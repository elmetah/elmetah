MPQ    �    h�  h                                                                                 ��B=[��5{��k>��IG29�~�H|1Qƞ���\x�u�h�
G�4R5u�}gp��7�j4)Tp�a܌�l�3���q;F,- ��M�(p|���л���� �LEy�ΪIT#P������l�6��*5�l��_	�r;RH��`ZlkOu�ckP�ő	���FDs1��)P�QU~S�9}���8�e޴�x"���V9�v���};�G16�I/Q�L���J�+�BW �,=��nҶ'eC���u�7���s�K
�~�(�x�6�S��og��'���	�h!��#RԌ\gev�"��&���ۊI�&�-h���E�c����g�g�J�5j�H��1i�7�:%�i��a-_d���VM�o �-�
�t�G|�(���֜:D�����h"M�!�+=�P���L̈́��='L���Z�f쳒���-"B�
_q�s%Ր]�J�NT<�c���קMf��ې}����l5r�
��ጰ]�1�{C�W�4�A(��L$T�㓟P<q+Pi>o����^^d�GI��ή���C���6�-@3�*�<�U}l?�᧦J�P�.q]5Ɵ�S&D���"�� !/ J����k	s�I��A~Ӆc �6�����^!]5#���w�y�Y@X(�2ih��W!����-AW�� �""XA^�c�x�+;Qc����~��!G��yN�C{&�!}�-�*;C/� V��U��!��b�Oa�1Ee����@H/�s��r�g�H�C�76�O#�Tr�F;)�S�
aC�E������1����[��7�V�Q�(�L�%o��i'3R�	RD��z���T0�eO�F��]��v�m))EzE��������tub��q�̄��Y�v�r��ZP�m���Ҿ��z�����G����	�f��t*C���E�G�=�����W���S汖���u�����1`M4�`�H�\n��� ����"���h�;�����lR+�\
�d���N���ؿL���HQ��(�ٓ.��h;/l("��><�&=�m�����B*�%U8��4%Qt��~぀��y5涛�XnYu�*�C3Y������"��6�����$�{���>|)��e��r�{LZ�����E�­c�g#�}	
%B �{,��YU��Q��+s	%"F�;%֬1��,ϫ�J��/�i����ixlxƨ�g\�,ł�O=�K��AgE2eX�n(�����;:<s&��ծr@�p�#�"�S΀12Fx)f�K|ա퍱ڭn�	0M�ʞ@_�юA
���9�P���?�p�ca�|瀷��
���F�\p�$�`],
K�����E��7ټyS�+x��	�)��#�;��Ip�>�p��Uj�>7ƴPG��+�(d�q�ŌuL'��jΏ7f�6�Ju�T����8#*���(�� ��P԰*g���F�$R`�yB�Π�A��l��U�W ���p��6���\ ?R���dM=��ŋlg��ٺr����[X���Hú����� ]q��p��l/=t�����������/ܦ�7bxL�K�/W��ᝣ���\�Ɇ�!(W�#5!%6�ѝ��<?M�F�ܗ�΋�}̐>��U��Mn5��H�d8D&<������Lj⫗_�~t[�:!��i�o����ӷ�-�+4�퀰ʕ�i4�6M@u�M�䰇jN�R�8äU3"s8A���t�� d1'K�o�i���a�b�2lVj�<ҋ�A�*�ܕ����y��������ww��V�?��M�\iB�=�~��-d`K�������{���ߘ���+cA��A��9�n�[��E.h���������+�coG�Q�������`��+O��Px%K��)X�Jf6V�R���)#�s�[?HR����c����а;���8D%�3�y�n���K#|�参�!Gy��)\�g���78�g('kp�i)��>�q��c!���".ow��<�0�]3��U�U����h�����n�8�����3���{�8�LO�n�g�pb����h��؋�*,��s�]����z$�w�_��eZ<�}��ӓ)�B�m�DȀ��|�Y��e~�]�������A���8r��O�Z8/?H���1��MXl�0��=�>��5��y��?�ON㳢�U�9���cs���i�x��EOBX�aT'\����ۡ��♃;w��W؎�V�J�O�yNP����>x�҉�D�Z�5��������
�;'�(z�r����ek06�q酻Fq}�E�0�	#,Fe{���y���qS�g�{�f՜"�ZQJ�c�-Ld��+(�_I�8~e�Xh�2|~���]^����zRKH���t,=��[��,�8��h�_o�1m�dsԄ�Q��YI+��kN��>h����')N�ǬZH�	�a����gZ�p��>_�#��]F+5�k�׺�*�n�f�q!s�43o�Tk��$��0�"�ܛ��K���)A�!�DC)U9P��xzZ�_�3��WLI�9��̟�H�Pi7Fpx��$O��"��~�>�xk����C<C����d\�����`u#����`���A�v�F�q��m�xw�//��y6d#���d ����1m����Y���66�x��!Ś`T�j�j�}Kpo���2��y�	E������'=���[Ƽת�r����I�OY&(K���[u|'���3)��yX�EP�����_ob��B���I�:�N�'׬���U�y>hn��dX32�+�]�?8��ڙ]�逊�
��Z{����#�'�DDߡ=���hTwYQ�~�s�$��S�y#�7f>�<�¹�u��Q������-��@BY~<��@�UB:��8�ڦͣ�-�v`�V2��,a�ܡ��#g�#�T��,��J�ѱ������:�m��eeb�b���)M��Iku:���v�����參��qa+1Y��{�n'N�T�
�,9��MZ~����q_}/K��,Ծo�b~͊^�E����kfe:�<�v���%JAjC(<{�4��>{����\�R[���9��C1���S���&$c����^IL!���g?��I��ܖ��X���GA�Y���z�B�:tN���	a.�-�S�CD�mF�����83ZOF�	
`�+����c����2��/�?ف�!�hƴ�h0��puo}�����K��n��I`&F�`���Y�"+	����T�����2zdM��釞{�)�) ����D�����W�_���{)
��Ɍ~��mӉ��I�U0\�\�o��'¥��zY�����pq�/�\e��ux�,t���i��Iz�Q���B0���jX@�,T7Y�r�$���|z(d����U�ϪN-�<��*=G�\����ַr*�y�]�C͡�\�=�fIP�EKL(%�����������n�m(Ɔ?`B�C_q��,0\N��;T�ibU<��ָj줧��'7�}��c�r��~���O]YN%{�X��«���(��*$��}�Z�qF��i��0��Y�^��E��I�1������^T���.�nG�׏�Ux�_�<�J�o�I+H5A�2S���jH�p� ���=P�k�`*I�$ A�?c�F�6/+��2�6!XC��Y�wR�Y[�A��Sh���W\o��^-<0Y�{��"�[�^��,1W�+��ec`]Ŝ�����q�C6��!�bAT�;�͔ʋQ��ˋ �䰛O'L1`�J�M�v@#?/R%�1{u;_��G���H�6��^�(�DA;d:���2��@� �s�)�2F�L4���i���rk?���#�G��o۷&'�8	mV���,���OP�2e��ۜ!���(o�`w��(l�ٜ���u�tj�l���G�1q%�	C]���?�f�� G�zUN��!jG�8��;s�`Tt�y��p�[�U�=������WhP�Zf���T��0���܈���M�lO`�\�&K˻���˿�H���4�ֿ�R��k�W���5�שKk��lNL]	��#X	�cet�ύ��/�$�����A��m@MZ��-�}%�8�4�x~�M�2��fy���y�An�mM*?C�Y���ܟ���Ց�
$t!��G�y�D�e���.�7Z�'��E�EXvc�|���u
��� �?Rt{��Yp��Q sQs��FZ����1������n�i��7��Q
x��Kg���m={jߜe]2 "�nC��x��;��sa��I���k���LS���1M2)�՚KW4o(�*�H�z	+��%�_�@A%��Դ:�Pl��?�J1��M�wg��/
rM�F�e���8�7K�an��I�������Y+3�~	2��S-#�aQ���R��g���kPL��7�5b����{(?���+Hu�T��zK���f���A�e����s��b��#e��÷\��Ȕ�������f�ٟ���T����@�r:���aW{	%�� 񦏌�l�� ^\� *�M��ņ��g+i�-�c��ͥ�fÕu���]l�p��l��0۞#3�C!�/���ߐ}���b���F��/����`#��	\T'��4>�^��%�4���(�?��N��� Φ�}G9���Bӈ!�5]��H��PDqSb�`ʑ��T��]'�r~��:�r4i
ӧ��+��7�Hڢ4D,Ӱ��/�����=�u�Qw?4�j	��S��U���s���&���$ _�y`խ�*�Mi{�ag7҃ВV���mR�A֨c�7ob�د�y�V�<4ڈ��w�����̚M��.�ݨ�B��j~��-��K^�7��wl�u�����V�c��CA"M9$([�Q�.��E�%���լ��6�oa2Q
-��;��`��$OH%���y�%�Ǆ���
VŚT7��#�.�[z^���;�^��U�;ִ�7�z��3[�%�Ӷ��k���z���bG4��)w�L�C��8�x�'��a���9�4�3jI�K.��ݖ�����30ⶕ����Z|�\���O��S�2�v���޶;����m�i�g<�Inν�G�SN��;����]%���u��w��� ��W�<��'��n���Wmi�Ā~:.|k���cg�x���6L���~K��`�r����UV�?�� ���T�h�elkR����3�y*�5N%@��(O��ݢ�ip�+�t�nR��K�� �E��XIYT��yÓ����F+��tλ������JY[6yI��dJ��?ѱ��rD�Q���F��p :����'p�z\'g�6Ce����L����Hs'�0��,����V�y��qΨ�Vn�fB{":��QE��+1�K���zk)��+�3}��m,t�e�]Yv*�>��R�%���=f��[ǀ�W�R�
+jSa��s�e�Q��I�mk) �>>.P�"M)IF����u9a�����p^�_�����>�5�w��q*�eif�?��C3Jm�k5p�͜"������K�M2)\�!���Cn!t7$�I�UtП��hWV�9��<�!�H�g�7�bw�A^��ӯ�.�r8>�2�}
X��C~�=	���9�-�#����'f�mve���� ��6�h��w�6/q/CQ�"�Z�P ̪gBm�[�'�����3H��q�����g�r	�	}�U����l����J����]����={�� ��C����|O�	��W����|��)�BZ紌�E�����_�p������~���%��j��T�U��|hi��d�l����Z4r�U����ϞE�Z=�����'S��\-�����T�#��YŻ�ZyLPҕt�V7�ͦ�ώU�݋�u]�������4-P�0@=�<_ëH���&�U@����v�^�2'UFa����@�ށ{�oie,J�稬�җk��w�m���r�b��'��kM�+kP 4�d��4��Y!�BU�a,�#Y](�{�߱N���
@#9��ר�;�h/�q4�-�׻��-o����%�yE������d:���vN�%��C�
{נ��d5����K�[|�]9��1m�S�Mt&_��`?,D4��_hIg�ͰI9D�b�XjǣG|�����`����u�N4�������SS&���'����v�3�B�F	�cB+��̄�A��{"���?���!�SA���@0��RBN�}����_���fH�&ax��L�j��E+D�<���G�����8�Ss�_g᤭����B�3������C_��,6>�����ϐH��D�U�q��W  o���`�����P�T�K;_j��edwx�l>t+�Y�M�/ˉ�̊���(���j�W��'_*7�����?8ї�dy����u?��6-9�� �G2��b;�������-���fۗ�s=MTlP���L��?���!�� ߑ����H�)�Fp2B4�wq�+P�G�Ǒ�����<�u�E"�þH�B�}��lay�rl�	��6]Ԋ�{��j��	�>�Q(��d$
 ��
�qa�i4^A�{��^��}&JI��s�i�}�K�h�yC���Y��P��sw�r��Us|���%J~���d�5�� Sܽ���3�6�' �����kn�I��At��c���6j�{�͎�!Sq��PG�w��Yv�C�(��hc��W����L�-7)�����"�^����U�+Ƕ
cQ��7������/��C�c(!������;� �)m�&m	���?)O�`�1{'���g@�;B/��n����+�����6���#�,;���@$�;�8��Fk���g{��B�D/A� <��Y��B��o6�'��	����p���{���e�M���W�l�f���{����,%۴lT�\uQ�!�g�+�u
���a<�$KR�c	����[z��<��r�G5w7���`�S�t ���K�ߐ�%=F�l��	@W�뺪m���2�������Y��R�Mj��`���\$��v�@��ݡË��񯕖� Ra�.�RQ�<'��dh��� EL�@���~}��g鍖BD/"AF�On�\[Hm��8��r�ø$�%�g�8�a4ۿ��ĥ����y+a �T2�nυA*�biY��z�JO]�N�A�އ�$��s��B܏��I�ߤe��6���Z�p˖٥0E�i*c�O�&�e��ԓt��I{�vQY��	Q�!�s� aF�!V[w1�k%�a�\�@�'i!��_K�x|�Tg�2�Ÿ8=v�����52��n^���m;���s� ��俼�f�)�`�YSDJq1h>$)e�K2�,c"��㑓	&�꧀g�_:��A@�F�/�PG�e?����Zfrl�n�f
-�F� �''��K҆�������/��+��z	M`_�Å#���8 ��tJ��ѡ���7<�;}I0��(��&�wu����uL&��i�mo�AT�Jz��=oz#���^pҘ���K���+�9�+����/$����9@��c,W�BF������)� ����[�	Ms��Ł�gt�غ�c��������pL��-4P]�e�pz#�l���Y{��.�B��1�Ӻ/��r�b����A�/��WC��Z)\Ϥ)��aUǙ��%lE���?
��RSM����}�����9����5�8IH�`ED̠���+ң�BqX�ME�~���:Wti,�LX�q���c�!4��1��Z����lNu�u����j��~�noPU
fCs��9�a��Q�� Z����Ћ�#�i0L�a�+܃�S�V��9mA�b�ߒh�����y�+�sb���w-͎�u�M�Fp�8��B>}!~#HH-ZU6K9���������v��V0c�5 A=��9���[��6.ް��������~o�&�Q%����w`�nO�P��I%���߂���BV���g\#�	s[����Z�YḚ̂Q�;��	RN�:r�36eQ�SԬ�m,�8�CG�I�)�3Z���u8��"'��\�����44���1�I�8.�7E�5��悁3k9앋��ld��,�s���n���-����ٚJ�dqyg�I1)֔G���0��m��F.�]��f�pTuwE����_�r~��yU��I��)]m$y�y�r|���\��ɓX���ĳ����;r���P��?����jc5ك|[l������״��5�z���1O��u�_�FoJ��`}��)���RE��#XmT���NG��ܛ�y�Q�fI�%�J��yDn m�ϴ��l9D�;��ٱ�* �џ� N�'˹�z���#�ea�S�'�[���)Y0�SS,��H�7y�*�qI���1�mfK"�:Q@�a��*�����S.i���b�����R=�]TA	���R���<=ᘷ[�`4������L�e�l#9sJfQ2�CI!��k��>yQ���j)D���b;G`ia*��]3p9�_.�ҽ�W�5���p�l*s|�f�-!i�+3%N4kpl��7��vI�Q\oKT�?)w��!��C����>RҮ7�P6����W�9ǆ�̕h�Hl�Q7�tj�ܷBԯO[�-Ώ>궀���|��CV7��ͱ�ԑ�����#f������S��|
��/���	�c�.wx�/,�PlN��$	 ��$R@�m-���1�6q���P��[Ő'��B��DǞ}�[���Ǌ#��y�(A�؄���*�2JY���y�1�O�����;|ԉ��z����E�����T�_%��������F��0-I��~��9�BU2�hd�Dd��ӡ���uP��и�˟~��[�Z��̉��O'�-��=s�͋TTm��4����x�l �och7})���}�u�Eē����7��-�3@8/i<]9���m2���	�Ї~��-�v���2�G8a�H&�Ty��2ՙ�1�,�kp��u�C��O��m�ع�nbd�M�	k+��=��X�wV�|���aGG>Y؉A{�p�N4�O
�V89;(�G��#�qOQ&%�ŀ�+mo�����{wEM��!�D:F֮v*%@~C���{K�<�tnI��EL�(�[7369�E�1�V�S��-&�ݾ����?<���o�g���I�8܌�XE�G���9��Y��0'�0NO�����k��sSa�)�E����3��y�3yK�9fb	 ��+���s�$�P��T�y {?O�!�^Ĵ�E%0�(�}GO}������8�G���!g0&|n4��F��[�+���L���ط�������@���=֡m�}���U�����_@�i�r���|��t�#1��J^�UC�
�R��of��a^���!���;�&%:�#�e�CWx��t_����;�JmA�Gp���$Q���Jj����"��7z���Ѳtd�W���0� r,-�aD���
G�a��$��B��o�|������;F=�a�PקHL��T�n�ҙ߃��wY��#4����B��q~���R�L	U���o<|�@� NO��m&k}�M
���r'�X�2�e]O�{�|L�q�=^(��$eaR�Ж�q|�i���Vg�^[��I���������Rx�W���D�����Un4u��m�J95��57��S����F[S��o8 �r���k:��I!ϡA�c�VQ6�1Q�h�n!N�$��TFw�CKY�h-죃�h>�Wҋ_����-2Bk�14M"S��^�P�'t�+��?c��n�ҏ����ԊC�2S!�3C7�;ԙ�C݆���Y���s���vO���1����Cԣ@�/ȃ��g���T�x�O�t�61d���;ڮ!��5Ѱ6�̬)dc&�����񆌳ɞ���L�"���=�"o�� 'd�Q	����7�|X��p�e 5���2��8?ҞZ���]��ۏ\(0Hnu����b@���oD�r��?s/��4X�q|ؾ��z��V���G���=S��f�t�F8�&=8���$=��K��EW��Г��1��&Z峒J���Mt�`��y\Ӱ�1L��~C�>����K�L�8R��I�M#f�8���u����LS������ى��pz���/}}؂
6��w[m6r���d���QB%&<8�ɢ46'��=�њiy�Nכ/�:n
�i*u��Y������Z�	p���$ő���������zO^e}�b�S/ZL���%�EN��c�B��a�4�N�L=���{]jCY�a:Q��s��XF�zA��g1}�Kϼ�U��KCi&w&��d�xW#g���S$4=q��R��2�[ny�nc7;�|�s�o����a����S���1�j�)��KR�����~S$	!̓����_�аA[�DԪ�P"(F?35�4��m�˷�`�
�_FG��l�#KUbӭ�X���x�����+��	hM�T�#��n�s��M������Y7����!4��]�(�00aXu�pmL�H�S�A�����Š��e�#�a���H`�q>�a�[�_�T��ٕFi�
��QoY��|~��3W1 6]�ܡ}�b� ���MW��|�gύ(��P�7������KCC�h�]B pupl@�����I�%��ӕ��7P�bIz]�<��/h���F��)��\JB�ز���ԍ%�����+?^L�����%�}=ꚛ�݁����5��nH�D'ϳ�ە�Fۉ��u�(�~%��:�ݫi ���*�,_á~�4:	���S�Ѓ��u�����bj���u�U�/s��e���Y� U������
iK=�a]@2����V�G�?>A�<���ܗN�y��2�V��\(wh����M��-�eB�L�~>]-���K��B���L���Ј����cr� AXJ�9�[f{�.��[71�+=�<Klox0Q@G��18�`�aO��ح!�u%��g�:H�{X�V���-��#g`[�ꚽ��q�T���B/;L��m��HJ3v��]��{	�����G�Л)����9�V8��''U�:� �/�o�������.��݌���~K3����&q%�������.i�:#�l���>��, ��H�_nag����o"f�I3���H���E][׆�k�w�U�ʖ���������$��d��m���t@s|!r���ɮMG�,]k�~�P�B�;r����K��?Y���%,zٞ\9la�9�Hp��f^5�𴭯Z�O_\��0���a:(�d���'0�)soE ��X�T8V6�	&�ے4��G�A�`C�J���y?-�Ȁ��o�ϱ#HD����-�e�w������*'&��z��Ķ>.Ze�����������Jg0��%,W�ћ6�y��q�=���Sf��"p�1Q;�J�>J+���Ή�&����V������4]O,���a�R|��#�p=\�u[}`������9�I`�T~��s��QM�I��qk�U&>���X��)?(xǽ��aE�+�؍�pl�_i���.��5��p�ː*.��f<���i3 O,k�����I{���ܬR�K�)�~�!|�;C��*�eT�IF�KƟD�W}Ϧ9�j���HG��7��Q�w1�P������>�W�sO-��`C�t��s�@��	,��f�#!L�{i�cQ��)��'fq�BN��^$wӶ1/����y�Pm� �:2��^mȰ��z#K��>)ک&r�������%�}�&���ˌ"�8�:�-�3�u�Scd�yj�m���CD\�z��Oj0�Y���3.�|�������*ULE!�`��ï_��!�s�4����������V�t3aU�Mh_ di?��\5���V�Kxb�z-+���eZL����6'	Қ��l/�貖T�B�Y|�Ѓ����j37wLV�E�����uS��[���r6�-���@3�x<�3�������ϴ�K(��u�'v��2]Zaʮ2��3�T���m,@W�bb��~�X��R�m�	^v�bk��(�M@k�%�x�GAPs-�҃�ab�YS�{x!�NoY�
v��9���^�����qj�f�P���|o4���[:�Ez߮�|z:�hvEVz%�'�C��x{�{������]�m$	[�9���1c��S���&�ʾ�H�:d]���gp�@I7����GX a2G�c���^Lx��y��?NjT-�z�t��S�횵�Lr�����P�34tUT��	{�|+�ŏ�B�]����}m����z?
=!�O�w�0����`�}U#����q���(�ܥ&����B �6ԝ+������b�����Cm~����A��9�U�ָ����G�ɵ&_���Ǥ��h���y�������U�T��MJ�o�?~��@��~z�a��/%�he�0,x�L�t�	h��IN�e/���u��٩�6�j)����v7j$��Uz��!5dod��xr�[͙-o$]��<G�67�����M��D�ԍ@���=���P҈�L9��)������??��順�2�Bj��qyc�A~���K��L9<��7���,�9��*$}����r��k�M1�]�ch{����C�	t��(�C�$�⌓�Cq�``i*ͦ�1�^J���gI��C��L�����|��ᐆ��ݨ�/Uij�ME%J������5�US�������l ���N�3k��I<�Aj�3cl$6��z���!I-���w�BY�X��w�h~�WJ:�Q7--{�ό�7"'�^�+����+}�c�[��m������	Cg!"!�����);�R�~�T�\������[�OM4J1�i
ľ�,@��/c��o���ا�sg�/�*6L ���p�;�N�vg��1_ݬ�h��r��iL�����#�q��r��8�Yo��'�	�L.�f��W�aq~e�<���-�"�W�Y �.�����jlLkSu�l�]��+�R�b���Z���Y���L7��)�z&�h��t^G뷶����ҙCt݋�����=|8C����Wy����O
��;9�m[���"pM�'�`�$�\�ك������\ço��%R�ټ�H=�ii��ѹ��jL��ȴ,6���E�����=/��j�������m�4��xvj�.��%�0�8�Q�4��]�~����d�y!\:�
��nE�*�Y�Le� ����m��$�|�o���*I���ex�j?1;Zbv��9EɐWc�Uӛ�`x���&�Ps{~�Y��rQ��
su\�F�����1x�����iA���U��x2�wgHN��/�=l�;߭ &2Q?�n�L���L;��ss�����\9����S��T1��p)	��K�x�6O�5-	ḧ6�^_�oAv���%*�P��6?n����2h�Ƿ$@6
�M�F!%4�ҝɿ�K�T�SP��#'��+db?	�Z���#cAu��v�o8��m+]�"7�w�� ��X�(Л��3u�� �k�n��'���$X��S�@���z�#3ƅ�A�}���A
�7�op������ΌKt�C���{�uW�̽�����Zb�� �A����M�%y�w4�g*oX�^];�R,��x�H�&Z����o]ݸ�pp��l��g�ϊB�d����	�pv¦rM�b���7p/�6���h{�D.b\��|؍��|%������?���Ȏ�����}��Q�a��9��5.lH���D������aR��8�~���~`�:���i�=9���"z��+84���x�^�U����$u��P~�j:Q;����U s��A��Ҹ��L P�q�V�[�ifN�a�tԃ���VV8I>fgA�69�H��	~[y��D�R��k˘w�A�ի!	M˰g��u�B�<�~Y��-P�K�`�}��粏��[�gU�c-EAsp9��[A@�.TQ����f�����o3Q[1䬘&`f��O�𭼑z%�"Ǖ-e6��V3���?#B�[+a��P2��O�|�fR;�s�Tr0?�3��XZ�G·>�v����Gew�)��d8ik�'W�o�շ��*�D=B��^.��3�.�����3�Gӕ�ﵨ��H�m/^�%	񤎷������g�J��2��Z��gM� �EO=����U�t1��h�]�+?�f_w�<��Q���i�o���ɰ�cm:�
�o�/||�%�����b�����YvK�}J�rQ�o�FpL?�$d��#ٹ\�l���膻��*5s5�c���O��\��d��|%��ݷ�jE=�dL E���X%�T����$���h��o�ܻ��'J*>�y:H#?��*}u�>ΞD��M��������P^�����'�lz�ʶY�eW."�ݤ�2�`D��0�t,��ղy+9�q?����kIf��K"M�Q6��X�|��ˑ�$ԇ��{y����L�]J7��O��R7_*�>im=י�[X�|��F��1�[u�Cs���Qhk�I2�k� >�@���):�C��F�xTa`?]�S4�p��_�(����5�[��&|D*�	�f+j�_��3�o�k�Ĝ�m���e�iKʒ�)��#!���C�qg%�*��twFK��8W8<t9�nűW�H"l�72�,��U
�I����K> u���!jf8C��s��g�ʡ3�>��#��c�Ug��n�x���b��ݽ��Y��w.y/��8��Ѥ��� ]���kmc�U�uQA��+��d�_"Mņn����-��%}��S�����}����f�N>���a4�bG:ƨ<X���V�u�O�s�F �N��|G���L��e�<E��c��R_�[Z�.�z�!	Ν&6t������SUh�GhZjd�����[���d��W<�U�@���5Z�މ���'d�bߍ����`TcCU�����9t��e#`7�;ފ �z�.��u��6�R˭��-!x`@.�D<N̫A;��'���_�P��vL`�2���a�4�
y�����!�,�bF�=�	���*���m�Z��cCb�愞C�M~�k������I
� j�)�s	Aa}��Yά�{S�qN�E�
%9��׹�􏙄�q���=���\oo���{Eu���k�:��v`
�%6_BC��{�}Pݪ�������@F[�b�9�c�1�;PS^c�&���1�$5���p�hg+�IRw܂jX���G-��o�	_���c�q�N��{���O�S�`�{�����+�/�3�o�	�-�+q���}�C�Z°�x��/��?��!'���0fZ�}�����[Ǘ�{,��&���ս����+��K�T�D��6���3�9����b����)?��c����Ŀ�_�c�g<K�u,�j�������Uy���Ho��@���u[��;���X �ee5=�x��t�J�Ԅ����=�ۮ�2�q�]j�^�@�7��(�!����d����S�ϖH[-
N��AIGC,뚓�%�#�ԅe L���U�H(G=ݥP͉6L���������b�mF�ٿ����!BfQqt/c��R��V���*<r>[��/��t3��M}�[�r|�r�C�h��]E {����~��;(٥;$���F}q�Ĩi������^��?N�*I�%f�z���|u�������av�ZK��Cb4Ud���<�J��Q��S�5-��Sm�����.�� �ؔ��'k�W�IW�cA�}cG�F6����!D�ǿa�Hw>�Y�h�왊�h� $WH(����7-(�m���"ɪ�^
'�+X�YcE���R��y�@?�C"0�!��-:�;�+|���������חP*RO��1�:��9�@�g,/>b���U��b��.m_��"6g�\�R�K@�;P�o��ݰ,�i�ߌ��14��D�|� �\��^ ��X/�3#-oG5['�7�	������m2B<��eVd���H�}��Ɔ̫V�.�E���~u"�W�X�,��������u#���� �'��`�z��r��%�GF�6���A����t�����(U�AM�=�R���W�}~�FA#�8���=��H�j�o�M;�=`�k�\5 ˧ܩ:��4Â㓖�\�R2��C'pM��ו~�
��LI��ȏ�z�O.����y�/3V���%}���m,�S�I�i�%\ET8���4�U�9؁Oey��I��h�n��V*��Y׿��[f���/�H$	�2�Jz|�e����es�N�.�Z�
b�*��EDT�cf�d���/��u�/k�3�{ӱ�Yܗ�Q�`sP:�FF��,Y]1s���r!(�q�fi\�����:x�g���ŉ[:=g&���>2��n���d��;��	sM�|յ#��W���q1�Suh�1�"�)��QK���ڴ6�	Z���&_kp1A�)�Ԡd�P�7?����j@}c�_�?�
^8kF<g���W����K��������P�@�e+�	����W#>!���Q%�E������'L7mx�1��xtO(�&5��uSK)�f�����ⷰ����ͻM��ΰ�#Q$��/ZĘ�$��ј��^�ً����fA��GC��c��v��W�wY��4��X�J �͙���MDS�r��g�ph��K�m�������
�]x)pkj l��$ۊB��?ױ���KX���jb㈑2\�/�_爫��_�z\@ݨ�h���J�%=3W���w?1�\��.}3՛<-�t.�5ɨAH��KD�H��Lm*�|���kt�ލ{~�R�:(�i��a]�*�������40f��SO9��BH�=@�u��\��jj������~U{"@sΫ'�"�� Kb��ι���i�xaS�y��V��٬�A�P�ߣח��y�(�FZ�wޫ	�F��Mƕ�I�IBoL^~t�-˴�K��ヸ�������ȷ���c襍A��9�9�[%	.���&T�����o�7>Qv�~�'0`Aa*O4�[�W�W%�h���2I�DV1��#j�#Z�[f��돈�J�o���Y;��n���U�3Ƕ4����RΪ�q��I{�G >�)�r�/s�8D�B'����p��%�����j�z@�.�r�݂�j�w�O3���\����bE���������b�nz�ޢ�q�<��Uȥg�~�Z�2X�?�O���5]����a�wVD������ȵ�����;�m�b�jƨ|׶�덚�����"�>�4^���-7r��Az?�E��0��|�lW 2�aNm�e#�5�;
���OM����Eޗ0��ZLg�E���EeEV��XYQT�s�C̡_ޙ������+�J��Wy56~���&߱Y�=Dw���|5ԯ��?�Tǅ�K�'�u�zH:��t�e�}+���$�m�����0��>,+�y�vyF��q�Rk��UOf�"��Q1W���襧7a���3������͇Y-T�#�c]Eb��VTR�4��Y�1=R�U[3���C ��o��Vk�4��s{(AQ���I��&k�v>*�����)5��s|�da{�����?p�w6_�y�da�5��iׁ� *��fF����i3��,k!!����	N�b�K��)�н!rC�Cp]t`���nA<,��o=W��%9�X��?H�77mk����t��`�^��>;���i3AMCOC���&��Y״���#�q�P�Y��S��V��xM��TCw�[-/]&���F^� 8J=��m����p��G9�k�8��B���-��A}R,y���s������W"�i���I��=5���嵂y�i�p}�O � �V�iZ�|����z��砝�EW�����_6�R��9��<�#���{�n���U{�hU�d����ޕ��d۩AW��0�F�1Z�Z����<y'�z*�H,��a�Tލ���l}�F����`3F7-K����$�I�uI�������6-�_�@)`�<n�O���%�+*c�A��+��v�K^2��a����e�d��;��I,6���x���p� �
m�˚,�mb���^�(M�-k�WX�}r��/�N �.0a��~YIn�{.�N�Q.
���9�������T6@q����I��s�o��d͑�Epc��2}$:w,�v{ޥ%��FCo8�{����EKV����#}�[h*�9#g1YޅS9U�&K����R0���E^g�XaIm!��W�X�z�Ghޕ�
W����A~aOqN�^��p;�*U�STy����͢Ċ��3�%N���	q�g+L���������T�s�ԇ�y�?��!B@~�mQ0A�|.��}�>���8�X���R��&���83f��E�+0]���^�ȕ	��q3�������g`�.�8�&\J���z_Q�a"����	�����c��l�U��CowHc�L`���ĭ6;˷�+VS�e�i�xĬ@tphM�E���Y���ۉ�뮬5j_�ϙ˳7 ٶ��V����dee��.5����p-�	��2G�A��N~��>kC��ە���ۃ�u=�J�PȪ�L�&�����0mI��l����X�2uDB�>�qo��4d�}-%���D<���������>�>}�K�'rXuޮ�C�]��{e ӳ�fm��(�'�$vE����q�HYi ������^�q`��eI�r��x�7���?}E��<��(����U_(�T�Jj�$�Э�5�p�SH1j�����޺ ���\Zkk�Ir>qA`f�c"޹6V���99!?i㿼<�w�-\Y�[���hϣW�&L���Z-#M��B��"�N�^%B���C+3.?c=N_ţ�����ԛ�C�^�!���9;e$���ʒ����㗫�OÇ1�+HĴ�"@jp/y�V�8\��<����7��`�6���叱�&�8;�̈́��*��'�r�:ѺW�������+y�V�5�����.��o���'��	��s�\���w�
e����اH�ϫ2�H��nM� ���\u��o�S�:��_���d�ѐ�7�Owg�оG��z\�t����G�x6�n�?�`�tjW��;�|��=�)z����W/������S�"��^e�#ݚ�>�0M���`��X\�Fj�b!��U�%��}�]߈���yR�v��>Y��,t�P4�%11L�^,�jZ����{m���v'/��;Mc���m�,�.�8ä��%�y_8��#4G����ہ"Y�y���en�&*F!wY�R@��Xԯ:ə�J�L$�.��%"R��o{�KsenR�KsZ}ӱ�Ef�E�75cA�e��[��HX;|�{�2Y�b�Q��s+8�F�F|�9�1n{h�͔�,�niw9��Kq�x�Zg����$�=b��c=2���n�nI�P\;\ps�}��P���R-����cS0]�1Ԯ])��MK��O���OX�	kw��x�_&��A��o��8P��G?�%��_^Ǔ��^�
C'FW����I�K��ߥ���6��1	+�m	��+��#!s�$M���-ό���7(���i���(����u�*�a���YH�r\Q�t�6����#�5څʒ�����r������l��[���gd�dƊy��q��WB�92��--���^ ay1�G�EM�"��m�cg��X���?���1�nnQ����=`]��pf�lQ'��E����;u�&Z���6b��-�@/y��C��z�;\�ڀ�CU�ǅ�%؂͝�7�?o�8�>J(�-�(}�c$��:ӯ��5dc�H�ذD8ó�
��R�.�U����~ְV:��#i�φ�y�]
t��o4�D$�.���˫��Чu�E���j�N���G�U�K�sZv
�M����� F�k'݋��ei�Шa�=��T�V��t�A���������py,C�����!	Jw6p�� M��O爛�B*|%~�$�-F�5K�Sw��!��������Ժc�`�A� �9v�[�)Z.�qt�,�����Mڵo�}�Q�ޔ䢹`�Oo=��%����KX��jVL��U�#���[�������E�^��.;}?���?&�u3����Y���/�l����G�$b)�k ���8�X'�YS�?H� z���iS�5��.C�����R2�3W�
��Lߨ����#�S_���ږ���eU���f���e�P%g{�5s�ڔ���*u��2#�],5x�\4�w�kY���[�fеeK�ӵc�4|mpb|�e��|2	��H8��������Z�f1��03r�r��<̃?j���VF���Cl�c��<�נ1�5U����Op�1�a�E޲[���"� ���^>E��X��TIp��:���,u�et�Ҭ��P�J`u�y0*`��Ϡ��t�$D�Ǐ�W��b�k/��5W'7��z������eM��BH���zob0�g�,h)�4u>yaǖq5���_ef7\�"A�Q,׮�Oh��˺����!�z�P��}N�ۧ]@���R�*��t��=�x[ �~{��
��Q�4�λs6�Q�{�IIckpF>e���)��)0k���|FLpPa�%��I�p�-�_�o����5���ܲ�*_fa&U�+3�5k\�ͣ����rܽ��K@�)�)�!��CKiQ��S�2�<~i�U�"W�u�93ף́��Hعc7����H^I ����L�>V���&��CB�&�D ~��1���#R4k0j[��	.�����p����O�lw�]�/t1آ٤�� ;>M�m���k�f}��C�S���|5�㮐00 }}����A�3,x�k�bل�C�ľ��C��������k�O{Z��0� �|	:��U�!��q:E�X��З_�����S�WK���ϻINQ�%q�U�A�hP~Zdzk�Ӎ㳱� ���v4��<�lD�Z�Љ���'���|�9�TY�Р&���SJ�[c�7�zN�v���d�Du�[�����#׹-Wgn@$[<����DT�F�f���q��$v�V�2.Rqa�����c��5%���E,��̨�2_�/�*���m�\3��bP>�y+AMt�Kk��I�)ʻ�� '[ *���v�a��9Y�O�{	��N ~�
Ge�9�$�o�0�q���v�N[�o����,6�EkU 獮�:2��v���%,.�CJ�&{7�4���J��yz�~��[#�9(m1ԠGSg�&�R7�g�+��&�sg��'I���xe�X�7qG�6}�����䞿�0�MpN�q��x�SM�浱L7�����刪3e���&�	�T�+'�#��kl����n����z?;!]�!��?00`/il }&�����Ɨ���"�&膽ճlS�ǮJ+k�ڍ�������T�6����)<��B1Q�ibL������3�_�V݅D�9�N�`��l,�6�U��	�>)wo�����j�ĵ��PS˒G��bek�;x���t�Gp� J^��5��3F�d�Ԯ��@j��Q�vl7{�[��Jd�}�	����-@,����G�vs�	_��Yc��[�ˣen�۾�=TؤP��LJ���Zy��KP8�c�|��ˌ�mF�B;7[qj'�R��8$�W�<hA&������|���}���(�or�=����];�X{@l���M�E� (���$�&}��	q��qi�����^�cu�I���0����O� Ϲ��Ȑ���%��y�UZT��^��J% ��'�5#.�S#��2���=� ���_��k&�jI��FA�nUc��|6����Գ�!:7ۿ��w�fY����xh�fqW�D��"�u-�`ϝU�"?�^@}�.�+��cxw��>K��b�����C��g!:�#�;@=�/���-�����+�'.O~a-1=S�/�@Eσ/���ӂ��6�����`ż6��L�
1���;���G�ʰ"N���5�������r�}�p��ԊY����)#�o�36'P7	c���ͳ�$�1�e�ݽ�+3b!Ҋ�"p�
�U��[�5�uX�_�N%�<E����ѫS���"���'X��,2z��n���/G����)��#�{t�`�𒔲߷/�=Mҹ��u.W��v��n&�ni��=��M{�ygMq�`�Y\�}�S�pb��*
s�8�M�8k�Rh�&�9������;�@�0L?6�E!Է�R=Wq�}��/�"���M��V�m"<ǋ	l8��F�%��8��14�^����=�y�Dl���nn��*���Y�H�kү�&Z�e�$��� �w��2Z��9*eiЫP��Z8�e�`fE:;�cNכMk������a��{Iy4YNMQj1sV�F��b:�1i���(({��i����
\xÆ�g�gJſ!=]�}߾��2�|�n�/Z5V;7��s�l���y�Mׄ�'�S�q�1�Zp)z�Ky�����	��G��_��A�7�Ԗ9*P��h?�_��y�Yd�5�^
�mFrK����ZZ�<KA��$�d���ؼ���+�#e	�A���5#�@j�_h��{�kḏ�n2�7����T�n�(a��M13u�#�\1�����-(�Qͱz��|x#�fe눘�`{�ͣ�G&����&فL4�v�7�=���˨�l6�W����G�HF��N� <E����MzQ�h�3g;�(��C�������÷^��T��]�%pa�+l���� w����}�|��#}b���(l�/Ԝ����ɕ\�\6��"���n�%s���|��?ʕ���W��Hz�})�?�������\5�=uH��D�*��~O��ɉ��#���~/_:^4<i�ȧ�*�.���4&C��	˞�5]�s��u�	xa��jk�$��ͻUq�s5����/X�n A`������i�A!aI҃�/�wV�E��A��K�Y'R�:l�yG�x�a��׊wT���|��M�����b/B���~�k-��K���.׮�h���E�x��c^;�A�R|9�A[�N�.2�ǕW�W/����od�\Q��r�z�`���O�/��ə%�TǦ�1g[:Vg�|a�#�/u[܃U�!��@J�wC�;8���Ͳ��F3}�;���g�I���
G�+�)J��%��8�}'FӅ����a��U0���CW.,�6�x���-��3��d��+x�̦R�~��X��J��X�0c�i��Q���K��g^�����";�5}tG��m0I]����W|Pw��ʂ�����cӐ�OPL�m�ɀ`��|�{���s�b|��B���.T�r"��7�i?Ŝ(��v�
�lM����*��_j5�@��>{O˽\����ͦ��P���^����E�F�X� vT�c1���B�G�(��mx�����L��J�@�y+i�4:�[�����SDm��2���QlX!���?'��_z�2���ie�|��n�[��HQ0�<H,��F��t
y|��q��t�x��fr��"�Q'w����V��� ���U����|�YS�];i�`�Rh@���p=H�f[�����/��y�L����s�IXQ�3�I��kKA�>�s#��
�)+l��)��a��!���/p�$_U|����B5�_��7��*έf|�^�L3l��k�9��>���(��l/K��)���!h\YC&���B�ҵ�e7�����WiB59N;W���H���7�w��W����,�D�>q�_Yi�0C}��߄m��)�O�O#%K�Q�O��	K�ǃ�����JkRw?�)/���ǉ�<ϗ �وy �m4�6�f�L���Yڕ<en���Hg��k�V}�W��Q�����&?'ٟϘ�?���p
�Y�-���ױf��O���E���|����0w��fGE�Խ�ڿ�_�f��_M��r����o�$���`p$U9(,hK8�d�dD�H���� �7�R��(#��N]Z�F���&�'u��߾kI�T��TԂ��{ �����ې�V��7��6�1��~u?1&��v�^�p-�	@v<$]�r
ǉa2�7ꬣ���v��2��a����	8�@�s��],,E��2�j�X�V��m���tCb���~aM�YvkrCˣdn�#����{%ݗa�=Y?Q�{�$cN[ʜ
�8-9�]����n����q��:��k�)7�o %'��t�Efg~����:�:v��q%�œC%&�{rD��{~���V|��U�[��9C�1O��S&�����v&D7��t�g\^I�����X��Gޮ��@68�Wy���j�N���f��D�S�:��L7)��)%�@��3 W���K	g+���.���+c��i��@�z?�K
!xvʹcNQ0�=r��}�e	��wp������&�.�l�7�+����%�:���l��N�j-)�D��ᆨ#e֤4�\i����?_ ��Z��TY��ی\jK��q�sUJ�u�9^co-�H���7�7/�����m�r̽�e#qx��jt&G��4��w�����?��"��j����	A�7���A"/�9�d[���Ԙ�Gz�-�n1�壙GT�G��_�t{م���@�5��z/=P�L~L�?��fS/��T�jQ��7FB�OqeSs�kg��:��&E�<��͸gr��%��tx9}����xrΘa��Ջ]���{��/U!��(ʋO$,(8�w6"q��i+���9b^6v~`DI�l�狱쟭<��~�sJ����C@�P�UU�V���J�B7��5��S�*ߋm����U �����@�k�`�I�(�AV��c�-�6��j�oN�!5%��rwwo�YYX�
�8h�I@W��.����-����-�"���^[ؒ���+�)�c��9�ق����0�Q�DCS�!UR4���;v�jB��Ȳ4����aU<O9[1n�Ī:I@ �g/�C�n�0�P��?��J`6��`��[܌_;����mu�3����� ��	�[���f�d� Ϣ)%��$�OoX��'��	*UY�RYÐp�ge'��ݸY�<:�E�V�(��O*����W��u�v'�I^넗JN�N�����E��bP���1z�=a���mGW����=��>�ItwS�mz�����=���QW�/�w5�ܕ�B�����M6~`} \F3Q�ؤ\���z����7�s"R���42^o��ƴ'�[��L�-l� � ��`[�x�/D�����;����m�~���G��%-C>8���4�I�j�O�X��y��v��n1�@*|�NY���l����^���$z������큄�edn$��+Z��}�{�-E�^�c�ป�Y�U6t�	��l�{�Y-Y�Q}ثsᓠF���Z�1dòσ۔���ji�9�A�.x�o�g4l��Z�h=Xö��2=&�n �9�; �s�{�Ն�t�H����S���1
'�)�a�KTLP��.څ�	u&���~_�O�A��4�ԧPiy�?Z���;F�Tgз��V
��F��y����5S�K|`��.���7�Q&+P��	���uW#π������:�᳅���7�:`:���(<���wu$�W�Џ�h��["���,A0�_�#�>� d����P�(�e� �����]��Qɺ�x�芯���g��W������cƄ�tk 1��\�M���c�_g�4ٺJ�����e�d�
Ò����!]Iߺp\��l ]ۻ)��5�� �ܽ��^��bP�#$�//TP�3�ɰV�\�55������%��wm?%x������c_v}�T'�͔��%�H5�8�H�TD��}7���҈�$�ݫo�~L��:��Li���n���q~�X�4�af��)�A�E�R�u��/�K�j&�e�tU���s�����>�� <�d�G^�i���aĆV�
�VBu��@}A�^
ߴ�ߗ�PybZ��r��ƻw�����M�(�ZG�B�;�~�Ҿ-<4~K[g΃i���S����v���@c6@Aߤ�9l�[���.@��b}m�2�/�oiRQ�8�Z`�зO��(�%���6"l�V�0��#�ʒ[z&��ho�;�1���Y;�Vy��-Y$3X()F<#�#��b���ZM�GQRp)4H���WR8�n�'CR�AF{�h��e���.G�r���Jo3�䒕-*i��xc�ٴ��X����Z�a�S����g�F?/g�Ӡ�����#��u�8��]�]b��R�wgz�=p��׵[��k}:���m��΀[�{|����9�5����7����W�i�'r���2�+? Z*�����%�(l�J���1��O5�ϭ��O&���s������W�����P�E'��X��2T�v�ð_t�b��[�������J�,�y&�h�x�䴱��D�p��G���"����iA'�Q�zy�Ƕ�ʱeC,ЃI`_�Å�ҷ0�1�,�d����y�նq+�˓S��f�F�"w?�Q"7���N�hb�7�*l�0��
~����X]6�����>R#vꎪ]0=�![�?Γ����@|\G�E��s�
�Q��I�k&�6>���_xw)&�KǄ�F��\a̋s�?�p[��_�-7�5��5�K�גiu*դ�f�b�K�43G3Vk��V��[����o�scK�Y�)<=!�C�{
��Poe2b��T�W$/�9i�r�w��H���7�#�~q���q?���>�q��ګ���5C��*�z	���Ak����#�f����$*�i��N�ʪI��EN�w��/�o:��� ��&��m�52�aI��X!��PU/�"�r|�d���ܤ}#��z�Ҍ�<#���oٺ��Ѻ���ξƔ�G�J�2�a�vO1�� A��R|��h�pu�QzE(p����	_GU��=�՝�[��u^�gU�.�hFd0~��M���������w���x�ZS������'���y;�oV�TO-�V�w��M\��o�Q#�7>9?��i�ƚ�_u�&>����˙7\-��\@��<�Y�-�}�|�Ł�*���,�v8��2d��a��V�vα���%�,�^,����u��&����m��X=e�b�����Mj0�kM�ܣ�l�N���>�@Ń_dRa�(Y�rv{�u�N�6b
},�9�Ċ�%m��Iq�'�/>�3�o[�F�bӣEa�X�Cq�:��hv�t%"}�C ��{����H���S��4�;[�A�9^ 1ʅoS���&�L��m!���;�g!I�߼�n�-Xg�GG���z���R����:N�݆��G���S�ݽ��A��Ň0ě�83�2���	��2+�#�i�e����d�1����?���!�A���|~0�;E߾�}\F���k6�i�}ꃿ&�rթ?��}��+�I:��1���rx�
�}%� �_'��m������������',_b�:SO��o��V�#EJ����<U�Y�4��o�Ż�}	�R�0�y�'�H@���e��>x���t�f�v?����Y�)q��B7�]��j0}}�,71X����F�Tc�d��X��jςu�-vт��YG�A|���֏� �Q.����4��=�S�P���L �T�аΙ�v.�Y�7�EW���H%Bq��q`�[7YǮq��AS�<^ġ�Bsѧ`��}���ޕAr�ZI���k]1��{����j|9{��(�m$�Iӓ2�!q��i����x�^q�{���I�����T�h/�6M���ɐͽ F��ݯ47UP$X�Z�J��v�!|B5	wS��የ,W�sm� �$Y��tk�N�I��IA�߽c���6E9�
	Y!03_��D�w*8�Y3���h`LW4�M�X��-xD�S&M"���^vS�	�,+��Oc�)��t����ԬdC��!p�� ;�������c�����p���
O�t�18�A�%�N@��/*�w�	0���է�� ����6���� �_�;�;<}�}?��8u�K^�0d�$�s�h�+A#�J�X��ab���o���'�b	EgȜ�X����(Rde�Bxݳ���6�� �8੽ ��۱���k@u��ǈDč��o=�	w���i����듽���x�z-�K��)�G�	7���R�Yyt}���H�P�-�E=�����M�W@��2������r���L���M���`x�T\���˓e����� ����H���/R�R&�/���@ׁ���v�gL5E.���;��L���s-�/��H�l�.�5�mᡋ��g�U�%��8��!4X3T�%���s7>y�?�Q�nl��*��Y�ˋ��kB���;	$����ٳ�Q�� e_,ydZ������.E0��cғ
��g�������{���YH�Q�f2s���F22���i1_��ޮN�]�^i�����-xyx�go����I�=S�+�t�!2��1ngP^.;�Ӄs9�8�!���C����Sa��1%�)p��K/�� I� }c	*���G_W/dA��cԌ��PD��?����2�O�ط�|o
J#4F����w��jK�c�Z���ZQ���s+��	
|��VD#��H���9���pᮛu$��7Y�D:�U�d"�(����wu�A��R�ߏj�S��=7aͧ'm�:ț#=)O������B��ڌ�3��V=�w�"�,*�γx��J���bJWS<c ��~��D�c �<�����M�,�^>�g�i�}u��@��d��m�?�ʓo]��pW�'lb��vaY��;�1ӷͦ�Fb�5��/�+6�t�5��pn\,���;�6��%�1��r��?�z��o���~d�}�ڛ�L��`;�55S	H��DI>�8���0��y��JYl~���:�Ui���"+���ɡ 3~4����D�|����B�u����j�J�+:�Ug��s�@���"�c� 7�48�ǋإi��a?[u��n�V}T�E_A��$��M��U?y}�����wʔ\ղ�xM�i��KB[˓~�Y-��tK6!��������C�.�c�PA��9�O�[��m.{���;�-��^�@o��Q╇�[O`��1O �R�Î<%���\��ݜ�V�[��#�� [R�k�WFW�6�-��;�����33�E�]�¾0O�]Q��(�G��)Of�9<8��'~~���h����f�&.b���n̶��3���H���jФ4����V�+��N�����ގ͕���F�A��g0�F������+��J5���]����MlSw¡:���c/e׵���F:U��6mA!��VR�|C���y�C�P�G��w�=㶤�rXr�-��?{7����M�@=wlC�3��٨�Q�5&RV���ZO��2���]���FF������jBE�g	X�hTZ�o�k�I�}w�����c�Ύ�|tJ18�y!GG�ֹ��/��s�Dc�����c��j�Wox�ݳ�'H�Pz4MA��be����$S�Y]�K��0�FB,y<��eԮy�q����.=f���"�yQ��`��#��R���������E.v叢�]1N����R�˄��j=>̧[��*�/M��۞�B����sg��Q��I~ۡk�V>�
��^)!���=}S)a�n���TPp6R_��x�Ѓ"5�W�����*���f�0��O{3"�nk҇�t�����H�θVKq�)4��!^�0C�L�L����=�-J�f5W�;�9�c���ܗHi��7YtÕ���gk��RJTi>� ��U���]C�J����y��e#�<�x6�E�?�ֵE�����@QRw�$&/I%)rB�2�e ���&�mj��\����2��]�r��Ϲ�?y}��f}���uc��D�8���<��%[�5:��,�������G��\MTO��g�����2�|z���戧献}E�+�����_�c����W�K������9����~UoU�hA�d��*Ӿ�f�2�Ʃ-��˜濞ÑZ�I�����'+LK�4+���=NT����1A�2�H$��L��7��g���5Ƶ��u5<�}n��ԗ{-(>h@E<ڱݫ��x��^!�-������vs82�iya����ѳ����<�G*G,"|��#(�������m����ub�1�ʄ�M�&�k(�~����T����1|<��a\Y5�{���N���
@K9�K�׀s+�@=�q����\��N�o�3:��Q
E\���:c_{v�n�%�T�CۓE{�h2ݱ1���p�쏮y[T��9y_�1E��S�\&7�d�8d��L�7#ug��SI�	J��M`XB.aGT�k�v�u�b��0MN��\]a��S��'��l������3���ƛ	]�N+�����v��an��_CI��Z�?l�!�,=�Y˷0�Y���}�F5������>��&9�	�$�#�X�(+.x�[����Q��e��� ��z���|Qa�,�����p���t_���d��������V i'���U����/(�o��.�8��m)���_��#
�B�ue<\�x��tܥ��1j��\���60��������j˔'��6�7��o�m��o�idQ�x���Ͻ�-T���/qG
��:� ֪�̉���nQ�o��=%AhP�nEL[h껋|���5��F'� ͉�z�B�q[`c"��iȉ�\�<<ٵ���ϧ� ���}�.�9��rD<����]���{�o=���%�W(�o)$�N���q9�,i��S�^��lUsI��V�Aj��#��Q<�iϜ���-����J94UK���o�&JV(چ<V5�&�S�������� ԇ��p��kW\�IޒwALH�c���6B�[���!+a�(2�w��AYN��� �}h;o.Wo_����-q�Ϯ>8"p^���ɒ+��uc)�d��t��N��P#C�Yr!�>G�ii;�G�J���ɮ��m��O���1S0%ĠC�@�ڟ/e>�����䂧�+Y���S6�H��{o��
G;w�b�13�]n��"1C�:�?4���~��J��_����so�o'�=�	`�ߜHΧy��c�e]
�ݮ�DQ,һ��S��{�7یk��6�u)�?�?J�M����g����;��n8��3O�z�X.��z�Gz7�Za�tl�t���#�w�hsQ=�	��iuW�F���"�濣5��$ϳ�`=�*�#MB�`s��\��8�N�1��]�o6��~���R91��*a�2�<Ϋ��A�L�|\��5�v�.�ӗ�n��/��ۂ',%�4��m�cዚ��Ð�%c�}8�!4�z���S���XyM��,��n��6*��Y����"bM�& 4���-$pи��ʏ�<��y`eZ
�aeZi6ږ�&E�c�f̛�������;Ur��{z�TYc�pQs�s�o�Fmk�3�h1Z�m�9���C�i�QY�7�XxT�bg�ԛŐ�=N!�����2��.n63ˢ;ȧ*st��ռ�r�>���8`pSpa1@)�`wK
*�;tWڻ=	��ŧX�_/;A��iGP�+?�Y��q?�J�}�F�
��FÑ����$��HK�Ӟ�������'��+��	%Izk��#�`0�z�L�7����7\�U������(���cHuZ���M���	��^KuX��".���#x��6���dP��%Tx������������܊��U�]��W��2b��Q����� �h��3��MK���Y��gLWں�I����:�ZLt�H���F�]�tpR�l����1�й�q��E�Ӓ������b��ۑ�3/�"<�/�����\��دH��qg!%D؝m�?ۜܒ*AEΙ��}��Z��$=ӛ5ЍH�P�D�����v������%�@~�i1:/�Ui�s�$��IY��;.>4��ذ�����DS�u��rr�j��ӦF DU�1�s�ݫ9��)߉ 2͚��닽qCiU;a�O����cV�S���A����j���kzLy�sU��؈��w���M+�M����p�B{k~� �-2)�K�e�߶_�>�����QGc��A�q9b%�[c}.�2D꘬�}Hܷ��o��	Q���{U`��O[*c�^!R%٦�Ƿ-_��V��N�C#d`[��$��C7�1��̈T�;i�*g<�3���	�Y�4�Xͬ�$�G��)j�h��:R8���'�ʋ�w͎�֢�fCw�!�4.} ������3Csk�c�S��|���7�K2��F'�30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�ڜ4�y^�*г�j���&|f~o,KN��xslЗH�S��ޣaQ(��OU8p��ӳ�ę^�|�ΡZ���%C�A�R�n�X���<���.���R��_@n^��g���+�¦���,t�_�_��t��T�(�gџ�l�0����G�KA�����tf,�8��'��J}����/rĞA�ɢ��`��F�qX�ߌ�����a����:��дd��-��q��!���7'c����~ZX�ox���\b� ���y�1Mfߖ�E2Gb.�S��^'��I�d�0�s�fz�={���|Y@�.����su@��_7ᢈ^.�)W�{p� �H�>��~νU��M�ز�����
�y�Q��]�����U�-j|@�'[vv&&�/&��΂|�S8G}(;�^f�&�<4�~]��X/�\�4�Iށέm�<�	�▴�����G������X͎0	��h�ٺ)��An�l�jǲz0��{Ո�᫶��S�� �� 9D�1A؋=��c�lR����U<��-�e�
��Im�g95K�^���(��jc��K����52�� n��e����z�1��8K|�j�|��;s|/�������`�D��K	�p+	�THˀ`�o�FRD+'��
8i��1V��05�Q��wExu��O��VGc�Y��leykD9|l��[���0^�mO��x���I�k�����T��ݺ|Eo�E0~���x�;H�WH
��i��������EC��
����v��(d�i������F�7$�z�$��Iy�,��;M=<� ;�$��qGU���n�L� �μ;,���ѧⰾ�]���t��[���1����>V`��y�J�^�}^�����e�kbt��'����ඟ>�u��>٤X^8%H
��ɭ����]�&�4�,Ԙ�r��p�$�:��$ˮ����r�� c}~9�Ǉ���c:2��|�Ll���[r˔�����٫،���,}܃�a�%"�5l�f9܃�&�%
���AO&�la	-�8��3�D�5�;;'�<���1<��rV )4���\H�i��y Z;І��ڽn���L�e�D�V;�H4]m����)�9˯բm�a����R�sd��J����p�\֢�h�E�r�A�Sނ���-F���">��_�A^vӀ���W��36���sM��H��~Cmh1)V��%��w�ɮ����Hqw�nۣ@m�7rVE0�;��h�zF�饋�U��Q���ѥ�(	�������.�.}@V�2{5��X��B4S��/
Q��T�}/B~4
O��NRjWף�ؤ{�
Yg�o}�?�����J�d#�	�r�KWܑ�\j*���4h1��D�^�d喂	�����	N�6��L=��C�1�3�vM	�XYg��X�ʖ�����ᩣ�w�г�s��\M�˹��GC�k����]���J��%�&�2��==�ժl�Q	hr��SZ������둷i������F@�r�st�%C��<�)#3j��������G����N5C�P=~�"lIZXM�|o�q�^�e8=u�&X��?�әI�t�0�k�f��*Ms��t��&���De#8!4VW�����H�!'�s$����~��v�O%lM{�Ǝ���ұ��%I�6��q^���gԻE�\Mk�*?���+6�'�!S���?-�?>2 �a����4�ǜU#>'��-,��y�n�=��0!���4����E�$3��#l]����'N?��F"/���9RGt�,N�ܪpE��s����朿8���(y�떦�u�`4�:-�W�Ƶ@�_�9�`���56zo��ĸ�B���#�G�ûDz=�ԇH�,���>��Z�@�B[4����T����G/���> ��k��UI��gl�˅� �&i���*=����hAr=y.gB)���wzW���i��6�4�	;&r�S�C�D������T�sLS�'3��P�ݞ���C7�"t���\T0�Uv��^f�P��}u�*��2A��>k���/�������_�2��f�|ex�q���(���P�� +[���}%��A�!��c0TI?c����"њ�L����y��F��w�hu���^�!�H�^�yc�2����"���O��'�d^6�*C�tp	я�j���Y�v˫h�e0���'���ە�{'�n;�` 2�z�nJ2���7R� �v�(�n�pJBT�W��V84i_~�e�,n*⪣w'd$r���l�;L���_j�dzб">�����9��e��T)l:h��d�H��������A�'�ۭ9�~�w%5���<�b	������Rq�%��6���w�� �H9�ػj
��Ơe�|�$����0��.1�0 p%qEw0���e���z�JQ[g��k����߿�4������n�H˩zMZb�� ��WG,+�+��b�����df-� ��v��X�Y��ųxb\���,�y?	2f�W9E=�.!��)�y�t���(s����~{2�|d��.���,@�0�_���I>�)]d{g� ��ͩ��I��U��ؖcL���O�����-y��j������,�U�<�5�'F�|&qY�/ѭ����1�(וGHI��h2��R�<�u]�8/.�e4�f�9l����D	��FE9<9e��ci2�;�E�s��A��A�<	�WNާf��Z�ް����*x���!{��X���;�|�)�P�>�Q㜑Eh<"�5%���1i�������d��?)��I��B�T�J,�[+�ؽ�����u���5��">�X_�Jt�d� M�\re�#V}��@�ŕ�Ηgcќ]-��l��(p�7q�2�(Ѥ�!I��P6]R(jr����_��1q/p�� �CC�]��a�KՖLa�3����&��_../��iX��y��_�K��R�Zܤ��\�$N%��f�X>��}�����I[ʲ����#H%x�3s�d˟�i��ƀF��/��)<eħ��c���1-�Vy���4��Q��������k����G��7���}(�Lfsw����S�4���5⫒�*N�G�N����f��Kl�xLK�AQ#���ca��߳�	8�u9lY.�R[o���0Κ�V��Z��N�RAN����@Ck4��0ʍ��;R�-�_�^K/g��褒�[^/��,M�J�Xt���>�g*�~lzT�#>�� �xA[�i��t�q�P�*�V���n�!/+�\A�] ��o$�x��	8e�i���W���A�K�(����h0��h�玀m7�X,����+��6��e(M�AM�Vx��[I�����c�����T=��O��Cp��"M4϶�Psk��P8���:�b�Z3�!ܼ�5�:��ϳɽ�0]o!�)!`�2��X�jP�7�v`c�U��na}�M���6��b��ǩ�r��!�{�x�vi|���߄���6N	�$Hw�~�6a���u�#x�Ѕ���9\u>�%\3 f��XI�}w�O��I����J/��� %O�k�6���o�8��^���_p�q����wF���t�c���-�m���U_
Q�)�k1���������g�k����}S[�f��Vǭ�<�U~b$���v*��ǳ���2^f�[MK�,�x��ܗ�����<�a�0���Ƨ8����~�=�č1�5�E���h��3��R�Ǳ�j<���sg��͞R��p_'fP^y��g�	��4�>��x,����Ct��|��vg���l�~蹮y���A�'JQy�t������
m�6���,�/)A����~y�o+xoI�f΅�l�B���J���(j=�9	�����lm���,v���v �68�7(X�TM`2޺Ťj�5��t�c�ad�9�{ϕ�N�ƍcHρ�*P�Ȓ��S� ���]3�������<��~H5�[��!2�s`�AZ���xj�t�܁�o��XYn,�JM Q6e�S��dϩ�y��2�{�~w��0݃\sY��;�6�,�%!H��gq8���l�1�dR��y����F���],�Ξ�����õ��:"�R�9H�u��$��]��"ƚ�/�`.+�7��Ը܂s�UO-d��2���DGp�e֦7x�<�[G�%���<����D���,��Մ�.K��@��6�0�V5���;��b�g�%�2��񌞜�V�32#���O�[S��幙���~�p_��=�\��6�?�Q�mz��&?�	�Ȋ�Ȟ����R8�y3%x����n���E��Ŗ���� ��hR寷�d(l��j�6�����՟᷽�m�Z�0��y:�:��ͥQ��W>_d�����Kg���y�Cm��K�:���nS_n�T,�������ʤ�K7��`�rL�&�S�rsح#ڥĿ�d���-�Jn�l`�����|-Q6�R�;p����;-b����d#��jd�z��uź�n=�̍�k���3�5;��v:Y\`O�M@��;p���ԥߋ� � �Ʌ�]|nG7��}��*��&�ٓ�*1�2�*���̊ns�S� �ʑ؟��`�ϵJi�̩�1�@l\�P�̷����?�a�Eȵ	*�q�cZr��܇�"���v<�OB�ZE��gL8�f?og3�7�"O,E�6�4c��/��|e�{����o-�t�*b���m ��I��k
.�|�e�!�z�R������r�s7�f�Iг�܊����sz�#"�J$I0�ֆ��dQ�W;�0WNK�v�#3����4�uK�4 ���a6�>�_]0%�4U����HM!�;l����k�O����Otϣ��΃���8B�X6澊$��n�����;"����$��׽9w�{�V)S��h#E�&��r߮�����ƛwv�:1U�m�>Mr��Kı�9y��Ә��myp���ђ��c�>
[�#UqPUjZoe��Nܤ9�H����9Lݶ���]eG�ӦpU��.���*N�[�y�E���ӆ��ez��*�"�7k�q68�?zqj�����U)W��^�����LT��m��?秝D�K�vbqЮ��aZ�)��L~S��J ��P&�%f�� 1�&k�+^�S��X�j�SB��b�%ʦ�b6�����<%��B ��m�XS6�5,xGC�E���A��͜G��� T�%׹����oR Z���;��ͷ�l������7s�\ P�+2&��%1���	na�|�ta=��&Ea���欙v7u�L�kDk�7PCsp}�ta��&���ݑ8N��W{\��!�!4��sѐ���Ž.����\M�\Ύ�N��?��2���(q�ڷ�TV���}�MC�w��e��8��'w�a�>���,�?�a���.���|4_��U(Qq'L��,��y������]���g�4�ڄ�����pN���BW��GlerF�o��3�kR�S������O����s��U�+�ؿYb���������"�*`���-	*z�?5�mX���&���*�Wvzz��lB���#s�|��-=z
Iۇ��
��{ҏ����BHԬ�S�?T$+��d�����e�Us1�
;X��% ;�Si�ۧ*
���h�MA��.Ì4��;��Q�W��i��k���;�z��`�%C��D�ƶ�����6y9�' =�P@��,ȧC�D��o>M��2�T�_��}Y^鎑P.��u����ŋ�A��E�+׋���FN��d��%��г|�)T�xK6��v�L���)�[�7��V�%����:�����I,N������@���JP˩S�%�$K�u�^.���K[Ѧ=��O�bf�"C��z�t��^#��C�t�p6-��j����ۋYѷ�)20Ψo���*�U���Hl��;R���[݇��Jߞ,�.O6?[�� ����J�DWT�VE�_+���y |Ϧ+w�ݘ$��z���Gl]f��o_��dǷ!���k�o9%a7���+l����B��ZH�����w�'�9�'N~v���A�I����[CK��%߫�=��c
�D;� � ��j"�>���r�e��/$^R��]��.��d ��%E��ֲhSp��z�W�[����Ͳ�r~�K��)��ǜ��HJvz:kߌ�Ì� +|a�<�W���[���M-Uc��X,~V��i�b)��n!�yL��f7\�E��.�䏶���;���sQ�[��lK{�/�|��}.�ZC2�@�_�����m�)j��{�% �;�͖����d�U�%��0?R�\�ŭ��qbIhyJ�⵱��TE�UgYԤ~'�e&~�/~&�&S�/�G�nQ��oE�~?i<�Ug]�cZ/�Y�4D��&a��\Z\	0̽�Ӣ�M�(�%/����򻗀sv@'JR�:���\����A�>�����3y����{Lv�J( <qH�2��g����I�
6��&��l����_h�q� �>�Cq�����K3FiLi�����}m�\�/���X�4�SY�K����x���H\(��%o��f6�VX�`}�Qs�U��Iy,����J�vz�%b@�ꩩ
�B&��\�A�dn(��a�P���`c$e��/�-P�9�nK�RXQ�!����+����-����H�L�}F�`fQlJ�`S�ْ6��e��pJ*�l���0K�%��f�~K��Ax�5?�_������a(`,�M��8�WJJ��gU�D��θq���l�fz�R���u�!Z��&�ɍ�4R�_�@�^�4/gs����[r9K�_,�!3�v+t�����.�g���l�C�)k��FA����K�t];�|N���t
��L%/���A������H-���J<����;�����(��i��(��\�lJ��P�mw,).c���6���(+M��e�X��֮��ԯjcG��Lg��!������)�P����18�g�6���39�ܚ������Y&�N��!��`�������jnٖ�T~���En���M�G6����������9�{������I����x6,�����H�Әg�")���#1!���`3�t�A�P�G�ѯ�]?���5��Mt�/f�"�R��,w)���.��>]�"9e/���.E��7&3\������uO��E!��kD,eE��7r�<u��xEg����$U҈�D�V�G��֠G�!C����~���`C�V�v��r3bQ�븸��,���:�������3���$��EI;���pRh�=��8����dP�����l�<id�����n$R�s�3�A������	���	�9a����` ~�~R[g��ȯKd;χ���	��!ѩ�tl�X���f0�O�yn:����dQT>��T�Nj�H�g���ym�keK�����bmS���Td�#_�놠q��k7)�\`�O�ڝ�S3�ؠ3+��Wdre�-�9�n"��`�@���:�$�TQ)6b��!�H�k-u0����7F�����;V��&�F�!j̠�sk obiy�5n^N�IOY�W/� "��N�j����Gm�@���Ψ��y8n����a��=&�����/21���z��*Qn� �S�vڀ�o��?SȢd�i�UƻĈ�@_�E����jٿ��,���)�Ȉ����Z����lU"-�)*�b�Z�g-ufr��o�y{�*�"�R����4v��Ӣj�|8�8�*�]o��Ft����l� ��KI��
x�e|��L!���2���c]���7c]�I�@�O�H�j.���q#�z$<!��ٿs���jA-.CK0*ω�R�#Ʋy��h�u��{4ӈe�t��>�T�0�j�U'
-!�0��5kyO�������ʰ�vI�ζL��	�X)���m��!���;;��w�LW"��P��n�)�_�h�(z�9i�rR�J�ԉ�BNv���U���>a�7�kT1��X���j�����'u�>B���� >]<I#%iPh�So�MG�!/97p��7��,��	~��3eZ�k�����_T�ͷ�*�׵�l���8ܑ�9��e�>�*=m�7>;�6kw�?���I	��]W��q�s��'^L'M�m�N+?z��DŐ͑��E�a�u�o�ڜ��LQ2��}�ޗ/������l�J��~:;^D��+��j���7��z�P�h=��R���	 �$ ��-���x:�NE�(��cͯ~���4 'Z�%
�������b�)Z��=;j��� �'���u�����L����(v�7ZTxY��߀l�c�)9�F�4��Χf���� �\]�8b�X��JBW	��X��Yrs�F�%��N�� o̴(�s�j��лS���k�[�X\�`b����8 �N�?}�h`O�	P�[j�รw�0A2l�;�5u��v�"�h���������0�Y�!m�/��
�5x�����$� ����zV�oJQ'k�r�+ɗs��J�=|g�r�I�a`��҈��aɥ��Rg�}�ְ�
���	v�& �$^�ؙ�.�1p�z�<:8[E�z��ĵT�v�bb[y�� FO�wڭЧO?q��1�+I�H�˲�f������Y������J���b�I����*ӿX��*�v����n�3���y�칡��n����	�ŤHWX��{��R����F|io��V��s5)�h�S�����oc�����kP��l@�g��Nd�0j�Ov�x_!m�Uk)5�Y�ͽ��P|Ѫ�E<+톧�x�[$��.�
�1tiz<p��M�?�EO��
;���ac����}%�R� 7���i���_,,���M��f&q$�D�qS��'|2�X'X�Zoe,��>�3h�	���
�օ�牝����>�ލ˅�J��Ӊ�Ԧo9��ےk��P��p'B��;]��J��X�(%
��Y g��Q!���S�@}�`��r���Ѱ`�:�q�����g�re�o�~ų{��R���:>1g��ELx���� �� d�E���^O���3�&�lh�|a�~�"U��2J9hш&�$i���LO���a����J3�&Q����;30<<}���=zH��P 5%;��H��>�� ;�i�f6���)�LR1�ׁ)V�bH@��mL���5��9W��y������Z���)�V晔��N�p2m�����:g�M�Sj�!��L7�G)�.�}�<-Aj䚀Fm�c/슿xz����^���E m�ٞV�>P�Js`ɺS�(ݛTQHNPȣL������VQ6	;](h�3��u���a�\Qz�����(��w���=��}n}L[��!�����ըC�B�ءm�j
]����s}gkB
��O���N�X�W�X�0Tt
eQ*o	�l�b�i��}h����R	y�6]��m*��Lb�\������SF����R0D�u~���4��c�s�5�����!a�蔫��{�۾T`�I]-�����ֵ	���"'�蚂�2!z���-�:B$Pe#����Z9z&	]�QTĆ�ď461�Y`B���opT�3:�0���������:��i��&��TЅ W��iv�A*&,��(�A��P.__'���G;�W)�im�~��J;/�e�|�CO�)DIf�{�Z�����k'm\P�6��Ho�C���ȋ��`�$T�45?��^�P��Gu�>�a��A��Ǚ&��/��s��L��h�����Ŗ�xg̚�o�h;���[�{��U%�L�jYV���Iȃ�7�"�cS��G��өo�B��Egu9��^�?V��&�B&$�K����"9z#���h��7�^���C��p����� *��7@Y�O���k0�������q؇��Y�W��iHݣ��J{-ͩJ��� ��y}�7XJ+�RW�#xVav�_�h���k(�wВQ$;J�Ol�U"�	ru_T*Od��,��4�����9����ʪ.lC{/�@��}��7��n�!'*<`9�8�~���>��e[7R��w�r;-�����4�`�* �MX�bjS☸�e'ޗ$zw	���.�� y#%E����
��z^%w[.d�4g�ժ���+־E}�8LH40	z֭ZߨŨ� ��+��������ժaǭ|��io
��XH�d����bE��
�yh8fӦ E�U�.�0̏ҢZ�=t���X!s��0�{{V8|͂K.�S�_#�@���_�=�R�)���{d(J ����2�?��U!�LCL��# � ��'cy'�=�Q���p�PU�3���'Oɿ&��./�ݰBa�� G�sR�ug����<(��]�P/w��4`\e����x�.	�P��/�n<B$s�	�΄a���f��U]���d�	cy�N�����Z����E��)��{_����F�e'��Y:k�z����bh�"�5��z��'D�tI���Ԑ����郬�g'���J�&q+AZ����z�0�&��^���k�i��J��8��=I\;7�����hž֌��%S��8���w}(K�qy��2����H�I!��6�M���G�p�_s"<q���	DaC��O3�K��Lʋ�,|^��^&(_�/�:X�PS����K�:����静q�\3y2%��Wf�XXG�}5��@��IĄϲ�C���g%͸t�t/�mDP�����,�y��ᵲ�����G�pCc�Dj�-�	!�Y�m��Q�^��)ٖ�0�T�W#s�%�Ϟ7�}�FIf�>H�k{X��_������z�*w�ڳ��pg�f���K���x��*������a��u�8~_8R�G���E���+�΃��F��eSR�J��:p�̝I�1�����gR�?V_%b�^7{�g^��q�	�j��,7��A�t��S�g��gsT�l�?���bn����A$H����t�R
� M9:��U���3q/��As�͆�v���ӄ-�E��RE΃� �v�r��4�I(�Q����
��Pћm�!�,4.���r6vֽ(V�M �C��!K2��QcR����\��w��L���K'����P�_܂ғ�r�+��3�����c�;����ԙ��!0$`�~@�!x&j9���w�~�kn�z�M^�o6cV:����X�h�p�~{���z����+��6�<��H@�g�Xt�ה�1����K���y��=c���@]�31��`�8����"msD�w�Hꢊ5��;�]U/"w@/�}.�;7s�N�ꊈ�O������@�6%�DE�peЗ�7��<��o�#C&��{d�!��S�D�1���֋l��l���>F
��j[�@�Vs�t�9H�b�#p��J�׫��.R��^��}cbϙ�$�����?�����p�-2=�>���t����,��$9�Ǻ��:��=O�R6];3�`��b�Ɗ�ݝ�������� �۪R�1�өcd�
��3��4Ւͬ���_eܤVna�_U0�$wyl�1:��v��!|Q���>ݯ����g�qys���IzK���ʈ 5S�W�Tj���4$�+�+��7�`��e�S����٥��d}ˬ-ean��`����C*��2Qt���9�i�S�-�����K�b�S�(�G���稗��<�,8��d�k빧�u5�,!9Cr]�YZژ��`̢��`禹�$|���ƅ�LnE��3C�%�&�7r�(W2�ໆK��@�nq�8S�#H�H���[�����ii�	��g@�BN#I�ua�j�%֟��ȳk��/?2Z�K@���"�ڇ4���ͪ(Z�a6gJ��f��Uo�{��uU�"M{���A44ᦂ�mWM|ckΝ�4�o�BVt����� ���Iw6�
Cb�|�!��6�NY���Թ*,�޹)�0!n;�?���z
k������1\՛k?y�:Sg����r��������Iw�Uֆ�6w�$4�� j�5%բ'�<�/Ej�E�K�b��O+j�N�~bl���n�K�8�j�je6��Q�p0�p����\��9�H���������H����#(eY��h�c��o �l�*`Ӥ����w�-�X�e��*p�7���6
�y?������@�癀W�3�p�أ֙iL��rm���?��\D$��ENЀ���0��{�HL/��n��X[�X/<��@���}��^#74��A�j�S����wC榏)ڋ�������Ѿ� H�֡*��!�x��E$�D�ͮ�k�W �C%�`�)�)����Z;q�;��	��t�4�4ۼ�.Χ=g(զOZ��o�hgl���5��՞�駒�F��h���-8�Y���QB6����/Y"F���%��'�o뚁�ro��ź�S�9�ҊI�[ ��\"���l�W�  ���?\R�h�`	更[���T�o�l��5t�}v��9h����U���b�Y(���nS�)��5wS��`j�1t�Ap_�N�#	+®��'����*��s�h)��,=����I!�ta��Ӡ����`>�`g��ʝ�uyO����%tvy�C^��ם|.ص�9��:�R��Ӯ���v�)�[��P���.�V��f�Oq#�KêC�H�+����v���{T޿M���|��qt�b)����*%�:$`��"�b+Ҍo�=�n��
w�;��j�*:>~��b><0��۝�a��mr�}�w�|ǔn�TҪgQN+3��v��)J8�� ����m�G?�NQ��M�Z��#	�[��Q+C(I,��v�	�s�H������8����@+�^m�d�}V�
<���O!eF�8t!r]����%sJ)E��%[�s�"+��e��z���;c����`lQ�5e���h拉��C�n��d����t���q:1��Np"'���1ZzĨ�ͻ쑎�|~�
�]�6�F93I�D�w��V��L��H^
����=�qZ�F��+itQX�'Fw����ESvA�I�}��3x�������md0>�ԙ��K���-2�^������N�۪��m�2�?r�>> ��Gc��Ȯ������_�J2��A�R��T���u09GX��Ld�ʙI�����!y���}T��:m��KԌ�x���S/,�,ɪK�{��9t�:���[g8)م�Q+Zj����}T�<J�ͻ�FP�~8rS|]��ʣ�)��B�#\isx=��cpʣ4u�x�������o8"`N�q�3����g��#�C��3�b�"���|Z���1�,p�$�)�zzC����G��L�}~:��]�)_F7���t�pi6�����F�@
~	̓z_#����F���+'�Xh�wٹ��CjA�൓�j�q'C��;n�R��m�~��k��1Ÿ��2-�*�9�����h��m��_2N�W?p�>�dG�޽�������_�}�	T����T�|u�G�o�L��)�G�(ؠ��!��⽵T���� Գ�{z��^���r���}!&�hf�I~���rA9���7�<1��3�����*�#��������=퀯;�M���˫��gKE	5W-%26�&���_�b��C�x��
	��h���ך��2�b��6�0�k�bzb:��t^'��~�0�*�*ꇯ�����׽�>@�撉4��J�*����a%-�N-��-=�@dwà�K0�ο�2[�K�&4c=��d��
r����K(��G�k�p��'Oc��_�]�G�vt�=]�~�I9p����F�_�a�%1��
,��ǵ=�1�����p��Z<���y?b�ť�/����#R�{k $��E׌�ٞ���i>�4�qYF�����$r�ɹI�N����e�~9=��KA���6{{ä�B�
G�F�����~ub�c(y���`� ��Y'�ywo��rP|��bXH�9ɥ������O,��M�ji�o����2Ѫ��a��5j��<w��v+o[�z� h2�2�����#�DY����~X��>��"��&��e���F���/Y��*�����1�ɷ�'w�I����'�GD}�Y朏���{+�����ܼ3��.4��	��5f�P%�}w��;�@A���K��3��e�
���|D��[�)�N|��@`_e
�CҲ�1s�8��-{����O��W��߭<��Ϧ���h��Қ��Z�B籬���K:�������L��S-�$�9�͚xaj������)�.��2M��"ex*�N�������[}׉���!����z����N�r3Y=�`����p���^I�j>��37 	�����u�[!�n4U�^9'�6�:l/��Y���B���eu �P:2�YG�rPF��O�?Д�'H@RgK������,�\��q}|��O%P�Tұ�xX��5�)����X\V�t@�R��.�+E��G�)A�=ni����0z�z�� FU(�u^�v%Ȩ_��')\`t��D]��|��wxMUĭ��:�ݒ�+��X75Ӷ���7�~�j�z
K;5bݽSԢ|(W�l^�h ķ�38�ijSy��� ]|�?�/��M���٢��)���S	l��HS���UR�B��o�ik�,V4Ҏ5%������F`�kvacBjV��k̋�l<b�� 2J�n0�	Ox��8isUk�W/�U��o�-|�cE�ܜ���@x-\���>J
/AXiv;��~�s�;=�E�[�
72t�y]b#;�e���(��?k7���䎒�Ѹ,=�yM�}���$���q�SȰ#�H��3�V�,Gi�/,���؍�����R�l���[g3>ޯ���tJ�����Ԣ^����k�I!����l4��>����L��cX�9x%��E�U�m�Mk��1y���\�r8l�Ѭ�:�������H=�raC~��~�g�,�����:�3�YL�.@��Ổ�D�5߇aN�w٢�Hdy�a"̵"Q�w��Θ9d��&G����`��LO���a��Ŧ�@t31²�9�;��e<y� i��$� ��b76HV�����;XAP�b�P�0LNs�S�V��vH��{mH��ڱ�}9Sî��S]��/6�A���l�ҡ�数���p.x.��(��?�ɴSf"�k�Ο�����@A�
�<n�����ݐ�Eء�юxY�m�\V9!ٷF��6��ɖ��6J n��O���V�Ԛ;{��h>am�q]���1QQv��Y��(��.�1Դ�'�}�D���:�+	�դ��B�&��i��
��*��Y�}�"B�[O*��N��KW_���,�Y
�#�o�zĠ�X/d����]Wd�y\�}���b��4��1�#�5�dm_=	����վk���	yO��1LB"v��b�)��F:�R��v0��P�M�k���;�^����vֹZ������/ge]}s���\���&M"�=q�0���
	���r,ͦS�ψ�`:Ϊ�㍷�y������D@�5�r`�׭�Ą��"#�i��Z���]��y*�Hr�7yP�����Z�TI�h�q�ń^+��=�y�&��R��8������@�k_g)�'�sKD't�*&D�H��_8�z%W6�J�<Qu!��'s�N�=��X����MD��O!��Z����j	���q���ػ�0�M��tkR)�u�_�'R|�yc���I�?�ߗ���Y���4z��U�Ta''`�,yP*ڸ�H���ۭ4Ɣٕ�%Ƭ����'2�[CM�����F�nB�NjVR���۴���24���1s��q��]p�����a�s����e�`���-� \��Q��Ae����G�Z�}z����L��B#<�#n5�KBz�脇�'�G�b�s���B�f�N�.Tj��ώל	���͙�0���EK��S�# 6�i5F�*�iۜ�tA���.����v�F�W��i,rT���;������C��ID9��z����L���'��P[F�nkC��Ȫo��_��T��o�h?^��4PI�uv��⠬PA#ܪ��4�~5�i\+�F���>>�K�{� �x�}ܪn��G������[��r	[�%Q������C�I����/�"~��_��kT�ά̖�l(uX�^�2������Ք?�'�}@�"�$f��� ���$^�"�C���p���%� ��YL ʫ�90	f����P	^��Y���꨸����;"J��/�i͝ڠ-�����XJ�gWo�V��Y_�mഩ/jWPw��S$���ä��lx��hؑ_�\�dL����K�f@9���i\l� �g��~ �V-��m�A'	)�9G��~1GK�Sz�ğ:��d���qΫ�b�ؾ�{���m :��`������V�����!������[͒�E����81l��,h���CH��z��$ߙŻ�1��+�Y��)�%�F;��>����	�X9-��E�bvVw�[��yل9fdF0EW�.{�a��d��Nt�%[(s>���r��{�|~5z.g\�PFp@�6?_�����"�)�Ӻ{��@ �eR�Ae��5�U���}�ˈI�g�}^���y��5�"2��a�U��^!�-'�T�&�Q/��_��vX�̒G���B�ˁ�<y�A]�m�/�4�j����ib\	�վ�`�<�1���i�h�5�ޖ&����l*	t�N���]PKZ0+�fg�D�\��{Ptv��$ǖ����m��[/�vPFhV�5m����)��Q>���8:XZ�W����n��J�7�+2�c������Q�w�<��0H��p$r�J�D��ɾ\L#^�=a��8�z�/�ؗA�"�w5u��
�(
8�q�_�2��j�:��I��_67���R�A��_dp�q	�^�:�5C�?����K�wLL{���������9�/�G�X"f-�O��Kh�^�tR4�jǄ\$��%���f2�=X��}�����VRIu�Y�I�r��%�Giꥠ���ۤ�(���NQ�`����fÔāS]c �}h�-Ll���l NgQjw��9>٧�ۚ�4TR<��#ƞȼP}B*�f͘y�\��r��ɫ�T�*��Q�(�`�!l�fqg�K��`x&-=�[�X�	�Ca$����1�8���������?$δ���g�r�bL�R�n�����1�"kq��F�Rw_v@^�B�g�d���g�[�0,'M�r�Mt�ܕ�x|g7l���}���fA5���"�t�������p���I/��sA���'�\/s�D�N�8k�T;���:���@�eL�(a���hHo�̃���m��s,%�Y�5i6�2�(���M�0��h�WQ�PxRcCߩ��>��t1ǝ8&Ƽ cϐ^�P��Q�P���c�}�<��35�k�9��Ը"ύJ��J�F!I�`�=�2)jjT�М��Nn;8�MD64�����<�i
�u{;o��+��k�Q��}�6�����9HQ�3g���(<�1^��XMp����%єͳk]�S��	(ːV�[�+�"�3��(���s�2��~�]f��"5:/5�,.Ab77�����A<�[��Oܚ�����g��D�� eA�$7���<q����T��h��N҄�/D8�Q�C��0���2����I�d�V�Y�㊴�bM�4�+�-��k[v��%:��E���[�_A��v�pN�+=xuf������;����u'8sۊ� ���R3��B�s�ˊ�f7�<k�5���#�8 z�WR׻u�ē%d�2�
^ڬ�E��S���-c�I��W��0�o8y}�:���S�QX>ny �{�[+g��y�H���&KJ����\�Sn"/T�����8�<oc7%+G`���aS���؜ظ���dn9R-v�on�i`4ȅ���noQ%Ӻ
"�D��-�?���\��$������؈�(��²�h���(k����5j�&�0�*Y+�E���u���	f+W�ù<�/�/�;ns��%��U�&�i�y��2�������&nB�1S�vh�Yo=��.a�3]i���@�@[k���f\�{���TZ�f���ZL�˵E"~��%�-��]Z�v�g�s�fn��ovO�&�*"w����4�ڭӞ�|�疝&;|o/t�V
�nM ���I��*
t��|_�!�7a����`��A�Y7_��I_,��K��ٚ�\�#1�$8Z��U����A*��0�V�N#Bx-����u�64�,����>��0t]mU�h��!�c�a�ku/\�;�¾������β�F�GG�X%�Ǌ���#r�7�|;�(���`cS�������j��)"��h̀b����rN4��55���8Zv~gU��>ݏE�g���tl(�X.�(���Y%�����>��a#��P仞o�옝�C93�ŋ��(�H݅�,��Be�:\����S����aE*]���h�%���5?e	�K*9��7�Q6g]o?�01���_�$�~W�IT���L�8m�pD?��D�!��E�a�]]S/�ژv�L���y7B�MO��î��h]�����^@���@�j*�󳑃�%���>�du��QHC��&" +=�����psx6��Ea�����+r�� � %��&�C�^n8Zx`;f̰�F���#6��� u����:�G(roEZ������ln������������/K��~���u�8^�`�ZBS ��ԡ�Yn9ZF��g%��dχo�������#S�Ɛ��m[Q�\��U0~;�4�� /��?y�hܽ	L�8[��PZ���jl�25�2Kv��hb$#����_�GY�
�«��L5���}�U�� ��\Wx������+��B��)����Ùk�����X���Sϖv��������XI9���ٍ�AhA�ۖ4;�F=�C�wM�p�܎�r)�<�h�&�Y�rr6��{ΉT�v��&Uۆ|>��㟋�\�'�1>��*1�X̋^�-���>}Y0#(�3P��vo��ƘA�w9W�{�WcL+�)�O����ez�1���p��,���(�*m9�����X9O�Y�>e�cB*]6�7^(46�/?-@�������p�W��|��ߣSLGZ�m �?�y
D�	R��lYЁ����nڼ�QLq_�񝪛޷$׽�1���9Hy���^d~�KCj/�D�Wͪ�8��p�ҋ��)���'�I� ���#n�8^xZtE&����C��� G�t%*-
�����JZ�};��A����G �O̞�̧�%(���Zt�����l����x�fVi����3�W���O�|�8��:��lBw��x�5Y��F9��%�85x�o��	��
p��iS;!g��[��\��ԊF�XB ӳ�?�+h�|a	pi�[����<,�P�yl̜/5�\�vL-hG�քC�FzY��8�O^*�*�~5��z��1�=�sD�Z ���SYG�'����K�is,,��=�3�=��Ba�Ŭ��I�遮����X�Ɵ����*gw�� �v�c��D?�����.�h��dJ:X�Ú}|�Սv���[�� k
������<Xq�2h�K��H�$�����9�ʞ�� �H�5����db�����^�*�\�;XO���ebl
oT~ nH�w�����%*����<Q%�޼>��~쥈��w��G|�60��-���Qo<��׊)�B���$�t�2�Nf?$2Q�����#j�f�/�+�7�,L����1{�I����{��~8r.�H+}԰%�\}7w�<�2�p��FSU{8�v]�8�Ƥ)�y�s���CE�ʦJ����	ּU�ߒ3�`�Ȓ����f��WC%��d�>�$ߟ���9�1ד�p#㭹�m@zF�V�.�R�g�~]o�]s/FD.�E$��$��싩�2
A�����N�2�-F��	+j2X�:w�����A]�Z�2������W��&�m���m'��@�{�I2P�G������R%۫ �m@�2Q�m?��>�1G�x�oi���_�;e��ҫ��TD��u��ZG���L%쨙*����P�!����c�T�R���3��
�Ux3�ߪ!�T2f�Ju�X��rݎ��Ɛ\�����N���e��)��&3�>������/���2�*M�%L�F�
��H�od��-��I����$b}��CխNӚk�5�:ի��P����0~��b]��?�tG"��༓���탱��x����@�����J��_�-��a��NP=�-��nZw����N��[x�s���fc`odO��U9�����(�-G�CpE����c��%��~ӵY�	t���= �u~��6pS�>������ay���ཐ��ְ=�)�����1�S�7�#��t�ʨ�$/�]���<@{��$SIE��s�"��Ni!�𨴎���Y�$����|h��q��AQ~�Oߎ	I񃲕6`D���Bf<��i�Z̅9�~X�cki��3�[�8Iؼ_Fy:�ˢ��P�c+E
^�N'��e7���ز;�k�j��)�9�2��{���ؽ�j�ՍwY�v��[�=� �Y]2d4��7�D�[;����ӈ�����.K�X`��đ�Ş�Y���Ю�����1�ZC�t��ń槥�G��pY����m+KêR��3��4,*������K�� �V�e�@�@���}3k_��(E��`�DI2;�QN6�@�}>e͊��
�1�9՚��R{�ڮ����Z{c��ޒ�0�)hI���>���mN��D�K=���!{�C<$�;���9�J_xEz��/�c�
l��sdB��O��u7e��N�O�����5A�R`�v�0�7���S��B*�N���3�|`~6�����V�IS�n��tl �l��k$'�O��u�v��q����������:�㎙�)������]vuÒm:5HG8u�F��KO�+���+��g�����ó�A�\1�
}?hOH�TU�*�[�B�5�)-��0�\k�:���u*�͙M�'��e)�nl���U��z{&xZ�ٱ���\'"�K9-�*7J�Bg��Wp�����U����~=�5���g<q��5�d���[3�4j���K~��`���.�ϒЮ+�X��G8V1j6'}�k|<�-2bİ�y嫭��A�"�{v	O�H�����RϜK�ҭ�i.�8VW�5����G�I�9ߩ�n#�c��hⷀ�k�{l����g����0���O�x��g,�dk������Rt�|��E[[ц�#x�՝�^o
RY!i�W��a}�~�[En��
:���� ��^_ʠ�ұ7�r��1�/�Ա�,�M��;���$~�q�fC�f&�wd��YP�,��(��;��Ir�&S1�5�1��v���a>�N��dQ`JdR��(���%���"Fk-��6�$�o&8����~�麃X'u�%n@(�"���@��v\����r[6��/�<:e­�kn��`grd�KNn�~���Oè#��:�E&�GV�L�E�������Ƶ�젇���,"م�-�Z^a���"T���̋9'��&j�|5������[���MHn�8�*R/!S�X��~���bKȷ���[���\��V%KS f�X�¡}��1��I� o��a)���]%>'H�lE���cKQ��P���t��M@#hB��Uc��}�Y-���J\��B�Qʾ[�zlI�"M����3]����(C}�ef-@=Ǽ���nq�M�s�L��*H
e��yܴ�tf�n K�&x������h�iO]a���)A.8c��&V��Lכֿ �A�@��ǹ���O�R{n�KA��9��r��e�Rp�_���^��gO����V�T���,��~��1�tg�j�8<�gd:�l�㗹݈Z��x!A��& �t9)k�*����z/�(��/%��A��_�oRS�ƃ��rrr����7]��i�m�a�Ѧ��c\�_ܩҺ`��;>u\�{^&����S хE6CS���"���[�.��X^B��C�ap�H�)�Ҹ��YP�!�t��0C���)�Tم'R������l�+���J>\��m�[^���΅z��J��jW��V��_����X���w�!&$~~�è"6l��Ѝl��_�d���.�U�j`�9���mq�lF<v�T��Zd����'1�9��u~5`'A�ي�	�ix����rv��.=�B+��hD ����dá����e���$]��<D�.�(* |��E�Ǫ�$�{z��[�u�w�X�x=g����D-����HW\4zY^�ߋ�O�c~+;L��,��8%t�pC$̌��X+�#��6ob�m^��Wy�@Df���E�gX.-�;��ɴ��wy�Ġs�}�d�{>C]|�.}�B}B@�KX_N�׈UL�)�3�{'(e �͵���>�U�?l��������oF�:�yJg4��v��S��U���I�'R�&��?/��e?��4��G�f7��g�=3�<+�)]uCj/:)�4����E���[�=	3�����<E����h��G�h��*��إO�ͽL	��Nj �T�Zq�����V�����{B������8��\_��ݧ �ah��|51�����㽷�6�����a�L��*�����J8�+$Lt��G)��J�)gd�� g�._!�UJ�U5��b�\~ڪ���{�����!��s�{��;��x�{(��mq�(�2-����I�Tt6i��L���<_V��q;�Ƕ��C�����w�K�3L�t�������k�/3�-X�g��A��K�x��Nt�R�\j�%�'f��*XJ�}�Ű���I�S�����d5A%Y�����p����﨤��#B�;���ĳvVc�!�z�->���[�Y�Q�����ٷ���U�"���k��:�}�n�fk'�N8�@��_>߫�0�*���ZZ����f#��K��xX�O��%���Qaz����8u��x�7��h�����&f���#�TB�RM�^�]�OC��
Ѝ���R���_(^�
_g!��0e�g�M,�,Yܻ��;�t��*���g6�l�1�/�,��H8Ag�2�t��8��E�����/��zR�/��
A�L���@Xw&�6-kD����������G�L�׷�(��ZX�ڱ�s��mC�],���7w6�`(Yj�M����D~?�mc5j���'T�\���O6�Ʈ�D��P�p�=��U:�n�i3����Ȉ��>�Ͽ�Լ��!�a�`}lȩd"�j��8܂�}���-nm��M�0Y6�fU���
��)����{�"��U���`�0�k6Z��q�H�̾gR1�ځ�1�ӑ���~���X1]�2�{э�xs���"0�������%����]]�%H"�5E/��.3j7�n��=����O��k�󃮛���DH�ee3>)7�{|<�O��rT�ݛX�=B��T�D�j�5%�N򘵏-��H��׽V��YVK��<�_b?0��f^��&�@�}��������<2#��_�3�[�\p�Q�=*��׉���N���'ku*-���F�`�R���3�L�ť\G�aN+��@[�'39�U�5 ���R�޷�șd��|�/�7�����"J�y��	�0�vCy�r�:�%���L�Q�A�>��p��g���y�?T����K�*-��^HS�b*T�Q���t�$nx�7�Z�`��MȧS�Q�ql�E��d`�M-���n�8`��f���;���xQ�	��Z��6�-#m��n��ef���GT�
e�t}� �N��k��g��75\7=���6�Y�,(���`�{ݡ		�.�!�aN$���#n��wϸ�~�븇&k3w�+�#2��I�8�c.Zn�q�S�2���9�aJ��мKi̳˻r�m@͏ѯ2�X~���o��B�:ȶ����ZL�/�=��"0:��Z���Z&6gM!f`@o�1��h"Э����:4$�Y� |f'ڝq'oEAt��Z� { ��SI���
��|�0l!ӥ����Z-,����7Q:�I�����H:��6�#c/�$�x���X����e0X���@��#t���M�u�3X4����"�:>eA�0&�U���5��!T&��9kgVd�m��0EfϤ�Τ�y��X��a��K���i�;&�V~Y�)�G�u��]��R6�;�?�٥�iji�.�Wc �ң�a�L9�HmEEi?e�D�cb���tгl�i)��n�{Lc�����)b���{�~6�f�^���=N�ja�&��\���R.�b'$��p��g����O� �n��ݞ���x��E�+dF_�A�%^�� 9�%\�,�<,��4�EZ��;��k�\���J����ɞ�y�P��(H�aZf_Ϳ4�ql(�l����X���Q1ǧ��ج]���n6"8��ށv�B)!��j�*Y��zF��%z�L�Ŵo�U��=Ƹ��S-��=�[3`\��$ƪ��`� E��?OuhrE	�P�[��������B�ml�̡5��v�P�h�ᡍ~��uelY��n�A""�\�n5
*s�S��/��v�$r�������\'���Խh�s�T���=�P���8�tMar- $�}���	�S�M��+�(1���|K���0v�#�v���j�.�'���G�:�(���ć�v���[˛^��;��I�uй��qօ�ý��Hy���U�&փ�<��޲Eu�'sI�$5pb =�q�R*��m�'K�b<oF׃nz�twJ��T�*I����x<��WېQʄ�ꥺCHw(2||:�����Q�
�U�ɇ7)�� ���&��@C�??Q@���M̐#\|p�F��+V��,�R���)��{´�O8��8q��z��+�$����})A�<�:��]F28���F)<�k+����]�lG����x
�\n$
L`xi3>���*�8�%Eh�
tK�Q�MھX�M�>(�+��7����+E��m,��MB}�fI$L�nq,�� �v�q!���J,$a�Ѭ�y��^|�`~��炬����>�0�޹Jʕ�"4%�_Ԇs8�k���0G�����]�z]%���Xa]�%�/��RS��Q��"����d�7�rUY�iXh:ߋI�d���pr���d�~>ҧ�I@x]��:�ȟi�L��q� v�y`������~���R�n��Ra��a���"�.Ԕkw�9��,&d$�O�e�jU�O�_a.̖���h3�D�:+Q;̸L<6/�������G NR�tp_H3�#�~��;u/��{��s�LK���V�rH���m����Γ59�]�RJ����әk�81��~��)i�qdp���r���c^�f�S�D��H�EKE��e��{GAC��X�|������"١���{�m��uV�>�Cn��ӭMP�����:���>=�|x�V*��;xA�hۖ���Fװ�B�Q��f�vLq(N8��nh���JC}eǂ������!�B��a�&{
6���)�}0ܬBC�@O�NWcnW|����7
>u_ozF��ۻ���d�C]�wW���\�k�����1�?1�`��ҠdJ��	����6��{_��1u�Lx:1���vsL�����G6of�3����.�ha�ش��X$%�՟����z+��4�]�����4�J �&�����p=���M�	��ir�_xS������M��4����!"��h<@X��ry�8תKQ�a�@#����7��� ��jF��UP�;��G�eZ�)����q�^H^y=��&=�P��l�nM�DX}k<���/C5shϳtY6&��$Ɍ�8FLWs���V!,?s�ZN��ŵV���M�b��F�7�3�*���q�[%�L�����M;-}�1�G0�'one�6��$7�?�x�솷��|;4W<�U $�'D,�dy�$��
U�2�ה�4�J����)Z�h7��J����dK�F�q�+�YR�
��7��"�F�s�c%�#����u��[���6����`yl�-"��60�e.��W����Q�
�z���	�B�j�#k���{)zVQ��<B�Ħ�������'B@�I�K�yT�s��g��0;�����Mu
�|Q�"G 3M�i��*�̜`H�Aw�O.�����)/W�iɒ߮�H�;��ٺX4�C��}D��B��m��مsqg�'�)mP8���$�Cܮ��g疕��9T�&��#�^���P&� u�(�m�A��D�#\��{=d��A&�ġ��Ȯ��!�jxC�Ȫ�.De̼!4[��{�J�%�5����I$~A��ѿ���t�Hf�K�.���u�^�Ս���PўÚ|��ZJ$"j#���f�l�I^ӦC��yp.+r�be-��7�Yɒ��c�0�!��瀌�Mr��@��3�����7��,J�P��&@�7kl��.���sJ��WL\5V=�V_#(�q���.�w�d�$� ���YlU*P���]_��Cd������c�69?����l�������t��������'F{9�}~n������A�;���S������,��[���<� �����H����e�TT$V�T�U
�.�� �g�E|�R�`�p�Uz�7[�Q퐀����v�C�!i�ǔ�H��z2\�߄?��|V�+t���4o������	���E��[��X$M����b!r�f-�yD7�f/F:E���.돮TV��aL����sIR���o�{בY|�)�.��D;��@�>�_�򙈮i�)b��{��. �T͎��Λ0U�;�(j�Tح�w�Z��y�P�aB�L��U�����'�Q|&v[|/v�ݰ\��W[G͕���uW�v�<��]�Fr/ӛ�4<s����T�	(J����<���h�!��"�`�햱�v�ƾ\	� N�C�h�(Z���p���on�����{;�����A��2R�V��A(�h��5
d���������M��C~�ţ���BQ�o�J��+-�ۂ��V;"���/�:1���~[���JY�u��&\�����ƤC�uŚ.3�yĜ��K�Q�(�0)q�u%2f�ܤE��I�6�6=�������_O$�qT%��,6C����f�uKzVL�����N��|�8�/lhX-�A��s�K3b�П��߭\��%6;�f��;X�Q�}���k�I��ϲ�M��]g.%)�&�Pl�����n�����L��,��5��4�����c�ޥs�7-�	<����y�Q�����)��:2�0��]3��j����}m�fXJ�G%��YE��MG��&�*S�Q��Jc�L�f�F�K���xqٗ^r�E�a�D%��M�8.]Q)M��'h�IC�_Ǵ�r*y��ՖR�7�G�(P��u��jWR�$=_��^g�1��c[@X�F�V,r�����t�O�CxWg��ql�N��M����8A�9'k�t�
v�t�y�囀��S��/�a~A�v��E0g#���dY� \c����<'��5�����(l����!f���,4m�,�t�P��6RG&(��M�h���1��߂�/�c.���z���Ǩ���'G��[RFP�����c�NAՔ��C3��+�!�t�?�X�>�ua!��$`v\1�}3j�����|�Z0nb�M:w�6�����y���!��L��{F���{W�6x����63Ћ�3�H�͊g�UZ�3-{1�0郧�:�*��W�����]����s�al��UH"�.�Sܴ���&˾� ]�8="��/@N8.��7mf���� ��&>O�`���-�vWD�^e���7R��<�㥉}(����bD�/�DC:(��'����HM���_��K
�VO<���!b�S����U��m���Ճ����܋�uL}�j������Xx�py��=��Ъ��++0��=��'�"�b��R��3�V�ž������G4Z������ �ƤRbi����dX��,b���}͈xC�� ޤ2u���A+0�R	y��	:��K���Qsrf>9��Ǣ��!Xg��dyϣ'��zKU�i�d�S9+�TF�a*O��m�-��7�j�`�A�ASzi�����լdYM�-�=n�S�`D?�# �k��QP/���?R�/��-<������������_��;X�M+����gY�k�Z��ُ5�t���-9��Y��s���]��񢴑8b?v���6���ͅ��n�4Uϱ%�S�&�7��K�2��>���� �n�z�S~1[������P��)��iE,h�,�@�
���^�Q�����{�������Z��Q�Y�v�[���;d�p��3w�
�#��@τ�'3�;4����
�D�i%ȘN�)�@��*ew�}ҿ%1 ���a){wU�+!҄�>�z/��<�����hs M����/�!��Kg��g`�u��W�ȜM9B\�x�(���4����ə����mEe% iN+_���L��n���T�YŔ����l�~N��3F��`h�m���e�eI�*"��� ����Փ$���,ujh���Ҕ�+�Zͣ��:y�@����_��`u�Τ:_7G�S�FQ��O�L��A@y���g8]�ų)��\�P�}��7O2U[TX��ŎO��;�)�t���\�0d����_���ß/�x��r�9)ί�n������z%�Mw�󵔶l�V��,�5���T3-Il������$62U!?���2����۩&5@B����B]�j8�K(���J����x�9-Y�ը����_8�ej��@ϰV|&4�\�;�_��U���+����	��H@�ߑ�8�R����<ܞi��rVA�5�'T��f�#��֘��c���a��k�x$l��0�e7�0s��O?8�xdf�֏�k����ڽ�[�|���EE�?���@x����Lx1
<�&i#�q��.x�(e�EX�~
d	GA\�ʸ/H���.^���[7�[���x��l,
3�M2����$<�q�Q���a�s����,�Oќ�?��v��P"���;�r����C->���XJ���<w�Og�c�uk��-� ǰ��?���j���{XQS�%���B3���6�Z��.���rEA��Y>�:�/�������qr�H����~.lه9�M|�:}ß�z+L��`����il��~V[�n��B���֘Q�)a��0"~lT�[s9�;�&T�?;��Z��O�Qa�����3��A�*��;�`4<&������n� >rYd��H#���n>;e�)�[�cY�L;Zd���V� �H���m�eھ�9 h(�B��y��Ùg�(/S�:�c���>p�y$�b,����V�%S�2Z�8�v;oT�����A3?���?�l`������.�u�����m�-V�R��3 y��}�@�L��!��)��Նz�l��Vw;h�Oh�V��O���Q��ţf��(>n��^\l���m}Uw���r����ϰB�א��!
&�+�ɋ�} |B3]�O�)hNG=�Wl!���J
.I�o��v�p��XZdx�{�g��Wq��\�
m����!��1����Pd:��	�D��&���kU��!)�<�01�hqv��'9����_N(#w:��Ҵ�X�G����H�6��ܹǂ��R��
]ʌ	|���:p�&z�|��B=ޒ��/	���ry�NS��3��ժ�rp���D���X�� B@H��ris�ך=�QA#����'���;J������W
HP�U�7��Z����ֵqi^8�P=���&-�m�   �  �  �  )  p*  �5  @A  �L  6X  �c  �m  �t  �~  `�  ��  �  P�  ��  զ  N�  ��  '�  |�  ��  1�  x�  ��  �  L�  ��  e�  '�  �   K � (  �( 0 �6 /= pC �D  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr�	p>!��L�>P^�x�#\`yq�~�tD{���O(dG6â�ߘ<����F�N�B6��~�'.>I��]�(��d_�R>`��	&D��3$l��� ��'y��T"`/"�	�|az�H?X̴Y��ǘ^�B| �e �x�@�?	hlHG �*&���ɵ@�<A&��H�'�T)r��u����`��/T�i�'�S�č��F�P�+ 8x20��ĺ�y��Y8#N�P��1�P	�BL��'�)�s�Y�1~"AۇlX<�XAL<��8h�B��.z��s��N�@�}�'fvM$��E�d^� jSG�>l%��ρY7H03�,D�������b�]S�lZ�r�̹�'i��1�	��~=Xc@ѯMb����ėL��Մ��?�Ox��W���`�~�p�B��>eBV��H�Yw�^�]�*�x� �nN}��/!D�����^����b��WL����O�B���J�l�٧�QM�H�R�ϘB)&��$:��«z��u;!L��;-�Eaș!��5z�y���6G!���.Q��G{*��\�Ǭʓ��-W��S�ə�"O^���.ONA+F��6[� j���%|O0`� �B�v�ڍq�ڂ�x��i�ўʧ`.Z��y��V�k����=y����&j$�y���^9la��&^r�8Ql����)�O�yA�B��6-�Kd�+�j���yrj�8tE�Q���T�*�2����y� G�g�j)"q� �O>&ݚg��,�yb�D�#ˌa�E��^02}RgN���'|z#=%?�j�a�/>o��rw���b��}�S� D�DjF��$o�`t
�H��,�n��1�>��p<�R�� ��x�h�&RI�$��`�<)Ǡ]�S���C�g]wh(x�ԟ4*	�)�d�p篆%%Æa��*`��H��Es��:u��n+���ᑧ y���A�^89�`�<�0��%kwL1��9MV���&̟f��CƸǬ5�ȓ��q:��Ϭc����U�� ���԰�&]/+�d<sF��4�.��ȓ׀)��[�A���Ȕ!d�(U���Ҡ؄�P��3�ǶnO�B�I�'F!�6�@��$ZB*�!Q��B��7s���$�p��� !+ց?��B�IWL����C��sT� q� Եa�B�	�23���BK�8Uzuq1�S���C�)� j��Q/�9�1u�M�I��Xq4"O�����	_��K�	��7���"O��L kމ����-u��Z`�'A�p�<iڒA�Z��N@W���H�n�<�`kÌf(����B�"�j`�"��<Q왻Z���z�䛫b(h9`�@�v�<��4W�̅RQiQ2Ć�k��Ui�<yW!R#b�H%B�̟�`�.��M�<!@�s��@�B���$����L�<A�}��D���^F?�5�p�RK�<�3��-6�&�i&+��
��XGjAD�<��F�a�<:�B!|��aE��i�<��c]!ؼ,��&�06�ݱ��i�<10m���(C�I��8�	w/{�<�3n�'�$={a��;�\��3�	B�<a���zsҥ��F]5g��(i���v�<����~9zBd��W�.��!�o�<�擰a���N?W�t�e��f�<!4)��%9g��7iC���W�Z^�<Q7�'+�𛅏�6?:P��V�<Qt�t�T<Jb��Xd,�3"�k�<��a�?pY��Ht
�*T���Kt�Q�<Yv�H6�\xa P**�Hh#�n@T�<1�
ס�ΡS���)
ֆ�I�!�z�<AE���)4�1χ(U���p$_z�<iա@6��$�9V$0�q"�r�<Qt�]%L�4�2RF�]�jq�M�m�<�Se��\gX0���r�T$�6��p�<ɓ蝟Wp��2T�a��F�<ٖgE��(
@\��2G\�<ī�}ߖ�I�E�l�`�[PK�}�<�%��{�\t� ��>D��� w�<�c!H�Kھ|&�Up�!B�q%�C��CWx� �i���-���
�B�Lu�u�4�R�i��#Q.p�zB䉾^5k�)�T�p1�3L��>^B�	�U��a���=n(��3��i&B䉺k�����Īsx`y%o�'x��B䉦*I�ӁRZt��rD�<U5�B�I�Y�ș��#|�(
�� l�hB�	'���+ρ!AVy�N9}rhB�I5���۳Vm*�b�E~�B�I����U'Ѐh�^��-�B��_�Di:rcʸs�6DY�+T�O�C�ɩNQ$|2g��E��P�a�im�B�ɭQq����S�)���sE�9SzB�*�ع#́����;��â�NB�	&��
nLo��LXg�I2^B�	;����#�����e�KO�B�;i����55�R�Sd���xB�I�E+`�A��Z��h�'��C�I�q�Ґ����/~�Da#֬��0�rC�I-�H�(�ѾSJ�ҤJɂ$XrC�I	���w@�4�>0�BL�\�TC�ɚ@�B�� �� 1�I�K�)� B��T�@-�4OW?;7�ơCI�C䉄Bq�Abe"P�'&�	���	=fC�	3/&)9��]� (���Q�G�B�I;p�i�OӤ-�&��c��q�
C�I�4(��];y`�M`�/�8�B�I�o���3 �X�-"��G��C䉷s.`�B�S٦	9TΎ�8\B�Ie�θbu��:P0��'F7u�ZB䉃>Tb�"�ɏ%�P�āc6B�)� |��V'�4�H�P��-]�(U��"O^�3���h2j5�F��o�6hp"OL,�2��9<ct�AބM��A	�"O${)�+3�y��*��U�D8�"OJy���C�H�쨰1�
U��-��'���'�B�'��'���'���'���%u&q+G���'��Y0��'���'oB�'���'c"�'�"�'�z9Yq��*g�Hr�F�A�^�ʕ�'(��'WB�'�B�'h��'�2�'b��yQ�H.&�*`�`�I=�\��'���'!��'���'��'���'�>9Q�� ���g���l���'z��'��'���'���'�B�'t�H�r�P�7 ˔�G�VC
�a�',�'}�'�r�'B�'��'F��s���L
p���M�,\���'/��'�2�'���'��'���'Z��ql
�lr��D�":��I1��'���'-B�'�R�'a��'�b�'���a˖�c��X{����TJ:X���'I��'!��'���'b��'@"�'G�@u���\H93B�p?����'X��'8��'H��'�R�'5R�'V�H5�-r�,�C�$Xd0���'l��'��'x��'D��'RR�'b<$� '�<3�)�� H8mxv�'m��'��'��'���'B��'c���Č��Z�b䡈5'�iCu�'�2�'e"�'�b�'p�hӮ���O�x`E@�a��B@���EЀ��Gy��'w�)�3?�B�i�!�B#�g�̥�T���$����?��<��mA����4�B��m�����?5"���M[�O瓩�jH?�0��[��<`����B�^%�2"/�I̟ �'��>�"6��Q�
%�QI��/�T-Cr�Z<�MC�a̓��O
�6=���#J=Lkܽ@t��=�J|�@��Od�d�Pէ�O�1 w�i{��ܒبg��
`.U�p���[�h������=ͧ�?I��)X%8dyKT �Q�"i�<�-OR�O��m�N� b���W9�A��>e�x���'Q��T}�I�@�I�<��O�9#"�%%�|SG��j��Щ�����	�i�,�C�:�6i�R�Z��(BU�D(����/�l������ry"^� �)��<� ���u�"L�MZd"%ώ�<�S�i�ށ��O��n^�S�;eպ|H�bk��vR`%:� n�����|�ɾ���lm~2=��,�S�U�H9'!��jX�ђ6ƷVjڠk"�'�<TS�' �i>y�ڟ���֟��I�f8l|�Gꐝd���vL�$[|*5�'3�6��U�~���O��$�|����?)�ɐ��h�.)�T�ZG��#��IӟH��x�i>}�	��,��aó$.���4eЁ25�c�P>?4�hoZ^~�`�B�����?�����<�/O\1�R�@�c�  
R�̴yIrd�ҋ�O,�D�Oj�d�O ���<���i������'O���O%�Pȫ������ti��'Zr�|��'���ҟ���џ� ���`P��d�M���g�zF�lZ�<���_�p:`?��'����w�����E
&O�-�bM�:7����'\�'�b�'�2�'g�>���%Ƒ&��|*U�ߦ}k`�B�e�Ol�D�O~ow���͟��ܴ��)�$����d��Yk�f��f}+I>i���?�'{(�1�޴����2$Y�Fß7���h�2Tk�Sq���-o:����䓯���Oh���O���A�r�>�Y�S2� ���ӄr��9� ��"A\�mK�f%�3g���'���O:���c�t�eӎG�|��%���yB�'�:��?��O{���,Z�N�!�F��^����-e<H���ýjw���I�?�� �':(�I�[Ij扂�<�Y�K��7�&�[B&7W� t��͟�����d�i>u�I꟤�'O�6-����yHcG�^� ���}�(}*RI�<���?�,Ot��<��.:aK�l�>}kҠ{1��:�����?Y��#�M��'hNY}�Ԩ���Մ
5k�*�N��"�M	c���<Y���?���?���?�*��HRwm̆B�� [��Ú@��U��򦭉b�ڟp�I�%?�	�M�;:0��KNn�� ���	�4]#��?�I>�|r���MC�'<*���e.�(0��;AQ9�'\6 ��������|�Y��ȟ�YV�PT���IF���D}�U��؟���ߟx�	Cy�~Ӽez�M�O��O� b���C�i0Lu 9h�(�I���OZ����Gy��m�E�T*�FL"��&?ѰK�)Y7�AD�׊��\5���
�?�@��W��d�S"�$2μ�1�$���?���?���?!����O�]���Αf;�\�q��6)���r��Ov|lڭJU1��ԟ���4���y׉¡ ��"C�_�;���Q��_��y�'d��'׼i��i�iݱP���?5Z��o���À�0Il�������'M�I�(�	ӟ���ӟ��ɷ`<0�kZ�HK���%�wJ`�'�7� �8H����O���t�	�O:��>	8��0D�B4[ΚDZ�陸m�<��'���4���$�OR@��B�nl�A��hH)"�XP�h����6��<iA� )�����?�eW�<�*O�ۗ,��e9�i�EMZ4y@w��O4�D�O>�D�O�x `#�<�V�i(�28�>�Z�V�(����UFUh�U��'�d7�1�d�Ob��'���'2 ���z���@a,V!�U�-/.��i���O�5Т����s������ 5��;B@�8�㤍�o�,�'5O.��O���OV�$�O��?yS�'���&"��F�*�t)
t��������\h�4iÊ��'�?9��i�'��]c1iL4���[4�S�M>j��3�|2�'��O:J!s¼i��i�5b��
 	�P��^'?� ��k��0:����d�'8�Iٟt�IꟌ�Ɂ}:0ٹ&�Αo��h�2"O--F�D�I۟\�'�6-�6����O,��|z��}�Bh���k�kCM�z~b)�>i���?�O>�O
.|W��?�@nFe&� ���#qQ�MrĲ��4��X���`��O�A�1���Lc���$m�x�i���O8���O
���O1�:�EH�fLӸ�b,���6�j!zv!R���'M�`w�D� ��O��$׆l4�؞�|��U	�UYr�d�O�����c��Ӻ�6Z��U	�<� o�r�a1�d�)+�
	R��</O����O���O���O~˧b44IWc�G���u��'m�b��iq��h��'�2�'(��mz�a{ �K$9,�K儇K��8�m֟��I|�)擊�6]l�<� .J~?"a�i+�^D����<���&���D4����4��&�%���S3��a!��Nv�D�O���O|˓G����J9~��'7��.wTH��`�z`�
���O2Y�'���'r�'-��Z��@:7�8y@���Y"���O�9��Z:?�pD�%�:�?�%��OM��Er
�)��?~mB�OF�d�O�d�OJ�}z�ZG���S����(�&�y���=�6�޵>���'u�6-'�iށ����>"�xb�I�k�2�B��{�P��ߟ��I�c�LnZ|~B��L�R|��w���%�3�T`Q��688y��|�^�����p�	��	��\{OJ�18������Z��-��xy��t������O��D�Oj�?��KEk�,A� �V��
���%ȟ���OJ������	/HcJ`���R̔���ȟ�3�ԲףG�����'7Έs��Ο�Ӗ�|�[�l�h���`�<��e�ҟx�����	$���By�d��ԣ���O����o�<Yy�����ۘ@y��Od��O���|�)O����O���1u�:lJ�k��1Ϥ���#��@��kr�@�	ǟ, ���c�TU�4��Vy��Or��?�la�P+��[ڬ9U%Ǵ�y��'�r�'i��'����ǚz����b��tÌ\1u���P�p��?�i!<):�OO"|��OR��*�gx<(@+�L>)���$�O��+�x��ش��8T�|���P�y�Zˀd/�%CG�@��?1��(�Ġ<1��ɮ;3����K�Ha�5�ML+�O(�lZ8������	v�D�U)D�p�1]2<�Cċ���EB}B�'�b�|ʟ葑��:����W#�Ce>H��TzHP2E遯y*���|�a)�O�I>��i�`q�\+Q�P�k��I�`/���?���?���?�|j,O�oڂ$�9Ŏ�E,���cX��8dޟ�����M#�rd�>Y��M��3ꖙ�\lI򄅐L1ֈ���?q���M��O �:g悯�2I?I��Eށu��Bh?KH��#�k��'���'�2�'O��'�哢O�a�œ�]Yz��O�<��4m��)O �$��8F�O��d��]	
�lM�5�Қk����VNR}����쟤%��S��L�	��~�lZ�<����7s/�z�dH�C�*����<9�A |I���z��~y��'��"v|Xe�j��~����kN)k8r�'��'���M�q�?�?a���?�v�H
}ˎ�Іm��z	�ѣQoU���'����?�����z#$,XU�E��bx���4[�'�}���@�t�����~B�'�00�� �z�,FE�m�e Z�<���R:|! =��R(�< Cp�A�?���i���U�'
��n�z��]�D�f,��+H�62��UMב3�\����Iݟ���d�ɦ��'t~U�5��a��lݎJIjl��∞%��T�	�?QcK�<)O��������O����O��!`��9���G@�,�&pHv�<��i��՘�S���u���'�R�B�Hxt�U�_}�(���0y�I����P�i>��	 �Gh�7}��l*PA�+n��(@Т�U���o�[~� ��"iV���䓶�d$4����ʂ8d�*q��C�Ah$���O���O��4�,˓@����4���¨��ـ�@F�HoR�1r�xӞ⟘B�O��$�<��H�R�V IEG������V�3B�	Qܴ���[	P:�8:�'@���n�+��̲�L^�HN�I����2���+�OX�	���,I�2)�FȾ�(`(�Oz�D�O�Imڿ +�+\�Ɯ|"��.)p�I�A�U8����(J�'X����� }c�V��L��O�=oR�<���;9d��YPz�G�oV��4�D�<1��?����?9�-	��4!��_�>5����?�����D^֦A��Lğh��ğ��O���QA
�4�ҁ�ӌP�C��U��O���'���'�ɧ�I �%�R=c����0j����=D� ��-�7Wv8[S���ӹo��|�	�P��x7N��G�9��'սC�^��Iϟ�������)�FyR/m�������p��L���ِ|�0
��Q޼�$�O4mZ�aC�Iݟ ���Y�d��A3��֎#�;�ȟ��I�I��)lZZ~�#�#w��=�SJ�� <�*�+T;0���ZR4M�%��7O@˓�?���?i���?����)�)����f_0fn{6d7ElH@lZ#���I͟X��Z�͟h�������5?���:3-
TNd�SĎ�?�����Ş&�}�ش�yR#L	e�Ό(G�\�]��A0�Y��y�L�r��)��Z�'���֟���b�&HQ�/\v�J`8��;L���П���?�@D�'�6M/U$���O��䍤G�FqZ�OV`�����i���D�<���(����H�?q��Ҥnk���I)�}Q"! �<���HшѩF�<|3.O<���'�?	���O����|NT�ǯ�S�"�Ba�៼������	��G�t�'��`D��1O��}QE��V�ѹ�'�(7�"�n����4���ɝ�w���S��3C��(�?O\���O���;N��7M0?i�LV((��)C'�y��7RVJUrF�H$<$LT�H>i.O�)�Ov���O��$�O� ����
?�USɋ�uZ~�2a�<!ּi~���'Zr�'��O[�N͡I�F���iY�I�"��c��/)*���?���ŞM�zJ�}��ՙ��P�T�w^�M[�OB	"T ���~��|R_��Q$M*;�0Q5�@�~;0e�t�����I՟��ҟ�dyr�t��c�!�O*kP/�S!�t����R�@���O�$mZY�QG��ݟ$�'��-�j �C���`懀��`P$�+Ư��������}N��Px���eာ>� � �G�CB�2�`����ǟ��Ißd�	���2�f�9oI�`jD�g��;�Α����O}m�,�����0Qܴ��`�Ũ��-;d���f#�|�t1JN>����?�'#.i�4���3P1̈�EH	[\���ٺ)W�kU��(�~�|�V�����,��ПH*a����l	���@�Լb���d��Zy��n�6@Ԉ�<1����ɑ>��)HV����AwE
,/��I���D�O��<��?Ś�JĘZg�͓����r�����i�D���w��%ʥ<ͧC>��Y�?˘A��E�9b(Y�f��%��D�	����I˟��i>A�Iןh�'L6�"\m�pK2/��v���S"�wC0�����O`��Ȧ�$�������O�5�s���F<��@�]���Ps��O���@4/�07u� �Ie�x$9�ܟtʓ7����Ď�5I-N[F��(0#��Γ��D�Od���O��$�O0�d�|�g�H�D�T)YW�+�t�rV��;_���%�B�'���d�'�7=��� H��m�@"�	�K&���Od�D$��	��nR7�e��!èΥ8�<�᠏"""d*�g�T�s�	�!t��Ey�'M�� 7M�
w#`�K�!$Q��'���'{剏�MC2Ȃ��?���?����o"(�Q��`m<E������'U���?������̙�$��hoM�RV��'<@��D����Ȅ�~��'�5��Y$e|�1jҨ|�L���'�6�z�cC�
>��œrN�!�b�'q�6Mv�j���O�TlZ_�Ӽ��È�L�Z�ɂ*F?:A���	�<Q���?q�6��Xܴ���яn�uQ�O_�hŋ�4C̊�Yo�x� ��E�cyr��(P�X�Ba"���S�
��jy����,	������	_�'6-�w�	� tJHؤ�����	9�S���Ɵd$�b>u�ėNK��g(�5�e��n�b�lZ���S�WCa0�' �'��IupR��֜~��� �^���I�x��̟"eߦ
��L�'w�6�@;C�����3Yؔ�B��@{�:���-A��DZ����Icy��'g�듖?1*OP�iۣV�h�Z��(��ғM�`��7|���ɝPL�9���O���'v��wz|�x�f���4�L�e���6Dz���I��(��埤��П��:t�N j�91D�ǘ�(����?��?q#�i����ȟ��o�X�	�@�8��¹(w�H�e�Q3T�'����ş�S�J`oZQ~/Гl6�mZD)�-R<\
��(���"�g?�J>)O����O����O~�#��� Ls�ib�B�(��)e�O��d�<���'Uf`���?������xdTp�Hʀ�8P�Y�<i�ɤ����O���&��?���f�`)SC� |*��f��X8X!���2?���|�M�Oj���n/R�Γ]@�Ȑ,�HW|(C��_�o|��@��?��?��S�$U���?�M�G���(=��QҪ1�f�@���Q���*O>�$ �d�Orʓ�?y�-��X�P�ߡR��#�a��?���%Dm#�4�y��'S	����9O�Z�N�{f�!��fM S�$�v>O�d�O����Ob���OV���O@ʧ
ծT�f|6Be�� E�-�M�Ҹi�HJ�!�3�b�'���O�'J�wb0���P�\��s&��2,���'X���i>M�	��%���� W\U{���5R�)���B�̓f�8���O�@`N>�+O���O��+@	
.(����a \�T����`�O0���OP�$�<��i��X8�Z����1%ؘ�9��=z��]���J.<�?Q�Y�h���T&�sDQlW�x�d`+uh>,��!?���ȲlD�8@ڴ��OȊP���?!Ъ��Z!�4�ϪsK�l�%�=�?���?����?���I�O��r���GNU�� r^�HWM�ON�nڵ\�I�| ݴ���yG���H��	�м�!^2�y��'�"�'�vIPE�i*��4/G���ܟ� 2eab�D�:`�* _�`Uj�:�$�<����?	��?!��?!"��7/[ }���X�KyJ��i�0��D��M�q�F��P��ԟ�'?U�IB�R�q�*�7kHQ8f2�!R�O|���O��O1�bt1���W�(�&�ϗg�qP�K� Ak.� �!�<�J�J
�ĕ�����19 aJ`GX	,\^U���N�h��?Y���?ͧ���Yæ=A����p��K�h�p����0r�����+Y���޴��'v���?����?��n��xݞ͋�T� o�Ueh �r�L��4��D��\4�������P�s�痎Y�bD\�.]�髒7O|���O����O�$�O.�?1)��\Q�5AU��l��i����ӟ���џ��4�@yͧ�?ad�iv�'k�ઁ�QB%T��$+H6f��i:2�|"�'��O���$�i���+�j�A��U\r��(S5c�%J��$���6���<�'�?���?�����	>�$J�-G�2IZ$�[ �?����ę�əńןD��˟8�OA �@i_�v�ToZC(��y�O���'H�'�ɧ��@�C 4A�LY7bu TH4��~���&�N�x�us�����*�BLM@�h��h�'�*���Q���=�� ��͟��	��0�)�wy�%q��5� "d��]��$����IĘ��z�*؛���u}b�'6�PI�#bNT�r�(Y%Z����b�'=�.�������������<��e�� m��(A�z����i��<�(O����O��d�O����OH�'�2]�!u<!3 Ϡ5��
��'��dA��?Y��䧁?1���yǕ�v�x��@�6-��"��z���'ɧ�OV�y���i��F�vF2�I^�E���Z���X��t�̟xqB�|b^���؟hS���8-���a�GQ_Z;'D���	۟��JcyRO`�x�!�C���Ofayd�1Ht��aD�r�"��O
˓�?�+O����O��O�uA�LA��<SA��z���2O��$�1(zP$W:2$˓�Ba��O|���9�XĨ�G!�n<���ι6��dP��?���?����h���_�U@<@���d��=qbm t�������
S��d�I��M+��w������R�Dl�xQ�x$�s�'	��'C�=˛v���ݮl ��SLRQ�B�]�Xz PJ	�>�蒕|BZ�`�I��<�I��|�Ip�"�9k�(� �-�5x���sy��i� ayR/�O����O�����dV`���"]�H鰁��
m��\�'i��'Vɧ�O�b<�g�6��ġErR�iH�L��C�J��c]�@�$�64�Bf�g�wyN�xà=B@.��e`����EY7h��'�b�'�O��� �M{�n^��?	�L�_�N����81�7N��?�c�i�Od��'�r�'����$��} ���yC��z��0ۈ�(�i��ɦ#�l|�tٟ�����"��M�TW�9���ω�|�D�O���O��d�O��d3���[��Jtj݉(��i��@ϸ|�8��I៰�ɕ�M��*_�|2�s_���|"+[er����S�dQ���@!��'�V�؉�A�æ��'��=P6��:V�T��FD�Vy���K	;����	�Q�'���şl���x�ə����2�K;|%��#,Դ�����'� 6mCw���O����|�,حm�� u�2�	��ZI~R&�>���?�N>�O�@x�d��}�@����+�.���
O<�|���G��i>����'�&�x�Ŧ�.@^��$���G�B�S`�Пp�I؟@���b>ݕ'�7�M\�PA�p��`z������M}!�F��O���V��9�?��_���	�=�p�y�'=��� /�!l�����؟T��		ئ9�uw"<���/�syb�A;u�Ii����2�L��l���y_�x�����	�������O���+<���'Y"M�<LP�KjӚ5ӑ��O���O������Ħ�ݏE�:�rdȲ+b�av	F(��	�$'�b>e��Ǐ��y�:Ī��`کE�R ��J݄qߜ�Γ!
&��䫥��&�|�'���':a�%WY� ��D�_~� �`��'B�'=b^�H	�4\S�Q���?�Rf��@*��Tc�J�m޻��b���>����?YM>�f
��F&赛��"�
�Qp�e~��?�(�ّ� �E��O�,��A��I�	�N�`�q���!�$m����'l�]��ɟ���0�	E�Ӷ4��П �����H7�`��Hl�%N��J�4PV�Xp��?���?	-O�9�����@	���Y��Ԭb��jW4O��d�O��$E4�6�b�p��O��R��}2���3@��r
��"�Q�� :�$�<���?����?Y���?i����(�L�b���.��"�!���$�1�E"؟$�	ן�$?!��F��r@�=|�)�Qo�d�T��Oh�D�O��O1�qq1���wҩR��a��hiW�˪��	�&�<9��V�$�L�d�����S9_�,���)U��LM�4"�#pTv�D�O`�d�O��4�d�c˛Fd�*�h�T�D�S̷3����W���y��h�㟤[�O|���O���H
NT(f��4Iv@�)ʂ>EΑئ�iӲ�(�	 b2ʧ��;&K�'.�t��Cō1��K����<����?)��?	��?!�����X���?���K�%ſBEb�'�Os�
(�F8�$��ަ�'���K�d���c�	J�^`Vy���@�I����i>5��A��=�'�D�
� ~�($j
�k���RK,V�e�aՋ�~�|�Z�D��۟X�	�ɷAk�N��b�8REZE�T֟���LyB�|��u���<A�����yR���O�Tr� ��8t�I���O|�$,��?Y�W�c�����9*�ʬKȥ~�H�q��������t��o?1O>��h�bB�AaTAT*z��$1Ш��?)���?���?�|�.On@oڿ*�L��������l�;
J��!�Dܟ�	(�Mc���>�OF}Y�����p'�"Ob�����?!�́��M��ODe�J��O{�q��g��n�f�J��c#.�x�'R�'��5H6��'���'��O���7L�e>jֈL�Z����N`�V��l�O�D�OT�'�?Y���?ͻ9	,�+�̺ p��r�..6��<����?IJ>ͧ�?i��9ɐ���4�y2N�0�;���+w"���ɖ�y"��C�ȴ�����4����A ,;acɏ���c&�ۍ[����O���O��5���C�Xu��'�b���̩�aM�S4p����¦U�O�h�'I��'6�'32�҄��v�`Px�.3e����O^���fޜW��7-�^�S89��D�O♚���)LR����dR�i�^]T�I�����OB���Ox��?��b��<��%|�(�"�n�|d��Y	s�i�I;�MV)���d����'���i�55�Kw��ɰ�If6�)��|�����4�	�	lEn��<y�>��+6a�Rp��CO9o��,��%WO`L37oJ�����4�
�D�O����OV�d�
x�^� ��c�H�x$m��[�˓\��#�i �������mH�h�t���p��oW�?�������	}�)擷MO�����W�8]*�ݽRv�S���b��{�r욷��O�YM>�/OH��sD�/מ�
�MM�R�z�)�O ��On�D�O�)�<�S�iJ��'����{�<� C�R  ך!T�'��6�3������O.���O�� �f�x
�KEN2��H׳x`��ݴ���"�M�qџ�����nC�更�TJ�.9i�5�� ���d�O�id��O�$�O���O1�(H�jS�E���*m��T���O4��O�o�6.p�����X�	`�?dL�˵��(��Ȓu�N�{��H$���	Пd�	�W�h�lZ�<�����Jjܼ;8���#��/vF�!a�K�a���������9OۢQ���E&�h^8����MsE���?����?)�b���̄ |�,�U���7�`(枟\[�OB�$�OH�O�ӧ0P`"��2��m�ȏv	nyZ �;\P�n���4�����'�'DLɓ�n�b��kp'HA����'��'r���O)�I �M��X�2��tp�O�D��@A�^(9�����?᧴i/�Oz�'��I�9��y�T	V�5��(ʿF���'$��A�i�I&i޴
֟��9��`�ELJ%w�F=���	΢a��M�kЌ�g�פk��� !���< Z�NO/c������ҁ�QO '5��q�s D���,�dP�,�O�`-��!ǀV�rGÌ
������3��@D���ܢ=ظp�f�R�����Ak��b��]:C�cr�)��Χ�H�W�٨)��Y��U�����i�!}-�D���14"�1a�ău=�q�$�D �������`�8a
Qu���š��%r-���Íi���&�.O�4�΄3�tt �&��sZ�)	C߄/��5o�ß�������S���<�ӌ�'(5p�K
���4Bڑ֛�Vc��|2U>�?qR�^6xܶ��!�I9Y#pH�S̈T��'=2�'{6,X&�>�)O��d��XCMT%�*�x"l���Za91�1�Ɂ	{t%����ϟ��I5Q*�$I��Z��x 0�D28q �h�4�?��.
k��Ly��'�ɧ5(�5^ �Հa�.&��b�ʞ���ď)x��O����OR�d�<�"� ���Ԓ6�3]
�q��W *5��Zv]���'���|��'�"`˛+��$��Z/�dͳ���Z�2)�y�'�b�'��I�U7h�ИO
V���!��hi�y��J�8�4$��4����O��Of���O��$���ز*�)�h�A�=ʠ�)�Ⱦ>���?)���Ą:�̌�O��*�#0.��v��Z�+S*X�]��7��O(�Oh���Ot�3EI1�I�	�DL����-3$�c��6V�6M�O��D�<qG�:!��͟`���?��ˊ	S򢌪��(Gex�j%D�3�ē�?q�X ��x�����d�������[�8%R��G��	�M�)O�B��N����I̟�I�?��Ok�s�����׻v��vL4V�v�'|�o
�B�|b��[�9��ȋ���<#V��e웶�ċy5D7m�O��D�O���_h}R\�ٗ.�m4�H����'?�ER^hX�4j䤨�2���OFm��Jw�4P#�����5�E��-��ǟ ��_����O6ʓ�?1�'�xҗ�Y��rebG8i��8X�}R���'�2�'�I�n���Je���t�\)$0L=�6-�O<)9�n�B}�S�|�	P�i��{r��\��%@��N �>��U8�䓫?����?�-O�a�Ε.PX�L:���̩�D��y����'!����%��������s�]��12C,� X��E�3�H�:ł,$���	����Icy���7#-���>���;ƢY:In8���i��6��<y��䓖?q��:d�'G��ʥ�k�j�@4�ڰr��٘�O����O���<���l���̟���Ϡg����&�L�f �� ȗ�M���䓿?��M[���{
�  �{%��=d|��LB!���i���'��	�{Y��L|r���1#��11͖,Q%��@e��'���'R��'���yZw\^%�A��� ���U�[Cђ`*�4��d��nZ���i�Ov�)�a~��҇_Z|����QT�y�I���M�(O����OR�%>�%?7-�	�bTʁ,��J9 �#�=w�6� J��7M�O
�d�O��)r�i>�h�B� |!<���Ŷ4�@X�Q�-�M��?�����S��'��_�O��ˀ�B�&���$MV�7-�O��d�OF J��q�i>��Io?)�$� +
�T��,��G��u+������\�I-������Ia?��hՇ-\�{�č��@Q�ɂƦ���5:*���'4���'�>��U��j5J��"���$"�$�5b�1OP�$�<i��P*6�Z��V$8�j$�M�Z�@DϏ)���Ot�$9��Ο �7�p���`�Ud�H$��1p��o�1��c���I}y2�'4��՟2�&dٵK?�d��&B�$6F��վi�R�'P�O�$�<)"�Lަ��Gb7휘q� <Snm��<���O�ʓ�?��l�����Ox�ڐ��G��D�cW
p�V�kۦ��?����䈵�'��tq��55���P�^,+���4�?1���DEsj5%>]���?ט�U��]�c�O�j�T��0!Jf(O�˓�?�����<��>8��χ�\�f�q�<Ǆ4�'?���(�B�'�2�'��X���4?�NY��V]w��BdF�8_�6��O�˓L�:ExJ|�^uV�1д���đ�@�4k��ƌڢ��'�'4�d\��:V��tM ,26���L�,�;�]�\kFN:�S�'�?^0
��%O*d��,��mږK�>�nϟ��I֟,��,߽���|R���?��#
�I���3�"I��P�.�P����'s2Y�0ʯ��ʧ�?��'T��5��Wk��X��Z�h~�� �4�?�������A�����|����5k5j�H0��a���'��:f�=?A��?�����D�'QQ�ڄE5S?p��@��\�R8��a�	���j�IryZw��� ��ה%�ͳ�"�JdI�4�?�+O����O���<����X*�ə ~Q�QbZx��x�"DPi�������ןL�'�[>��I�(���c��ޔ�@�7#������O����O��?QWKV��i���Rt�C*aD���Uo�T���w�L� ��IyB����Q�Nဉܽi�� 	#-Ʉ��8n�����	QyB�ؤAO��'�?A���5dC�c�&tI���:n�xr��<I��	�t��ӟ��f
l�,'�D��
�rw$k�X��'�+�<�mnyb<Y�6�Of��O��)�P}Zw��f�ԋ'��uzu"�&I��4�?q��Z���ϓ��ϸO����7'ӂ-HiEa�{�R�[۴��`R��iZB�'���OR����đ?P�]�4���Ղ���!�r�m��*�I�Ж'�� �Dص?����Řd�4��G�ӪR��l�ݟ8��ƟxGi����ĸ<����~"`ұ7�lx�B*I|��c�̓��M3�����سt��?E�I�`��h��1��B�K
r��1h���o���X��BI��d�<����D�Ok�C�Ә|��Ժ7�1��+O"O �I�6$(�I��|�	ȟ��	ܟЗ'�4�rf�� a�t#sE���0$F&��gNN듯��O���?9��?�pC�e�����|dhQᛀL�͓���O��D�Oh�r\��S0����ڂ2,!��4
t��r�i\�	ȟ�']R�'!Ҫ�0�y�%(	A�u�3iX�(%<��n�-s�7m�OT���O��D�<����f���ޟ�7��}ͦ|	g�OD�t!� !�Mk���$�O*���O�X����sӤu����\)X�Mǂ|]�\ˤ�iLB�'��	���믟���O������%^�T�85�jJ0�X���Y}��'R��'�l,�'�U����0(8��ň.�:tq ��5�֩nZeyB�p�7��O:���O����u}Zw�X���'<}�!1��:\$|��۴�?��)%Q�}�s��}Jq"�%[�D�uKƞ:d"'+¦A�v���M����?A��R\�t�'q,��� �X8"b��d&���Et��0��2ON���<I��T�'>�%3���^�Hࢋ?5��Hq@dӞ���O^�dʋ1���'^�̟|��,m˄iP�3�TY��N�2 "Xl�cyr�'D��yʟ��D�O��ж�H<arm�I���CYl�LlZɟ̨!���$�<������Ok�/;i��q���[�@Tk��ɧ~����{y��'��'��5���^^u ��P�d��<1�	�Jvvu�'��Iʟ��'�2�'(�[�@4P|��`�o��I�
�dr:���'	�I���Iş �'@<�A��s>=�`,38��S�+'�HdR�sӜ��?!/O��$�OJ���2��Y4m�Y��*L/(�tͺ�A-@\Jn�`��㟴�	Iy�^�MR`�'�?����m��ĸt�vD#�bK�9Ϟ�mZ�Ԕ'Z��'�rJH��y�U>7������EY`g��[r�;i]���'O\�,��%�8��)�O��d�6ԪC,�H���Dh�f��i�� �P}��'Rb�'s2qٝ'��s����;�=@�"�#oo����a�J�2�l`y2�����6��O��O&�I�S}Zw�X����Hn��Pd�5w^�޴�?��0�����?/Oz�>� ��D��
� |�0�S�T�u b�izpR�}�@�$�O��D�����'���.:�(�!�ˆ0�VA��͞^��(b޴*b�͓�?�+O�?���ü�6�Z�kБ��W3}��H�ݴ�?����?i0+5��Imy��'y����/����Ӝ<��,S�"6z��f�'�"�'�*����	�O�d�O��� �]�vab�c�&G ݈y��k�馽�I�^���O���?�.O����N�Z�� #lDt8�LK$U?���RW�
��c����՟�������ky�.B��Y�<=*�(��f�`qp�>)O���<���?1��'�N��$�̛`O��`΋93&��Z�K�<.O���O�d�<1��ܩ1����
Â`�Q)�|r08`�@G Z���Q�d��Oy��'?��'�$�'�}�aNQ>P����W`�O���SQ�s�����OX���O��.�<�k�[?��I9E��z%aC4o�,���-q)9��4�?.Oj���O��$�R��$�|n�����xg�*~�FГ�EܷYnD7��O��d�<�������l���?=㳈U�*�ԑG"�
<Q��L	����O����Ov��A8O���<1�O}�̉�(�:"x`)p��3$�]k�4��$35�m���������S ����X!֌�!??pt{Q��g�:�ط�i���'b��'�r\���}B�ؗv�Rt@En�#�0�qA�ަia*�:�M���?�����Q�,�'����S�4��H��˯^�|� -x���
W4O����<�����'Z:M�g�,	5 ΤZ�r��'I��'�#��'v<�����O��	��yqG�[M#$�V�L]@6��O��$�O�p	�:O��ݟ���ٟ|�W%ʛ=ň���az-J2����Ms�����a\�@�'N�U�D�i���e�
"d^鰧�h�6���>Q����<����?����?	����Ċ6 �>�%K�,x�p��;Q�Z���^�Iן0��]�	ן4�I)y�@��%k��5���)A���Y�p	��$������Iڟ��'�z ˱Jt>e�$N�9�M��m�M�6KD��>a���?M>i��?� ���~f�%���'h��D-��K�������O��$�O��\z��0���4��2��])֬��KXP�ԭ��:�6m�O��Ov�D�O�]C�;O��'F�mB��̚B�-p�N�%M��#�4�?�������,%>M�	�?-B�#2ĨX�R,"��x�bK�ē�?��x �������4��!=�D]#&倥D��e�/��M;,O����Y��)A����d��n��'ĔKPb�5z�%�֏�p��!��4�?��q�Z(�����OP�����
0%F�ӥm}pqP�43���a�i�b�'b�O�*b���Qǐ�{�5s7���.�������M���W�<�J>َ�D�'�����N'�p�눣0�:��b�q�����Op��XS<=&���I��<��4���t�^ }_>
d\��-�ڦ�'�41��~��?A��?����K�0�ׁ�}!�6TP�6�'���4�#���O6�D"��ƪ b���{�tY����wLӨ���m\�<Q��?1O~��kO�on$D�Rć�e�@0xf�ɪG�\P8іx��'�b�|��'�B��T�F�X3 �<w���1c��[��Qڥ�' �I͟D����'KDm�e�~>q#&�G�}T���H�4*VT8	�c�>����?9J>���?Y����<��C�$>�V�!�훹+�f�����I3��ȟ���H�'��:�:�Ϭ	��y벦�5y����*7?��`l��'�l�����D�ß�O<��qEM�a6��gŀFq�l�B�i��'��IfG�@�J|r����1$��J�iBh8��R>��>�+Ob��6�i݁跨��v	��b���opr ��e���O�9���O(���O�蟔��á��L�N��.ϻ#DxAr�L�9��Iy2$�-�O�O����VB}�vH���jZҼ)�4�&DP��iw��'nb�O�����Z�q�Dh��i�S�$�{g��4�@�lZȟdE{��|��'���OԪ;ߞe�G���`C�!qӶ�D�O"��3C)�����O:�əw2��G懫i>,�fۚg�`Ҏ��d��ߟ��	����Ҝ������ک|6v�(Ea
��M���8~bX�-OP��OR�|"gG����BV�ϔt����k�*s\�O�`B���l�	ß��	ny��-[%`����Xt �;�jC�����m6���O����O����5K����X3�C�#�>�{p�!Yxc��������I˟@���f����0�|��pm�-ALQ��� �4��m��@���\$�D��qy� �'�M�@�'ҠLsG�0YV�
�&�X}�'���'h�	�ȕN|ڃ!ԃ����+�mS@�a��3����'��'g��'9�ˊ}�,1%^�C�%O?k�H�	�LA��M����?�/O�M����D�۟��5e �j��//`�
�+ي��݀J<���?�%N[C�'4��X�'H���0���Sd4�S���hO��T���Ŭ�0�MK�T?A�I�?�(�O2��,L�;:̨PD��q�8'�i�"�'s�����"�S'ㄵ�M�)�6� c끉/�p6m��	�V�m����	������?]Jl9�&$ Q0�+Z���ٴ5���Gx���O��1�,]�Ę2���^ː=i'������؟��	�S$P�L<9���?!�'��J�g�C\�M�7f�,z44��}�`���'�b�'1�+=� H=�H�.�p�+uMJQ T�i�r�\���c���	}�i��Kg�ħ(/�P��.6�(���>i�	�b��?���?/O�8�5��u�&�`�S�`��a�e�C
!3ް�>�����?��T.�]B�iL�M�$��a��vA�����\yܓ7�$���/v�k��	�5ڰT��i�p�4,�+Zh!��m��1c�2_�<�%$VqO����R(� L��@�P�i2d��`�I-
ǆI ģFF��C�^�+<Cp|PB������ 4{���G@	:*]��s�4m8G�&w����H-T��=8���4vF@Q[���1D�ڄ��j����'�X	v�0���-C�d���O��B,��2r-P� ����kP����zDV,��������O��C�x����%[P�����tS>�y)ǎy�X����;�����e7}r��R��q�	��7mZ�'N����A+G����s��"E�>�<�a� ��O��hem3}�BA��?���h���d̦0���Bq��2�$K��\
S~!�d�~�b�21��"$��ʀ⋸Mfax�)ғ�0�#��'c.���گ/�|y Q�D��ȟ S���(Ko����џ@�	����65�����W��!�
�U� �b�Ŗ~殍a�
�t!��v�g� s쨴L�HA��Y#LS�:�j�3%�zl�����q� �2�3�d@"/ yK�ȏ��p��M�.1�b�D6?!֩����`�'���҇T�MA��Y&!��m
����'���ز�Κ�hb��axp)��O��Gzʟ��ں}hVNءM���"2�!9(��+Kj�~Z���?���?aV��4�$�O��;E�y���Ӷ^����#Ԛn�E�W�S�>�7	�� Ta{��=���S�t���$�AY��p���N�ID�=lO�����Ŧ%*�1��t
t�c�+�+r�'�ў��?�&��,��I � �
�v�K$�^�<)q�Z�� �jÏo؜�w��C�}��	OyrČ�,� ��?��m�b�p!ԯ��B������?)�Nk����?Y�O2��G��9m�h#����q�0������O���� ?��x���*G�hqѳg�n{>�	�TҪ�e�,;���y�gI�l�j�񄀔�r�'��A����4��%c�+m��5hc���I0}>���_!���h3�S�BNC����M�6II/)�ty&��$���'fQ�<9*O��3�i���u������O���I�'D<�8�.�(E��[�Ék����'�B�ӧOV6�5���|�'P�Mx��S�2rl
�d�g��qO�Ы� D ��F8>���t�6pN���t�Z���A���.�)ŗ>�4��֟�I,�M�����O �X���:;!Fa;�$Q�6��'���֟ ����+�dE:a�R�S��ѱL<�1� �%c�x�i��7��O��mZʟ�{r- �-z�ԈV�O�4i����<�M���?��)�b�s�D �?A���?����DI�!!����B�Әc�Nh����8͘'���
ϓeJ�bff�F(��d�� F�4�=	��[x���ԅm��ݨ�O��ܩ@����L����)�3�	1VS���7��������H�!��TU�4'�Tʎ乇)̗E�����HO��(���{���pէ�+È��Ĉ�A��e�r���,}����O0�d�O�����?�����H�3d9�qȑ<��9J�g��9��EksD.��}BAߘM��hɓ���<Eɠ��`զ�JgO
��}Bo
U�|�	��u�P��V<)��Q���?y���?�*O&�$2��N�x���Ϸ�
��었�C�I4J4��Q�ޱ}��<Rf+�JFzb����O������CS��I
(�vՑ��<�T�Q�JY�8QZ��Iٟ��UCUٟ�	�|7���j[-`���0�$�A�l��X�t��� A���x2I!V&��LƗ����0F��Ç'B;	��rѮˬCrT���ߞ�2�'��I,$#2��''Ƚ�L9�@`
�I�c� ��	*Q �(٢�<r١�+�\�vC�ɕ�M�1i�0����B�^�:$ Z�M��<9*O��"�/�v}��'n��.:k���	>m���0��%7l�@`�β!�>���ɟ��`¯7*��*���&^�8$��S��\>��g�%Z�R�`�mN.J��	�<�'�r��oߐHu�]�B�|ۑ>��gH�;&b����NM0o��`�%1}e��?���h�X���=�pu�Q헓^v~���fN���C�I�eyV�ۣJC>JMp��.fSaxBM ғ2>��c/_-_���HCHv�n�!òiv�'_�E�(�:y(p�'���'�R�e�Q��ʖ����@�݉NdP����GE�m�H��	%	J��C>��2⎨~b�\`��8<O��K�F�6Y������G�M�ua=�����|�Њ	�^��7垏g)��Чe[��y
� << ��D�jK���,l��� 7��ؙ���ӮG�n�I��:V��{�dE�a����m5���	꟤��̟�A_w�R�'���:(�L��*I+!�)�0���0O&�sħD6
4HЦ�y|tа�ȧo!���6
]�1C�#B.�h@���
 n 3��'�B�|��'�����:=H^����V�V�IQ��I�Y!�d�
[%�1��.j��H+��"]1O@��'e��
��b�O�D�,��=3 �E���)I
ɄE���D�Oj�2��O��db>}JC�0T�F�H�.G�~⪍�F�h��r�&rjXด�د�p<!׬�A��P�A2U���҆8�
%R�ǹ\�3T�i �x�(��?����D��ҝ�Ć��1�JA�kݴXd1OF���R�KtN�8`Ӑ;�2Cv�T�*G!�d����I�C�0�0P�wjH%َ}�W�b��E{��)@�u8�x���\=�9�tk�")�!��0h�F̓���b�H�sDJ��zx!�d@�WĒ�qˈ�H�h�����5ht!��3z (�+�J&RuԴ��$�(_y!�ĐY�y��3V�:�E�Oj!򄈨;��0 ��g2�r�b�4*�!򤝀7�8� �d��q`K^�!��ņ	�.8��`Ӕ*t�Р4`X�3�!�Ě�-�ӗ��nj�0���T]!�dS18��m��_�s�@i����-	G!�dϩ7L���+��R�㗆A�B!��*u��t�k��zW�:!�D�*MC���� �b/��r����!��K�Y�rq7�o�,EbA��;y�!�]�}�dX˒l�0)��,8����!򄄁p�\ي�W�O��<b�$�!�dA�AV$i�I,EU��)_	_�!�[Ze�i�E�m�8{�V��!�
� ��aK�'Ez9�FiϔO�!��ٽ&�^e�b܉}T
�Q�+D�!��/���80���@�)�F�.q�!�"T��8J�IM�I)65˱@̷�!�۹]��i���Q�P|���d�U!�ܩu���f��<Q�(XP�I.x!�]�2}���̋�C�6�"��Y!�!L� �7�C(i�4�3.�Y!�dZ�lr���E?l�p�d�Z	E!�D̘z�;�޽oTp�i& T��!�䓣GN ��䊟5|�@B�R�!��1�|a)��Q-(�v�h�(:BO!�/�tų�aY�g���SH�9k!��N�8K ��[N�"p&� �!���3����NN�ut���増�=!�D�W!��J�ƣd҈+�L�-s�!���:U��5 �H�98g�X��(L
!!�� *=:��H�n��p��U|w!�$�P�̸��	+�y)T CbU!�dO$�*�[hZ-�,A��1'�!�Ăk�x�)�o�<֌�VPc�!��NPցXE�رE�z�mߐ�!�$�{����/ldp�o�F�!� �~���͖*Q\�0�!/�)�!�ʜu7���ŠM�\���.�	(�!�d
��9��G�2p �gٲ\!��,x�ʤ� nO�N������ȥ6Z!��.Vڒ`�Bgߵ#���a��A!�ӲnĦ�����$�h��5�!��P��h�ٍW��ړ�Y�F�!�M� �@B� ޓ��9An!�$*]�99��Y�q�VŅf!��=&<-B��&��̣�c��^P!�� H�! d�� w�hk��^Ej(��"O��Q-̾�$���-*�E��"O�y)��R:ʢ��#j��;"O�E�f�K�7]v(����C�� JT"O`a���أR	� ��U�<��ܨa"Ov����Н�h�*FHē�R��e"O�h��H�}5�л&�݁S����U"OZ!QU ə�d���K�/[�|��s"Oh�ab 30�x��w�ޤM�%�F"O�%HҩFt*��Й��Q"OΝ[W�W�L��(6j�'X.�C�"O��ɤ
��D�� z�	���`Ad"O�MA"+�A]��b�B�C�K�"OT�##-&#М����{���&�'��i{�収m���Y�j� ��]y��W�B��4^������]E��)��	�C�`��&C��>���^�&G�px���T�>a3�
N'V����V*������:��g"r��:s�܌@���4�Q��/Ĺ�ff��S���Y��Pp��g$�e�e
�7��B��λ_�z��ȓR���g�����ZB͝T7���O|�5��?�~dW�G�`,$��E�6TF'͡MZ����6���	t2��-��3\ԡ��C�$"��X
ci׀.88�M�z�dI f��E~���i4j��%+�1�b�:� �r�t���
]��Z3+�gi0���5+�FI�>@��8p��!XX��Y��v�աk����v8����o�Dr��(a�^�af8�)�>ѓMG/�*,sC�YL9���q0B.U�L��/��P
r��$,U6O��E��0H|���DH�,8���M���䞮&Wܐ��V<W�(  6.H���	�Q�l����B��@����$���~��;:�a���$���c��5y���D�^!1O���@�0��L�!/
_���Z�����'�ܭa��6#.����J�o����b�A�?G$�(�\�K�υ�a^�'�}��N�x��Kd���x����ϗMn����B��fX؋�����O�pC�_\���ϫ �6���D<s<d�PCc�?	�a�9̄�1�K-u�Fa2���K�'����ƈ�{rH�aŊM�/`�c��n쌙�����K�j�a��]�f����(�$MY`�R� n��">i�$@�@d��!̼��~�<ݘD� �%���C`�|��Z%gL*Z�� �@璮#��(�f� LLĻ3�d� �Ź7k�K�.�86a��2�1O( ��ML��Pa��>ga u��-�)bք�*3��8	��0:�B�
�-ڄP��+��b-� ��f*xt��ئE5?�(Ҋ�0=�0n�6m��v��_���e�n?c ��3|4��ROU�mKvh�D�V�'Tآ�7*�����:y����'�@ʖ�;�P�.p��e�(��D�{@�DxܓO�Z 8m�Fx�;F�@��T̼a���H�#W� �B%��I��A�,z��J�' �=�"#h$�c�<�&+,(��$`��W�.T}  !�I9w-��*�dM?R 4I���Ģ>1S�J�F���!AP�tll�DI\7��h���1�Jq{�.�i�������(o��D��i�Y���8LOfY��EK�-���2�N�:���@�OLo7�ꅩ7�?J�fX��M[�m}��0�J��h``���=H�S�J�S!�DR�",����ʙ���㠊�+�$d(�J��਽	�Z;
�1O���JJ"xͲf2�<�TK�:5��� �Wx�b��';�\��KA1����$�B,�6 *� ��\��<�<)�(��v�=7A�(�,5�6g@�1�k"&TZbh�bǒ�F�x�F}2���b�RĢQ(��k�,�i��q!�A�K>���Aŋq��93@�;B�t���S��T��gA}��� ��Cȕ���T��a�a���ZƦ?R.B)
Sm�L��TҁӪadJ�ce�dI9X�B�Bpns�R��gE>q!�{󄜈%=th�A�?:�Z�s�̘�L�ȈZ�K��Yt^��C�T>#�1O^��G�DcG�� 1�H�`�ß� �����:�����'qbb�h�;f�1b.�1G�n�;p)իMZ��<9t!ŋ�Z�c"E Fa2q��\̓A���(6�ܰ28i�lb�(|G}�'�&��X�8h�d+"H(}@'�qH�Se�4`�j +DK�t�Ji���u��Lb��4T���	{���� �=9�F�K����z牍Z����7dU�d����3;#����yKFc���dX�O:��tg_,�.P�\ �dH�P�:�"~F���P��AOM>Ĵ`�S��8`�t�ORH���Y�H�RI���9O��;?�X{����L��"�^��L�'�1�2�'�&m���&s����%��:ƜS� ���'�ƝQ�(�F�Hl0�g�a��S�:Id���D�TK�[����J��8��L{����L���Y����
p��3� e*2�7���Q`,&���2#�A�b�Z�s�;P���`B
.s"��T?��$�E�D���Qi�">��%q�s�������*�R�O�D�x��Q?��?!���$�.��������k�In���ڠ)d����	O$�Z�UI�5V����м]�E0%�� ���ɬG��CD��k]v(Q�F�L�">��@�3<��u�ۮC�j�ju����r@X�8(�����!�hxE�B�<A���c���RV* K�r�YP� �<9Bf]%%� ��"W�E�
qA����h��HJ�L�\��08 ��!'d�i#W"O ��C<S�l��5�S �(��#
i0�11�F;C:2u�B<��g���6,�G�_�
��|��,�L�\͆ȓj�QŏfA�B�� �3q�EѦ-����$���{�,�_�"!"b��rU�l�E�3�hO`!Ip��Hƈ��b�L5j�v`´�JB�X�YҸ�*�ѷiF��j��B�<���+��1�M��oX���6��Ħ�g��fB�H���ZYFp�$��OQ>ט!E�z��Ǎ�e�mˤ�#�$B�	�)�,aP���0c�䩁��3.5ܐ�v�&�?1�C�:8��<�V˽~J�E(�I�R[H�P�[9��0��=�����7E� 	Vb�W�L��`��3v�B�҇�E��zA�DL��<a%T��=�S�ѭ/��. �I������ܓ�`�
g��n|sf��0�0M�*#��͖���؂2�2����~�<!�"H�&���,�QaFm�Nr�� �d�OI"�n�f����)��y'n�4-`��ːoV�/��aW����y�Lȴ��t�h��;�(1˂&ʓ���5�hP`�]�g���ҩ�C⟠���<�1�a�<cLx%KV�/LO�2f�f<$)��]8n9�D�?�u���4H|����冣�4��tKI5>)H��DY�jHu�\��#�X"\I1O��'�H����D`q���A�Z~��DX�s���:2��Sg50X�Q�daKO�<��E�T��4c���]7r�1�i�.��!I3$_F�na�q+8w�Vy�bM�PˉOf2���w�h(�v�X`p��I�%����
�'�be���W�^4�ą�=W�&0�6!W
�>�9��T#�H�q�b.�bd���7^c�Xa�7&��`� =�:\:�<lO ���C���Ѡ{ր��G�	�lzV�Կ%��I�}\��Ѱ��d؞p�'��uh� S��	�H��H9�ɴ�XpK���L�O���R#�	_�$$�4K>���'�跖�1$�L��'�
qF(�[d��p	��OQI��3?��ӛCR:�Y�/��6�[���P�<��,$C�0�ԡ�(�ܑ+V$Fh�aq��!�:��1(�&����!;=��4��H�az򃈭z�X�A�ST?!6$��Ԡ2�M��ԡ3��^�<!���>C���x�&ͣL�L	c@$�A̓�( �(�3b��~%���p&քYذ�bQm�D�<9��Wy�$���<��LH�73�@s��0}�#������/_2�1�D[�~q�%i#L�&7��B�ɡw�D8{�׵Ey��P��B�y�C��B�\X��'��`ѫU�w� i�ՀU�B���ӓP��i�&V��hK~�s���,.8+��ξ��C��-a�x4�aE�n�|�ʍ3mrb�|�ƕ)S�����7Cj��adHKx�Y�3�ʜ7��C�	XXJ�F�Y�ʡ�R�[�6"����L��T?����F��O����9"��Y�S�{��ء�"O`Ȼ���4�2E����/gP�����;�<`J�&KDX�P� �Jg$���	0e��X�d,D�<Z��x�D3 �Q,%�J�F�)D�X�ˑ*)0:Т�Хd�z�qU�$D���Cl�T�Vĩ�s_��(U>D�x��@Z�q~HJ��O6G8|+�:D�h �
�(Wƽcb���d����3D�8�6͎1W<�{`K1�xxE3D�X����	&�8�r0�
0r���Pa$D��؅PWƶ���ʏ7����#D��B&N��y�}�pM�r�~(� =D��9gKO�z%��/G7\��c�O D�H�s(9x���beGk�J��5#D�hS�G�2q��A�=N�J�cL!D�� ��sB�^���yDU� '��s�"O(�,A��h�4��@�d@2"O�3+)u`�Pᣃ��Ҵ:""Onq��L�;RY����Y�"հs"O �6-�6u�Pp���_��:4��"OIcэ�6_�B�"�mɑClB-@"O����u&���vW7Ee�E�"O�(�V��h�@a0�x}ztp$"Od��$Ř�G�f('�\�YX�a9r"O~��Q+K�&�z�Yģ�)/G��e"OZ�Q���U!����@�3V�kA"O<(˶�Xx!��ă��*�t�"O<�.�4k=�`	P�Q0g`2*Of=Jf)�Y�vug)3T�U��'��*@��$?�T�Wj�R���q�'_�H�eD�<��ř4J��I{U��'񐕛u)�?���{d���O��Y��'�M�*��F¬��sa��^*�*�'+ u&����y�DV4��5�
�'��1��)иKj�"���>����	�'{T(Ar�:><�F�K9�Y��'Jia��B�z���:�/��$��'�<�X��S�NA�0�(U����'��d���G�[��E�2#OH�m��'�z5����?5��j�ŰA�r�Q�'M�P�N̪v���f$:��p�',�T�6`��3��!�v�:�͸�'U���,G��Y#�� 6�����'QZ!���D�4<�(����-K����'@��v��"z� fR-9�~�Y�'�jqj�G;L0�����"O���
�'&=��M�wzb��P����R
�'R$�6_Eb63��Fˢl�	�'��Hb"O(nlhzU�Q+�lI	�'�pe�v�IU� <D��ya���'��쩐r^��b�^����c�'�*%5JT���N&r����� &�yb��w�-Xq��h�D�1���yN��W�1�O��bZ%���ybJߨ����& �r4HIK&L[��y���^������bły�%�˱�yŗ�C$�,i�/��% �ÈA/�yr@�c;��I��&�"${#���y���sN�۷�J0tD�r @��y2邇�,k��+|m*�
���y⯍+|
�Bi��"�i�ѢG��y�'Ȩ�t`�@�r{İ�m���yRn2ŀ�a��Z2j�z%��(�y" �b96E �닼c3P��tǌ��y���&8���6�73�Z`($E*�yr�6U&�y�n��(��=+FŇ���>��OL �xC2Q�3ժ7N��蓨.D��PoFP�Jf��/!�pY�(D� �wM�3ˈ�0mʘy�d]`*$D�l('_�\���F���R�骁�#D��H��U������Zw��ӵb?D��ȰgO'���&�L�+���Q`<D�x�U���ITDX���n͢1�u�9D�8A�)� g�p�@
Ji����6D���D-}�|�)�k�F��De�2D�#F�Ϩ
l�5S�AR�2 (�5D�<���**
Z)c[�W�ؽ�`�>D�(Z`I�j�v�Ȧ*�?���2�:D��(A�v݂PZ7꟪!������6D�� � ��<|��%.�2C��\�"O��)Q
�l5��p�ź����F"O������JB]hS���ԬѴ"O�I�#BJ�d���9vYX$"OH	H���%� �����$&z��"O�J�J�[|DL���Y���"O4e:�+���Qz���(l�ly�"OxY	tn�A�a�1�T;di9b�"OXi�e����A�F	f���V"O�mqf��,�p6��
0RLyq�"O�-cE�?rf9pk��c?�@�"O>�At�	�4 �Y	£�28�nm)#"O�J�.��L�q�O��dX�H5"O� ��ƭo�0m�C�C"Rt�L�"Od؂�5{�a�d¦9n$��v"O2Y�!##�\)@�B�kU���p"O�$�Ζ8t.�i��ӁtCN�qA"O�a(�)�!=f�]�5�Op��k�"OJ�b�ˈ���7�4c$l;!"O�at�B�F��	��/\�OHZ�J�N���������E����/'#&�i���yR&H�+"�BeCL� x�B"ˁ�y�b�!T��욤�����Q[�Py"kĎG$���s��%5�{�Nz�<Y"���-�r%8��Z�u�h�ꤤnx� Dxb�00R���DG��e�"5�yr&ĿK:3`ݢRT�iC�c��y��G'[�j�j���L�ym�&�y��'�NL� +��A�<��'�0�y��O�+�Vl�k�Ks�9ar�M!�y�@��|��o�x�N��P�ִ�y��A�KN��� \��W��y�ؙ2(<S�"	fZ^<*'�֏�M��'�3`o��oQ�����+��m1�'�i{3���%d�
E�
����'~N�0qL�0A�!��@�'ln��	�'q�eY��W�*��dPq��W�`	�'��8���S�LR\0�D-V�.8�'Ѧe��3GP"�f�S�6ʺ�[�'��`�qɄ�R�F] �ě)q�|��'7,4	�HҫA��q��⇿ P(p�'e�����'>��L�a��8$>�\x�'T�3&Ǜ%�hhI��!��d��'���Q��N��'.��m��'����gJk\�a�/�z�P	�'�idh\�x�ĭȆ��@հ�'z�Q"@�H� X���e�B ��'�z]�!]H�	2��!V�̀��'�@ 0��E�F���釠b ����x��I�(�����YZ,�u����y"E��y+ܔê�5K��|h�����y�,~�����Z]�x������'�ў�O�����Lf��a
��P�b�4�P�'��(�ZM�����Bhc�'H�ظrJ˴|�	"��˸c�,qj��:O
��գ�:���$g3,�4j�"O|e��nKiʚ=�;I��� U"O�Q�@�V;&dxxY������'l��`��H�6&��1�/W	i	�DzB�'_�ܨ5�A�b�;4B��T�{���2��e��i� ��"���L��`"O���c�& ��P m�Kv�
�"O�8���." �8�E�>]k^Lt"ODa�ȃDy8�q1�X,Q:-i"O� �����M&~�NLR�)�,O2}	#*O�x�W��j�αP�!Up\I)�'٢`j��4�+T�O!Q���		�'u`1�Ck�8F�.�8Fl�D*�Z��6�S����j�\���߫T�t�Rӌ�
�yb	D�j��!F��S��r��ɬ�y���#�l���M�x}�ħߠ�y�F�{&�d�Gi[KAB���D��y�3h���'oA�J�<�bް�yR��"^��xǖ�G�ly��˽�y�NQ�:�p�ch�%=��ݻA�̤�y�/&-��`�`N�@��xpm���yB��0���!O�1����*��y�+��r�P�!����%��h����y2� d��T[R���$��DC ��yR	�#+��h �-�� *�i%┷�yo�x鸠�ri^�L4�G�.�y�f\t��F�9|N����AZ��y���MCt��Ȍ{�Ne!��R��y҄�|D����J�i���5�U8�y�O�\X%�b�17@�a��yB���L�)�f��2���	�y�H�o������6�)��P��y⡂ryXi&���4�d$��Y��y��JC�D�IfգyF�($IL-�yB���r��3�[>�$ЖN��y������ۢh��F��Qp�Ț/�y�DD�JITp�������y%�Ǘ�y2%<L�J)���I2b�'�y��ԣg���R��-)7� �����0?�*O���g��@R�H /=Qot�"OZ�Y�ҹ�����ɱY�`(!w"O�a�e�Qݕ��P�{��83&�G�<Y�dξ���� �X� ���[�͐E�<���	0)v����A,S�ċP-�j�<��?��PW��lܬ���GL�<�1	ߴ$.P�DO0hb|��*X_�<�����ZvD�Q3���.� �U�<��+K�iߎ�x�e �w��!�ɖE�<Y��ڒk��m{�oޟU��d��u�<!
��V���!�J�z�h�#��Y�<Qa �9&b���λ_�d���V�<鑋E�n�x�q�K�%���0��	R�<����o*��5�ȅKn8ѱMR�<�'nƉJ␩��|�b�)��r�<9��D�Z�KcBżFތ)���t�<��M�v	4�b�B�D�rQieMMv�<��M�=����nB�vu���Ee�r�<AdC�~�h\H�"�4��8��En�< )�$:�E�ĨWZPxK��B^�<!�3�Z���%{Y��2G*A�<QtD[��DT�N�h>�S�X|�<���X��6�ܘ4� �3#��{�<�jF�1��p��P9#�
_�<!���T�9A"�7Bz$� V��A�<���Flᮨk2N�f]�P0f��h�<)��5\�j {�S�fm2Q��fCf�<��ݸ<2�9��.D(.(��X�L�c�<���P�pxE�٫g�B�В�`�<�⫝��@ź�Kר-t"�!%�^g�<9큮!��Ja�էB�\)�`�<�J%1�0)rM��U?z�Іs�<15�s�q��'�X�
c�<��:~���j�UIj��uU[�<� ��@�����2�(�W����"Odѱ�l�4u��A"'E�E�¸G"Ox��DF�3d�0�£]<	 �xC"Of�y�c�:,Y����$�	i�T�be"O��X��4���â�(�(�
"Oڬ��ˋy�nl1�/�S�F�p"Oje�a,��U����JB���#"O>�bF��G��+�B�+aƼ1�"O�Q1�&AnZM��V�]�A"O�$JքؽP���a�@��s�&h��"O�E��KS�L���eo�-�D0C�"Oj	࢟�T��ʦD�/x�2"OB��T��7U�]�$�<x}�"O�� �X�W�D���t��'"On��O�pO�t�UI��%�[�V"Of0 �XO�"�G�K�0�F*O��q�逑z��X ���4Y���'<�4�!�%h�Z4;�L�<WَL�'e�QA�녋b͘�`�Y+S��ē�'R`LP��è%�V���f�=q
�'(����hL�zuv��V����`��	�'8�8�oM8n��tk��T69��
�'���z�H�4H&4h���K+)����'���B�f� ���i� \ĸs�'�����˄!Ξ���Z�$��
�'E�Qdq!Dh�G"
fdQ
�'k&IJ��ܢ+��<�d;��]s�' :�P�E��v�����@oM�5r�'��sD�#/pds#�/c+�	+�'��Q�m� cH���bE�$-���'R�*F��GR�����0d��'v6��0莥-���@"��w����'m*��O�=-�xA�A�h����'!`p�v�U((��%Hg Q178����'*�X8�Ƅ?a�`��F�/6�`(�	�'F2�c�͛7�*1Z�	����	�'HL-0�Nٙ]�Le�o�i4m�	�'�L��֪�4~�nu"r♐��r	�'8,��c��4{<�����A[	�'^@,�B�F�"����@����x*�'�����ĢPb^�٠f��h��1�'O�#R�2@{��k𡏳�*�P�'��U�fN� ����j=u:����'vz����p�P]��M�?x��c�'�I�&A�=�8�I��5��(�'wX�dl��n̜ Ǧ�}´��'�d1��`
�̌�F*݄p~�i�
�'u�r���)jdc�o�|F�	�'`��陾Db6��5��ml����'iV�R��ܚljpň�âW��I�'�$�;Alݴw4�G� b�9P�'Uzq�M_4)j��vG4i+����' ��TO�0B&Y�����e����'m�u�u.��_,��h�pَM��'���r�+�G-:�O��9�p���'ppQ�k�[b�	�MZ�r�'UȔRh��d�$M��b��v$��'%��g[�j�rIP K
����'f�[�_�G6��"7Ϧ(&���'�Xq��T�`���v-�--.p�'U��DN����3/�O_�i;�'�~�ض�yZ��I�c�22@�t�'�4���;u�h��+�!0nf�'�x��LܝL� �H��$�"�K��� �qY!��!.6��]%J��""O��)rF��8@h����Ϣ��� �"OX �����Yd���	�/��ѓ"On	C�su��U�7}m�"OҤ,וl�F�!���W�L��e"O�A�iX��[��R�Xk�}�<�1���EG(\���̓<�TE���U{�<	�(��e�ƴk�G�8j�p�F�t�<�#隿q�h���u���Ze@Np�<n�%^y���C�N*���AF�
B�<�Q/^&	� �Y��$�\U�Zv�<i�T�g ��:���#IoZ}�"K�p�<��iQ�=Y0���>��Q��Gp�<�A��j>�����Q42�Fa
 B�T�<�"�J<��{/B�U8��ׇS�<Q��0X=�S0+�*�+��N�<��l2[$�n�-"�B�Ka��M�<�cGУE۔$�TL�d�tHs��
H�<�v	��<��Ţ���O�6�� �G}�<���57,D��G�`V�mj"��|�<դצsm���AO�og�,*�D�q�<���&Zm��X�Á�>���+�A�R�<�d�72��u(��_e�e�P��P�<a���~�hڇ�@� 0�]#�I�<9�mZ1j6Q`��_�H��ʅ��@�<��bͪh�⭸� :càQ�Q��S�<QK#,/�� �B�55��D��	O�<YQ�C�VT��!dgX�XS���K�<IFˆ�@ۚY�p-8[�� I�<�ǏڂZ���i��Y�U��P�c^P�<�C/�&4���
�Vy2Uz�s�<���VZl8��_0���S�<Y5e�
&)B�.�5{9��\N�<�B���T]*�S���u�TB���s�<�c�۱a�p��&EV�[H�����u�<�U�_����
n�(S��E���Wu�<)Ef�?��5������ ��q�<��LX�\�V	d��
Plxs��x�<�qj�.I�D�,�2W��u �Gu�<!�m	2�X�1sk۰�2�+�WG�<�N#�F913��Yw ��w��y�<�r��oު�ґk\ P,mzծu�<Y��h>����Y�r}"�bKo�<�O_tA8�K1�߿a&�tҕO�A�<�f�9k��JǊ�"Y��Y���U�<�Ќ�;b�[&�.��T���l�<�E�	��|H���U�&�a�#�T�<��K8M$�h1mȗn� ��u�<�6���'�L$�1
)v��u*�o�<)3n�W��:ňM�A��k��s�<YV�BК�j &A����R$�n�<a��2&�%k� ٧���P�L�g�<iCl�,-sb���^%YjY�ï�}�<a�)�Onu"Vk]�UP��2hu�<a��K�|T�� Sֈ-�7%�m�<�e��!�h��Tۗ*Ɍi{#o�`�<�JQ�*=��@R�ks��jS�B�<��BŲBT�:���A�X��J�}�<3�C�.1�� iD'��E�w�<E,�G�@�wLJ$SĘx*#GJ�<iԩ[�t0ѹ�׹o��mr��[�<q�,�p���g�2.\�n]�<!͞	;I�|@T7%}��a��<�GK��)��y+��C�����R�<� :��榆�;�jHÀB�&��lI�"O���m�uz��"�"(��H�"O�h)1��G@ ���A©A�6�B"O]bb�,{l�	[���¹	�"O^��7��qB*9)�/�%(+�I�"O�M��ʊ�d\9��Pp�d��"O��$-Εi������H^��C"O�Ԑ%NQ��@�CeRL�j�"OB�8�/�Cpz�K����2�{�"O�@���&�X�r`f[�|�x�P�"Oz�1bi�Oo��ðĊ���e:�"O����]�|�҂�?�2�2#"Oft�P���Z�Q��Z<�(�b�"O�,
�j�|*@y��J�qg8q"O ��$�?�\��hMOt	7"O.�hHm��:�i�{C��"Oji��%ӞF��t�ӛ13���"O@!���?[2p��@��Jx�"O4P�c X+��;�٘d�̐�"O���B-^b��̓V&1\L�"O��c�ł�2��� `jmZ�̂�"O�q(���hS��s�	�n2Ir&"O�0Z�%
�z�jϐ�6O���W"O�� f�5�P��ş�(<P%X�"OP�SS&�4b]bѫcW�5<�dI�"O��p� �d ]�B!��p+Vmj'"O���錵|�8rb`&��c�"O���3��73���`M�33S�)YS�'�ў"~�e-=OUn5���9g��=�!#���D'�S�O�<����f��%!ƍΙ!��r���'����łA�fP����>9��)
�'e&�F�:Q��Q�$���h�	�'i��ˁ&Q!Ox�%�F*��kR�,A
�'��<��OU�f!��k�@�1��I��'�H� �&x�V�֗��L>I����> Z���K0�4LC���,�!��S(��95�x���k#N݅K!��\��h�������mÑ��O"i �*NC���YƎY�x�̭�G"O2H�Q�:���[g#ü[���0 "O>���7
�樘4�ώ�0���"O�Aё@N�l�Z��v-�J(-J�"Op��NU� Zn��"�_�<�`��"O�͡à�mˌ-xc�S�L��ɠ�'0!�ĝ�H�*�ŕ�L4j�-� q�'�ў�>�scS)��q´��%�i���,D���סI(,��{7�֙K j	˔,D�L�S"�6uL@��@ur@��-D��%�>x�q��Њ�<���`7��c��@hs��
M#�����	M�R+2#6��]���¢U�<@�0��/8.�A�/D�@�2���V{��?53�	�C�Od�=E��4Ojq��� ����ـ�*#��lX�"O��(�d?ތh�JxizW"O�c�H����Uj
وv���R"O����%	���p4�Ս3�ZH��Y��F{��IF l�<L�g"��:K�ܻW���da!��8�N��j�
6�8�F�](>!�ݺK�JՋD���*<$������]�z���$��B�`���>{��a�ڝ�y⭍ 
)�Qɓ�\��t���yr(� 0�v����B�7�y���l�P�c���Vi��
bF���yr��� �eFU�\AqKH��x� |ɉ5�I�ba�zI�6>���"O����'@�!,���'�l( &"O�A:wn�2I�*��0��$������!LO���Nڍ2M��7�(Nh�y�"O����蝆iP"��8dŢ�"O4��)X8�ZV�X)I
��Q�'�I�w3�1rԠ�P���FǄ�p�B�	\,�}X���<$�}���҈U�y�ɇebb��J�l��@��߅=eh�O��=�y�L݊6�J��1�*�>��G��yB���"̎� Bϊ>"FL�����yr £@%���v�oi< ��y.@P�Ȑc[5e�X5�f���yRLW#\���AP �Y����k��x�'An�H���Ϫ�`��0�؅h!�דc@ +3jB�y���pr(,,�!�GEQ�l*�"�F���42�!�$ƳpC��I󡔃n qd�M0F�!��N�d�:xe+����+�h�G�!�Na�����X�P�ʃ ĀY�!�DL t���#��4X��z� ��$���;O�zU��EL��g�2���Y&"O��c̔�e�ڬ�&L=,B�4�$�<YO>�˟v�b-< ��+4h�J_��C6"O�$���
+1��D�7��Vb��"O�)rŊ��-�8���G�h ��"O`u���g�*-0�HU�xfI�"O� G��$ꤔH�GZ$eP�1"O����n+V��zT�:X&]���	J�0、�zVE��%�"n�⼘5�8D��0g�3L��%�G�d��e��!��������F#(xa"h���'�P-0�f��q�kЧ8Qo���'�X���a�#6Tp�fTB�t	��x��'7&��qB�ѓp2|��Z �yLK�%6�|[�
L<kXZ�@�h��yb�рa8�����0�h�S�yR�>z�.i"i��u�|��C���y�I��AJ:pRr��Q���y掅7�NU��gQj�8<�^.�yRş�^ώ��@AE�f�<��(��y�,n9�����,Q����!���xBI�(���S5�@9i��� �N�'&�!��"N���D;���� NG�!�$_�l|����LZ�+c�=`��@��u�`��7E9B��Bֹ͚��ȓU�\�W�sC���c�m����'nd�[�'�rQ��쒎g�����'�!a�O0�|�c�G/[�9��"�'.�e�r ��t%��,��D�s���'@��&�Asq!�f��
2�	���?��*��.uX���O���"O8:g�܀� ���+��1�h�"O�U�7O��JܮLZW�B���"O�᧧I��qv��8�r� "O��ʁ���T��WiȍQ͎� ��0LO��:��k��!s��>M�j$c'"O��qK�����C�D�<{x���"O�����ػ8�H��އ%pX$r"O<��A�1�
1�l��XQ���"O6�J3/Iej�8��Қ#?��u"O����mΛ�)���� ��"O���R�O�@�6<����
>	�a�"O,xyAk�2��v��)!��}� "O� xɳ׮�͖ш0o	�F8�"O����
O��f��V.��lX�҃"O��BQa��HHb�,{��x;�"O��{Ӆ��wz�[��f[�D�"O(k��"òHC`�=����"O �r��(K���Q4Ꚓ!�N�Ӵ"ORM{�eҌ ��8'�D�X $��"O��:A�^�X�\9�߄aj�80e"O�j���D��a�ӦH�H�ޱR�"O�\!c蛂Aj��y�F�"�	�t"O���C!"����F �)�\"O��/3f�r@��΄��č��"O���hV�k�H�RX�v��� �|b�|r�7o�,�J%�ђL�-��Ȟ�BC�	�<��)�F�V�A��Pj�C�yY���4 \\|p !�@�!�B�1bsR��A�KMD�����n�B䉲���qR��h�L�=1(P���d�������=b6���V��ъ!,0|Otʓ�y�OӦ/F�:q�E�I-�Ȣ��&�y���}P��2R�
�A�4�04����y���(��H�AU�<�>�TE0�yBa6]��}PL�7Uu�O���y�MÖioT�5/;Q��yiJ8�yҀ��]C�i����7���*,O��y�J ����ߜn�q0�jд��3�S�O,�lނ��� ��v���'�b�AT3+È�aգ�����'�)�A��'`��B~�BA�
�'�(�C����)��p`�	�
�'�%!���.G�1`�K�b"��`�'���C�O1w$$�����8Y�*y`�'DB�aV��	�l�gϖ�>��99�'�B�{�ʟ{�D�&��5BCX� O>����iý,��æ[*9���#��.e!򄂯ń#sA�#�%b��!`�'+ў�>�! iD,k7���eM��cQA�@%4D����K�\�f�I�@�s;�C�$D����`�'^2��j@��s���"D��H�C�t�`�
�E��|�0XB��O��=E���E�Z��l��j�V'�u���:�!���.N�(�3��>���"0`��W�!�D�&r�� �J	)����sM��P�!�S3Jgz鐀&x�(�/U�1x!�d��Fؼ�Q�ߡI�*�����/{t!�dN�Cl��BD�$9~t�!�i-m!��*(�,�#f��Ja��C�_3:Y!�Ӄ+
H�A�BԿ!�D� ���WS!�\�+Zp2�l,v�z+�n�2$�!��$(�B�RSLΝs�Q7䁀��'�ў�>�8&/�2+�Liਖ਼3^�$u3��4D��[p&ٞn#ny��-�5T$u�f(D��#� E2�J��t���)�Y�(<D��V�[�ie�l�,R�AE2QJ�=D�TWiEff��zE�]�C�0��<�	d��k�ƟO�6S�ɝ�xK�![��9D�0���ɯh�#M����Ҫd�!��20�pgc��*C��$	�!�!�¤=��8 '
8l�13W��J!��?D�%#�oX	!$�82�Ζ<�!��,����$��Ya썡'S!���/C�,�'��'`I�'�иM#!�D/p�3 ��"3�j��tm��
!�o2��r�j${�6�D��u!�� =������!��@[��B���"LO���՚n2�lD�ҶXs�4� "O@{�@yrܥQ,ɺWkt)�"O�!#���8(BA�U
n��#��'_�d��Zy&�Y�(�P��dB��FS�!�dK�=�BP�'�@;_����*9S�!�D�+lT�"df��$xbń�!�W�	�T	J%J<"4x��,�k&!�$@�3�6H֏�� 2��`,#Vk!�ʃp;H�Pr�`S Z&�ջ5!�dH�H`�2��?4AP k&��3!�D�>���hׂv-.e�l�3!��'x���p���#z�jVAҎg`!�$�;1�R�����X��!p��M�9]ў��S3�2$)���Y�r]{1�$m~�B䉬~T(P��5L��`�FwhB��6?�~���ǾQЈ4#p�"�R�=9�'�d��C��,w�8S`�]�v�`M�ȓR����F�]NX�bVoߋ=y@u��y���B	Ӯ)�lt�F/PS�tX�ȓ�e %'�<tb��2�֊��Ą�,4ƭ��E��N�'iT
?BNԇ�>�����`R���h!m�Nz���?�zĭ�w��L�MU�^H���j Ys"�c0bѡf(ӕ"�؆�IH���́f��@9 G� ȓM�
��T�J��
A�ʛ�T0���s����R+�mD�
o��ȓ|��զ�!�h�G��z�5��3�&,�DJ�B@��� ���iO�	2L�S�,���cX�S�̇ȓrb"�T'a��\b��0#�~t��6<�(Qc�)G�j�I�k�� ��1���Kм	�q)�#;|��|%}�4�$̲a��ND�@���wp�y(�֊s���H
0���ȓ02�x�I��y�g�J_l�ȓK�`��ƀu�0���%$݇ȓGT��*JДI3iP3�`@��t_J�7�
�d�:�ǎ�{�bA�ȓ2��s4M��i�8eK�/���ȓ$�,��nW9 �����#�0���G{"�']JH���(��A��/"�&�)
�'�Ą8Bm#*p$-C��ճq2nb
�'��{狏W!��zD,jQ:r�'�vb,� b��4�V�c	���'lX�ȓ���P��3X䈰�'��p��b��(�q�ٛS�R���'h> "�>$��|��j�EP���'���`TfD�O	�A);	��'$D@���'�� ���7E�,r�'�f�Zh��7�����N�+*Nȝ��'����@��:�Dѓ�HYWδ1��'پh�(B�L���S�FwV���'T���'1Cc�0Y�IԞ)��F{��O ̹H�H�%fK�J�K:�P��'3����2`�d�lR�[�@Ap�'����7!���d*۹W��(�	�'5t���G%E{�a�@Ã:����'XB�;�C��`P���N�2�T���'=X{�BL�::�R3h2uz��
�'"���%"C̀ �����V�P�P
�'6�q0�d�JU��kD�� �v@a	�'��9�I�#}�>Dz�O�F{p8���� ^�1@�Q/w
@��7:9�6\4"O���AH�%;v�R�Y lێ�a6"O~�0i�	J�����f�2T�$�{q"OB�
�*�- �vP�(1�� I�"OT� �JҵZ!P(�B!ۻa��ٰ�"O�5��D�)*������!*�y
T�|��),6"�p��� .�q .�K�B��%Gc(���L� J��u�A+�6oÊC䉍d��������J⣖�vw�C�'�H�a)	�.���Z���h���=��PF]�"!+{H��۷GD��j��ȓiŲ�����K��H;*f䕅ȓ*�~�f��7;�@[e�j�ֱ��:h;�I�M�`[q-�h�}F{��'9V�q�dE7%"�"�)�?.T�H�'DP���̗n��(�5�C$�p9�':�ia̚�g��H�ݠ|+�Ku"O�����N0��B��<E3���'"O�T(e��3�f��*[�&D��"Ot����Hk���K�A��u�'�ў"~j��#jkʼg�S�T��ȡ�(��?9-O����g��j#�9�|,S�I�`����^��͢e�ĸ�F� ��ϕX��ȓeN�� %��, 8���܌��A��Q>��wK	w��U��dB��B��ȓ4�|۰+Zu��ݺP�åY��h�ʓ7�!�Ǫ�\�lQ �a];�@B�ɺU�L �ˑ7�2�a��5;'B���Y����&��`���᦯˚I��� D�2D�@.e���;R �?��)�6��	!�$�:ab�pW�6�]`Ձ�=m�!�]++��
C�Įn�<{&@ěo�!�d9=� D�&CM4)m���άg�!���@=Z���EU�A�F�t�!�$�	�Х(�!K�DOj�#�L�9�!�D�iPx͒�nթ1�	C��v�!��E�i���a�����YG�!�$KtN��V�O9#cfI��%��6�!�Č�o�:��%��78FJ\�é�!l�!���/3�	��_�T⭨�'��I !�B&k��	���2Y:�9gǞ!�D�q��Zw��'%�Z��e)V�!�D�7Q��À��'����EA�V�!�_�" ��)!JQ>S� %��F��/�!�F����U���R�kRN�!�ԛF��a勅�x?�U
��<�!�$	�J�;%���h���(X��ȓW��P�����-�*��cb�.�6��ȓp�IC��*&W\��ON�O��܄ȓ]��1�%�P#�x7bK8/6&X���R��Fġ�ihm�>4
�D{��O�mp3N2.�z�8'c|!�A	�'�HQ�6&8,ap�VCC�CfP���'��(���C� t"�h�;S�T��'Ħ�{�㉄Y|Ja{GC�Pw���'M��A䀨^/*13Ðys�eJ�'j��5�	347��;2J�5����'@"#��؈w��gJ,O,�p�'�]�S��>~���� ��XY���'���ɇl�?t$I��RJJ���'8�Ekf	�B�إCC?4o2���'݆�X�f�1��#5iC!+���
�'����n� |JI��苶�28�
�'M�*�&Ƕ�>ɑ3��0h���	��� �����_�In�����^)ON�R"O��`�N�5u�nE���J�0IZHAd"O��S�,�N<Y��C���04"O��������iӃč,%��9�"O4�ɗ��#6��K�bEY<�6�?D�D{���7 N��s�Re�Q�&�>D��*��5�I�oߝy�r���/D���D�'_�(�v�ް,�P���$,D�H��c� {�@<!��@�^�� ��>D�Th�ϖ0BZp�t��8 ����l)D�̡`i؈d�B�ײNhD��p�'D� K����@�z��H׹z%<9(5F$D�d�'.H�r�)3�U�1�i� D�0rd�1[w������M�f=D��Ge�Pr~��'�ĩGґ"ō/D��0��O/��a��-GB���� D��9#0e��c�nA�	$��/;D����L�:?� iV"8��Ex��8D�8�`N#2&�$[��I{�����4D�`��D�L)��@�C�NS��8f�8D�L�ᔂmz�l	V M�����;D��be$�����.F
d���1��;D��9v�S�+Dy`VK�!%z@�D�7�O`�.��q���P�I�$�@��Y|\)�w!w���J�cg&(�ȓ{6�<	3��`M�8K&`�,B������G��l��y2�	1u��Ȅ�mΰ�ϸv( ���+9�$��ȓb����� �%�x�x$ӤZ�f<�ȓN�� ��ͳ(^�Ю@�r��]��06"�@�.	��x�R�@��h�ȓc�f�!�*ߙi+��%�L#zP)�ȓ}+rX*��/)���H�'�d��ȓt>}����4����o�<rv���,0X���V��q�# <f����P���0n̍O����!޺9�0$�ȓ[?�LZcbT:WE|MsVF^�
5"%��9^��׃M6R7���p�h���a��q���_	D+��C��J=]����ȓb����OҊx�*dk׎=��E�_�,�|�H�9{�z�N(��x�F�N�<a��ͬ� ���ʮ>m(��Xt�<��\�>��!	 #�y�C�[�<��G�SވHkWił�쐺6��X�<I���<�=��cؾ�n3�`�S�<q*�m�~,3B�ٽ4�b�"\g�<Yd.G�G��+w�Y4
�\)H6Ϟax��GxaH;6����щ*/��u��,��y�%.m�<,ĉ��+P$�/@/�yroB"V��Ҧ��*�Z�����#�y�g4)?��Ʌ*�.)����0J��y
YTY�����8!4��g*��y�&��
�� �%7��a�F�D>�y����Up��o��{ޱ�s����>Q�Oj����Ʉ*����_dV���"OV`�%\G銌��/��Ye�B"O6�rwb�;�f8�(�S��d34"O����d�U������3c��iH�"O<lH��Xn�Q�,��-��9y'"O4<Y���9�U��_�b:����X}�<�a�B�������)Ų]�ŇƓR��0#`��Ӽ4@�@\(Q�*��'/�Ek�*e0�Yj��ˋBK����'4�Psd��<vX�G%�)@�~l���� hhSO�$��ЮM/
���"O���듅c�����ʁ�%"Oکע�<J��\*�����1Cv"Op5�6`]���C�� D�~�"O��Q�2�hI�A�e�F	 "O�`���B�d�sK�2|��y��"O��A�ʑr�q�$��	L*��"O�Xj�܀1���V=����"O�cS��%��|���&�x˧"OP,p���
�긪g�Z��~abC"O�y���e򐈠SLZ�3�:Р�"O
a�i�u���y�Ȏ���S"O>�A�_[4��S��=���T"O��;aH�h�|��eZ<��%"O��a�Nϥi� �3Q%�%D�D�)#"OD9Yq�':RAqVK�6��!`"O�e��K_ƄՓT)�*u�H�"O�s��I)�2�!J��^�(j�"O.M�R��/Q��հh�*~O,A{"O���p�@�K@�<��T�`��"O찠����6*��2���	7��)�"O� ���/��,.��E�!"O�8��ҼqN�	�r瀫:Il�1�"O���F
۶7,l�擽s70�"Ox�9�瘝' ak@f2'�)�2"Oڑ�U�%@�&�$5*4ݡ�"O y�SlӘx�N�S���P�"O�!�c�Ø9��"�l�,�|���"O<��6�m����JĨR�j�{#"Ot���[
O3�E�RDܛ-�F(Q�"O��LV+reH<H��Qخ�J�"O.	���
�`r��,VvR��"O� ��o4T�p�!ɺO��m� "OV�aUjHD��eF��$��$��"O8�"-�04��-��L�h��y��"O�k���q,`�U�H}
���"O�Հ�
��=Vj%�q		�
d~U�G"O�HБK�4�T��K�A�X@�3"O�A���˛@��e����/^��RD"O�d�����%�ebw#��Ĭ�b"Od�j%��KTذ����!H���ۄ"O@���"�@pV���S�4��|�R"O�$s�P���j�W����s "O\�:d��rȾx�1E@blLI؁"O|Bŧ��'��c�mQt�"OZM�&h�@<-2W�W�\BhiH#"Ol\�҉ƙ-��Ur��1�U�"O������x��1�c@�9Q(�\��"O��q�G�-x䐑H��<h�"O�5x�X"w��lS4�ֽj(�X�"Oh��o�%EU�I�&A�_�.lq�"Oذs��	ra�ǣ�>1v��6"O
I1�!��Y����a�� ,�4�x>��rM�P���A{�F���&.D�<B�H@M*$�D-��o}�)��.,D����=}���E�r���j�8D�̐�`Z�S�nt`C� �=dB$�QL5D���C�՞c��	0�ę�=4�y�%5D�##4G,X�h� "�mY� 4D��ʒD�R�<"��gb���/3D��pkT9/�D�2��k��9zF1D� �!eȿe�j%I��1Tku���.D�H17L�U^0�2B��0�4�㴧(D�L2#��$2��x���U�4�vB�)� �� h0@����A&�
AT���"O��Pf	ʏk.���  
0+944ɂ"OpK7*�sT�ѱq̐�.(�$��'!�ܐ��ݷPvh����<	f��U	%D�X��<��r`Y�]du���#D�\�lINz5���9��H�j"D�� �!�%�����!.$0���;D�p�E瓬/���:��X�"b���),D���lX�^��'�&#�&�:��5D��"�kɯ0&����#�8b>�Z�9<OD�$?�	n�Ȱ���S7�iC�(L,)�hC��sY��`�ʡk���0��
��B�I'4S�-�dg� T{\Z�̆8	<�B䉨t�<��f��y�1|2�C䉎p涰K���<}�A���A�C�C� t�H�����6At�p���^�C��,5gPhC�ϩ|�p5a�
.8��![E�=� 
/%d�3�Ԍ1k}�?Q
�
�N$��'ҍ[��)��A\��u��SO�`r7�	��fR�)P�0|���!�l�i�)���	��c�bą�C��膊�b(^hI4��]�ȓ(<�x�*A%�*`�HIi��y��-�QibE 
Ʃ	�
���Q�BѢ��4lZa
�#A���܅���L�T�,m����.�r��ȓk����S�385S�-:X/N��� -"�%��1e^i��%�f�* �ȓ<*( ��׎/W��(�Ɣ�2Pи�ȓ*�&0�	�s�x���G��t�8��2d.-�SW{�j�c턚WWj���f=`�@%T�[�>���VC'���Et��KB�za�H�h�4����ȓDqju�dNa�-4��\S&�ȓN�4q��
�w~�P�0퉓�l ��4�����'B�sd����ʊЄȓQ�h��B*���i�K�+T�Նȓq����U�Y�x)WNI�0.���ȓiB�X0����U��c�|�j|�ȓU�T�yp(Ҵ��l�"ɔzv��� ��신��1<�>��r�?�Z��ȓ.�,��dn�.��,y@�[.|͆ȓ�=��n��!�c��	�ȓJ�a�WY�rɁA,�S�6Y�ȓ$w������n����I�i�l�ȓ9Z�a��Iօ)\��BbfN�4����E�@��d�N.T:�}�E��$�^��ȓsv��I1��1Y��������ȓ,��m(s��.:��>��P��n��8��^,�4�rLޤb�ZB��t��9� V��x�Ɇ�n�B�2a¾YӔ��CY��ѢG$b�B�I�t� �C��W�ș�&H8=�HC�ɹ ФM�3�C+=���@�J�6��C�	�f��0v�ҏg�E�a���C�	=n �XR�똞]G�R�*N;�C�I'U�V!��CAY�D�
��L�hz�C�	 GS�LҰ�S�@���(p��0P6zC�I6F�fPB��2B��A1\$h�bC䉗�\�(�3}���E�)[�2C�ɾ�M����\��fH�)��Մ�g�x�@�[8w��E���
>f|�M��L���Q�&�)��1�-�>9'6݅ȓ/+�`�+����Hr��?� ���S�? 6m��Ç�^�H�R 	�k�Ҁ�d"O����<]q���qǈ�>�^��"O*	AԀ�4D�,Sл�����"O�]&��4����&d	�����"O�B��)H6��#��Цv�CC"O\��f���a�	����6"O�	P ע4z�𮊝)�}I"O`L;V�9{L�!�L�A0�"O�Hs Z10�� KULɏ7�ira"O�M��Ĭz���@ߴG"�p�"O"�铈ݟ��E�E[�k�@@�F"O6%bE*5R��ip
_��v�k"O�=����mw|(�(��^\���"O2��s�/t@B��?BE�1`�"O��hq�Bxu�#����~ pR"OiK�����:�e�L�F�S2"O8E�W�o(H%['�J�4oJ<��"Oz�A hG'��<#�%c��a�"O�4ˇ���*n�
�SJ�}:6"Ox5y��K9���QC�6P�	0�"O��*4$ZN"\�$ �b�	0�"OԈ���"�0��e\-Q0D�G"OD��O��T���"c]2W䶴�%"OԃK�$�\��!�>@��i/�y� ��LSB$84�����6�y"l�1�V�1�ɰ)���w�E��y�3iB<k��Ŭ)D�!ҵ((�yrς,\��y���� ��a5K���y��Ӎ9N�A FˈK<$��$	���yR��8V9��G�=�r����N��y���#QB��D�_�4�:P�-�yr  /�(��F L�3G~Xhb���y���fO�CR�^71�ʌ�$�$�y���
��Iq0��.�@ ��޵�yr �Nwl��G�)m��L�y�Z��T�7�O�(��C���yh�ȞT�غl~��A�ퟣ�y��ӱ=��@��=N8�t(UIH$�y�LG
�Zq��z��J����y2n�	o�Ŋ�����i����%�yB�ޒ98,y�kǰOݤ)"�%Ƥ�yr��v-�n߇`4\3Rm�*�y��	y�!r��^�!�ݢQ߸�yr]2}���T�Ķn4��@Q`�;�y�	O�"�����c}A�6�y��ߨsq��#�Y? d�1�M�y�)V�Dg��*�X� ���p�i�=�y���w_:8Q����u�B`�C���y2�q;����s-Xm�c���y�͖	���Jg喞:������Y�y�`�2J�.�*ƊV�,�\lI�&�y� CTTL��D��W%X:��Ά�y�披a����3�+K����գڪ�y�G-Q�x�ө�.?�\��W�y�H�	,&!єa 40�\���'��y�M�/{�0���A"8��˱���y��$w�ܸ�lP�P�N��O	��yA[誰�E�*E�P�!<�"C��-i�ȸ3�V i,Qo�"+��B�ɸ;�dp�͜��qsTF�+��B�I�g���A���0�����G�!�B�k�8	3�.Q�p���R��b�B�ɷ4����d/�EeN���&bB�	>Y�@3���B�>�'j��(B�)� rԩ����QsP���p�""O�!Y� K�c{`�U$�
�t��p"OJ$�R���Xt B ƽ�
e*f"O$Ejg�A��@9H��L(d)�4��"Oj�s�� '�F���ǁS��=@�"O,,�兊/�jI�@TTux�0"O��!th�a  0Q@�]Y]�"O"D:b$�lŦX �oR&WRD@"O0�P���z��0I�+NjH���"O.�a@h!�ܕ B�	e0`���"O�X�솤>J��W�ܠf:����"O����IW���8!p�Ϟ!-�9��"O�i�O�&
B� �'Y"����d"O.rc��!WÞ-���<1��j"OxDS��N���	GD���Z�q"O����j޿Q�$����=N�PY
�"Ot$2.Z�4��Az��;O�`AF"O`HqEoM�U�H亠�)!8T1�"O.�iJ�?�0�)sE�9 <�;�"O�`(ժˏ�T� &<� �S�"O�h�Q��	N�-U���;$�7�yrjڝ�6��Ȍl�8��l���y��a�ŋ�+��b킅��E��y��iM��*���G�DPQP��y�&ɘZ��z�L�*���ρ�y����^}[�慮W�"�H��yb�A7�*�:$k7S`$$`���#�yr!M�*:i&E�@����	-�y��P�_"�U�7��@����#��y��	N<�����5M���ŉ��y�V+Ჴb d�;/��H�BRG�<���J�G\:�cs L�t��P��^�<�B ��2�T�@+�ţ�'_2;�C�ɩ�ځz�m�
 Dy���۞.VlC�ɜyv2aH�i_4iG<mJ"��9Y�C�I�,��|q��%��R�"�8�/D��!r ӏZ�t����e2�k+D��H�E����̼*z�X$O&D��"����4���L�3G�*'%D�� �ҕN���Q�cݳ�r���>D�� D�FP!p��B1``i�>D�dI�e��.
J����%P����)D�d�T� �RJ��ア�2�����+D�,+B�@�%���T�W9^�<<��)D�`��˫x�(��dԗ��5q�()D�8X��L�_� ��EqA�dв(D�l��6M���Q�m������$D�4bB&��G���	�8��8�,$D�8H6aE�*,S�ș=�@�S�!D��b��B�kl���m��W���"G?D���5�ʞ-��MX%L� \:P���=D��S#bE�6
�� �%�� ��C�7D�4	EK�,ip�H9��Vi�pd�)D����'@:	q#��T�-q��Sw�(D���uF�-R-x�W�&��ts�'D��K�Ɏ�.tHզ�3�TI�m2T�Pq�AT�)�$��(G;C#���e"O��[���<N��ggH���̀"Oj�:����{��ग़�p�҂"O� ����T>��rař���{�"O���c�3UXn�w[*[)dEr�"OR<�C!O�3v-(4�Y7y|�)�"O0t9��M�K�NG:Q{�i"O�]Z��S�l�*�.�>�4�b"O� .����*��@ N�=K>��7"Ov�0r������^�1��"O�u[�J�G'���R�Ȧgs� �"O��3�Oѷ�~! f
T`�Es"O���s�(5���ֺ$��xr�"Ozx�բ@�HT9KU�F�D�"O����2!����/���X1"O"BC��r:}�P�Cd�|R"O���߃b��ɉ^�4�v�rs"O\�R(�"-���`նq��Q��"Ole�%��� �K��'&J�{7"Ojh�Pl�;-��%S -¯�`��"O(�@��<=��2�+�-E
u��"OX��i��"�C�̓#��H�"O`4�1���L�ʗ�[4X4@�3"O&}bj�5a p�#B�qɌ�� #!D�ȱ�Gz���I7t�4��D2D�\�G�<v,=8s�E9�
�Z1�1D�!��]�>s��Hv�e��$D� E�߷0�djLY�kڌ��e$D�@(Bh��X8�#�*����ad#D�,�a��*J]`�Hւ,Y���7�?D��S�On���c�Α]7腡�� D�lh��F���كN�=c���`"�#D���T�;W�\Q+�@fۤT���'D��@@+�'�^Y����#Dy�u;�9D�<�UCV�s�9`ү��N+�8@Ӡ,D�$ccG�'��`�SI�vК3,D��JK�#�(i�*K�~nV��@(D�hapϝ�D��µ	�+fN`��F�%D�x�`�^&v�Жj���Zk��"D�pR�h�
=|0���Y��a��=D��(�`}_�=H�'@(2 h��;D��۠?j��2b���%D�H�6ǂ	d�6��oB�Z#0U�W�%D�I5$�=>��<I3�_	ac��18D��h���)G�}���&k �5D�A�e �J��e�o��Q�� D��5�E*\��U+T�'. �)�=D���v�W�J��C`b��a�h=D��h�/
�t����)�Z���R֭<D�$��]�k�H��׍ߤ?���AE+9D�dI]rF�4��Y<d���O��!�D��Q|<���#W�bXi)VhͯH�!���&��9Y�!�Ա0˸o�!��ƄG��<����;:�E�I�T8!�k4� z���1B5��d&�o�!�!;'0�j@��5'�`Q�E�:B�!�dϯ#S���'�$>{�ݐb%2!z!��
��1H�FF�B`�,[&#� �!�ƨM����M��b�ys�S`!���i�:����#��j���!=I!�$Z-��d �w�\�����%�!�$�>S�%�C^��Ġ�!MP�K~!���S>�(��R���+"���#!�ă9!����� I�eeDY�7�!�d�j�K�g��(;���b�,�!��T�-�����_+��A	��!�$ݍ{�t��"厫aJ�Dł�9�!���&%�����_�|]l5��Lx�!�1A������S tH���N.�!�+|�hIH_�Op�hYv�n�!��ɲc��ݰ�Nވ.I�,�r!R�q!�$�n��Q�i\%�28�p#�=!�� hի4��7�x8Ã*=x"OT��e�>hتi�$Yx*�C�"O\��s�p�(���:�H(�"O��R�
�[��S��V�"O�PR�O��Lz�dh�	594$��"Or�c���,<H�E:w�۪$`a�"ONx��f��6lP`���()�|ف"O���(�;0�m1��	'<:��)"_�����<�2B-9���s����e���V�OX��O�����2:����eo_�T��2�"O��ી�I���s�X��tڦ�,\Ob|�t�T�)(�)���R"JDQ!�'ɱO�8rA�9H�����	Ϻ@�M"O�٢���o���x�h��*�<�b"O\}ؒ��l�Q��}���A"OP\��H�9.ѳ��H�C�| ��Ii�O��ed��[L\�M�@�x�	�'�8��wC��,�dE3DX�2'�Th
�'44׀A�>�(�n�A��0
�'��4��J��n�J�O�?�6�Y	�'�Z��AfZk��Xz�GL�Y����#OMA�n��ՙ���=�2�)�Z�X��I�80E��-��j�B��R����.lO��'��5"V���X��I]�V*4�
듍�����,T�A��+�L�"���|��1}J|�OT$ap �8��Ȑ�kD.X|�0Y��Iw���ɓ�~w�� ��^�x�f�h����M�����,�����!J�]مF	� ~�  �¥W����G{�x�l���[+R����s���-�X��=D���c��.�H����C���m���6F隍"G}��5�Aլ���)��:��-zE�-�p>�ܴ��dǪ\�L4���D
νȴ+�m��D�O���$� ?�ҝ������J�iX�qa|��|b��8���kP
­l��Z�o[(�y⫚�Z�=*�M	�8�r aZ-�y2�5K���xC�D��q1�
�y2�>/��	��Ɩ����ّ�yr��n��|��C&N*ƵZ"����?�" �OdU�C� �ɀ#⍍s7�9�"O.̚��N$.�b� ߪ'8A�&Z�|D{��i��!���V���CEC^4A�!�V8o��h��4��aR�a��:��d���=���ٟ- XI����c(6D�� N9T�!�d�.�%9d��!V�T�� �!���P���NآB\��E�j�axґ�$'���_�^�ha�i�<kk����j(D����'��� @��ϛ�6�����)D�l j�. P��#�m��(�R��(D���C8u�<@��eD< ����� 4���� a}*�hLW�6m  ����~�<����h#�q���[�eGt���C�S��i�0��h{*l{��{���8 �6�6"O�WN˔w��!CH�
�D�в��G���O���8�

'߮��CAؗ?�M�	�'��H� ��P� ��Fʚ+�Z	�'t}� ݼWw���ա�N���	�'j�8��U�K���˧�0`�@�'�T2� �E� ���n)C����L�R}�_��S�'~d4��\.Hq!V��!J�h�rs� "Ar�C�^C@���R�w2F���L�-���C؟̣�
X��6�e��<^��D�=LOV��$I'w�)�2�?T� <Q2�<Q�	p�'2�P�H�<.�l��c�.. l[�'�J%���j��Ӗ�O������� Xr��.C��{�bE�	��e�b�|�~zǥ~�����߭iY��'�ě /��;D�@���GEJ��&��n$#�8�	X?	���O��P1$���y��1*Z�����'�X����$�,�%��O/NY��'{$�Dy���S�w*��p�;Y��t�\��yRb�1��H�a�N��y�Sj���y2�\ 0�q5��d{�����	�8�1O�t��'i,-@��vt$�C �<?����\�$�8.\��aK@�3c���S�; x��^��$}J|�'N�dp0ۖ!���a��<rZI���HOډKtM}0�!�@X�Z� R!X�(���)�' ��9z�ƛW�Ti�	�i���z�r,:d�ЇW�0pjS7y�
����M#𧒟*�<#���,W��+4�TC�'�Q�$j��'v0�!��ҖmS����ʳ>34����D�O�#}2񏗙0�=�ē��H�1/����D#��?#<9E�Ѱe6��kL(|����Bk���'��Q� G �
�:e`D�`(Ru�dO��xr�6)뀵3$�M�t\�կ�%�0=�شj��'�P�N1`RHXE�ٰ �.W<D�4aѩQ$Bht�U��.?X��� 2LO(�(C���~�8�8Q&}��_�<Q��	!+v}{K�Is�M("�X̓�hO1�d��!���>y�3�\�⩺�"O<�A�i�f�Ң�l�0U� "O1B�m��;e$TZ �5_��T�"Ol����	�����_'q�q�"Ohx�À_�)Sɠ U�Bn"\)C"O4�;�]��0����>?���3 "O6�� &ʹ���3Ɲ�5NĈ"Olɒ5 �
���B�%�r4��JP"O��26�3\�b�.C�B$,���"O��pDO��	��Ś4��;n��Ɂ"OD�	AfO�h
�`�
���I�"O4�xA�ʔk�͚`ϗS�\��"O���J>Q������R*F��IS"O
��E�A�ay��Q�ϣd'�|d"O�ur�B���(�
5�@�1"Oܝ��n�ex�@+�bP5c<TA��"O^���ܼf�¤��A�" &�"O�\g�'D=ZQ��O�V�dH �[����ɸG�1R���< Y���g��}|>C䉳	d���
"w�
��7��C�	�<�r1 �O�_��y1�e�B�#<я��?�I��¹G��	�+�&_֕x0%3D�p���d��іǖ�B��L�X��I5�hO�>�ï�e}�U�bJ�i��()�@;�O��y�m}�]���5"GRX�cIP�y��* o���$j�m�Si ���<!���� (�r��L���sd!���^��d�e�۵V v}ӵe�ab!�D�9w^�4 �+7|!�FK��#1!򄀝#� �.��N����J
+��Ic��x�c(�)(<Txa	G.s�	P
3D�䩡�J�R4�ّ%_'K�b��@�1D�@�l��.H�C: �P`�C�9D��05ir
��� ��[���#D�k���xP*�� �M�eR�h��"D��a>{ڌ
�C
`�D�BD`!D��X�ɝ�u��$-�=�8��3D��*�*2���a�K�e��ٱi1D�03�)\02���o�%� 4S �.D�`Q�d�,���Kp��������!D�� f9���]�x�>x�"^!"MZ�Y""O�u@¯@�U	�j�lW?$��b�"OȍD��]�v����X7p�k�"O ����e���z8���"OԴu4w�z�A$A�Dl�0"v"O�������| 3F;@2=�#"O���i��_��a+q�5C�*t!��I����N4�yq��X4��Q��2y!���{�R���2^0c����!�7m�޼3f�	�:i�I�c!�$�!HW�D hH \��́g�̅L�!�DC�?/�����'.x��h�>�!�_�^��Ib�+���b��҃zz!��ՁAv�TAƆ;v��ӵ�6>�!�	��a7m"j~e��[�fT!�޲N�|QZuPF4`� ���K�!�Z��A�S  
T<H\���	u�!�Ų%�F���K�O<�e�`��8�!���L�� e�!-7Tq(v,�g�!򤍥lj�CK���08���z�!��]".צ��KZt����JY�!�Oj-�L2��3	/(�����A!�� r!,��w߾V�J'�< !�ē7�H�!T"}�"(ZE	%�!�dq+R��LS�LƐ$��Es!�ė�2Ӧ��C�����0mF�?e!�$�)�zx2�&�PQ��A�>{]!�$ߗ�T�r��\t�=c6ʑ�P*!��T9��� ߉~~�hr��2�!�d�S���(��gb�a��	^k!򄂆#��H ��V��88�E(@h!�d�.�X�� ���{¦M�eL!�D�/]�
q����9@�� G�L�n�!��^��\A�K��W�N1C�;�!��Ƃv���Ad��B�]Hu�Ѝx!��MY��6��+T9��ܐs^!���}>J�i�'n��u1��45@!�DS�|�R<1�ʆ�z��m�Q(!��4�r�ɵ�'j�4����.A!�_�8���YTD)J���a�;E'!��%�������i[�23���?�1O�J�kZ+8�V�"��XF&��F�'K����27�H;�̆�F!�$N�P�dD�d�D
��h)�D�!�d1+� Dk0*�|B�had�)�!�Dז��ʷ�X�0=�5SQ���|!�DʡTH�-�L[�n�lYы^�N`!�$1\�,l�`K;G� 1#��j�!�D^.(o�����V�#��}�&C� N!����~���6G�8��d����!���=�lJ&J��?u�h�d�K�;�!�$T�!D.]{�K�x(�9RM��!�Ï��Q��e�;gǲ��c� �!��+ai捻��ȞT�&]�ç�	
�!��(��m��G�6B� `�݅4�!���;,�F8��+����d�Y�!� �"x�u)��D�4�#��Ĺ�!�y�JI��&N+}���D�߇�!�ųjz (�,�u�٢��c!�N�\hD�B��.b�l�5�W� k!�dP	s;b��҉D�u���m߁SG!�$ټ7���Au��>���+� '!�D�0sdhz�D�B�rIy��Y#�!��ޑ4����V�Ð1��;�o�)|M!�ĕ1%k[�2T�l��V�ݠl�!�� �se��0�B� pJ�^����"OVH��)�"�X�c��_ �8}��"O�����b�f �g�0�"O�Y�'��0�s��1A��9��"O:,pEk�>b��X�4�U�.��"O���-��C��s�a�`��9�"O<m��h6.?����W�H* �%"OP����6R�$[bݦ
nʥ�r"Oh\��$��2 �nH�%G�� "O��Q1�K,h����clO�=D���"OZ� �` fI^��ЎR1orH,2r"O�@���'x�=���J�~z��ô"O�x��8>&�Y�j�Lo��"OV�X�`
����9�}!"OJ�1f�S�z�N|��
��K@iX�"O��@��Ѷ�׉S/KIX�yV"O�%��kHg�2h�h�XPҶ"O�p�䅧-�qI��H�Y�<5cu"OF��Q+O$z��`��{��P'"O�Pp�OC1���q+�,@�"O�U��BQ�JY�-XU�Ȋy��"Oj�"¼Ee ���I8\�H1 "OH�	V*
n�P����?gDT`�A"O@	�傅
�lIhp;QH�
""O����.�;�r�c���D(��"O$��	J�y��!�'e�	y$�EQ"O�	�*E�v���z����9��U"OJ�w�\�Va,�P�#�^f�5�"OxP����m���� /n��d"O���Ւ.	�C�`�0_�I�"O&��u�SS�����@�D�1�%"OJM�aR�p�\m��uaR%I5�%D�@��NԮI8�,I�N� �%D��� N<)9��9�VpI�d�<)� ʔ2@��S	ӓS��x���u�,;��N�a��e��ɝU�)�$jR�~�y��p�b]�U,ĤK3|a�Ovŉ[�#��x.�&C4
��,/Q�,٢��+g��b(�g�FjT���	d-�$B'p�U�ȓC5���$���G���;5O��!�\8t�	,K��*$�J�Q��)���F�_&8"~dr�/ܧA�,�a=D��;`
��4�1/)� ���⤟�`e�@��`y)t��]X�(�#X
�ā��+�`3�9�O�+� +a��;
5Ӱ�2R���3�.h��Џ^�tC�	aB��ᔬ�?6��dZ`"�T�.�<Y�	�gN���4L�>��O�j����шw��{���u�ԍ�'�"!ခ��o����d>d]1i,�QX}^��S��?�"�<���nΞV�*q��.�A�<A���3׮���F���EȡN}?�V�6}ش�%��<�®�"Bl�K���>]��C"OVX�@�'.R�H4�K$.��6G�*;�DͺG
�_�B�	�u���#kU���ԗ ��=Ib�ĝ��pȌ�iҗc�B�p�kf��A�#���B'!�dû'�l��f��J�Ti��i�r�Q��k��	l�>�X�M�)���h�d�y��h*�<�V⑒p����$V t��@�d]�K���13��Fq��I�Q�d�-���t&�$#����n�^���y$�D(`颅дb�CC�I�H�6xrŭ�UΥ��M��B^���.C'W�^Q@U�[�:��q�;�>lZ�m�D�I�?qbխB���M� R�"ljP�#��+�ax/��`qC�i ���ï�l�aE$�t��eJ����X&N��4B�TB��8�j�榵�'q���v��qj��֓4�$���$�U2��M �	�f\�h'	��7�@��d�-O ��E	t���P#�ȅ[N�n��m떝�$͜�(�	�@˥O���ܧj�Š����0=�"��;��R!�H�
ߠ8���V4-��I��M�~������.�hu��ʘ�	9�i]�m]Ma5k�R�$���ȏd���IN;,�THo$�OB��B!	=h��(�"?ڼ�����#dҌ��V�� &D�!�M
�OR-Bvm�<h��8��\���D�2i��q{�� �Q��-d�E�F�C�bMd:�ɟ��=��)ڐ/�=��*{^h�)�I��\ڲi���K�`CkܼQ�(�u-;Tl=��Z���$		�nӬ��"�)�	c,��"4mD�2�	󄪋�g��˓����L�(-o��;�d��>�U3�M��i�2��bfX�pI�ם�36�b*
�)v䄈����-�牬$������	*�x���9;�����)�n�@+�e���o��B��e���,�p]Ҡ�v~��)�O�b�8��g����ӬW�Z+���P��9u���`�`�U�x��DU.W�N@�ƇI�J&��7J�rĘX�����mp�̂❱{� q0g�	�9�ם������ś�%*&�C�.�B}�%��C�9��+��D�;���6`���'(�&1�%M5Y8xI��->�>�����'P�h�u�{��i>��ڭ����N<QQ�U�ʥu$��!�T9�b�ry���������H�T?�B�`ވh���5/#����%Տ>��r�a؞���>TJ͈���/���I�pɢ�)����>���#@�&d�$�O���'���H��Q&?��g@���c��^�aV`���"G0P�5�u��F�T`��X��<�U��m.�$��5]���'4bV���
�As�'	���[w]<��/�/��O�Z��@JO�>Q��	͸F��-(A�$A�p��c?����I^V��1aӢ�,J�\9��I+,��0�i����O�qr�"8uNduQ��N����W�0��ME2S.�#��>E��J<6J�*�&�/V��g/̾��D�54Y@��N=z`ayR��#�^#��ܦ|B��*۱Tp:�'�(�T�f���~B�Z�Up4��+��x(���<
߶#p��$N����I>Q��0DUGD�Ii���I�h��O@iYd�ĉ(,������<d�>āH̥E&�Jr~Jџ`�p�"4�%�@���Ї 鲉�"]_�X�2�	�y��Pê��v�5��
��<��$[�aB�h�?��)�'

�1[ %�8<Z$j�X�Ct�!��xT�Y1r�Y�����'�[ rċO>	�^Y%z��|�<y֌��Iܲ	��Y���u�v��{(<a�U�Q��i*��T�
Sry�L�,lF%�?���e�'-hF�9���,8�P�b!D�<Q��:P4|��K��R�$��!D�H���+άdO#f�v�1��-D��s��QB��h��]�ipH�5f(D� �u/�)N� I�B'e!Ftеd'D�̳�b��$�"1Q	[�X�*����0D����͑R�T��UiR�X�RL���/D��Bg�Q�
S�\*�e���:̚'�+D��{O��s�dda���39uؔц*<D�d(砏�i�Դco��;h�zV:D��Y�"L�|��L!FAX }i6��t"D�$A$@�6�D��$�8���dI%D���� �:�����Sߌ ���$D�옔�\�%o�0[�K�|��@�@A!D��ңaP�f� ��UH5[�xs>D�P����*pjx��/�l�+7?D��ҲlĽ&�H5��}�\ɸT�.D����n�,��4��EĦL����#,D��(�,^1`�h�AMI���"9D����b!���"@I��ِ�4D�4�U�&~���S��-����&D�(k��
8s-Xe�Ic�q�5�&D�h�Å7`��`E@75�Fu*1#vӺ�I�&8��>�b��J*���낹9jj$���B���U��46�A��O�|9t�P�A|�L�3LM�o] �)s"O�e��E�(�TB��f9����x�(�#�z)%��6MZ�D�Dgjam�O&��zI�$�q��'?�s��#V� Q�௛�/��@٥��e͔=z�*�O�!���H߸��C|�"^$(U.ػ��Ć>N�VΊzy��P� <�r!���c㠤���K�7��	�DJ�Vg)�Q��, 9㶼P��4O 0S�-�f��Y7G�!��"SN�Y7 G�9���S靲k�!�D�/8���Y�#/���ό-����GZ(�k^<t)�e�5=�Q>{��*^�x�K"�T�q���k 8D����0��pP�L�?�ukW�<U5��K��H�D��̢�#��r�ʓ��b�����N�~X^@�an�o)|���=�O����.� ��
� ��Vظ�f�A���vJ̯
�z�*ď?l�h��'H�T�c� b���Ň6[H����dNz�2T�U�E%�@q��^� ��\�U�~�f����	�A�r��(D����\
O0��s� ��S������<YO]+zZ�Z�N�-��	�Bӌ���{�n��~}D��ë�(�ɉ�"O*����T����0��˛`�j�ax�Z=)�ʛ�H��!&��s��OI1O��*/K�y�X��m�;h���;A�'e��s�X'Zi�A�`�e�hT�4K�8\o�Q�%��b��,F�N�az�a�0?�j�;3K�2I�D�����O�гE/-a4\��E��>�d  �O _����I&{F<�0�P�F4�B�I�[���nV�"X�#	L� _~�iF�7&S�Y��8�U z�ģ|B���/Wh}����Kx9;@C	C�<it�i��PJg���1V:0�Bl��C;���vl
$ut*�C��-�8��|�<��&Z)�T�q&�6~<1k��E(<a#-T�/&�:�[�=��A9���ur�r��¨@�u�S����=�F�q��]
G�K,(����K|8� �GI<,8��0��-�D�mZ�'߆9�$"^*vV4�8�ϑ=��B�	�c{�T0�i�pUv����j��O���U!=���F,��h�@�Y�����ĚS�2@O�hJ�"O24*�b��R���WhK�q"�(��G�##/�"M��AF�/�g~��P-bѐ��X�F��}�Pꚭ�y�)�8A>�����">
�{3�S��M+ �'0����K:w�̴��.A�	����dV4z�!�D����m�.��"�cB��!򤒋z�m+�j��D�����NJ!�D/j�PIr�ةc������p6!�4(np�q�B20U�5�w�D!��2�8�a�͎eM��!��z�!�D�8;r����(��a`B��!���-	������3�����B?b!�d˓I�`pJ�M�'�4ȒLܹ`f!�D�>=�͡���ktp������cu!�"��p����g �Pf �]�!�d��c��E����*�"��p�i�!�$�`y^��$
�s��#t�HZ�!��ȫg��ce_ݖpU�Ʈm!��hѲB#�,R�0x�3+�!�Ğ%���fHժT� ��BA�m�!��
?+h� 㪔�R6�6!H�!�$ϼA��w璅�lE0�a_�!�$Q�ir����R
H���#၅��!���|瞤( �DX7��G�+�!�¤>� ЗEW7_5.!
V�ۗT�!�$�2z��;��E���
HH�c�!�D!n&5R�'�i�g��!���r��
��G�n��y�À�!���c::���^�'�t�@��	|�!�d�/S�f����l�"�����(�!�Dz��XJ�d�8j��U��e��a�!��"'-�A��K���0V�U�*_!��)�����ŉ
.�$�3���!��K�dSB4�ӏ�w�&���b֧9!���V\�P+�)ŋRt�V��_%!�*x��5S�g�~K*%Rנh!�D��^>���:�$�� �$�!�ʔ��r��	:�B���� �!��I�e� ԑ��G�Xu�k�+�!�D���z}Zӫ��H�XA!��ҞnJ!�DO�'�5�DF�O���`@(0u\!�"[�2`�7^���a凁5&!��A�I}@�Z��*[�`<s`Ǉt&!�D�� ��p�/��]��ijd��4<�!�US�,�1�����遵�N�Mr!�� 3���&�q$�(�nCT
!�� ��1��Ύw�b��QFD5s�B���"O>Q���o�yqW�Ŀ�>l"O((�����˗OŜB��A��"OFe˒��*v�<�8,�.���g"Ot[�6Tj��e&Q�xɊP�0"O`|B���><��V5-D`��"O�p��A�2AA2����A6a��ۢ"O�� �`� O@�
D��;:�b��"Ot��,@�3kP���jZ��B"O��`��F��L  ��)~�;4"O�EꂉJ�M��&LA�!��#�"O�L�%�_wנ%����F��<"�"O��+�X!M���K��P�d���"ON]�e��4u2�q�G�ٰd��xY�"O&��׊L*C>�mA�(w��1R�"O���(݄}0�Ͳ�%M�/�v��"O0�{��T
T�$hU�.$�V�a�"O"�j�+I�8r�8Y����J�z�1�"O���e� 15����
�r"O���+\�\�(��Q2I��yz"O�8K�D�2f� q��J�D��"O���o�<���(��سB��""O��������΋�S�=K4"O^��7�}�]�E-Պ$*\�	q"O�!�3N��"4��C�J�!b�$b"O,X��#Iy��È�$mW�%CC"Od�B��Z��麴$A%J$ �c�"O��̔�M���Q�Mח/L0�P#"ODؙq&�D��D3��HM��!"Oġ��i��QG �ӅT9 *Y:2"OK������7k�X�`'��yB��8�r����D��`� ���yB��+�����ٔ
j���g��-�yRo��26~��FH�	�� b����yb�-V*8؉2+\������/�y�*��W������֭L聑 ��	�y���Evi� ��*
B�@ ���y�jɨ&�*h�C����+PGY1���H`T�� LOZI�l�\|	�c�P�9�|�;��'rT�h'J*#��� �f�f��T�h�:=v�+�`�Mh<9 �=�T�$���*�"_]�'.��	Pc׊:�@�4�	X�j��R�<>�j�z� ̕$~!�DA��HݲŢ���t�Wa��f���A�U/^&�u��+�wy���'�����¡[�F1�EHQ"�-r�'��c�ɇY�a��ǅ|�V�'<N�:@�	(82:�+��'�V�I�gdQ̤Z%C	vxHM[�$E��A����a\��(�//D��t�Y153�Q9�`��x"�[6C�,��4v��l���aZQ�$8��j��iz�Z�9 :�F!O$`����gI^979��ȓn�|���o\<+�$XT�O�3�<�L�l���s�˃GW�)����L��i]�pCD�����:D�\#G�)�n�S�Q6o�-(a���HQ$�\e��e�5(IX��a��J�R�J��H,{�괠UD �On�I�2��0{���98�\qp�����i���<��x�"�nf��s��ۮ�!A�˒��hO4��R�g�^"|��*ۃM欤	p��*ֶ���kb�<�G�	3։)��P ��\D�'e�#�X�O�"y�AQ�%TH��2������(O�X1�KK�=�nǼ2B�Xդ&Nn�8�HT�<!��WHBi�L>%>� 1��)���'/��d�������a�^� �C�	(�E�h��1��YccFE�~ވs4`��l�r��45aZh�G��8F
Q�f��N���?M�hZ��L���
:f\�2���  axrj��]Pr�!�i&A� ۤ�~�i�jp0�" ��#R��i��d���������'`���hu:� �Dʹv���r� ;8\|S�f��zy剁A��H��՛ ����\�1J� `�N�X�!@o(��� ��)�*W�-�墧��OPv���O�xa�>��i�
ӓ\� �ˆ1�f����#���᥉�x(+-_����\�V��1۟N������~�؂D�F��8A��2pzP� �h���֒E��!���w���c�V(� ���a��w�l� �nκ=�v�����*i\�!��V�u��˫OTAې��R��=	)��e� Y�v��@&�L����$>M��z�����HSMӼfE�]b���"G� �s����F6PI�-]85�

 �tҴ=ADS��QV�"U
��)�	�=�	@)۔M�l� U� �8&˓mV8)�����X��υk
H�E0&N=I���F]���lB:�[�F����j�N�6�^��>7�t�[)t�&���(������WI(�0+��у9�؄n�>V��c	e�0瓘T \U��O*�<S�@��;�ޘb�J�e�$���J1�"2o��4d���Č3�tU0c!@/��	�C�^�(�y�GȆ7L�RL02 ��U�y������A��L���M?)�~�C�����Q@���5����!����'tM:��Y���M�@
R�0<]P�D�"UA��S0Nݕ��i>�r��t�d M<��LX*����xȜ��&FyB#�9g��p�F[�T?)0S.F�1��!4�:4q�@C�d�X�F�B�����D,)�	�j�"L��	�I��1�Ѵ^6$��#����!�L�@ЇA�4j	$�'?A�ǁ����dn�'lJ���cE���q�A5y��\[R�\��eg�!���P�ҐuR[�, E(Q*b�	40�'A�D�\w�P�������O+�]����d 	�鑍Q�Z)R��ңzL�q 䈧�ħg�f��f��>��Hc�&@�E{v/V�o����c�52��)��L�WbҢX���#�XH�0B�ʵ<��6ea8��H9}��)�*o � '�R׋��S�`�ѫOʁ��C�1��B�'��ȪP� �dSv��M����I.}�L�2�x�kg���'�ܥ����az�;1���Ӟ�"u��0�����'���з��.�QY�%�$~3r��baԻI�@M����U�	T4���L+�'i���`!�B��&�E��F҇�LF~ �X�S ZS����?5�P\q5�ժ�^C�I��x��R� ����D x�˓Kc���!�ӧ(�p%P�ɑ/e�v�T��-@H�p"O0��rJڃp4��2�&�$�f&#���&
�.�0F��dA��`D!Tk��p���
x��q��;U����Sg�oԄU@�,��x2%�	h���jS�H$[K�%�b���y���/"��eːQ+�
3%Ɍ�y2 �/t�̻�AQJ��8@4M
)�y� 3�,�l��Fa�0XNX	�'�<!k�C��!�5�I  ��]��'2��ǀK�V��{&��7$���	�'(8y��E3 ��a�`[	
�u
�'���+3V�����&0tb�y �']:Đ!��=~��I@��k�� 
�'��z�������b 
pl��':�@*LZ@is���
�n��'���[�n�,LV|\QdE�vȸ��'�:@��bԭy���s�ƤXY( �'z����*�<d�&��C�Q+dP<P
�'�~X#�׌U�:��FF� e���	�'E0�sN�h���S�L�a�'dv�Itn�v��P����2�%
�'�H�xA��\�	�q%Bq�	�'�T=�s�]�e�<�a�(1��-�'�4�e��R>��M�-�|Z�'S�F��b��h�F&_A�� �'iF]r��{�"��UM^�'��<��'u�8Xs ��cP�͹�hޞ��)��'���{�� =W�L���&E% fV[�'����ƿ?6� �M��.̉�'g��[� �)}���8�:4P���'�r��\,��V��~xj���4�y�&��;p@i�C&.G��}�Q��y��M�s�j��<�����޾�y�/��jlxZ�T�,�`o�y��?f�]��!q�
	��V��y���4N`��B�.Z�rB,��܄�y
� PtH��ӈEZ:��l t�J*O��B�ټ.����Y������'�]R�h�I��	�������'��(��E[D�n���cV��T��'C��q��59bJh93��VIn���'rep��(��A%KI����Qb\���>��:=�6�k���P��ȩT�[I�<��i�5B�Vk4g
��"���/�E�kv�c#a'���v���8.<���H�)S�	8E"O 8� �s��j'�;(M����@�gb}p �>	@?�gy�H�I�FI���)~Z��k��y��ńW�2ų�,�X����M;c�X\H�n�>ƾ���uf`ɡC�)�����ƴ�뉻g<	�DcD:3/��(��Hw捋"�tLi#"4"!򄊆5���8�d۟kˎEѵ����qO����C�	K^:���iT�
��s�XG�vY���E�w�!�$Ѽll��b� 8A����*���F��"�U�T�|�'sn��T%�h'T(2UA�b�옣�'"�  �N}�#�Vd�,��aZXJ�!Ԇ�0>iw���_1���ɑ1mT�Y�G\��xb4��sQ>�7O�rg��R��a���p0n��"O�e�u* ����a��@����C���=����%6�bF
�+��ɻ�n�K3J��@�ȓJ|x0�D�͠��ț��t�B)��ǇHEqO�}���&�9�F�$S$��5��7��ȓ4�ެTI����cf"Q��}��&�L��տ^�9�BAO�mB&�ȓo�H8J��@?v2�r@FCx�PԇȓsHȍ	��0%��A��,�v�B)��t̠�E���~���M_0Xl�����8Ӏ�/-Z>�*�bW�⨇��0-8&n��V�0,�l�R�Q�ȓ.UB�(Y�O(��A)�Y�ȓE��y ���%H�\�*T��p��ȓ;�1���@>@v�B���Z<�ȓ�� ���S�|�b���69������F�.j��0*��(T:���P�0��"6���9���u�hM��i���t)�����Ղժ3!�4���2�*��
�H�yBB@� /�|��;K�ɪ���}�\�@!`����0~����L�A�l[�m�%s|��ȓlWb�S�A\�t�kFNݕ	����s��} �f6�[%/�	���ȓ�n�x KڢE�As7��uL���!�H���-z<~p4�ZѤd�ȓF��t��lǇ����<y:p)��2�l��U$Y�yzT���{8�H��1}(��y�f�����VY�Q�<�	 �QV�mh#gS�z�n,�w�{̓l�H��Ө�t�LH�s.ҳ �D��ȓa{�:��ǟC�H��(�65&���/o��в�ӂ�A�3E5�6ń�NaTt�T�udX9"5��H�R�<�v��<Oڮ��`��(�8���C�<�,[�
P�l��"º.�v����x�<��$�cܪ\����6%}F����L�=mK�"<�'��	�T2R�2q��7kפ��^h�@T.�>����5k���I"rq����B�ɟ��$�L��<)LԬGM���W��2Ph@�d㓌B��I��)�&_�S�O+�jS�K;wn]����;�\D*�O�زD�)§r/�����56H���pc��I�dH�P��<E���\M��;�/dw�Y�1�ʛ{*M��ө_k�l����d̂1ؕLE�b&֣<!vB=�b� 6�RU^�2�j'��Ѡ�$��(O�Op�<���Q��h�d��~3�xH>�y��3� ZE!��*o�i�FT�p4p" ��>I�O�Y�S�dl�(6�6mC�aXA)��X@@M��"��`y�hTaA&
M�ĂM���6��L�����|j7) m�N<�� c&Z0��LR}b���o�;��4g됢�@B�		��) ���O�� �͔�%������1���t`��<�	�'(�QQ�..'n,�e@LW�d��@�r��b�f���de
v>M��隍�U���7ETtL��䏱WҼp�v���,��C�$~���'�H��t("c43�2�����	Z��rZ���0.�#�qOQ>řB��06J����8� ����OL�s���ڸ���"0�.��Z
�xIF)�\J�(&B�?ᰝ�=��'E�ɳ'�0E����iCt�Y4��4!���?�'�NA�`G(B~<e�V��a�&�	�'�<\�@��'|̠$H�ٗ`Q x	�'�N\i�+�4�&�����R�� ��'��D�߻�<����{�=Z�'�X�14��.4�<YR�N0+r�A��'�h���L�.I��A���D�'�R���'k8р�G�/�8)����A[�'m��G*��R@�!��J-{�'�!�b�כg�h���ƋS�H�	�'�[ H��5�9y��	4&�|z	�'�P����#�\����
&�֥K	�'r>�J��N�:���A ���h�	�';j�@!,D&���:AoG�Z����'N���pi��4���O��U���'��h���Mf4�⤭�8bT�S�'�~䉳��1n.n��$�`�.-j�'�x�c?$��@�ӈ�,U�t(c�'t���8n�Na�#�P�EO���
�'%(�;�H8�����
b���
�'����ɱ#�cw�݌X:Q8
�'�ܵÑ`�#g�4yuC��s�q�
�'�P���<X��9�D
��<�	�'�����N�"�b���@ ���(�'S�X§0R�9(�k	 k�i��'[((�2�kn������W,����'邼�7A��@c𕰥�Q�DXָR�'�Ab�M4�L�z�8g28�
�'V��� O5' h����X,4�@�2�'�xU����5#2HJ�㌈Zj��'��i�F�Vږ�JW"2�8%P�'�@��ǃ9W��ɶ��h��|�
�'z�M�dH@�}=�x�%ُY����	�'������=����e�T��D 	�'hyk�NY�hlT�!�D�IJ���'��	��J�)� 8˲	�{�$�'�>0vL� Q�H�Bu�
�zf:p �'"�0��\���h�$pJ�Y�'������T1��;���7V�i��'����+�n����͌��y��'v$���T�����~`�E
�'9>L�P�.z�E�����BDٺ�yB��|μA�嬜�� ��,F�yb�%-2���aE֣N�;�H��yD�n4~����?9:ԫ���y�-��{��4�
m��-��y�㐡16ʁ�æ0�U�����yr�-@����z����(F��yRř�B{�r#��&L\d�V�3�yB�ޝ)A���u��-�QxsI*�y�B���ҹ� I�\�<%c�!D��y�j�8@���a���\��A`dĽ�y��T�	t��{�ЄUy���Ǥ8�y�%,O�����I��L�7��'�y�N�8�B�"U���8H� ��V"�y
� xh�g�Xi����Pc���"O
�d	5E[ e�ý!O2P��"Olٰ��Y}ŋ��L�,���"O��spI�c�(��fD��
�(�8B"O�`�����N3NECp�ō1�
,��"O�i�uO��]zJC'��"]d=�"O8�8�œ���I��C b�ʝ�!"O(5��+> I�b[�
�*�p�"O����H�-s�mT�Hs���"OD���ʟ"A@ٔ��i,�z"O�A���0���'2\�Dإ"O�M�P(S���C�W�?�>��"O��� ��c��y$�<@v� [�"OqW�5^͢����QZj!��"OJ�ȳb�?�x�BB0{E�"O
�I%���.����5X�8�"O���C.H��Z��1 ޚw��1��"O$�(%���C���)��d���
3"O�,�s& +����9U�ܖ(�y҅ҏk%�D�dNI�SSJ��0�ȱ�y"l�2	mڄ�V_d �� �y��I+��b���h@�wD��y��^	@p��ғ� ���7�y(�@�R�"Ӣ!vp@��fJ��y�$ђ'�4�c �WŤXzk�y"L�G0���)�:��i�����y�NԤ7�{�i��d����0�՝�yB��:zX�xA��Zהa�P�$�yr�܆��)q��JY{�I��m
��y�D!2�̤��N=z`C֯K��yr�Z��y鐉9[��kUEM$�ybI�[�����;4*.�E��0�y�#�hy��s׀U���`� -�y2B�83���P"k�J��$z��A��y��'	�lې���@�l�����y�lх&��S�̅�2�ڤa��y��(X��[Y�����O�m��s׆(��̘(`��q'�SX���ȓ8�԰���f���n4�8p�ȓA�
H�enk[�(�eoO�[�乆��d��P �=Rݸ�g)V  en���x�U�"��	#�q�*=b� �ȓ�D�`�(ٌk��X1NB;d�ņ�Wb��E/��?�n!B�*I5�$!��H�r�%U!�:��α�Pu�ȓ1�H괉S�v&�,��	*-JY�ȓ1-X5IF�ې�pJl��k V�<q �Cu�r�:f��+O����S�<��,I#�r'��*SP\��PP�<QVLS�B�D����Nؠ����r�<q��ߜ*&��R��
�'z\y�/g�<!��۵�4 2��n4�Bq��h�<�RUX'ܽ30i�VO��ҡ{�<����*DZ��3�&�6���C'�\�<IQ�ܕn1* hfL�cَ����r�<��ܕjXTQU�ۃx&t�jŀ^Y�<���j���*Z�(�2h^�<���-�:�:��Q=jt�RR�[�<i�FՃ%�X�tn�?YD��b�AM�<�À�9wc�j"�B�.,N�:���E�<i MP�'��t�ufK+GX쐂,�A�<�tEҡ �4$��l�}l\���G�<V�߻��]�CBN�V�%ip��@�<9D#�9M'�q��'}`��7 �z�<� H C%�W3?rF���Q�l|#f"Ot��H�4z�
�ɐ��42pf���"O>4�%�ȅk��4Qt	D*��D�"O����^��!*� �3L�%+s"O\��*��)��Q*qIQ<q"O0�Ѐ�g`�Z���YKn��S"Oz���
.cв��@�C$/�=P�"O�qBuI�<&�N�)���o��\�p"O
�F � �Db׉�&�����"Oʜ�QC�#P���V.K5b�l@��"Oĵ��EC�E���΅,1p&�"O�e�v��.s
��rPǀ,"Tj�Q5"O5�C^� ��q34��2io�չ�"O��D �/��i'���M{���@*Oƭ�-�*�&a
W�!<��k�'�8e0�(ձB� ��f��	���'�yae�[�1X��T�X�4��')"%IT�Y��;SK�C�'���q�B�0I<�bsF	1}��+�'�>�Ɇ�A'/���P �кv�R��'�&��bMe:iÚhxq�	�'o�9Ҳ+L;$)6����޷b&�%�	�'���Ä�L�:+�x���ĕ`���"�'�t���c��k���UZ�n8��'�8����B�uI�|	 iU)&�\���'B�Dcg�4%z3R��qT|��'*]�Ao��8�����h�3K��h��'�̉����YC���B��DLRE �'��`h1��7��x"A�̊C&�s�'�� y�
[+C&�������U��'��I�AeɭH���J���
�T��'����������烽�p��yz���C7:R��@��ɀ����T|���t�a#B^�PM¦�}�<I"%[%G�:5jԋ��}���jM�<��$�	>^��8�D�K�b��3��K�<��+E��� t��&pJiyB��~�<9�Ꮢ=�� ���# �|���͟N�<Q$"IH�	�J�1�D�#��@�<��(\�'��Q�"О9Ĭ�r`Fs�<9�J`�����d�ht@'Fs�<aU$P �v��s/�H� �ekf�<�K��1S��s�Ǝq��Y��Mj�<����s���r��%^>𰙇��h�<���:�&�0�	 w��q	&E�d�<�Í�fq�]�� �V�Z,�3�G�<ar���&����������!��7�yRd��d��%��5`��y�G��p�`P9V�S�<�����y2��L
)�fJF�FZ�L��Q��y�{�\�T�R�@(���%�Y��y�k�,P���bI�g	2d�-��y�$Xk]$� �܅XA���U�J��y�S��mB�+L�M:屵���y"��u���a�E�	G�����Ґ�y��ۦ
;�P��N� #K��y�Ʉ*<�f�"A/\)CV�]��y�թh]%�"|�V��ugP �yr�t���'��u��PiԷ�y�n�4x���i�
~S�ukd)@>�yr�ԗe.��oޥs��٘���yBM̭����N��8t�#6	O��y2��� C��2.t$������yr�W� ��"�dA%����@��y
� ��fi�N�N��r�<d�a�B"O��r���'���E��VN "O��#�X�Y�`�!E�?YM`"�"OR�z��]�2
T{U#92,ؐ�"O|0�aJ"\�^ )���"w��"O��; �(@�Ax�A�"��tr�"O���ȅ�"R2nYJ"O�%�@Fޔ[�x�����l�,t��"OXt�"Ƃ�F��Cw��G��w"O&��PK� A^0I�A�)^x��"O�=9�-�	���v��{	F�S�"O�T�0f��D�d��O�"^&<r�"O<��/@7�P��5�;�݃"O��G]W�����.9M��M"�"Ol���   ��     K  �    �*  �5  _A  OM  �X  2d  Bo  
{  �  ��  �  �  ��  0�  F�  ��  ��  �  [�  ��  �  ��  
�  ��    x � [ �   U& q- >4 �: YC �L XS X[ �c 	k Uq �w �} d~  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR��D�J���ӳ] �K��F/]$	����kϊB��.p2:d�a�,��������=QÓh�D}*���\�<�{ĥ��1	bq�� U&�2�A˼m2��v��$&����
rdk�A�)!��T��ΣT�8��re�q���W4O ��Z���+�'�δ+Rh��Zc�,��D ��2�S��f��zA�QW1�ɢ�݈�yB�S��n�A��M)3|��
I�v6�=E��ULD�S��"�l�B�C�tgZH�ȓp�(8�6̎��.��7�(1�І�_�%�l�-�w�K����ȓ{��4���`��n+h,�ȓd�Y9`X�^�zQ0QN�GU�ȓP~�����+���
u����5)�ذ���
T
���A�N+���F���c�H�h�>�Io:[�M�ȓ���G���,�+�T�g�0��ȓvU�M	���}0�P;�/a�f��ȓi����P�C*r���� T/jt��ȓ7��0�R�#!�X\�4�c*)�ȓ#���H��&l��:�"?r�����na��جT�0��j3R��܇�Z�ڜ�B ��w7��1��X2���ȓY���K�K<�fX�&�VL	�ȓe˜,�ӨN�Tu2tX��ĭ[NrP�ȓ�x�1m�(H��dϰ:�����4x�M*O�����,�\��>�8� 'ְ%?�8�3��t�$(�ȓy_��Q`&��fut�@d@Ϊ>�-��qXXգ�
�?Q�����'����Q�հ <A\ ��j��#o�0��Z����-�;�`��q��-/ y��g�&]6HK�Q �/I�����"D����@�,c�vh��F�<��"�g3D����l�Z3���^2CG0D���Р� 'Ava���ƴ�V�1��/D��A��� &C�5��gļTzJ�7l-D���rF�+%�(:��_�Tl��7D�`)���6 e��@����B����+D���a"ϑ"���b�C[t�$��s�*D�pڳ�& �*��e�لF]y�U�&D�d1�-q���/�rߖ �&D����oH�B����w��JAn`�.(D��:�`
q~��Kq�^>2\��!T�XCe]��H�Z�@5h���2"O�M��4l�d�
׃��8�ndñ"O�1b�b4��-	c�σc�4��"OH�y���ov�y���D�s�jU�"O0<"�*��0@p��-b�
��"O>`��7`��ܱ� ˅8:3"O��S��=ǰ�Y%-��N���"O� &��'��=y�~���L����2@"OT�	���Q'�Q0JI)RXIw"O��KD�5�F��(N;( R"O��#R��39���(ٯi�4A�"Or�PVꜴ-c��e�؞
�����'B�'}B�'��'o�'���'
&p�k��8�5i��3O�AP3�'�R�'U��'�"�'.��'E��'�Ќ
a��R�`A!�D�K�^���')��'�"�'���'�r�'���''�y3���o��@3����3��'��'�b�'�"�'�b�'�b�'Bh�CQ�S��)en���K�'A��'+R�'�B�'�b�'���'ONI�GXt�"�J%Cۓ�8���'o�')��'D��'�B�'���'aV [c�]�DJ�)�����bD�'���'�R�'���'2��'���'��$��D��ߠ��4*Ol!6�'Q"�'�B�'�B�'�R�'���'_�	��e�,y5���U������'���'�"�'*"�'�2�'r�'������ė/*��;�)��c�u���'r�'���'\�'<��'�'�3P�)-X(�q�fA�����'��'�B�'���'n��'��'Ԕ9y�HG�<�����dݷ6�bLH��'��'WR�'2�'���'�2�'�F���+��: 4��e�e�~ ���'���'$"�'[B�'�NvӮ���O��	U�wY����^�!�Ȭ��xyB�'h�)�3?�i^�ik��M-gYV���#M�+g�����"����ڦ��?��<q�zXU�C��W>�B�b�7A�����?yt`E��Mk�O��S��J?�7�7eD�G���^�,ٕ�-��ş(�'��>-�C���
�o؄p�!u��M;�A���O$L7=�28�jS�	Y�lN1fXp��r#�O��D{�ק�O���ºiE�����\#�Q�I>)�PdN x&�$m����E�=�'�? 
�(��e$(���׎��<!(O��O�@mZ�?�"c��9��]�bKB陁*$��`��X���I���I�<�O�`e���̞���Q��٩2&�,��O��K�rf@Q���?Y�b�OTx��ꖂ��#���(:�|�q�a�<Q*O~��s�,�wfP�<\��o Ԁ!R�c��ڴ�b��'��7�&�i>9��ƚ�L>j$���S�����l���I�d��!\�`oi~R5�da�Sk���P#C
5i�E���&n��ꢘ|�U��ʟ��	Пh���|��� =!nJP�VkW� t�ەIAyrA�O.���'��'V��y��;���x�`H�IW��+����_I��DX�v�x�*�$���?��SgT8��	�^u�#C`�H�IS.�����542���7�2	��f'�'!��0�ڵ��$N0KWxAx`JVU6����?I��?���|j,O�n�<vHR��I,
�<��*̫4��+0ρ�C,,��	�MC�2�>�#�iN 7M�Ŧ�+@LAzGX�5N�i@�����+F�l��<!m��u��8g ������z���������"d�4�Y�E�0�%� ��<I���?���?i���?����,߬��dJ �L{k�p�4F[�5���'���f��1�6�t�d٦�$�({%��,OE�����&O�8�3
2�䓈?���|�E+���M��O��]wx�b!N)˦�����=�F� �G�O�t�*O��n�iy�OC�'���(M)�]�2(��J�&q ���"�'�剂�M��e~	�I�$��P���O;d�&�b�̡���.6����Y}
l��m�"���|b�'f�j�q۝��,�$�^R��|ɗ�.ъ`��ML~~�}�y��'h�i�'�wH�z�(�W#E�	�h�Iրt���'��'���tR��ݴ!�H���"e���C�
KI����i��?Y���F�'�'oh��?��o�g�����Aպ'x��""<�?A��i;z��D�iC�c>}��f͆�����j稄�I�|��e ��^@:P�)�M#*O��$�Op���Ol���O˧n��ӐgF�fC�
'K�'���ĵiʂ����'�"�'��O�ҡr��2�{%,J���c��0�� Cv�'P�fi;���(�D}��;OzaׇG ��ٸ7K��I�A�P2Ov 0R���?��Ĺ<��i��i>�I�iH��x�M�QyP!�r��>�*��	��D�I���'G:6-��f�$�O���ƣw��t��)=N� CӉ4h�,+�O�qm�M+��x��
�\�x�h˞]�l�M����іͫA�����I"�u�I̟����'���$Bڭ9\���G���].����'<r�'R�'	�>�]�d�p�����?ZZ\z��U�s���I������*���OL,oO�Ӽ#SG\�B�`���8qx8Y�R�<)���?��i�x���i���=�,1C�O��ףJ@5�����^�1㐅Py��oӲ��|*��?)���?��#���d�[=��P[�-A�it\��*Or o�2Z�E��֟\��_��֟�#�ڋx��R��)'�.�@E�[/���O���j�i>=�	�?"�O��>DaG��mdQ+ԧ\82�����-?�F�E�{e���^���Z�՗'�H��W�V��4�3�K�dY��S��',R�'�B���S��c�46�F����-@"mx1�+k6�����8I�D���8ћ6�d�ty��'���ehӒ	D��.-�`�ǣ�F�[F�Y*)�7�r���ɥw�(ut�O%��H����� �!��a<{�4��DL������7O����O����O��d�O��?�r#�T����憭V/��ٟ��	���ߴ7~��O�67�>��S�*��𢁓b��,9ԏU��2�O�4m��M�'�
�`ٴ�y���n��$Z�BT�r�L�R�^�A�|�7�X&H�)�u�O:��'�r�'�r�'̜u�c��2k�\�sgϝlE�U���'Q�T��ܴZr���?����i �W���z�l��̕Cv��;6�	����O��D,��?I�g Y�VQP�	!$ �q�LТ"EX�{`���4�֦���ĀSA?	O>	`k�	2���̰,�����)�?I��?	���?�|Z+O��o#��|� W#l�j�)\���a�GmN������MӎҪ�>���nm��*3M�~�x��*�m����?q����M��O�LS����zI?I�ê�(.��82� M|�5��k���'�'���'%��'�S��4��2(МE�`�f��'ވY۴M+z���
ش�?9H~ΓM��w44ѵF��]n��w��*n}|����'+Җ|���e��EY�4Or%�F��5d��wm��0,��1O�p:S#�.�~�|�[�@���kFD�QlΉ�!��EӠY/�۟��I��8�IPyB*~ӒaBG�O����O�P���.�(0��'���xrO1�������O��d%������Đ&��#Qꩩ�(_�V��I�(�``����+K~��`�������l�GM^#St�+6bϡe��9�I������IT��yg�W	t�� �	Q84Ś�Ķ[���f�zH�5#�O�������?�;�����üT�x�ʳ���p�r��Nӛ��s�b�oڄFz^�l��<I�:���������'ϫ~"����*'����t�K�����4���D�O����O��W�)�fŊg�r$�B�!&˓Yb�*�P�'�����'�riS���5>��i�dh�
F���h�>���?�H>ͧ�?�����	j��q�pi�:�֘;��A
@�X�'v"�0����R�|2]�H������L�{�RR�܅�@��������I���@y2�~�R�:��O�)c��Ĉ/YB�@�c�&l���O��l���$���O��d�O����,Pg~4;�� ��
œ�v�Y1G�?��3O����B+�*��L���?i���a�5N�6/Bif�!�H����|����x�I퟈�IO���D���8Yk�E*ƍU1b���?��G��f�X���$\ڦ&�� &�Ns����mO
D�&����I�I����i>E���Xʦ%�'.���K�CM\萗���4���O�X�������4� �d�O�$�`�4\�@2*d�2g%�O��d�O,�u������_O������O�rH@��b�Vy�Ř�'���j�Oĥ�'HR�'�ɧ���'���au
51���(��m�e��ϝVȌ}���i�rʓ�.�:�	\�	��`��=]zPY����"��I�L�	���)�S}y�moӮ+D�-z��tCݡ8^�h�2�хp@�	��M��2�>y��#�dls�l�,O
.�h7�Ԗv��(9���?9v	��MK�O� +%�ׂ��O:�ٚ�G�
�b��b�'����'~��˟�Iڟl���(�	l�4jͦ�����*ʹ^�����̑%�r6-&*U�����T��y�ǜ4�$�˧����:�s��&�b�'Qɧ�D�'b�䊥.$�f4O|�C�I��c���m��#�2O6�JJ8�~�|U����Q
�=�ʙ�s�EX���9���������4��Xy�e�&�����O��D�O!�Sd����q�c�SJD��0�����d¦���4J�'m���1 ?:p�� J\+�>�ڟ'J� G	,���������Hh�V����ҷ2 �E��lT�KNMXBИ'tF���O,�d�On�D1�'�?q�(ю��Qc3��"� ���]�?�ÿi�6|�g�'�ңq����1*%>h (��S��U��^�u��.�M�P�il�7MS.9/�7�m�8�	q��z��O1>�3��ѿ�ֱjp�D�)C��}�Ey�O�r�'#�'���̆-�*�I�gW���a��cД@�	��M+����?��?�K~
�	8 j-[Y֨[DRsO&u��P���ڴuB��)�4������X��t($�"X"@�Zv���(�a�R���c�Kt[��D�IQyR΋�\�p v�ͶIߪ���m�s���'�'��O�剨�MCBω��?�m�>l&�P!C�V�+�D� 4�Z��?D�ib�O���'7B�'~��Ob����C�x�@h=1���0%�i��ɡ-�� �ҟ䒟��/YV��1���9#�� ��6��d�O��$�O[l�ܟ<�	}���0Lbfd�>`8h6�ņo\fLB���?Y��C��6�����'�t6�1���X��X�V���1�]� A�F|ܹ%�`�ش��F�Oa��{�i}�D�OƱQ��9�CLׁ<�}�oD�X�,(;��'�t$�<����'��'r2�iW�ٜ�T0�GUc8���'{"R����4w�v�����?�����IU2v=|�Sbn\�����¸d��	���Z���Y�4����)J�����!+�˂��|T���5�JT��h �j�3��i>�0�'l��%� AF�����U�����.]ܟ���ПH���b>��'47-ц:z�b�N�(t���˅�r٪1���x�ߴ��'��듪?��ic}Dr�����^	�� ����?�e�ܗ�M��O��!֣B<��π �Y0�@_9B�&`7�&F����R1O���?���?A���?A����I=F-p[Ч��@���t-��o��n6Y5����ן��	S�Sן������e��#�6����@?)8�U����%�?������|
��?�6I�5�M+�'W�X��$ɒ;����"Ot��j�'K�����Xi?�I>�(Ox�D�O����-HrIn���(�g�O��d�O\���<d�i�x�	��'b"�'k: �`RM�9Q�A��9���'�'��듵?	���$.4��"�al�颥n
�6����?��旮f��-�ڴ$C�I�?#4�O���u��9a!�����]+׎��2@����O����O��;�'�?����jh	Q�ʪP-�YC '�?���i2�QU�')��s�.��]�W_h���+�-�}��=9��	ʟ��	ǟ@�!��٦�uwW�9�ɐ-�h�%`��mrr!a%!�|���Oz��?���?a��?��P|�!�0��P���`�ת��",O�l� �T=�I�P�IE�s�P�rN�8+�!��-�*=�*U�߁���OV��"��ɔ�7�(1t�4h>�vfI�*��]�U�n��0�'H��D��m?)N>.O԰[K��[D��R�PMrY�L�OH���O��D�O�	�<�t�iJd�@��'l,u#b�TB������,@p���'7-(�ɗ����O����O8��X9ci�-p�/�J��� ��/{�7mc�x�	>U}�!xڟ>˓���W���X�,�e�bYx���>��?!��?y��?)���O����/�\GZ�	Wl��b}�=��P�8�ɡ�MK�*N�|��
��f�|�4��\�Rm�k��i%��3]+�'�"�����38�F���4	�4�R+K�kYR��E��+!��H%��c?�H>1(O"���OT���Oܐ��`�:�0F��$k�C�����O�˓<��o�0<r�'d�S>���L7O��YY'�Բ4�H:2�:?)�^�H����|'���CD���$�r*�!�V�bo�=D���Y����Mr.O����"�~r�|�/�$*�`eH���
޸�@/2&�2�'�B�'����T����4qsz�a�#M8����M�Nb�(�`���D��Q�?�\���I ����4��*gr���	֟�q������Γ����4�	�<q�g*6�hD�	8! kW��<A+Oz���Of�D�OD���O�˧%_�M���ʀf�x�M�/K�d@аi挤��'1��'M��yR|���#
L޸�ъˢM�b�_� h.���O��O1��(�+x�4扁o��")��m�a�F V-OA��*�"�҆�O��OJ˓�?i��sH�+ѡ�B��ʅ��<��� ��?1��?Y+O�<m��(�h�Iڟ��'lHI!E�'42��h�c��n0�?Y�P�H�	ǟ�$�����T\�ą���+��M�Մ&?3C��3r�s�4��Od���?�D�5����+H�H�pM�,,��d�OP�$�O��2ڧ�?��P�|�@���G�}��`���׊�?�]8��������4���ygo�:XRQc�v�kWL� �yR�'���'�S��i���O9���,�����	-�}"u��r��C��(	��'��i>�������џ�I���`�&IT�]���J�|�ĕ'ـ7��"bU���O��3��1Z>�b�K�O�N�ѷiӊ��P��O�xn��M1�x�Of���ON���̘V�(�Fi��6Lv���\;,Τ��O���o�9�?�0�İ<�A��bA�G�2ʚ-��F�?9��?����?ͧ��d�]�w��͟ p$0q�e!�By*fM������4�?�J>�V�d�ߴ	��&�yӸ|��� �e�B�H�#���:u.�MӚ'V���E���8��dퟲ�.�5G��|x�oR���(���'X��'1��'�2�'�����Ӭ,*(\ahN�r�0��c�O<���OjLm�<�b�#՛�|�L�4҈;j�8=��Cw�ѩa��O�Yo�-�M�'�vLߴ��$��i��5
�<6�Ph0v� "o�uP���?1�/%��<ͧ�?���?Q�7?T�K�&�;��0%ꗧ�?I��������b��Jy��'���?#=�U���6v��v��&,t2�9n��֟��IT�)� K�3z��a�����"<�m:c��
��<S��*\�l����-�ȟ��A�|���M�T��ERĽ���24L�'#��'���T�d(޴h5�	r�T�%&bh�U��7V	��K0n�`~2�p�T��*�OR�䝖
� M�b*T�ʤ����8��O��Gi�P��ӟ`�D��T���<��G�YE2@��oXi��(�1��<�-O��$�O��D�O,���O4ʧi��cmC7Y�r���OV�|��i⵳i� ��'��'���y�Jr��Q�F|z��lS.<
Y�K�m�����O �O���O��DZc��7�{����%�+*_�,��`�$x�����%g������[��,��<ͧ�?Q�gW7F�~�R�C���LR� ��?���?�����$���	Bg�e���۟���e�A��E`���q��a��s?��ܟ���E�x�D�bM
�RGFxVa�4�ŗ��)b����\nZq�'[6���ş�2T��[�tиC��6'���[�@U埴��H�����G���'K~<k�M�J�VU���O5p?*�t�'��7��]^���O0�l�g�Ӽ۳�m�tP�I_�@���*��E�<���iT:7W��! cn^Ϧ���?a�-�*~H��B�? �H�"b�7q�敊�+ �1��*���<ͧ�?���?9���?�U(�zr*�Å���۶��K��d�Ʀ�@�wy��'��O����58��@�r��i�E+�33L�
]�v��x�$���?�Ӿ���B.l��-�ǣػ8=�O� =��u3Bq�tG�OR��M>�,O�ȉ�ڻ���Q�k,:��i"�"�OZ���OJ�d�O�I�<1'�iӤ,K�7� V`�s��X���@��KC�'Z�6�;�I���D��A��4n��6���2TO��x�̙�&�ԑa��i��I3gj��¥�O�q�N�N	%��tp7M��i�� �F+��}��$�Od���O���O���+��	~J(�����F�ǧO�r �	��l����M��f��$�ͦ�&��rb+X ���������u��#Zm�֟��i>���fB�Y�u�-X>0�@ňC�./� ��ÁGf���O�O���?����?I��2Z�L�[6�m�&Am���?,O2-oڬN������h��w��\w�R��D�Ng�$X@��"���R]}B�'�|ʟ��"EŬ?�NY�Ѭ�^h��xg*.RȠ� �}�~5����&MD?!L>ID�"�����⇯+b��A���(�?9��?	���?�|(OTMlZ�U&��I�#�\Mp���8$ㆁ[Xy��y�8�hp�O���<5k&AST��i����E��{���D�O�B�Ma����K"WM]����P����KC&�Ze#B+.HԵ�7�y�`�'���'���'���'N�ӟl�<�#v�\�=XH��G"[�,#v�X�48������?!���O~�6=���c,C�W�ذ)rG��	�P4QU�O2��-��I8O��6�~���� t�T��>6�z�{�p������A��d6�Ĵ<���?Ѧ"H�r$��h@H�}F �ɰ�?���?����ݦ)��K�ԟ��	��@�N�?(�H�P$I� 6����`�T��q���� ��l�	P��uS-D07ߠ���2Q���	���s�-s��n������z���'12O��nH�s��(�Ց 땩\�r�'"�'������R�eՓxJ	��"Skd�qh��$�438XH��?���i�O�!L����F�+����f!�C������ش+����$u��F��H����}��$�ު<�Z�bB��R٩��>a��&�̕����']B�'3��'Ė�� E�i���%jH�N��P�_�\��4=�h�h��?����?��C�2=�`0��NJ��ݡ�g�C���	�M���i\�O1�Z`QA��K�&�Ԁ�	_^`��J5[jI�䜟����Y)mrəD�	Sy�/g���h�"DU�Tը��Q�0��'2�' �O��	 �M�W��?Q�>�|�����$~���L��?!q�i��O��'��6M�Φ�8ڴT�Nh�׈�u{��A@&eZ��f����Ms�O��;X�@��6�S�ߙi��I?Qn�y!����crL%�'�|����ҟd�I���	����B蜑-�Ȕ�U���X�T���G8�?���?�G�iN
�O\b�|��O���nͮO��`�j��9�E�v�9�d�O����OD�QpӾ�Id� .�+��<+� {a�h��
��)pj��~�|�_�D�I��	��<#�T�th����/X��m:'�۟���_y��v�hmh���O����O$�'?�D�� n�x:|�1M����'�>�]���%~�(�'��=\� Ţ+��XӔjDv~)�У��N�D]*�i~�O�����R��'7@���J�?�ΘV��> �� ��'���'�"���O��	�M#A@�����,K�B� �7��*��5���?�Ƹi��O9�'�<7-96�݂��
�y�ȍ�W�Y�)�ҕoڷ�M�v�Ĥ�M;�O��Z���
��O?	��Z�\} �}���s�z�H�'yB�'���'3R�'��S�J�&���S�x���o�3�~�:޴_S�p�-O��$=�	�OJ�mz����-(�Q�Ņ�i�Hlx��6�M��irPO���i�%4�6�x��`�k�;lE�!J©���в'"v����ۤ&�B�Am�Idy�ObKJ�xh�5ɂ�N�EB�L��ÃK�B�'��'(�Ʌ�M;�L�"�?a���?a�,ɼ@�D��W�"M>�� �J���'\듀?����'�Йtn��ѥ��$z9`�' H�c��M�r踋���������'��"0�P(e:����m�j49"�'�b�'�2�'��>����a?dA�����k�FA0�z8�I��MCvkW��?��h��6�4�B��u���2Hr���@��
�4O���O��Ĉ 8O�6�b�8��
'���E�O���w��"I?�8��yɸ��ӗ56�O���|���?����?���,�� Q+7�8���o��\�~� )OZ�n�&�&��IȟT��X��J���)��<��y�C�C6/X�0�[�������$�b>�qqN$���0a�%S�ju�@%�h��SQ)5?���@,,���S*����!X<Q��R�����#IG�}BV��O\���O�4���rs��j̧�y�&��f��&E�E_6MK� _��y�)v� �8��O����O��d
�C �p1i<ul�ĪG@�o�^I�i����ş��;��*0��'��T�w��p�wOܾ�R�rǜ�}����'��'O2�'���'���Q�KЄ=�IUd\�BE"�S"��,����Mˡ��\~�h�@�O�$)�HD1rƸ=��A	���#H+���O��d�O��pӐ���HI2�1� ���g�	��䁡#��~�c���~"�|W��ğ�	Ο,��'�2b"�5���|��Pu�����	}yRӴ��������H��N�0B$5
$i	�1d�h�����$XR}��'O��|ʟ,D�E9�r��r��!�f�s��B�md*�"7jlӪ��|��J���'���&�K5
D�Q�G�q#>	�֬П �Iџ����b>q�',7���X�1qVG]U7��3��x5K���\�ߴ��'����?��H�5H�m��	C}�`U�M��?��Sip ��4��d�K[ry����őY�
����wH�w-!�y2X�������� ��ٟ��O�N%���'�J��d��'���+W�~�|����O����O|��|j�{K��w��Hj��K�(�F����V�p��ȳ��n��ymZ����|Z�'��eH[��M#�'�8�HA�W�!ʺ���hՍ=&��ɝ'�~�b�K����s�|2]���)���`%[��I�O��0�@�ߟ��	��L�I]ybnӠD)��O����O��"J�6H쐖$� T�q�.�I���D����ٴA�'*��f�Q( A�PN]�,C�'��҂�̅���R3����3��czV�$�*=�'G6^�:Al��qՀ�D�OP���O�$-ڧ�?�t�69h��A��8p���zA����?���i;��7�'.�zӦ�杹h$��i,��I S�gh��9�M�°i*�6���u�p7l�@��1^*�a��Ob$�1�@�ePj҃/�h{�mC�nL}�IRy�OLR�'l��'�b�~�@�fF�\�T�5NZ�)R�	��M���,�?���?QK~��N�<�A�mL�^l�! �B�>�x^�<�ڴ;���5��i_� T(���)�F����
�����o	�[��I2�0eie�'�ڡ'�l�'�li0j��.��p�ǋ̕R�N-xG�'���'�����Y�8�ٴ7��;�'Kb9�솂GCpI�*ܥauA{�\Λ��ds}��'c��'�nl��[� )f")Ee
9)��H�4�F<O�$J!e����'?����?]�ݮKAN��1�Q�E�j�'�3TZ��	���	ҟ �	⟬��Q�'M�� �� 8� T���,��}����?�����F�M)����'#X7�#��]�V��C�)��1��� ��M&�`�4^M�f�O/\���i���O�E���`��	d��1K� ���8��E�r�O���|���?��88�SMns��C��
�����?I/O��o�A��������ID�4��:F{�H
��ae�!��C���D�r}�|��mڜ���|��'<�^d�4\0Sq� �;���	��V�m��qRS��o~B�OǺ���_+�'N�}!�ƵG�6d!�*� )@P���'a"�'���O��I�M[���RdD�He�W��D�[��1t�2���?���ii�O ��'Kf6͏�o�6H�f�B��T �@�U���d�J@n���J�l��<����سt�����'<z|���O�DZ�Lz���(/zn���'������	۟��	S�4E+e��1�4Q'S��;B�K�0��6�ӝ/�����O��6���O�ymz�}���&yVٲgN�1&�n��G�ߟP��l�i>��I��{��AǦa�|�x�qf��7"k�T����[O0@�f6�|��&�O��M>�*O���OPLde�$v袭��f� _Gu����O����O�D�<� �i���r��'�2�'Q<�Pc-�9q5δBs�	����D�Z}b�'U2�|���X��W,Bv�ɀcL��y��'v~�#���s���O����?	��O�aCf�T!z\6|*�I�;K�X�i���O�����I��P�Ix��yG���$81V�4n� b�(�?bX�	h��ݨ���O���i�?ͻOC���たTx�����6��Γ�?9���?��#޾�M��'�ReYy6\�S$�	X�S�8w�ID,$@�l� U�|r\�����	�����şh3J�2!��;`'�[���p��gyB�j�l�!G'�O6���O���4�$>kp0�2��.A�P�@�P0����'�7����5�I<ͧ���'>O� ��N�5���8����W����a��A����'��eBRR���Z�	ȟ�}�T��7���(X���� �1�:Y	T�Oh��%���6�N*?���Or�I	�{ƌ�<��
�0:��!dO�)=�PI21k�6�?��?���?9A�A��e���h���`�ӗ1PEK��2�����5�����Γ�?!���<>b�2(�������
�Z097B� ?{~��-��0����O����O���O��d�O�Ygb[)O0L[��Ԋw`�����Y�saM�3���P��	�O��dX��%��e|�|
��n>1'�0�����`jb�T���=�C_v� �џT����0�	�|�t�l��<y��r�R0Ì�W���
�^*���&�Ȩ2�X����䓔?�O��'n�%�A�p�HV*�h�ڱʤ��3�|=��0��E�3�4�Dd[A����'WR	i� �Θ�C6����?�:���'��|����b�$�����r�y>��O�R���\8��gGs�0C��),d�`���ΑɛF�����:A�$:�dԁ'�bI���\��q�A#WT�.���O����O��	�<W�i���k�K��(���fM�����s��G46�r�'�7M?��6��d�Ϧiچ��\�	�&]�fl8勆�M���i%��z�iA��]E�m2��O��'p�ao��{*u JY��Γ���O��Oh���Oj�D�|B�DN9~Ar�ш�>N]C�K�E�F �%^#��'�����'�z7=�1#�@�:/������-�\������@ߴGo���O?�5�&�i��� ��c��8q� m���E�D��!7O�B�ї�?��h$�$�<ͧ�?)7�C���q(٥)��]����?���?����$Ѧ%���r�����hP"BF���(�W>s|�`�AOF�3n�I��(��|�=Xe�FmϫB��pQD�B�P�	�\*��#m�fDm�V~B�O�����?i0��m8�\�p�Z�L��?���?���?�����Ov�R
�-6�H�3� ��໅J�O�lZ7$�tv�6�4�L�	�N�

���#'^�O�����9O��$�O��D�%7�6m3?ɗ$� "~���z��C�c#�xs$�+ M'�`�����'[�'��<��\�퉌�`���jE�+���2�[�h۴U�ZX͓�?�����<6�c�n���V8���@ᕿIa����@�	E�i>U�i#����m�~�[ �-Hv���$>w�H�G�iY�I�����C�O�Ob�&565z�F�\I�V�_�( <����?��?a��|�(O
]o;et�2mQ$̚elƯ��0GK_�=1�I��M���k�>	���?	�o*t �l	%�*,��r0@����M3�O��p3��
�(���Μ�b����?H��X�W+V���O���O&���O��� ��=#`�9%üזA��G$~�~��ܟ��I�MK���O~*g�&�O�}� �Z
"U�x��N/"6P���?���O ���O�Ia�g�f������Y`*��8z\5W�=�h����On�Ov��|���?��!D`��٢_���W� {Ȭ�
���?�,OjinZ3I��	�����?���C��I' ��s�T1Q�\2�R�H��Iן��IF�i>��+Nv(����1���� ��EMzm���rߠ�m�g~��OI�e����n��`1-��9�&(R��k�H�����?����?��S�'���֦!����D�8 ���'EO�i��f�P���b�����b}��'g�A�b�9m��ku�ц%�ʼt�'hb풇Z���3O���ļ@�^��O?�	�J��@*v�S1&.-ʆI�/��	ey��'o��'���'��S>q0���wf�`�č�� ��|p����M�s	�?)��?�H~2�&���w���cu���N�)#�E� $��8	Q�'�|�Ozr�'�}øiS��]�K�0!�t�٩i�@4���3O6!�w����~2�|\�H�I���!��B��ẵ�m�~LW��П������IOyfh�n���%�Ot�$�O�	��Ǚ�dO�[A�E	r� X<����$�O�7��I�	$��;��L���;PH��4��������E̘DpmI�!?���?���d���?������0j�t��T��<�?A��?���?���9�>���ʌ'*܈ʒJ� c������OH0o�3Pe��ߟ0sݴ���y7�ԩ.(fxx�GGt^��'坯�~�i:r6�E��	�%PѦ���?�ЪD�%�r��U[���סR%�Z̨���h�fl�M>�(O�I�O�$�O����O��P�y"α �����(C��<!�i��Q!w�'���'��O�2�ώ#Ġ��$�ܧ���a
���	�6z�0D%��S�?��S0U�P��*� }�zaƆ�+h,42F/�8K�6�bW�Y�Tl�O^mL>�,O	b ☴K{�uo��3����Ak�O|�D�O��$�O�)�<��i�ց��'��b��E<x&�q�LB�BA �'�\6�/��<��$٦��4M �fOнF[�h1�ED�p�.��y����6�i_�	�X���O'q����xa��ônH����Ӌ~y�{�<O>�D�O���O����O��?�a"׏B��C#�J�Լz�J\۟�����|�ڴot��ϧ�?��i�'BL+.�� d0i�n\�Xea$���{ݴ�"d�W�M��'��!�r:�@���R�<�]�aBP�]���QeB�ş��c�|2R��ٟ �I؟,���Y�3����&c��-/lQZ�Ɵ���|yr-g�H����O����O$�'�T�*5��;½z�@�)j��P�'Xr�
���Nu�Z$��b��wfS�}�!�բP7�A �;j��Q3@Yk~�O�V��	�V:�'8���L�{j���Ș�S�81���'���'����O��ɞ�M3��D�4x�l<U{赢%(O7�� (���?���i��OB�'��f� �/���"�׶y��T��L�S&6�RЦ9�+���'��d����?}��6@����s�b=�7Ι{��|��9O�ʓ�?!��?!��?������׀;�P��	�@��|�q����EmZ�Mw�=��۟���m��79��w��Y�#?\r$:�)_�#
#��{�"�m���S�'9	:y��4�y2`C�_��Y���U`\��&�y�J]�I�Z��I'��'��i>��I�s��G"��*4�cX ���	П���ɟȔ'@7m_%`J���O����
PT��$> ��`�����c��4!�O\nZ�M���x��!�Vy8��K�Z��8����9��$�1��Īԫv61�$�9��s6���G(G����c�Cw�8d�'�*���O����Ox�D!ڧ�?�� �1��h{0,��W�:���ɛ7�?)�i�����'~"jb�@������p�53PHQV�]���I��M���iZ�7Y�[�7m>?��̝;�i^ �6y9d/;�h%P 1��l8I>q.O��O���OZ���OD��`C�q���jc�7�2|+%��<!�i��@���'"�'��O	r���_}����C�1
��$�[�-TJ��?Q����Ş	 � �vh�"E�H}���3S����~��͖']�$���WT?�O>�+OFysR�ѾZ �|҄����}k �Od���O
���O�)�<1��i��	�'ζ�e*P)b�x�ćW�b!�'�7�,�ɫ���O���O�쩂��1E7d� '��̨�k�._�W��6�(?��nź(z��|��;"��S �#fLJ�(Sg�%|IB�̓�?���?���?�����Ox0IّCL�J����A��R&*\˝'<B�'Q�6M��Y���+�M�J>��	�~���
�/t�M�@������?���|z�ʇ�M3�O��qA�/M��))�m�oq�t��G(�����'b�'s�i>��Iʟ�����za�A
!�P�$i�<5��I��P�'KV6���{���d�O��$�|b�ǂ+6M@�ꔥw.�R⡟_~���>Q��?IH>�O�~�cG��('�\� ��SE������)v.D �Q���4�x�(����O⽋��L+h��yx �N�S�P��1��Oz�$�O��D�O�ɗ�*2����<�ջiI �C���H���*b��::uF�X�䘥�y��'hҗ|�Oo�I��[�F��!���K�R� �@��H͟�����m��<��iCε!ɖ(��9O�Hr/��"���f�Dta54O.˓�?9��?����?�����iA� ��)�3�F�x�v�蓆;��o�.��ϟX���?іO=r��yǤS0?X'�	�k�����j�*,r�'�I՟�џ ���
Ml��<yc͎��"j��د*�,$k#��<a���!V+��	[�ky�O<��ʶT��u�r�^7Cb���Em�*$2�'��'��	��M#��ѡ�?���?�U�R�+���)ԍ�5�,�ȓ��'���?)����:@A��*���#��^�J �'&lT' �8𽐉�t@ҟ��1�'��H���p���L���yٓ�'T�'���'��>���w�pw�����ȿ.�d4V��ӟ�ݴm$�'�7� �i�U:%G�v�@R���o�&� �m����ȟ����7�pMl�R~���	Bi�''��g�KC��@e�}ߌ�{J>Q-O�)�O���O|���O\��s(П^���oQ�8g���ν<	��i[�0C�'���'���X>���|��`�����.��C K�/��ѯO��D�OƒO��OT����wa��aJ�?ĺ�ړ(�8L8�9�D�s���8q�p{$�'즍%� �'����Pg[4�A����6����'r�'R����U�L�޴*](t���Z�����љSU0��N�;�:��� ����'��'P드?!��?	�	�==(I�Ao�:�04�aaG4UkƬ��4�y��'q,��V�S�?y��O��i��NՓ����@��0�
�rᘱ+�6O�$�O ���O���O��?-�a��F��1aG�E������K�h�IӟH�޴8�>}ͧ�?�@�iUW��%H�%�8s�n�}9�IQ�	����	ßT ��W⦩ϓ�?�K��8�
�X�B	�2D�`B��i�`���O ��I>)+O���O����O�y�ǌ�]��Wg��
���s��O~���<I�i��1k��'0��'H�x���Y�fH&"֒�����5u��eF��͟���^�i>����*���z��5$r��f��|�����/Y�	�r�oڒ����LI��'F�'\�xO�4�U���J<M
t�'���'n����OX�ɇ�Jd̟�7��5!/?������O	���������۴��'����?9��JnU
�'��f�G���?���J��E9�4����Ur�g�?��'����2�<QB$9���wW�Dk�'��	��t�I�0��ޟh��[��lӺQإ���H�.nz�B,'f��7m�z���O���8���O$�nz�	��O��{l�	��HJ���@Ɨ8�M�b�i��O1�6�q KvӘ�E%!`��f������<O��r���?1�-���<ͧ�?yeB���@�R�]� L;1�B��?���?i����d��h1��ß�����(KR�� e�1��
S���)AL�p��'��8�Mc�i�rO���:�VD�&�ѓh-�Q�v�����FЇVG�ܡP�6擀TM��ן��D4\TvBN&��9f'���������	��`F���'�VA�'��wP�Ac��cښ�ˤ�';6��-w>�$�O@�n�N�Ӽs��ܫG�u
��C���B���<y���?)��O6� ܴ����B�:���?����5o�Bupv�B�/w�}h��	M�IGyR�'���'Q��'y��ƿ|�ܡ�H��h�@!�����3�MCtG
�?���?AL~��	]:0u��j�HD
�b�\�	�U�T�I��'�b>����ۭ?`���W� ��Yib �sT��l����J�'ƙ��'l�'��z \�AT��e��b�4I�d�	����ğ��i>-�'Q�6��Z���� ��ɁA�C+j�w�R�[���dZަ9�?�W���	ş�ݏw�(Т�D�p��T�R�C��:7��U�'v�
 �F]�H~��;����d��}�F�qcU5�J�ϓ�?a���?����?1���O"����F�r�H�hIъ3YR@��'���'հ7�J��i�Oęn�t�I<0\0:�Ř"�p�3�)<	9��'�,�	��S�'$vml�R~Zwz\�h�ϫJ�H��B( )4�x�c�F��D-�d�<Y��)o�mё��܀��b�-�OЄoZ��M��֟t��K��@1l�r�b�����8rM�����Ox}r�'��|ʟ� h�N��K��(���p7��pLP�1�qG
c�v�����H{?9I>q�a�=@ l���
�b�8BmWx<i��i|�ʀȝ!5��`�$�-�d`�(�$����5�4��'I��?1w�M�sn����̀�l�@���4�?!�5l���ݴ����P�{���?�'c9��R=��T �?��c�'��It�� 
�I�}#��
��T	���M36���?���?��d`l��>r(U�g��K�����.SN@���Of�O1�j\��be�x�	�+EI�@�l	��E�� �0DB�'����P?YL>)/O˓LԼ��(a^�C��8����	/�MS��>�?	��?�U��?7ɖ<�D�	��9�t����'�J��?������Bc\�H%��7#�22���ABH~�o�VQ,����iR<���\b�'���c*pdk�&�Q�ntxL۬�y��Qo���;񂗦UB�h�T��Y�Rls�N-#���O��d��?�;V�p9�ǪU2�cG��PQΓ�?!���?�D��?�Ms�O�J�T�ov�)Ŋ�V ���T�Q7%RZ�%���'xџ؛�J�	�r����$�Q�6?��i�椛p�'���'���=Ѷg��uZ1��i�6�&�9
VS}��'[�|��$�B&8��xG˓#VFt컑��?kH-��i���}U Y"(���&��'{�X�4��&`jl4s�n��`�j)��UY��Gb�+>m��S��/t(�aV`D#�rCz��⟐��Oh���O��ƞ؜���(� Y@��ŝ#Dl`�j���v� ���?E'?��]''z^9`���<��iׇ:_~6��C��DQQ
�j���j���%/R�q�cB՟����Dc�4*�H�O��6�:�d�L�}�ą�7�,��E��o�p�O����O�)ˀ39Z7-6?��{��-�C�&kU�9�6H�{}|�C�����~��|]����ǟd�	����f`@�M�L�M�Y�|�¤T�d�ILy�'b�Z�"@�Ol�D�Oxʧ1�+$ωΑIw�\�*��4�'n�:��6�}��%��'$���WM���,(���E�ehr�]� ��zŌ~~�O!���|��'�\%(���+�܍�w`/,�1��'Yr�'e��OV�I+�M��`ȲE6�yJ�eW<���S��<(C���?1ұip�O*|�'G(7혙07x�ISgLz{J��Ea��i��m-�M���C�M3�ObّWG����M?�1wCkn��b�͝Y>���`�s�$�'v�'O��'^r�'B�� �V��f(֖M3�ԃp�H�[QRa���V������?������?1W��yG��9�3��j��]B������7��֦��M<�|ଞ��M��'� �I��Q�pwjp"�`����t��'lY	������|�V����H��U�c��Z&JX�3dX��J���������jy��u�>]�7��OX�D�O���k�,O.(pe � �l��)�Ɏ��d��� ش��'���[0��<}�A��P�i�����O�d[@oS�����C���?�C��O�#���*_
�ٔ-\+��"��O���O����Oآ}��"q��s/�z�6Y�1#�@���x����O��k4�'�6m&�iީk�����[g�W0$L�=�gc�p��47ꛖLiӜ��n�L�fJ����/���P[s#�g~<�6m�74 L=����4�<�D�O����Ov��8':tє ��NVy
F��3���%�6� �0���'���'��QD/�+�P�80�M�wjP}�6�>���i#�6M�j�)�O59�ʂL|��� m�ڹh�@���N�ڬ�����O��PH>�)O�M�#&�.'�bݘwO3�ڕ{f��O8���OV�$�O�<Ac�iu�H���'���FRZ���lʤO0� p�'�h6+��8���AԦa�ش��$��n{R`˗R8W�tAQO=���P��i��	<Mo`��O�q����8����-p������Y-\����O����O��d�O��� ��Hx~�d��$&�
PD	=ߚ��I��P�ɻ�M�&�|"��K�V�|2�R5	�]���9dp��዇�X�(�Ot��g��i�'>�6- ?�e)�����l�oF	+�I\������O>��N>�)O�I�O����O�����X�ti��K��<">�3�`�O��Ľ<��iB@ӂ�'���'�S6F,� �K	'T'd2�aA21�.�g��I�Mˣ�i=�O�ӂx;�9I��+o�����Vb�9��ht�&1�f!4?�'-�0�D@(��q,H��P�� $O>u�(�X0����?I���?�Ş���ߦiWNK%G\�8�풒��ܓ�քʶX��ɟT��4��'Fb�i'�f�R7C.V$�"�՞y�1ǬXf(7�Dʦu*&�ݦ1�'#R����
�?)��<�"��Zª\�o#�P��9O��?����?���?i���	�}�� ��a�	(������M�~�Tm��@_>`��ڟ��	Q�Sڟ�X����Ū��t�t賑iM&��� CU��rݴT���c3��	ݦT(7�c���#��/0�)���?�B���"m��A���R([��Dy�O�
	e�Υ�.�g���S�/���'���'��	��Mc�γ�?����?��#L�G�^�j�mĶs+��c����'.��w��֌{�ޥ$�� ��"�T#ԡ�K�$���CQ뗐9\�8V	$��;�����C��?���p�8sP"�C׈�ϟl�I���	���E�D�'�:�Ꮾ;�z���A
�(>I0�'XZ6'�8���OX}l�T�Ӽ�n�WI$���T��p��â�<y��i�6m���Uc�)�ަY�'&�1�a��?�"Y�f���p�2Uߐ�y��J>�.O�i�O$���ON�$�O����(X�/��ŚW�Bk9B�!�<a5�ir��!�'.��'��X��勯��H�@S*�T�1�k}�r��,l����Ş5���C��;J "�,ɥ+,,-���hd�p�'RX�X��K�T�T�|�^�0�능R�������72̞i��H ş`����	ß�cyR�f�Y5��O
��p�ۆ|Yp����4W�V�ۆ��OelZO��h�	��M[Ծi�7��!H����1�ɣ'a"�#�D�3��E�|�"�ͦ	�6H�@�>9���;uvɁr���F�'��lrϓ�?)���?q���?!����O���ԑY���lW��X�e�'���'��7͙�|����O�5l�b�"T���.�K���6Q^y0J>Y��Mϧ=S\���4��dp
��p�H�TA!� .�*5�6��c���?��1�D�<�'�?���?)���l.����-
0��2��.�?����\릡��o|��Iǟ��Ox"�`B�݁-���I@.FZ���x�O���'|��'ɧ��	�/ =S�Ǐ�V�в�lř�����F�J�7�>?ͧ	�:��B�	�1�$	���#3&�a���{�R��ğ��Iݟ��)�SKyr+f�n$h��ްT_�E�0-2�L���ַT*���M���>���Zщ	��UD�!ke.��6���H��?A�Κ7�M��O�@�
Q�O��]��!�%fz!YE�
��	�'�I�L����Iϟ����I]AD���ΠR�bD�w��U�p7�B=����O\�3�9O��oz޵Q�]$5�f�Qa�o��
!�T�D�IZ�)�ӛR3:1l��<Y�ϖ�L�̃�o8]~�����<�@ż:����h��\y�O�rM��NcD,h�/e���X�h�1D���'UB�'��I�M����<����?�d�;y
���/1�ؐ0�Hǚ��'���?������D����Q�l�&��J����'���ؒ�8�f����~2�'��U��]"��a�J�M�L%q	�'�bܑ��c ة�/�-��ڕ�'�|7�&JB��D�OF�l�p�ӼSlS#I�Р�[=wU�e��<���?���6� ڴ�����U�uC�?�"��;z4�	6B�w%|�I�Yy��� !�z��uc�2����{�X�D^��Nؑ�I�����s�' ��u@T�V3K���c���
	��\���	��X$�b>�CDΈ��aFU�dt�93�"la�0n�*��)_�e�'�'���;#�l��LP�tr���e,%��������{�!����ޫ9�W+�9Qb!�#'����	��M��r�>A��?ͻ�0���U��(pÉ�~Oz�"�+��Mc�O�=��JG���4��4�wU����.�#{�|�PlK2��,iu�'���'���'��'!"���Mx&ђ�'�̘��P�>�X�� ď�&���#�'	��'X6���Iw��O��� ��øvXЁ˒hʆC�$tr�lr�t�p*�Sv^�D�O��d�O�\�d#|�L��꟨�@�k�8�Ώ/�tiWi�]|h������%��)���?I�&jl�@V	U�#	be��BW�{V)67j�x���N�����S)������?��)�f�wM��
�F>'nnm�J�PjZ<x�'�66M�@�D�O��$S���i�|J���uC"Nאu�B�G�g(03LS���]��4������'��'a�S!�-x��9VǄ�9�L�$�'���'l���T�'�2S����4[i��C��ݒ'EV8�Sˎ�R�����<i���?�I>ͧ��D�O�� <.0)��͟�fL\u��K�O����H�d7�g��I.8\�Z��[@��'�(\ˀ�V7J��y��BǨ�ja��'N�	ʟh���(�I�����q�4�$! |	�`�(-�*��q�ʍ�7MMS���O<����ʧ�?!�Ӽ�v�\cH�� s@�;>EMU4�?1������O��Ol��԰fv(6mt�s#�H� �ȹCNY"�Rlg{���g�;��D+�$�<ͧ�?����ms���(Nc�x0�b���?����?I����[Ȧq�A���������*�Ä$��IZA��R�>ɉ�Wi�	՟��'R"�'_�֟p��b�G��m�5/��R�:)��4���Z�b������)�'I��,�(d�����\�c����o�0h�|I�cO �i���*�?�N�#M�;&�l@9G�D��� [�m�:|�,���J�E���(3,���)rf��/E��Hɱ^
CP��cj�)q�&,����o�u��� �.��ɲ���%Qʨ�Ї�S!8��,y��-S��3~�<���q����9���!d怨�䇳Q�*4n�8�88���<&���RB�|�YR$��_�L����)7�̊4g�SN�`Z�͛!���93 ȧ^_�����	�K#��R� mr�c���c,p�# �&]�Ā�E*b�ZQ���Ŧ��K�h[�}r�'�ɧ5����2�a�c�� ��l�e���d��771O��D�O��D�<eK�;.�h婵hՖ>RΘ��he�����x2�'JB�|"U���`(�/{�8��L!	w�K4��n��b�@��埄��Cy��
h��S�|����d�)
�i�i&Tꓥ?�������^-p�)� x���@7
4�課�ׯS�� P����ӟT��Dy�lҁ]���~=�g�K�3��]X�F����c��u��z�xy2`ә��'>tu���E]��[�l��&̫�4�?�����d��-�jT%>����?����B :]BcGS�Y���arN������0	-��L������ȯS�P�B/��{��npy"�Z�z	j6-Nh�d�'���&?)e���1[�`"��C6%��ɨ'�ئ��'2\����I'H��p��A�� �!�����fo�N��7��O
�$�O�)|�G�Lh��\54S�`�폪-���ҷi�:�ȗ�4�1O����: � %��&@ ���h��wDPm��������,���8�ē�?Y��~2�	6�,��	=b0Y��lX��'n�J�yB�'��'�p��)HD��"�X*W�`K�
b�0�D#j��'�t�����'���}��fb��j6���$0���x�@��<I��?A����L�_����J�o�=��[�>�PgL�Q��?�L>I.O> 9�͞�#�Up�K���!�����h�1O����O��D�<i����rH�i[�X��@�*_�i�0(��+�=!0��ڟL��f�Zy�����$�6���˕��HO�L��X�+����(�	��X�'qK��)�i��}@hC�r�~���_�P�6<n�\&�h�'*V���}rL�=���p%�����@B$̑�MS���?9���?��$���I�OF��q���E�v��YU�8Ã�5v�'z��''�Z����	�	�xR�l�&�.5r���Qr�&�'RCD�F���'��'=�$�'�Zc��j��50��	�%�VF�۴�?��0*a8!%w�S�'t4@�Kf��6�����Y*��-m�'?L�Iß4���\�ş0�Ir�do�7���/ �4��2Ӻ?�J�ξ�Gx����'?��Iū|-�l�rK���t�!��m����Oj�D]H$����i�O��	�Orݒ��E�(-�4)�!۝[$X-��d�T�Sǟ ���D��H�3)<P	���%���*6�ʀ�M�} �T��'�2�|Zc�\pEʶ���DH2C�C�OUe���O ���O�˓c��Ivd\�Uy�ř=~�p �& @� $��jy��'"�'���'���r�[�5�T�Ƞ*��ݺaK��4�bY���	ߟ,��ey� �*����<��Q��>?�XDPB��p|�7M�<����䓧?���5��1��'v��h��^sy�4�@�C6Q��O����O����<i%M��r�Sԟ�hQ.�)XѰ<����&�"@���Z��M;����?1�D�zd����	' O6%3�ӦE40�8��%r>6��O����<���]�S��S̟����?�-&I�0����xo*��6F�;��1$�P��� �-�Z����%�R �#E(R, n��憶�M�)O��Hc�O�=��Ο��I�?�ҭOk�3=v%���[�#�jI�6K��_S�v�'�2���O��>����q�0	�/)�|�3�i�p�Q�	����	�����?ڮO�˓mh��3��3\����
3(���x²i��<����/��ߟ|��/��G�l�u����vI��a�Ms���?9���(��Q�h�'���OѱB*@vfUp�/8�t��U�dF'Ux�O|���OB��
)Mͤ���O�.if,�Yq�>�ʴn�ԟ�s����<��������'G5X3�}��g���Yr%Ob}�b�7��'	��'�B]��'aP%v�aj��_��Ha`�Cauy�O8ʓ�?�K>���?�'��=a���!��Z�H@�W�f��bI>��?����D"aJ�'�ZY�GfN�~fJ��#�=��0�'qR�'B�	�����4�'�,D���E�yc��@���w����>���?����dϫdh��%>uqqb�8��LGG$7!4U{v-��M������4�z��?��_�~��P�b��(��p�U��+�M����?�)Ol��ӯ��S矸�s���'A�jT�k��DqcrU9uE�>�����O|�D%�9O�n~��([���h �p�7�&N$��_�,�G�C �M�ER?%���?��O�)H�iؤ ~�c�X$U� �iH��ӟ��I�ħ�����ES�����^�d�c�tӊ����I�L�I�?�ZN<ͧ.��x`&	�F4@��D-X&_��a�G�i~j�0�'��[�$?�f��q�O�q|�1��k�%!&�L鷹ib��'D���)��)�L���7��D���)LW�H����0��'|ƔP'0�ҟl��#Q��AH�Q�Qy�kדM\�m��h����ayB�~ڌb�@�{鮍�P��RE�&�G"B��(5�4g��H̓�?i.O��$�?�"9s΁69�ty���
w�]:�
�<��?a���'�����b�
}��A;n�\Dy@d�	Em	0�B��'!rP���	�E��'v�"q��n��x�"�FA�:�m���I��?��O2|'iBЦ��c�#�H�U��MP4:rJ&���Ojʓ�?9�j�,���O�T"�Xl$
���S	F4�!�ʦ�?���?A��0���'��Yv� 2`\�(y��<ID%Ђ�b�V���<A�8�B(�,�L���O���Ɩ(Óa�<n���j�
�,�n��%�x��'X�A�g�̑k�y��� r�HCݛg����i�=Nځ��i�剓!��tk�4b@��X�S���A�H�I[��P�Fu���7)�Y����k�ޟ4HI|M~n,u��� A?ͤyS����<6�Y�d�OD��O��	�<�O���T,�	�N��T��8k0$HZ�dcӸ�sd�k1O>5�ɶq@�i� ��*Z�����4f]�%�۴�?9���?A��pw�����'��d�9
�H3��;S�q�?_��F�'h�I�
�������O��d�OB(�1=b�9#���E�r�s$�ަ���*	|ց�I<ͧ�?O>�����'\v~xД�LmPD�'��e�"�'O�	��X��ǟ8�'>�(�m�}n2#U���*V��w�߲5O���On��<Y���?1`c^�	a"$�v+F�[���бK��G�����d�O����<���qF���a2��PBE�u�Y�Ug��M����?����'r 4�"��޴g��;T �T��T#���7��X'�T��Xy��'����V>��	�v�va��M�B,Y��M�ai-�MˊR�'X�ȍ�7M� I<鄬T77�a2)��_��"u+����Ο@�' ��A��+�i�O���Ƅ��e��� ק/���j��x�]��Z�c�럔$?9��]7"`��Z\杘�*�j���m@y�n߲U�6�X��'��D�/?�c�W�z+B�rTf E��Z�Hmoy��"5[�B*�	+��i(T�NӞd|b&8 ��CڴG�0hB��i�'�r�O@�O��-�����G�NQ^4��"[�sò�l�&;Z�A����`�'���y��'�Z�A��+iRLI� �
l��&e�6�D�O0�$�q5
�$��S���K1�# A��+ܮ���ʛdn�nП̗'�t�3c��~��?����?Q�$W��u"`ʅ�8����B�P�6����'\�Xs��6�4�8�D3����eY%��*�$FDҗ�v]�X� � ��x�'��'��Q���V��2�0�gh�O��XP�P�˝Y��͟��Ik�MyB�[�oe�0��eN0�a�F'�e1�T���'u�ݟ���ğЕ'lZ�[�n>-і�e"X��ᎠWw�9c��>9���?�K>1+OΡ����O�0`ǉ(y����GjPb9.�*��n}�'���'V剒3H�QK|b"jX���qT��6�r�"���w:���'��'��I�f��	^�����z]jXP�̕Q�Ù�\0��'SZ� �O_<��)�O�����[`���C��}�ǂ�=�H�HE}"�'���'����O�˓��TM&�Z {¨�v�}�%fU��M�+O��cW���Iݟ$�I�?���O�.M�CGJ!�o�i/<l9�ٟY��f�'���y�[���It�'j��P̭	��Dh"ϼ6��]nZ�By�Ȣݴ�?���?��'%��	^y��&K*8%C���-��?6�6-S���O ˓��O"�3u��y��,J��Q�働.��6M�O����O�8xօ�]}�\�h��]?���L,zJ����b��4�\ۦ���iyr�ߕ�yʟD�d�O���L�lv����bD�z�B9j�Tm��Fo�6��$�<	�����Ok�J�9�meA�R��h�0�١��If��Ɵ���ҟ��I�l�'34a�-�Iv�M��CS%�����-V&����D�Ojʓ�?y���?QU��%#,�+ �n����\�c�`�ϓ�?	���?)��?�-O�x��E�|��F� W�$�0!dR�uͦ9;�����'�\����ğ���	>�P�A'��!�E1\�"m��M[s���4�?����?����P*�fM�O�Zc�eP�U9bѐ����$��4�?�/O���Or�$D3�<}�<�LQ��E�n��S��ʋ�M���?a/O�@�f@�H�D�'�b�O�@�C\���X�"ġ]��t��a�>����?)��q������9O2�#^��ei�
��݀�@K��7M�<y2�B
=ٛ��'���'��$H�>��O�r�{F�W -KD�JVA'=~t]nΟ��I�G6����$4�ӵp�pr
��e� ��P��0�7��%fN4l������X��8����<�aY�S�EBY(/��3A`��Eʛ���/�y��''�	i�'�?��g��U@��B;I�})TՔw%�F�'@��'�(E�r��>A*O����������o%�7�
1����@�h�<���<����<�O�b�' ���R8t��%d��d��Q�F�'���a C�>Y-O2�d�<Q���$(�jTu�$�D)D�Z9"�g�v}+Ҭ�y��'z�'��'��I�"���/ƍNCXx{�֮B�d�ea���ĺ<�������Ot��O�lC��I6mF����Cf���3��+0t��O>���O����O�ʓF�~�y�:��}�gM�h9���C�����i��	ޟ�'��'y�b�(�y�	N�6:�B��lF��連`Nt6m�Oz���OR��<!B/UB ��џ�X�x� uQ�eYW�8���蔞Q�86��O�ʓ�?q���?�����<I,��nQ�P@`�ʎ19D,�Ĉ6�M3��?�)OB5°�]N�$�'��Ot ���G�w^�Q��~5�Q����>���?���lny���9O��Ӟ e~-�Q�W��Hk��]�Pt�6��<�T�G� �V�'lB�'�����>��n���ɐ.|Xt�@�Ep0��m�ԟ4��81����^��Kܧ9�v���ձ�.����K�Aa8\m��7���!޴�?����?��L���Wy2�O�����dYP�R�3�
h�6��c��d�O����O�Rh:� |�{Mݳ4�q �		���0q��i�"�'R�ߕ&֒ꓴ��O���5���t�ƍU���Ԏx��6m�<9��N\��S���'�R�'��`;Aߟ�����$�����f� ���>#�n��'��	񟐖'�Zc[Ԥ���{�-[�\�v�(��OZ��>Oh���O���O6��<I��<%�T�R�� Lq^��mt\N̓�Y�@�'�Z�D��П ��n���ɳ�d�f²E3�z�r�t� �'\R�''�P���c����TE^�>5�ȱ�J�/ ���@��"�M�)O��Ĥ<����?���`�~`̓}����9Ak������L}��'���'!�0=(V�詟R��J&n[x0��A�5����ܗ$�lZןė'�2�'\��[ �y^>7�Ғ���k��� /��#!�H�6o���'8�U�P��fI0����OJ���r�SS��=��Xc�/�"�Q[c)�[}��'`��'�Z{�'L�'Z�i9�hq�����<[����+(e��6W� P� _��M����?���J�[�֝=[2��)��l���V!?�7M�O:��ѡ'��$�O�ʓ��ONDՋ��B{�~	cBn˿j����4F�X�W�i�r�'E��O����Y<K2�`s ��e7�R�­P�`o�o$�	cy��'e��$�V�Hj�엘*0UrV�,��hoП��I某�!�V���'��O`��  �==�b�bqG�	���:�i�'�D��)�O|�D�O8�d�٪d ��/ng ���ƦA�I�K$ޑ�M<���?�M>�10�b1��)�I��I�%΂N
���'E2�k&�|B�'
��'p�I<Ay`�s�	I .�Ԙ�v%Z���!����'�2Q���	ß(���7��C�I�6��}�&.+�,�w"`���'���'��O�-�2
~>!�jR�e^�XS��ݳ&�̩�3H�>����?9O>���?�U��?I5i�;a���I%,@/鰙����d��	�@�	� �'阄��L=��ا!�f�	[8b'��21!�Y�w�ŦI��E��L�	�JUHu�I|��:*�!��D�"��*���3ܛV�'BT���r%/��'�?�'"�Ј�'���R�kB�( ��������Op���O|xR0O.�O��|��y�⍙i�x��D�X��@7��<1���$OǛF�~J��2C���q�E%:xHe��K�N
�k��rӜ�$�O�Y =OX�O|�>MX"���ڴZ���ᅔ(m77���-+�m���|��̟��S����?��oX��s�R9iuHS���S�m��t�]��h�Ix���?��)��8Y�%�̓R��a�b��Pk�f�'��'�����-��O"���xa�/��a���Z��m �L)��=A�\0'���������.��&���)��=���W>TfE��4�?�P̒�[p�'/"�'�ɧ5���K~8S��U�> 6)���D
���H1t�P���<���?����
3�&���g0F�yQ�:go��:C��m��?iO>1���?�UcQ*e�>yIS
ЂGd��$���n�B����d�O`�d�O���Zȡ;�La(�BU�hrR� d˺[v̙SZ�P�IП�&�T�	П���~��C�.ʔ��Cf@��*!�Yx�EN ����O����O �L��I�b��%�/l��$B%{Uv೔��2RT�7�?���D�O��'@r�i�֏!�E�#d�4gx��H޴�?y���䍥_9,9'>A���?�؇{0���@&��Դ�xfc��'g����a
���᠅�4�䠸"�i��I�����49��S�� ��$��k.hQa��LX�MJ$g�Cz�	Hyr�'��O�O֞X8��,hi
�$O8�l9�ݴ!�jqBR�i��'2�O�LO�I�!R�f�kT�Q�i�p���)^��'�����O$���ǜh:�L���K8r�]Ѷ�<7M�O����O���OR}�V�T�	[?qEF��L�ls���{�@1A3mЦ��Iҟ��I�&��)����?���q�f��p.X�&��2P%��X-��1��i��Z�������O���?��4R�9	aL��a4,�kb��u����'�6�ɚ'�B�'���'��s�l��j��:��4j�Z;��(qN�pQ�)��O�ʓ�?�.O����O ��>�8�C�ػ<n�c���!s 8O���?����'lA4s�<��Ȋ�܋����Ee�4"���C�iZ�I���'[��'�B��y��"�|M�W�֚8�b�{U@O�8qX��?����?�+O
��g�L���'�|mHd*�^�`�q�C�a�ȤQҠvӎ��<q��?1��7����?q��!�X��4��4r�͐�fڥgW�2�i���'��I4X���������O2����FAqC �F�N0	 �Z�:��'b�'�RF���yRP>�	b�#�ܲ9 �U�5\�a�i�ߦ��']~l�B�l�f���O
��򟘐էu'\-N��L;��S��}�C�'�M���?1����	eyB�'rq���(�YK��`h`���zr^��P�i�����Es�H���O8���Ne�'��/�`JU�ܪK`�����?t:޴td4Γ�?(O�?��	�T��i)�-
�(0��b 
P�4�$�Cݴ�?���?��狄��	fyB�'�DC6,r����^9q�blb�n	0R����'A�	*0�^�)���?i��,r6���**�P��̕0Aư���i�B��=
`�듾��O���?�1!80��b�
i�h�0gǌ�ZC�p�'� 4��'e��'b�'�B�'IBg)� ���K��	ކ����a��������Ĥ<������?��'�VX")%���vOw��t�ܴ~4���'"�'�R�?������|JQ��qv��t��n�ԓv���A��֟��I՟��?���~r�K�Qx؀a�k����'����$�OZ��Ob��O,P2�O����O���A W��kVcI �<��M�����u�I۟��'�Ƶ�N<���5u���s&iZ;�X�@զ=����H�I�$���K��T������I�?���O��'�k�l���@[��ē�?�)OF����i��j 
Z�X�b��� H4e�cj�B˓/f�ɕ�ih���?9�� ��ɞ�`4JvM�-]f�k�O'd�OQsG"$�I�?O4N����)ď��'�ƕ��i�H�p@�'���'�2�O�S�$l,e���:2�����;W�օ�6�fa�uGx����'��A��J�@C��`I�:%�����o�Z�D�O.���)�*��>a��~�� )��8��x�"����8��'��Mq�y�'�r�'� ���%J�1��G��0��sMeӠ�D�y7��>�����k��Nyʐ�)�
;E~�q�Q}b�:��'4b�'�[��iW�ȅ~�6l2wG�:�
��#�K�����O<	��?�O>���?����k!đb�HX:�4���U&��<���?����D9H���̧Q��9�
��WZP�gL�<h����?I����?A��\�'}Hm�0
�8>�ME�vi��ɫOD�$�On�D�<�G	̢��OZ"`S�eA�g��D
�,*Uf$K Kb�~��;�$�O|���O���Ձa'p�E^�G^�c��iR�'��	q|��J|2����e�#:��Z�&Mwj P�c�.��'���'������T?cg�؞(x�u`�o��UT"��� q�N˓W�h�%�i[맽?��'-���/2��"�M�������rk>7m�OR���2}�b?A8"%X"�d[��4^u��n��G$Ӧ!��ן ���?�xJ<Q��	�L=J2��L*X��	��Ai�q��iQ�!C���S�$��ЂK)�xA�O�"�MocD�M���?���yb���tV�x�'�"�O�����%s��"��S�v�ⲵi���'�����yʟt���O
���jQ�5��i�:�$��D�v d�oZ���2�LG+��D�<Q���d�OkL�v�.0&뗏<���g��':�	Ӡ���0�I����	H��'��ቇ*E.5㰘V���Ԋ��w�F�xPT꓎���O���?����?���S1��qP7hT*�JY�g�S	W�vU̓�?���?i���?/O�kE��|:F�_�T:%?��9c��0�n�}yb�'����������B`��k���>�B���d`���E��	�M���?)���?1)O
�1���r���5�b�"6�����J;<T $�M������O��d�O��X0O8�wD��{��L?B���"CK���ir�'��I�w �j��|���O���;pllm���3�4L`��X5MUD�'Q��'�R
��yB�'�ICJ���7"��$�6f�
P�bKզ��'
,�[��x����O��D��קu��"6
R]�	�({4������M[��?�%���<�M>��$�χG�H� �³l0�f�[��MkĈY)qc�V�'l�'E���>9+OH<��i60j�����0^�P���O�����f�L%� D�d������cF�)c}� 9уɒ2Д]@(:D�l��b����$�CF�>�X�� *$�OƄ�傊+ʈ�u�!���f��7Z�\ #p#��Q��i���ΡwT�C4J?�hy���l����=N��@��&��}�����N�T0��ѲZ:��� \x��5�Jif�Kd ��!5h` ��R'��p�ԸN������X
9��l˧��7f���)%kzEd�2��'���'�҅���'��i�@4��0`	�>Z:�m����Q�Q	U�mE�Q��.9j�$��h�N�'F�bH�(�4� �<����LT�
z�l���SIu�7-ժ3pACag�U>�#� �� r2�'�D��/$n��ʵE�A����I{�'@V�ӷ/�}��D05�Q+Z�x��'�����#D��G�	K�m��'�V꓾򤊆8����'#�R>]�t���:���Va��&ű&a׍H@�Iڟ��IC}�y��E�	�1�G��?�Od��i�Î�$��ɚ��۷HF�\i���v	h�� �Hy�v&7�i�����M� ����S�Er,�GyR�Һ�?�����O��!rw�P��)�hq:"(��<!	�_�zHb��jlxC�P�1�rx���-�ēJq��q��#N�d�!�ܪb��H���W���Ip�D��3&��'��-$�xS�]8F�� /7ɒl�a�,5~,A���	h}*�"b>��
4��9�@��<M�Lœ�(��[� ��HV�=��T҅�ا����O���T�� 8�0 2��.l\�Mh�dٽOU��D�OL�S�D�	),�AC��� �#YIY� B
�'���s�	Y4"�\M u.X3+��0���HO���cAX���J�s���BJ#S;�����(��D�@פ���@�����[w�r�'�h�8�oXP����A��?�Q��'� �	�	&>�d���\M8��   ��A�"x�X�$׾*�H�f �*�@�r�C�6h�92cD�9U���=W�.��L�v�
���.����	-{�ԁ��ޟ���t�'i"Z�H�vMZ��&Ee�;�4Z�":O��=��(�'%��P�]])�9`G�"��&�'^ɧ�)$�I�`�iSi��u�8� �92�tC�	�GJh�r�g��1OjRsGQ7zB�I�b�`u�#��[m4�Ȇo�+�C�	��|��	� V�N;V��^�B��6�-P����a�2�j#UqpB�	H>FU8�3��&L��HB�ɬY{��
qNZ�$��A���c�C�ɘ_����"�?U���e��9BʄC䉳^������K�ѫ��XkbtC䉝#Ę��vU�:�b\yl"!6LC�I�EOz�1����:�L�Y��a>C�I�ua�p��7G�h P!H2݅>D�`Q���J�A��K+�6@��&D��ɗ��
�&L�0��>  ر�*O�a(�M<*�v	��
���B"O���p+��2�q�D�_�m�� �"O�����O"
eniA@���xp�"O�I;�a�+y��z����$@c"O��s��ʕ$X �����d �iɡ"ON���i
7-f��:%�4J�$	�s"O�e�%.��A�b��K�`�B��"O�͋��L�,�r�	
T2%���"O��H�[�C��يQh	y�ui�"OX��8]��	6�KEp��"O��'�з?`�k7�	2[��h 
�'��U")�5�.�;s�ռ{1���'{.9CĄF�w�hA�]8�<,h�'�M����q�d� )C4L�N\K�'���l�%�j �[�n{��	�'펬�G�z��@g�d��`��'��p����=3��< ��C&Eq�y��'�(q�%(�N��X��r�����'/J�J�	<+^&!��E,R�|���'�QP�N$&Q0`0�n�45�L�h�'9@��gJ&\��d��Dۆ;��1�'��#&	��<�0D�S��:SV1��'��h����Jj��2C�,�D��'�<�[4߇���s��W$��`	�'�z��pM��+�rI��MY��>m��'����Ά�m5�S��3xԀ�'�A� ���h���"�@�'�F�2b 8W�<5�Q*����'���&F�akb0BΝ��y��'��[G!R�>�1�*�
q��I��'7,4{�G�
G��*)�#�LJ�<9
U�|hN�9��	*� ���+�|�<�U��T��������]���Sz�<�����w��P�ӥ3�-q���y�<ɣ��2�1��	��֥Rv�<Q6��4����TUNk�1x�ct�<��M'>o4Ș3%ڕb1����+@q�<	'F	�`^`	� �D��*Q�j�<��#ȏZ�F�wgA�dFDKg�<�g�I,IjY#�n >�� ǈ�W�<q���\o�� ��F,ܽ����U�<����%x�*�q��`�h�k�<iF��3k�9;B��B�`Kt �e�<����{e�x�wIL�C$����ώe�<!��ƳH8�i# 7���
��NH�<	˞�Yɰ�0���i9:�0L�G�<� �����

ufpS�ȡ	j=�!"O��{2,O*h��q����3�l|��"O:��
��Ox��!R� �v<rQ�"OҐ�B� ю�"D$��v�$�"O�h[A�ԥ*�FQ�Q�_�I
���"O��IU�@�#�f��V:-�p-
�"OH�(��{�H{0A�Ɍ���"O���"D89v�	8�j�	���R�"Op�ЅbZ6k9�+���������
Y �E��i�d8|�2�#V��%��`���y��E�
����T@L���(�5�~�憤�D�=E��oY�{��I���>Z`y����yH�$�Qiȶ>�.�Ȅ���ɒiu�}��'�4�� ��@RC��D@5x�TU���
>g{d�	bH!:*xкTI����B䉆D^������`Jv�׽&i�"?arJ��#n>��&OȊHW�`H2���5Q�+.D�����ۚ@�\�R��J� ~<��uf,D�h�C�G�T�����FhP�d7D�h��N�/�lS�c�=�J�Q�,1D�(�J��N��a1�UH��{�%<D���F�:�Bd��a?E���ps�4D�t�g��1E�:ใ,.HB�Q
��.D� J�:M�2؉5B�.v�tI8b��O؁���)�'r`}�&��*$d�yZ U�OH��a���$A�x�(�
Q��8aZ�Q�J9[�h����?I�	�/�|���*޵��O��S&e�8u�Z
���i �:EM�`�6�G�D�t)�y�M�d�kL�`q<��P@�Q��l c��77>�K��C]�V-2��N���z�M���Ѵ�6\�u��D|�=qdĆ+v�(���MWh��Ua!�_!����0�Y(K� DJ���T�7aϱT�\a�*,�2�)�Ջb6\��?,��)j��'�L�h�iҷ{5�������:�?���Q0~�P �2kF�QB�ER�jދ@%�'��d�$�Ծ��Ϙ'k��פl�"L�6��j��N��<��+�(k�3d�V����d�4'��;Ì�'aq����Z�a�$�e�[�7�H\R��'�4��a�K�wD�Ay����K:r\��b��e�P��b�7��ٸ�򄝏2b|�qb��a��I����2�NQ/,R�fK��fV�=�)�##̡QЃ�TE�ؤ�����&�;M,8�@��[6��x0���<�7l7�Tp��@ ���2�Է[�h<�E�' ��@�� n�H|����3D�?!���W�q�8��Q?5LH���l��'b�(А
 �Ϙ'�D�iV����3�K�d����F)���y���;7?T�I�@N�*�3�I*Um����	ʕ=��`Y��Dd\L|��@���|��,<O\\�a�P�M�}�cF�>�1:��C0ML,H�A�P�f�w�I�z��zA�B2ID<�j�����?TVR��ʎ�I���G{��)g�~9j���T����O?�V언�p��Ӽ��U�C!=?1�l�}0딇Cx>PT�ۦ\h�c�&D����pf��O�M�e�Ff�B�IbI+'�|����&?�����|3��� ���y"���J��u �ڼ�@(���	$bx�	}���*J�8t�N!��(OBP�+DD��B�L��h#��ˆ�'+����(� E?�Y���xA��Z&s�@BF�G�t�X��'n*�H��͚N1p< �#�
n�����$��$�er��C,\�q��ɰ'�ӉSE:L���N�\q�"O��EI�Qu]�#�-3���x%�'��]P����Z�r�0�O?QR0�K�I�X�x���Re`�*�
�V�<	���%9�XRmV�w��貣-_Qy�AI�]%޸�Þ��p<q� `�=��m
�q��E�4<a~�A��P�_��p�ƃT�`�"�HR��5�4� ����*��r�ra��R&j6��	A,�ѓ�� 24����FK)�����F!���e��a�1�X!/����U��������
\i�ᓡH�Й�NG4u3�/@sȖB��1')��`���5DΐU��,�6�tb�T��$�Ye�x����G��,1�#�+6XhB��U��x�薔�����F��}4�$(!(� H�*�e�I(<��@IAA����o�ڳ��B��'�'�qO� f�E^�
�(q�r� 1zn�%R�"O6$#Viś��e�c(��֙�<*Ð7h�qO>�3g엏S�n�q��.|��0��,/D�tiA/�V�Q��`�l�\�#.�	�,q\��'j������ +��R���Ѻ
�'ꢰ���^�J�@��S搨�(�+!��S
OV0����}(D�����{���!c
x)�ՏR��OA�9HAl�\b��J'��	�',5�t���ORV���N�
��A��i�NPE�8}r��Z�O��)���q����'�?u7�a�M�2��OD9`�a�`����A�Ih��g��hǯ�>q���X�'e���,b4p�$l��m�d�q��A�Y.>I�!�E�}済 *��k�X׌#K��%qm�#b�"��Va�=y����-sp��'
@^IhJģj�Y�4�
�p�셔��<{����m�p�'�y�)�3n�lT��#�3GӲ�1��y�1�
A��#4���R��v��x磈 4ʨ1�Bg��L�
�i�O��SB��7z�d�'%N`�1����вgL�B�lC�rE��� ��;��=뇪M@:�Ի���!�x�����hZ��Z�{�,�f��X�,J�k�&s�
��q%��Q̤X�l7�{��3J�E�ջ�U�h�R-`�cA�kĥXҍ@4?nT�W�a\8)�"O*���j�K�*��������ҽmV����[Kj�9���*\*6��<��>�.�/CȨ���� �����L)az�'���dL+er��r��I�N�z�cuj�@5� �ͱ[�9��_)v�^��]h�Z��4���`sㅏyВO.�I��Dy�����
]������ڲ֢�H~��i�1�j�Ӄ��:��J��K
?�zqZ�ψ�C�]��
(�8��E��E{�Ii5��%QY���ψB��\�aP�`�d�AT�V��hkʧN%IF�Ob�1�d]8���s�$Q:rJ��"N#V5�1m�-�f��,�11�r�� HRd{f���X�gj~�@�A��(��d� ۰
&F� 5�P�A�C^v��C� ��	SE]�p���8�m�8@[�"N0�9�D���
�n8)`u�#h���L��'+�t��6��UK�~�1A<I;P1����e� B�e�5Y�����Gc��hYD4�X�')��Q2������-��} �Iώ;�5Ä��w�"E�R�����O �k�)+�R�N4ɒIS�Fu�P���ABÏ(r~�ŊqgL'j���B�8d��� ��'`����N�49 �ղJ�zE�FA�Y����$M�1 ZL�t�W�d������).Z48��ĐWjeK��Yn��ªʧQjd .T�QЀ���'/@C��S�qT(G��'^Mn �wB`�H�K���j���8�``�R���V����݀FbF�	��C(W�a�pN�>7~,C��
U�%IhQu�ʑ)CK�,>��SQ�K�t��S��V|��ǀQ�	�hA<(Z��<i挤:(��+˭N%�(�/�~x��B+ʯJ-�Ӑ#��2��i�p���w�<��B�/x�� ��/J�9�G�1#���R����!L֘�:�C3	 � �<��b9�	���ܴV=��ZS�P%`6!�'!��.c���`��#�*��*�U`.C�	�:ˮI�T�ת��N�6t� C�I-Vi`���~�Ybť_�R�C䉗@����hۨ)��8��"ڕ7�C��'*���3�_m��)ɇ�
#�C�	�q�8��\�y��MӲ
#J*�C�	J��l� ��-M��r�!Kg�C�"���׌W긨{7��$[o�C�(0�p-�Q쏿��HfDѩ%~C�	3��|����'.����b��5�C�I�WxrM�s��=n�6�����8y�>B�	�6�h���<�R���-Z/�B䉟M�����1|(�d�h�C�ɣ1T�(�i��L L�P0�Ӷ��C�ɄQ
J!z��O@�§��?�B������+s��� ��*^*C䉢8Gh�(B�
�NB�Do"(�X��zLD-;ɇ�f�y��q%�=�ȓO���W�X/1F"�0f�\��DՇȓz-ā��U����M%I΄�ȓ�0;�͟7&ʝ�g��z���:9�H��^�=?�1���P�a<�<��9�%1�-%wrBU�ӮB<O~����N��@��鏬#la�[h���̑@�<� n��Pu֩�5���E)%
e"O��������Ԥ�)@��C0"O�,�C59|�6��e�p%��"O4B�D4Co�œ�!�E�pŃ�"O"��3Μ�V ���/�{ 4ɠB"O�Ȣ�˩Qcb�X�#	1r�0�"O����/ ]����$�ψtR �c3"O������Rڨ���K�	C(��"Ox@Y7c5rJ(Y�VN�<r$� d"O�)���$R�����X8C����"O� pɎ+e	M�eYE`IS�"Od�:wꋁ-R%z 瞣?&�Щ"O!s��*g�"d@G�¢-"�( `"OV�8�HL!�j��6K
�Q�@2�"OX�"�aP�~,f��v	U����Q�"O`���	��pF��5�2î�h�"O�� ��צIVh)E)�
{�$�S"O@��"
ؠ	SL���%D�(��ɰ"Oj�����<�u�E�X��\�s0"O�K[�9��kY=3���6!�C_����`U�q�Fia�*Xu!� � ؎h���8A�������!򤑲qȆ�Q�A��"o�.I�!��٫6~����84�`.P5Y�!��їx���0)C/��Yyƍղf�!��=4Ӳ����+5��m1�,կdS!�ď�SSi�+�J%Ae��"?!�D��+%X�mͯZ4� fY6�!�D�,p|��k�+�(vˈ�+���4�!��<.@�Fm�P����r��fm!��M�!_����/-5��]���#Xb!�� '��p�����qk1�B� `!�d�6�r�FN�;sh�]!�D�%/�`��6��C��u�&��G�!�dL�+e�T��?J�� &A�k�!������cA � |�л�ŻGT!�$�#!��B�W�Byr�&��6N!�$GJ<��֢ėI��qD���_!�$�c��%qr`�!P6�,HV#
 G!�D@�yr��� N4g|q,�;>!�D�K܆��LV�/f8�MM# !�dԵ��p��.��XL�FA\�!�D��i�ٛ�$�)W�\b�\;V�!�dϻ �� 
6�N��8ɔ̜<p�!�dj����d�>H��\8憰An!�����%�UD��2���H�#"7�!򤑕&J	�֎��.t2ܐPI�#!�� Ű���UT��)�g�^�!�d����EPQ
�HRr��s�Rb�!�ГY�ݢ�'�l= <�ׯQ/@
!�� �,7�� &kѐ+=�󮀥y�!�$ԲR϶��엇{�8�% �CB!�d1�0E����i�x����:1!�$�{M��·"�?���a��/5/!��	�fa¤X��b�X�0)!��,����cȚ5�NLJFcgIc�'����p�|��&�^��ԑ�'� ���Y�p��FT-]��s�'�D����6P\P|�oŅO�  q�'���e(4��tī��IN��
�',e���X%���*�tR6Hr�'* �I#����oЃ?�<H2�'�Ƶ*6�T�G���^q���D�6D���u�ٶwg�1���2"z�Ѹ`�3D�� r������Sg*
�o��B�"Oģp���(
�b�n�s�4�(�"Orl@C�^�K-R3�䟴jʲ��"O�5h�'���ٲ��.㎜�R"OH-1��0_�X� �w��%;�"O|h�bN�$/�IG�W�W�j0"O:�A��Φ4�n�Y��O	1¡��"O�e��W=�Z�cw��6Q���J�"O����
�+F,XP�E��A�P`0"OVX�7.�*���*�(J\��u@�"OJ� ƯG�G?��D�t�9r3�
w�<iP�K�r���K�,ph���p�<�&�Pj\�l�S��c,�l�<�Ue�7g�je���C.r�y1`�c�<�bj�e,�`���N�=���H�Ʌbh<��kY�my�$ݰX�(��G��;�y�N�p�Tm�Ï�!S�&`�����yrd�D���H���@��3U��y�#_�pԜ��A��3�XM:�)���y��U9�.�#� H�����y"�ݱn(�Ϳb�>P{����yb���0��d�F���Y掔`�G�y���'1�� tIA�U�-X+��y`�m���
ef�8G��:ŉ"�y®X$9����ǍגKy0�������y��آ���`�W�B�V@*��]��yK�d��s�!ـfRx�����yr��Cw: �P�+r� ����y�o׾k���
��P)q�ļ[�M֑�y�^5;���r�N�b�T���ʔ �y�H���Ȝ���R%e�~D����yr�����D��7^[< ���S��y2L��
�+�>cɒ���^�y���G+P\�B��6+��A����y2 \�gn�E ࣓>*i܄�3EU��y���z�!d�6 ��pK���3�y�i�$����m��d�H-9!�8�y¬�3[���E;_Ρ0R�>�yR�6x���1�^U�<������y���&J�}�U�[,a�BA� T%�y�i߷;��`�-�}�Z��ͅ�Ps�%2k_�<��X)���|N���=�bT[�h)m���k4E��=��@-���Od�а�!mE�pH�ȓ\z��س��#���Hd�F�]�n��ȓ �jp���;JҪ����n���R��驢"J#Dm\Ѫl ^���ȓ!0Ty��R&�<���� lꡇȓ� �/�Sղ��aK�!�`�<)ŌCM)�<"��Yݴ�9#k�[�<�ƢNh.MC$�^,U[�H3�Wb�<yu�]�8HpTNB+- (�Z�W[�<�M݇X���r����s�8�
�*�P�<9��H���vO�J�q�	�I�<�s�K���@�K¬|"9� �M�<���%u�s����#�U�y�J�Vք��O[�A0�`�M�-�y���!F~�)#N�*=�Qr�n�y�K9{T
�b��O/"מ�6�J��yR"��F���a`hÍ)���%ۍ�y­;��Y�AG�x,�ٛ���y���]֪p��Y1XH' )�yM�<U	�#uJ�0M~�̀7�D��y�(7+������M�P窚�y
� �)���a�N83shQ�kܖ�c"O�y	3M٨9F��2H^�����"OxȊ��.�P���ݮ_ʰq[u"O�����E;�~��6�1`Ĳ�`"O <)��πa�p��!��o���#E"O�2Ǉ�gO��v
Jm1 �c�"OHɘtJE.% j���"K�|����"Op�R f�;S
�E:bб(��<��"O�xgP�7CJYA��ӄ>���hb"Oh\A�.V0{�E��${�}�u"O~9��(d�Тv!�U\ }8�"O�p�&��bS��4JR$O�xQ)f"O���#^-5�����<A��)�"O����55�������O>� �4"O�؄��[�
�D�ӟ.�E�"OZ��a�S���Bɛ�E9F	�S"O�`�
�?��[�"�-ú9�"Oz�ɇ16��u+�!i��}��"O��@oJi���%I�+8K&"O��P�I��8�$Jt�\�H�u��"OA��a��;ndx��L�{�v���"O���S�ߴA�ɢ�B (���"O�,:��׫-0���� �bw0�h�"O����#ߤW�h���\�Sp�1�"O��X�'��,����@��(n�q9�"O��G��
,P������sg�ظ3�'Mў��L��m�u�W�f0f�h��1D���0�&2DI3(�_�\PRa.򓞨��i���GR���$x%�B"OtӁl��zp���R����"O�p�)Y0 ���9)B��`"ON�
e�In���Y��ݥ3�HT��"O\�Xq`�. lh$�(T:/$��{p"O6�9���BN,�9�撾><�}X�"O���D��([����@%N\u*"O�2�D�)*9f�Z+Ysٰ�Ґ"O�����	}(`��u��r�Z6"O���"��'f*�#��_�{�굑"O��F��f�`-�X�4rp�ط�Ii�O�����
]j��ꢇ�5�$h��Ğ$S�ƞ%/猙���	?�]��!�"�i��
$#�H h�'9n����e��| [" j���1��
v�ن�D���e"�8rI��c/�L���Z'��z��ڈ>P:�j�j 9\l؇��8e�ТO4n|�������pϘ��ȓY�˥�L��z�	9pt�T�ȓl*����
�U7p}
%�� �4ч�H�@�`��2��9
��ExHԅ�l�f Wc�cd�E׊X�����]�>�X��
:�͒��M�D0�ȓPC�ԛ�cnX��D�99��ȓ%00�VO!w8E���+�+<D��;�+�*^��SC�}R Y��	3D��PD0�����(�+x� ���+$D��6
r�1��
N�Y4�6D�ؚQ�0Ȱ����3\rQЅ@4D��̚V�|5ْc�]\���'�1D�a�
�n���k"��+����0D��z0Z�6t�U{�bب 񆕱�3D���gH6�
��Ժ �'@0D�<��썄~~�X��CV~|��WD+D�$�R�
Aɮ�R�k�J�%D�Li4�	�X�R\�'�v��h�%D�� �,�����p��걧��}]f�K�"O�嬘`E	0�GY�H?���"Oh��Q�,5�����kO/��ҧ"O�l�a�I�2�d*1kԨ-���"OL|1T�ss�X��D-f����"O�3"eİ;����d��R�Ƶ�"O���5.؈��Z䌈ie$�A�"ORi�$Oے'İ�a�D�L�ʐ8�"O(L�Ś�%o�p���K.>��cG"O�)˕��kQ^�*�L�"��r@"O�̑fe����bs�@��L3�"OTI���<[N��a�CV& �F,�"O:y�Woݔ%��c����q)V"O8��nT�}�t{��_��"O�Jч'}�ƁK��#/��x��"O�����Z;d���Ϋg�1�!"ON�$	�C=�,���ϖ�a
"O��7e��61ްA��k�B�KC"Ov��� �̥K�H΂���!4"O�<��"��4ކ5.)c��=k "O�@�H�E�L���M� 9�fD"Oz-�� ]ar9�D̀)s�Ib�"O�����L.���!�����
F"Oʁ�#�L�
��)�	֍<�xm�!"O��B��̛Y�<D���D�H� �"O2)ЗIBZ������Ŕf�$��"O\aa�Gk���-�4Xޤbt"O�<(֫�	q(�%8�-� U�-J�"On<P�f�,H�jË.##�1i"O��',޴k�Dm�C��1�$�"O�MZ !��|<�PIE#e��*5"O��(`�?z4�d12jX%Q���"O>uY0�$�%p4ϝ�-�f�Q�"O-[��_;Y�dC%[- ���c�"O p9Q�Ft�]:7��Wmbt��"O�"��pt�x�����P8�H�"O�y�@ �0rTcֈ=Ldٔ"O̴�f�	,>��6�^���@��"O.�X�^u��P���*�(ti"O�X����)5Vd�q��t��X"O�9��ar�iGaV�f�z5�a"O(y��K}@��"cR{� ��"O6�ر��?+��k���;�B�X�"O����Z�/��)"��|�2H�C"OR��͇Nv��@J�|(d�"O.pq�����\-����Xf�i	S"O����)�(�T�`%
�]�U9u"O}Q0@�Hn9��@�<�N�YS"O��B���yE�+��(F�X0"O.�+�jD)x)oC>�X`+�"O,	�B�֧z�d K�Η�f��W"Ol@�����B��0��K�	�Pq"Oఠ��\$ � �k�r��"Oe�� �<K��y�b�E�-슸�2"O�QI��B�;�h��OP�K�,"�"Oحj4!L�O�����('�ْe"O����*Ю%K�gF<�ơZ�"O�	����i.H������z�ٖ"O�ʃJ��y �h��ڇ5-���#"Oz��ժ�y�8���2$�x��"Ox�H��A�?���y��Z0Z �P�"O�t�B&+T����Z���[�"OҨ+"��p���t)��J�"O���`h��W>��8AM��r$��"O� rP����\�Z�̃Y����%"O�m{4�Q�T|����^��i�e"OV���(�B�"i"W�ħ �~��"O�MJ�g�[ZQ���^Gb��"O"�acDۭY4�Q�+��vc��JF"O��ǆω^��B5@��GI��"Oh��E�LS�-��^$ �����"Odِ�M��+�8��6#ǽ]*����"Oک��N��Z�(�"3%�8"O|�شO[r��ٹW�Еd��[�"O�R֧B'D���d��ȸ"O~lb�G8X��!b@�0�.)`�"O�`ؕN۫Z���X� �~�n,xa"O���C'L��ɣe��\���"O�Œ,
"��Q�� ,�B�
�"OrpK�AC�&*ze1��W�~�PtR�"O���R㏡���C0$�+]@��""O���,	�*�PQש0d@PB�"Oh�S*�U�,�R�K�ifzx��"Or8���O1%�(�Y��	F_|��P"O
M��M��X�X�CG��#NF��"O����U�I�(���%N\��"O̪f�Z�su*�8ÃϡonL� "O�Y�A�	9Z8T�#��S��-{1"O� �nM2jW`�"�
q�#v"O$�5�[2w�%�k����Z�"O
٠�[9�JT9�oW�J�J��"O(��W��8�d����)O�~SQ"O���"Σ>�=����#��09r"O`Ȩ�eE0\�PE�����F"O�-��+ �.¸��c��E���:"O���	C�2����l��aq��b"OT�ʓ�
�Q:M��L�	"�"O:��������C�MԾ/�2��s"O�LJ�NW-#� �r�G&���97"O 鲨��m��ܸ��?:v�$��"Oa���Ѱ[�f`8�Na�K�"Of�3g.�?�����N�L��E"O�!�,��������9h1P"O4�Q�ǯyζ�s�iԕn�j��"O�u!1nN;����ȕ�L�u�G"Ot�Pd\�^�8���':~2�ݑq"O:E�B�uӂ�c	&��إ"O*�X��\^�D �͖.e���"O�d�����_�L�@����w+n,�"Ob��5�Җ����7޸0'�=:!"O8jC$I��8�ɛ�N�~��U"O��"W�Z<X��H7%�^)��"O�|�B&�Iֽ@d'�5��`#�"O6<���ڀ�^�a�TtB`��"O�Hh��6��Q ��tiF 9�"O@�B�Ȁ+8�A��Ҽ{Z��ye"O�T�Sg�?)�6�#�#����[�"OjD:c��W���%$O͖�ڥ"OJ+���e�4,)&D�(C(4��"O�Yh"f�R�f��䘟(��"O��{�L��*V��b�ħ�R�23"O̡3!�ُB�2]0s�]Fn��u"O�PgHA6F����',F�E�u"O�e�7�q���b� C%Uj�!g"O�Pb`�I?I�t�0��7QlHI��"O�����ڷ1x�!E�BR<̻�"O��d�_�k�<m�'��/?*��c"O����P\ެX�"_�Y6B}(�"O� 6�g�qRD����+��@"Onř���Xˡ/�K�8��"O���b��e�~�A"�
�K ��7"O���?/�9b�N�P1�p��'d%����r���Z�k0}�JH��'v��Qږ&�T ;󊛭g��'>"926oR�M�z�s�ꈵ_錥��'N�q�~ �|cC�PM,����'�`x8��7G�h��HN%He��r���hO?��O2u�T�R��W��9EOQw�<�r+� 0W�����\�:�<Z�e�G�<� +�(@��A��ȊE�D� w/�A�<��c���܋C��8N��Bb�z�<�@[�J��I%��D���"�x�<QR�P=	Ԑ�^+�z��B!�uy2�'����S�L1O���if�)G��}��"O`-�� ւC�h	����|��	ZT"O��C����r�)Ң� w���a"Ot��rd��)O$8���X��Tȡ"Op�c�ܠI&����T ��Xp�'�1O�̋��P:Uz�Yo1R�d�S$"O�d�'I�2|m��M�,N�D:%�'�!��r��
��$P��,�b�0&�!�1ajxc��Ǐf�jp1�K�w<!�DM*�r����t�<��@��M�!�DM�S�u�3�J�0` ����p�!�d �2y�d�-2L�������!�$Ԗ��8jB�Ⱦ?�ၥ�@�-��d��Vvd+b��7�M�����B��>v} ��Μi�~=;v�V�B�I:I88�M�g�|ي�eE�l��C�I�p�Z����<�*���cC�S�C�	 &��u���� Q�`�SI M@�B�I8 �p!a4���)��B����)�hC�x��(�z਱�E/˒ՄȓhJ4��J&�2t�F�(RBj���U��bM�*?����#c��Є�w_ �1b��:Yߊ �&��~V*0��A�����L��\����Kך'��(�ȓ	�0��N�-<wn�*��@���ȓ-��0� �05E��ʕ�^�=��p�ȓnC��L��Y`�?s)V0�ȓ7, �VA�*p�<ȕ�4_����	Z�'�lpkDU|l��f�*^��x�'[�ق�%��;�-3$V���Z�'��v�_'ikm!/��K��Ah�'�xd٣��*R�R�r�엪B� ��
�'�&<��m�C0���%��<�
�'J�-���!��`c�R�4�������*�'3�0�� '.B�@����ρE삭�ȓ1"�}�#�G�tDXqgB6g�Y�ȓE�"剧lE�Xt����Gb,ф�*�Vx(7C011��`���SYR��ȓB%D��BkU����4��`��eDLʔ.���j9��հ,��(��
@T�� ��ac̏4&��G�'>M��
 C]ȱyP�CU�� �:D���S/�z{HXrD�7mh�X�D&D�x6��`�N� �e��[K�%��e!D�t�H��#)I)ΑZ(���*D��Pd#�7Aa0����R� r�i3T���T͂�s�4]x�EO�sN�T9�"O�Ѣf��g���c�D:j����'�1O���܈d|�!�`�ua ��"O� �<��i��@ zQ-G;[����"OֵS�Ŗa��c��Z�8�2� "O��j�@�n���8�"WO�U�"OP�����6��ձ"���� g"O�����ȴ4s�;��D�C���"OA�ᝧ/�4�P`)��3""OTPٰȈ�4"NY�g�w{D1�"O��0�Z-[U�����"�0�"O*��R�9�rݫ��̊[�ċ�"O��{�r��r��[Mt���"O$�	R��J*b�� LV�#Ր��7"O����=FFp��=1N�B`"Oԉ0 �K*`����Q�CH���1��0LOԄȳ�^,�R胶�ğczT��`"O��X�@�~��9:��3�ؔ��"On0�
˜�:�Q�I�0'��% �"OL9�#(��l�ڝ��g�fY2�"O��ī��t% `�V�5�Ա��"O���W���)�!{��ĉjaT�a�"OT��t������U)�E��$?LOxY��S|�he��gFޑ+Q�'7!����#Z��Α>��y5"[�!�d�=B
8�qҏպ|���S���<�!�d���<��&ô0>Yk ��O�!��Ŀ��]� �΍ZZ֬�1��!�D�~�4���$B���w-u�!�\�XV��P�ʹ9)R%��.BS��'2�'[�	O�'��$���J���x��P�x(����h��ə"�xy	�ͭK���т�TC�I#����ɀ,u���%G�\JrB�I�>1���t�
�&h����
@�B�	%x����L-�&`j��^'�B�ɥj	��Y�PF�Ɇ�xLC�I�]�4��c	�I�`� �X�e4t�=�-Ox�?9�$ˋ�vD����[&|:��j���U�<I�L���HX�/���%�>m�nB�ɢV|����c�m(IL��C�I)o��jl�-���D
{��C䉋A�f��2�F9��p����C���1{é��=z��q2'��W��C�I"f�i�Cg�g��ٓG�60Z�O�d�OJ���O�#|��eL6"�0�l�_� ���_f�<��ٔ8�Q�4m�Z��KP�Ni�<��&O$a�ƹhdZ�?�����bK�<�WJ�{c������}&p�b�}�<Y�g�2ev%�rAS�0����|�<�c��YH����ק1g���	�|�<)c��V�UGS�{|���@T�x���O�bH����/��(��.
3����	�'>>�&J��z�脪Sg: K�k	�'�fU��+|CjXP 	eߦ1|B�	�v����Ԯwm���q �#l�C䉒|��k�ȍl�ذ󃟒��C�+[Έ���R<v����%K_�(��/�S�Og����a�m1z`�3�#B��Xqg"O̭҂W��L��c�B{j�2q"O��y$(���=�d�^(@^2�Z�V�F{��)C�r�����-�`E���ً@�!��òb���R��Hp%F J�O���!�D�ZY>hY�hא<��B<��'$a|"�DP�
)(F.�	\BP����'�ў`�'���R B�zZj #wO	Y��l��'K�h�҉�(�����bD"N�؝#�'�h(&��b:%�Ə��E������� �s�?>�����̄����e"O,uIE#������ۉA����"Oġ�Gm�! QQ�?GId��c"O�U��>?�TY���*�"hkq�d1�	ߟ��'�PaC���O,��a�h�Dl�
�'�x|�L�$�&)��ā�zm�u��'�|aSG��S����a�1<���[*O8���O���VA�uRL���yI�?�!�DE�{�4�t�Y�;|w(Ɋ�!�䎲i}�T ���2D)r	�+/>!�� o���Ȋ�����~�!�X����CpZ�5�$��X"D�!��ob�=Q�	|���6J�!�$��qr$�A`*5�ej/A�!�Ε*	��hç��,�̡�4��V!�$ۤ|�J}�3(�:y�=B�ه^!�ĎѨ�,Vm�.�"�11�O��d-���r��fz8� g 5�H���'�ўb>�'׸�R�)
:���L��h'(
�'�\u�1+Ģ;@��OY�Z����\�,%�T�'�9C�䎛i�b��q��
P��4"Ofx�HJ���A���ഴh&"OP�1��-cd��p�],��Ђ�"O��;�%I�)>h)6jE4d��@*s"O6p�3��+�b}T/�gs��3GOz�a��N�XA���^�S���9�	=D���Wk�Kv�L�h[/ ���9��hO��I;R�k��ūn�b:1� d�C�_rn����"F�z9�EfK0^�C�I���]��m��6��M��'��R ~C�?>��eB�ѰjS��	3�'C�ɒ&dR܊3o@1Q�����C�n���O������;$����q@)3�윰k�!��cy��A�-�5�)��*]��!�d�Pt����$Uz!rA��¸R�!�dۮ[p2%dB���x�� �!�ɧ<�$u���	6X4&+@0{!��V'!E�)�A��7c4�	��J J!��5/�;�c�� %xA��O��Y6!���!QVp���<����K'!�$؞jE~�q�ʷs3 ���C�n!�Ͻ-+�\�Bc�{��`��y�!��]%@��%@>h�ڜ[���"�!�d\2:v��&�H.C+X�Va���!�$��8*�Z���9�{���h�!�ׁ�0�H2&�F���1W�!�dK!`��A�DK�uѪ�a�nO-0*!�I-Fp�W���d��q�bcǓCm!��y�.� !i׹6�,\��!P�MY!��9�YJ3��-��fG�M!��Q/_��u���
0�x���:j7!��_�[��*��1r���rml�'�b�'2������;'+ �i:�L�
I��v�|͊T	T8gu�IU*D���ȓm����X�bQl�3��ղ%�(D�P�7劏�1vؘ���w�1D��Xp��"��p*�R$~kp��/D��YS"H-xh�����E�4%c�'D��[�G�0O��M���܍%��l�R�'��G����]�ܨ���H�\Q��͙\'nB�I�%�4�C�*ܿ,ؘm�P�M f�(��0?��l�5k
�z�!�o��19� _�<�S	ֻC��tY�oB�VB�sR��Dy��'w���'ܫ(7T@#Y=f&��x��� �U8�AŹ.�����A����"O:,H�(ԅ9��!��D�	���D�'��'�r�'�ў(����/z|JI��킛G��R&f�y�<� �� v�!�.�1��(2	~�<����U��4z��M�`�֌p᠐z�<0A�)"��2`��%; �ЅLv�<��'Q Y�p�˚%I@0=�G�s�<���ۯws ѐׄ_�!�a{��l�<1�,ĳG�D�C�A�q��E� B�]�'FaxR
Z�+e���@NԲD��y���,�yR���D����f�-{~��dA���'laz�a����ڷ��1!��l�S�
��y"�S0q�;���3l�1�#W:�yRHO���B1�î/���`R��y��9�J]����~���KC)��yR��6{Ӕ�)0/�I�h�R���y��X�in��U*�9����[5�y�M�/{�K������yRR26n�'��4�B屧�Y��y�ß7N�0yP�S=p�4Ӈ��y�ÊV�H�B��D���
g����y���0��9�M��C0�ҡ���yR�V�KmP�����:4Dj�Pb#���yRB>co�u˂�R�&(�0񢡃��yf
��.I��
�FY��C�(��<��D��t�\��r'[�N�����A�!�F�
�j,�GD�E��s%��9!��/:Pxm���K�f � V�Y�!���4.��j#H�q��5���GLg!���=Ǒ���/L�ճƍN>�Pyr�L3p�V���m��Jw�$� �y���E;2����J�F��T� ��<A��d]�<႔*B�P�h�����!�W.6��q��/$�
��@G� �!�䗾t�hz��W��J1`<2�!�dF�FX�g�"h��%��Ӑw!�D�	jeQ��I��"Y�sEY�n!� ��i����X9â�}P!�Es�T���Y\�� �"+s!���Wg�鈔��S������1c!��&B~!{Q�óQ8�����<!��	w�D�c�͆�*rP�s!��`�~��`ҜC)�����x�!��)=n!ҴnG�wo�]����<<�!��q�b����Mbnʸ�``ҼJ�'5a|��ǆ{>�$�V F�B ���,�y�D���������>o��jO�-��?i��:JŉŠޡ�Z��EなDL^���'�5�4'^4��p��LI�'(��'�J|Ka�0�����Q6u$��
�'-\���E|Xx𛖀�{05z�'��XA���bI��!.r��+�'��ڵ��?�
��Ua;jh��+�'+ܘ�@LۏJ�,��ANf���	���'p�>�I�t���s���2������X;9X�C䉺
4 �Х@�!��Y5��1_LC��v~��pt2F":��¼:LB�I�\�>�u�ӸGT��Kf�V&ʓ�hOQ>A3���ҕ  
�c"ΑKA6��+�S�'l�V�z�n��L����A�,�މF{��O-p	{��C�t�]�ѥË>���#���2OH��� nnZ����;�"OB%X5��T_��(����I�r%"O�P����h������xyr"O� �(tNB�VJ<Ӂ�F$j3�=1�"O0%����LӔY�N}��q�����O���*�'~%: (�ܵ1�H�ڧ��7T��UD{��OÎ���	�%T�1aɄ���0�'_����E&zJ�i�A��]��h�'t.8j�I�\ry���5Q�^� �'� �
 ��8;�^mkЬM�Ih��Q�'�y��K,�XA�n_�4�@� �'3�M��lL L�"��p�>.'����'�J9��'�x�k�fUxlN�*-O8�=�O��	�{�씨���*X&������B�	�
D^��X�M���`��� ӸB�	4$�Q���6Y�$��3R�*�~B�I.A^�s��@�J[��B�O�X�jB�I��ʹ��OK�|���QHdB�ɩ�6Az�d�(8B9��HU7Z�C�I�~_L�G(����*w֋�n���O��6��?E�<y"L(,~Ёakׄ�e�g�<	�ˋy�j@��C]�F�|ʄ��b�<ٗ�O
wi2XZpM�����΍a�<�wоZ���z�W�l;-LEh<��k�#E�$p�� WhHA�mP-�y�h�q�@�#l�S���U,^�yR�� ẽ��'6M8� �wh׊��'�az�f�c�B��Fg;I0��1a$����<�J>E��-�;vpQ����FQ��ٖ�y�̰B%H��W$�P��������y���;�L%�ƥ�K��(!M����x҃)g5�g;}���`� �vX�O�q���u�΅�v��B<b�'�ў�G|R��DD��!B	{aĎ��xX �c	�'�N��h_�Aj���cͅn���I����D>��ӧ8����Ӟ@�Pi2Q��3"�@�ȓj�,���U[��Ń,A� �ȓ��f�#'�2$��BH1µ��IR��+ԃG5L���hAf��ȓz���#g��a锱�W��,G��%�H�	D���'��P���6.p)B.����i�
�'4T��D�!�6A�h�L�"�'�<񡣢��M<b%As�0*Xe �' �ԛ6�T1d���A�M(T.>�#�'J�L��P!"�e�d焳yk����'_naaAbډX�P]#$��7D�-A�'���q�M1||ڳ�Ք'V޵X�'��5�
S���$���iIP�'�l�S5�		B����𦑍5F0���?1a�Y(Sr��D��W�iN��y�j��TB<��A���'
7jbj�ȓx<P����(���dԽi�L��ȓ!wj�b �X�!�j\����]0Z�GbZ���|z�F�"(������̏|�X����p�<�hO
)��L`���p���/�B�<��X)B��u��jܻr�ԙa�AB����
}�Ji�fM<^�$�b�<'fч�6X��c�<_�݋v뙒o0�ȓI>��#�A!"w
8r.�la�ȓjkԠp��T"��������]����P�k��^?i"(��� %l�"��+D�`��J�+P��4L���p�&7D�d���܄;`\l��K���) 6�'D�\k��R�t <h�$'Pb�mvA&D�����ԙ(O`X5��$��!c7D�d��� ��p"�/һ3�*e*!D���Ƈ��K�q��32��Y���<I���3� �I�� 	&J%��s�ݟP.�ѫC"Op��	8�`]K�&��5}��J�"O~��� ��:�dX�%�+Lֹ�"O�Ih�+̪3��D[ě:8r���"O�kK-_ 	���u-���!"OD"
���\q����7^Q�b"O��(J��I�<�b≲A��hr"O���I*#N8@"��1�[��"O��*��� e��u��,K�Te*1"OD�c)]<	���K�\v�س"Of�C�� l�#0/^�9jr8�"O �����(�FH���Y�����"O⥐�(��z�$��Y�G�0a5"Oҍ���2HZEpvL�~�hya"O��0��d�T��d��|���!�Z�����<Ȑ���זK��4a��݅5�>��0?yv�ox"80w�N���ㅂ��<�7k�?R8`eM�g�8HHs�g�<���ޕ&�N!�Aؖp�fP�g�<�ĬJ9>�<�הG��p����k�<��h�&������րy`��j�<1�,�!H��ȋ��e��^�<)�çj�f�I���!��XZb��o�<���AO��8��FThV\��h�<9p*ԤXgj��g��2.ҡ�,e�<�Ta�,<(1� �n����Ϗj�<aǃ_5phLrD)QtӌP�Ԥe�<Ѵ��?���
3�s$\j7�]`�<��-��.���_�|��IЁw�<�6M J�E��.J7tD�Q`q�<���/i����e����)adX�<i�o�>X�DPF�
&����TU�<բ�>0,)�f�	(�F!&bWw�<�P�յMք��p�z~P�0SMAw�<�J_65�
ic�*T1x�� �w��o�<�Į	N���h�N��)�ڑ���i�	hy�X�lD�d,FP��] ���$\�=X�З�y�!S��: �C�RN�L8���4�y2�B=��
�#�>ʅi �R��y���3��$4q($��oC$�y�-�Pf1�B�-�p����y��^j̖�q�������A�y�#O�V��Xr6W�%@CQJ����?����e�4 )JgA-n���g��y��s�N4�E�l� @9��Ƃ�yb�Ѓp����@g
j�n��CD��yB� 6����s`��y�t��C!K��y"� 06��W)�q�؍����yRN�3�BkCѰ��eO<�y"B٪ H�#3Ɋ�e���P$�]�y���>ltM�-V���s�ߢ�y�O̢O���P�S��ϡ�yK�i��q�F�\56}���S��.�y��d �(�R$)St�R�R�y��T"�x������\��y�޻0��1�6�Q�Npa j'�yR`	i��ȁ,%b8i��_��y��0�v�H`lV� ��sCG���=y�y��Z%�X��'k[�qQBtS�d_��y©$E�J�sa���A�&��y2ć�;�h�.�|(zY0�Cѧ�yb	S�*eʭsw��y�T�a��
�yb�пb��YO��oTrd�a���y��܎N�b�h���=f%���a�Ӳ��'!az
� �(Qq��5���WE��R���'`1OQ�q�֏z|�`��IQ�����"O<��U,�G���q#/�F��l�"OP�g6w1ܴЎ��|� j�"O�	;��I8x��xe�G9f���"O0I��$E�i�����G��ʟTF���ܫj����@f.9FL@��ˈ�y"���U�Bꞣ����uc��y�"�zk
�R�-�v�� ��y��= %p0Q�CA�iX��S�6�y�
6 xb�]	Z�A�R���y�dJ�"���q��V�f�I3�Ρ�y U�|��1�D��#��-[��K,��O�#~*�c���P�3� ������W�<�dO ]�\�ׁ� w(�A�FQx�|�'��Yk᠂3/ǖ(y̆2/.�B�',p�eD�U��c�&Dv{�@��'��0�2Ù"E(<=A�Àp�*��
�'C"P;�ҥa�ک9�
��B�	�'�8d�PC�Gv�z�f��G��A��'��u3���M-:(r�a
:+88�'�^e3ǭ�/)52�pgIZ2g%�
�'|��b���$	|�	��7m�B��
�'�p������Q)iֆrH���	�'6H��p*C	7�(p[�A�:d�d]�	�'J���F�P�,���!�I�T%�i�'�T��/�� �b�ү9z b��O�<��3�Z�3(�b ���"O�
�c܊X1�Q$G �aP"O(Qb`�/s�&8�E��[5�U["Ox����^%�0�cg��Ib�"O����bġvmvx�lD �b{"O� �SF��$����P	�v0ZH&"OTA���(/��m��C�B{F�1�"O���f)B6��dj�,�8n(�@�"O| H�E�p
�c�+^�H ��1�"O� s�f��a,b�B�,.A�<��"O�%I�)��%j��@�%�2$@�"O",�`�O��x�̉>&ՊQ��"O�xч��H�>�k]�#�n�3�"O � �%¯ex!��ĚX��9R�[��D{��ID#���Ȁ��l2T+�X�!�DW4��C&�./��w*?.�!��L$Z4j��Z�İ
I�G�!�D'y��q�d,GzD1�VH���!���t%��T]���R!�#b�!�D�v���a��J\qqO��v�!򤓋;�Sb"�\�䐨`��!��۫%Q�-�s��r�>��M-�!�DA�8�V�I�vnQ��Ã!��
c�p�@F�qY�%Ⱜѻ`�!�D��'Q�����c3����BVQh�C�ɺgE�`��
)X���F� 	tB�	�GZ*�� *��<n^E!צ��'�B�!A	�4���~�k��
5K�C�I.24-J�A��Z��x(��'D�8S�XctҡI���جc� D��4)���NM�5�VF��4��2D�P��i��Pq��΀�OJ�W w!�ãFB�@�2�"8�:�i�@V&J!�B,!U��
�"F�\��a����S�!�L6����Y��RI�`��!�d��B�*��2h�w�\فO��7�!�Dd�0ؑ�������o�3�!�� ��!.��(�8�G�}4��E"O��1���G"�P��D��Kq"O�a��C	!�.����&a9���v"ON���/e�t\��[�N��"O�u�䌓+�h��a�I=��c�"O2�i �
�d~�#Da��
�Lm	W"O��)�+��0�y��I�j
г��'�ў"~ҥ��A2����F�*	�A�����yR�M1-���2b���N;Q����y��� >leSWB��K��d�alP�y���-i�$����,K��!B��yR'�Yb�{�>0�I�)A�y�K��Z�:`�2B�8W;�IY�%�yB,�?_`"Ԡ���|;d�A���y�����6�2
Q�|h�)�)�y�	�
��U�E�6����W8�y�R45<�j�_(Xf|#a���yG�T���b��L y��M�ej
�yR@
3Nҝ�רW� Фux��	2�hOn���O�܄� w%���t�X�-�,�[%��2LO|=#�n�� S��Q�.A�k�\��"O�Mٴ���S?��)#^9x\�S"O`�Z��
bb|0�D֩~��P"O��	�;xf�Tz��Rf���h�"OV	{�#I TB&5�U	�.�7"O� �pፙ?�J��� � d�4"OĈ�RJ°�;���<�����"OFu��R?���fhva\ 2�"O�R��ˑm2��8���9`L�r"O,y"���X�q+T��<o58z�"O� L�ǌe��g�!B��)3"O���UBێ�^��"�Ȟ)@�
�"O�wݨ^
6؛�)�A���8��'���C�i>y���@�a�TXCᑿ>yR�'N��y� �b��p��GnS 5�v���y��U���]��.��l�&�Av(Z�yҥ#1?x�`2	&p��:FhJ��y���	�N}���G Y��bR��y��|���1�ou$r(�y�d��?�F�9R��z�d��ܣ��$:�S�On�K��;��-�g���K�M��'�<A�E<\���"�W�\���'UNe0)�'y�!�2B�'^x�b	�'bB9���B�v/>E��H��X�\H#�'Rz���hH0pn|a�!���Ȩ�'t��S�\'�q:D-�#"���
�'Θ4S4	#}r�y���;F�����hO?)R�$�B�CB"U&A�K��B�<�t)�[�b���^'k����X|y2�)�'�nu�cmH'8ߞ�a4�F�T�V4��C���k��58P`�I�S�,�P�ȓPB�DM&y���7�B�Ĕ��Bah-R5�Y�ArJɊsM�����ȓx�5����#p쬠�D�)�j���^)]�D��
$� ��4,̤Q֎=�ȓYK��I)�N~��/
;2�8��ȓ0%v��e�R�?���ㄟ+�P]��bF�qW傭vݴ!�7č?$&%��A{4\q��ڻO�Rp)�g�i�����&>|��G C��(�,�W|�a�ȓ%䵱Q=	
�(DoAC����,�\S�OtL�i��Ė����E���Â@�=~�Ad&Ȇk"X}&� F{��t鉑65�)KVi�S�aAEH�4Bh`����?)�Ʃ�?9��?a��z��y� ���c"�[����aΖ4A����"O0(�ee��BE�$ K.D?P�2"O�Y���όD8��(C��m͚8�w"O�8��$�s�Z���ٻ��`Rb"O~-2�(�9�yDC� @w� "O�;�o̗���jC@�nfV�b��'fў�|B�'Em���獜�$�ԮE7�d��۟L����->�m�I^~*���0�~��tH��!N<1�#���̙�ȓd:p�d���x��l�sx(���̚��T�QD!�� �wԎ}��:�¡:�FI�.�q$�� o=�<�ȓIٮ��	������ȓ�|���X�B?�d؆�HhĦ���_y"�|�����`E2�΅V�h�)�IEojC�I5��Jb/<;�CC�NP��C�ɫR�p�!%��!M�<��o`�~C�=���1�a�d��8�q�ZA$C�ɷ&�d�Hq��c��qCG�4<� C�I�I�Wj~$�`�զ�),�C�I�+�ƌ;a�
Ib<H��;Tm�C��o沠 ��!��[tc��2rXC�6󰐳v�Փs���颊�&�|C�I�'�@x�B��5��9���Z�d�B�I�v��D���h.ɣ%�6VoxB�I�*"D1��K�6�$I�P&�)AjhB�	�L�(����ò`����2�3~=tC�I��T�囅P����a��0~~B��j3���^yƤZ���$���	�'QR��&d�"�X�q,��2YD=y�'-�F�W%0���D(�}��:�'��J�
�1��QtKތ]>�R�'}�ะ�\�m�^a�3�K:�(	�'`<,y��I5xC(��"OH-r:X���'Y�M벥и�j�$�ҨV�NI0�'p6�(��PKd PC& H�z	�'�� I(Q����kw)? l@+�'>�Tac��*|P|��3)�5DX0���'�T�2�hުb|�&��H�>1��'f$��ӎU�%B"T�F���BF��'x}��ʷS��|k]�;I\��'g"1�G-�:\���O H
�'����E��?Va��S=,�L��	�'v6DIS���
�� ����(zc	�'||d�2�նh��k�L͏!����	�'�>�pk�K����Hgc��
�'����6�J�j�r�A�!�3�T	
�'�ıa3F�9�:9ZS:3~4[�'��r���|�bZ��	�|��'��2!��J��B�Ë�{s� ��'^d�H��ě0�hܪ���y��!��'���aD���,U���j�.} �'SX\ad&P4&�3��F�eن`�
�'�B(Ѵ��� ����7iA[N m�
�'���1a���E�>a�g��" dLe�
�'$ą�/��S�B�"7�pL��yr�ґe1dCC�.r�Х$A��y�L\�e!
�	\88���E�ϛ�y�aY��(U�Wa�:Aq0��@Ŕ�y�,�X�P�����8�x5	ѪK	�y���Q( ��Uj
���I����y��S[�2b�&`�T�4	
��y�%*y��s"Z�E�N�D%@��y҉ �����Q?=��Q"5����y�CN:n|	�eĭ!�P$Y��2�y
� &����Wj
����D�VQ	�"O��*�ˆhU^����	uO�<��"O�Y��(� `�U�h��04����"O��j$愗q�`9��V�(2�1�"O����/�0{Q�<��!`�����"O�S�/�%�Q	���l��"Ox�`�I�����JPs{�ݓ&"O6}c�oE�rDxr�߾}�&��"O�4��*�{��e�S(;�jP5"O�d� .�@�Bi选�.y�|��"O%��Ts��=���6Yv���"OrAEA�P�m�V�@�9rr�T"OjQxfLލ� �%�N�sbD� �"O>��	�8��H�������d"O���w�B�Č�D`��.ы"OR} �ڽV� ��O8-V�K�"O��T�<;Բ���dG�"O؈�cI^CZByJP$��b�@*#"O��a�ŋ<Vjz��Py|$pG"OR��u X�8}�Y�Ո�b����"O i��)�����IAF�R�j�"O>-�$��?6����Ɂ�g�BУ�"O��4� ?W�a�.w}lY
"O()�'ՎW��۶L�Rcp�е"OFmr�@F.ST���e�%U�|��"O���(W锨Ie��R�N��"O䌚�o^#��(*�㚜z�L9!"OD��D�P�V��%J�MR/�ޙ3"Ov��f�Ƽ4,��3��I���"O���SK�,F�!����g�
�YU"O���؋8��\A����5WrM#�"Oj���P;i HPJ7 .̥�6"O�y;��<e^���"��QT� �"OZ�8���W��\)ЎN,xP"O��rbo6wL�x���ҩ�0�Q�"O�tbV��^�f�Pc���f�J�XS"O
}3sNG�j������\���c�"O�ڱ�N	&i�4��U�{ҁʢ"O�����7N�v1�\�US�x�"Ox]P��H!7����:<�#�"O`Y�R�S�isz��υ���2�"OrdK`P2k�(8���q���r�"O@�+�hͳT�ik�.N����"O�A�pjԁc��k1̘�|x0���"O8-��
�p�0�j)0`�4r"O2mxRc�:#��QهG�+?a+�"O���K&\�8ڷՁ_#6�0B"O��6
�pP�E�L��Ho"O������MtVM����}��	�"O`���D�$��EF	�.p�@�"O&�h=ˈ�b%`G�
jH4%"O�� ��9\��If�Q1��P"O,4K�j�$�x|ӆ�,qE2hi�"Oj�0�����h}�"FS9���e"O.����ħO�B�����/}zr�"Ot�ȧ�F,^G���FA�-�e"O,ܑVI��F���zL�	�  AA"O�i��bT-8�J�ӡ�'�d�t"OV�+Ю�wZJ%P�i��M&�Hp"O���F����TbU.h��%"OFTb$</���a�F8R�
���"Of��Q1�Ȫ��3K��ҧ"O�	a��ф6Q�i�5)�8���"O^�BuC2'5llfW1H��s"O� Ԡ���ښE����N�0-&�"OTШ��#ZP�UB�ͪ 1�w"O(�{���t���'K�"�5;r"O̡��bG�d2�A
�9J��,:"O��z��0
����aJ�6&讌R�"O:��ӇE,ۣ"��p��\��"O��[�$l5FTPtc�g�¸;�"O(� ��h�Upb�[cz�j�"O,�¦�G�v�fx��YFDX "O�9b��\* X�F���T�H�"O�Diu�B�s �!�"�f��r"O�eH2l�*oY0]���QkP�j�"Of���PV�� �-vSX{t"O�%j�JI�Y.D��b_m6p9�d"O��BB�2[q�}�!��sDP!"O
�#NO���@Ѱ��9"���"O���m��3i0���E�� ,��"O���
�d��M��%W
�h�aD"ON(�RNV	H�ޙ�v�7�8�"Op0!��39�]P�D�*;�	XQ"Oll��ДvAf��A�G��Y�"O��e- /K�蚀���u�d�%"O�-�W!�z#�d�p�g!��\�z��m�2���l��&�!�D�p�j�C3K�-8�ޕ"!C�4�!���HN����`�;N�ީ��o2u!��̓7:ъ4	���
����A�*�!�$�f�ص@C� �phj�(�n�!��L6�J4��:&�]��]o�!�D��-1���2`�y���9E˿xt!�ą�QB��S�����`Q� *�!��Y#r��i��A
2�����ϔl!�$��D	Z��s.џ|�&�S�d��Bf!�ǭ\bb ����'t$���X$i�!��#sXm��)M�$"��d�� &!�V�]=�ēV�M�?"����
!�X-B��{E"͞���4	T�!��U�`�J�fű]8l�i�)�!��[Ha�@�T:b�Z����l�!���,\�p �U=1zX��B�;!��%��9į�Y@�c�C�;,!�M97Z�(8��4  �6��=%!��ώsed�*e�́{�@�QA`��J�!�$Y	q�� �9����G�ӥj!�ĝ�&�Z9�� ?Z�$�s�mO�!�d�� T�PiҧI�|��U��d�!�	�#lz$"5$�W||{g��6�!��Ds�D�3յ{X�h𗂄0$�!���.#>��"��BPG8��0�U3�!�$	�U�����(,4� ��\�m�!�Ւ}��Q�I�7l&̈�7�
6/!���)LBUǭX�/-�x�GG�c0!�DH��p�a��˛���V��f~!��׃�>ԣ�nD>@��vN!��G,C6�(�'K9O��D�P	!��D&RE����&�p�Y��T�i!�d�|A��5fI�1��ɐf��d�!���k}���b�/W��}�Ԏ�'=��Dy��'�������+5�mȱȕ[�ޱX	�'(��2O}��3V�_�S�4<3	�'��X�RS)B*E(1(Ԡ d�Y{�'aXp �Mܬ�a��A/0N9�
�'J�MD�X>_C�T�H4߶ Q�'00��f��0/�d���R���#���>ʓ��� `��B��)^�̴`���e4(�P�"Oڡ��ҁ[��l��²��X�pGyBj&�')K� q'Z�S��ŌLcH���(���jR)�sT��9"�A�4��4�ȓ�0qi�#�`S��[��*T�ȓ_�����DRTFX��{��pD{��'Tt�8Wl�6�X[p`F/�4��'�݁Ҍ�}��������?��*�QS�B��S͚�끠շ)st��'�ў"|*R��$���I�2@� �'��t�<�hʧb�H���?H�4[��px�Ex��� ���eϕ'e�E(e�x�#A
E^�A+�N�G�J�b�;�C䉎׊|���S�:S�k$ɖAS�#=Y��T?]Q�д=�vq��+^�/��Z@;D�x`��G�U�nآ���4.Q���E-c�b���S�L<q��!��h��,�>�li�,ȓ\L���	B}�IRrd��e�K���<�!
�3�yH��L�:���.�v}���\���O��~�Պ��A�d!�&�ܺL4�5��J�\�<1�
W�� �J��uB�D�2�U}��|B�*�g}"��,���z���j���i�>�yc�%xpI�F�6.X�D�'�M�	�'(���v��+�<oܭ|����"O&�2ǂѰg��bP�21{�I)�"O���v䓰i/\0dV2�,�h��I~�Ie��x�-�4���J�H��V���>XRC�	>;�� �d�A�'�0�	s��h��� 3m˄[ �� �'��0S�'Q��:A
��HҎ��RQ`}P�`�p�����>���9����#Lq����g�q�{�^�L�Po��9tH��P� B�΀�sY
=��I}�'�"����޷j�:53g��G�����>�#}�!�K&xpj�:��$4��0�JY��B8����eH8+A Ɇ�8�ژ�E��,��4����O=���U���0�M��a��@K���6�!�Q�r22͒ �ޅ4�Z�b��E��p�Ն�ɛNf����e����ِ�+7�C�	2poH���9q��uS҈3Z�yE{��9O�9����7:&`�n"c!����l7D��ڶE�b�:�
Q��XLn�lt�@���2Y5��9gG� |��y�ȅ6�
���<�� I����RŔ-I��H���ě��B�I,_뒰X��Y\��4�fg�&p~�B��g�i�/��l���q@e$2B�I�F�qC�/1�|��%Ԑ]�b�d��P�'��:�F�9���D�v�2@"�4Z��	W�'�iD�4�	IS��AeQ8E0��,���y��'Aܖ=��@��2eg������Bܓ���m��:}��q ��2s�igѩl\��0?����r�E�#A[�2c B��)��O|�[ v��&c]��@�υ�Y����I'��d�>Y��@�@����%Y��u��o[S�'���=�'C����H�*mL9i��!,:x�=������F��w�,	 � &
��Uoݞo\�0��-�q3,��L�c��0� Ȑ�y�?��9��V�<w>I��*t@�Xu ğ]�C��4R�� -��f����wǆ7��n��hO���D3��p!�;_�x���, �V���He����CCc��^!94�%:p1�>�����W��\�+r� G[�4!�K�1��'��3�)��U;�E�`ɃV-t�I��	j�!�$�.9�v9kC�H8	%f�bUo٨m��O�D2�`�IX5��J߂?�q�M�?)��B�)� Υ�&��+��94I�@��Q��"O@�Fa]�s�X���R.��$��"OF����KȾ�+�&�"u��tӂ�'����;#�.%�|Iۦˆ�ՀǦ!D�P�c�N�j�aaP�fF����G�>a���S3|.��*�/�$Q�0I�[6�"?)���PcR�mЀb�\� ��k\H�O���D�k���h%�9zl}���C!�D�;�V�[cFm䎑y��)!�D�i��@�˅>�x���N,xQ�`���/~B���v�ĉOIjA"C��f_��P���ȟ&�0���U��9�W ���v�Y��'�!��T�l�+�(�Y��r��+��D2��z��~��S;W�n)���O!m�	�E�A�ybM�V���2�E�gG��0%���yR�6g�YF'�-,�"iS��ީ�yBI�\�P�e@5&2\��0�y�h��ٓ�K�!�XTB�ᆫ�y2(��'\���"!���dH�$���w���O���CpD�ds�8�R�5<� ��'Y��z�A�\	��cl�N� 9�{2�>\Oxc%�B�#u�9��X�7J��G
O�7�I�(<���E_-xN�D�5���a�az�D��X�B<���tE0`˃���!�U�ØmAF��oB��"�!���2y���ʊA<�y�"�J�\�!���H�h�QV6o�n�	s���8�!�$U�9��xZS'�i�8���[�(�� ��ɔ���Fk2-(s�ŏe�t#�"O�i�� �+6��Ħ�%��Q0"O
�"��+^�*$�3l���"O� ��ː< ���#e� c��S�O��j���zJ�]r�g�?6���&-d�܆�ɲA��ā�τ8�tS�G#����$l��b�8с �7�
t��!^;+�jkfm?D�lH4�3k�i��iZ�#V�Sv�>D�T��+���U��&Z7Bf=[�<D���$B�~�<�$���p�H}K� :���<9�R�x\�,�!�� S^	:�G]x�'�Q?=� �Ӑ�P:��Β+�8�{��8D�ؠA��+'
d)pҁ�Y�>@X��<���'1����&N!g�r,A׍�8'`A���:lOFm��%W�r �)�u턣UQ����
OF6��7+�"�ؒ͛�=s��e�A`�!��M��� ����7o&�"!�Y5=��x��	�)*Ƞjv�	���Ό$O�>c�����)�ӇVz<ਖoE}��a$���2��B䉺2�@�"Jj��A��M-��+cDB�S����(q��H�g@�Җ�¡nB䉢'��d+l ��"H�s�K3=4z"
O���I$l<����[-lf8��'�:Da�S��y6���}��dX�'���R�2D�p�䢖1:��1#� R��!+1򓿨�>��V�Kň}���9Ex��Z�>O>��U��8 ��*��W�*j��z��Ëp���aAÐ8�P�*���p0��O����Ԟ!�0���"�<-��m8���fh���C䴟����'	�Sj�aʄƐ*6)�tJ�Y��B�I<'V����r( �(Eo].F���$?�S�O���:�I� (� ��(��
����4"O 8�ƩU7�L�����d��8s�"Op=pvMؑ*T�-�"f%w>���"O���V���_vVy�CE�9 �M!�"O�5����V:�;����$�4�qV"O� p���l͹l��y �M9���9�"O<U�� <&t����T�j�"O������}�e§�/x��0B�"Ov ��"�.<��V�G!>qqw"O�-"��|�P�0 �2X��"ObX�2�OȒ�;����#��,�"O:�"��8D|4����3����"O}����]���"ЧM�+�bғ"OZ	���ο~�J)pW���.��"O�0�d��W���rC��rx^��v"Oƨ�g�/,C����薓-Z��I�"O�\y�YmT B�	fQ��÷"O���j��8c( Bvd��q+R4rP"O(J�`����碚�U����"O��pSƊ7L���V;N��5�@"O8u�g��KΝ#",�:��3"O��-9O|L�qIC�R��]���yi�	���cQ>=�HXs")N��y҉��2̌�ό2�� �'���y�HܶK�̸#"O�-���kG��y�䎐o����6독 �R4� c?�y���-w`�J�[�Dը�E� �y"�#-�vE���*u������y���1�z���Je�2 �qʄ;�yR^�d2��p�T�VѪ�Dd�0�y�M�����+�%�A���y�h�%�����Y� �¡���R��y2H���SRbj��Ɵ��y�i	������J:�P��EV��yRj��h4<������p3 �5�y����F�`u�4�	���F���yR� �,N�4o
��H�/���0?��$�e�X��E	y�����a�	��,N�<N���8\��>:KP5�g��p�<���4� ���*�@�RӉm�<c��1E�h š�&Dʀ͢��Jj�<�t.�%0P~=��#(��E"ǆ�k�<�A.�f@�cBã>��k#�MH�<�0�٬���.ܳ>���I�b�<9��1BN��$�J�T��	���U�<i�� +���6��`�cT)e�<���I�d$I�h�I���02�Uf�<Q�X�,����'�(C�� �(P~�<A�	��J�Tn��+�)�m�t�<Yh�	[����%!�~�h�Bw�<9��\�;������X'��͒R�Pr�<��"k�H��ЭV�w��i��Zi�<�����@��%���=cX����VM�<9��Y4�I	c��X�\@�q�<I"���Fqaa��8� ���Vj�<ѡ3`5�T��__7���u&`�<qg�*Z	��"i�_7��S-�^�<!Ǎ��9טqh M��4S�g�Z�<a�jJ�:�V�§H�Xj|hH�kZW�<٧c�L���*�r6�-BL�<I�j� a&)�o{�4�D�a�<�C	��h�c�� o��`ƨu�<i�� U
h�[Q�L�h#D��1C
l�<�wƗ,�P���L���j�Ai�<yg�MH���	ط=����f�<Q�eڢ7���h�D��%ǖ��%(\a�<q��{�y1�$Z�@Z�zrC�k�<q%K�2|ؤp��&}��!�c�<iЮ3E$Q�q�*E�
yh��RE�<� J�uHb"�Q�ti�:+���"O��Q6��uN{&�%�M[�"On��!T.L���#5΃vz�т�"O����9c@	����'r�pz�"OL��B�G$<���#E�vǶ�ku"O��`�a��3�$yb�J���Y"O<)�)"uHvEbG(Z�v���"O�z�˙2��c��?,�Nm3c"O�4�RO�.Z���D�Xξ��"O�%h��ϴ[5��	��ɷ�B��"O�$�Aи?J,p�m̞m�F"O`X��D��'���5+�,~�J@�c"O�h1�DҚu���%�14�H���"Op�C"�ϗT�
���f�D���� "O8�ZN5��� ��Ir�"O~�;ꙻZ/���K6��Q'"O��07⎞U$=k�ˑ�k/F�c"O�� �B�:d�p���@(��'�\�a���8�Go�?w_�uzd�ӹ~d���-(D�����QP�<�0ҕ:���7L5�I�h��{����:�	@ /)n
���M2C�I�V=���*�7<`���D�@�1u�QܓU'�>�!�&t:�#Ǿ��K¡=`����ȓ�L9�-��Fiԙs�n�U�o��D��I��'H���ĎJN��W`�]#��(�<�����<�#��4f�*���»-#jXң �`�<1`��NZL�[����blF�
F�P����ׁ ��y9�A��6ml ����!KТ���xc	������%S+�~�N��w�@��h��D�;�z���K�7��i���:C!��B�&Y#e
R."����,N�_�!�ƳHu���N�	Ǥ�*"J� (!�ÁV*�Ȳ������jjqI	�'��Qc2(Ǖ��EVe�:]��A!�';��3l�	J:.�B�QWx��B�'s��XtdJ��#���v)��'�c�AK�O���8�Ǣ's����'���`$�L�\�N�0�lƦ68",*E)�G ���I�{��H�T�6\��`��,H{,���1n�>d��3}bBM�U�T��T��9������y2i'L�*$K�B.��� �~@�!X��$!��E	P�~�e/�JG����tiIȭq
bT`V���q6��ȓL�E(�gM w�T �a�>,�$]��'��<y�E:�䫒����9O�Tx�
�R�wG����ę�02��q�E �\��� �V��D�}0t͢c)G+:���hY�bX�#V�>�x��+O~ �%��[��p��4mbH�)��3>�
�� 	u��"=9E�75.μf��[	Ri���~2�k�Nx ���V)�@I80��Q�$K����i+�H̇�Iæ��&a�]j"萦O�G�h���,�8h�����h*���%�yh/6pL��#���Id˟)_�!"�K���BB��$MR�+vɔ;)\�܃g<d��%P�b�@��1T��D�A����(oV�0ż���ϣ}���  "U�Kz)��-@8�@��L�62�3(��ez���tG�A=�L�B��0��ּi2 թ��O����Ro���q	�E�N�1R4F��1��pS�X�+��Fy"MP/B��FA�4�����*)��ɑ���AQ��e^<PdF��\�Ⱥ��� "dl �e�A��xzǧ�4��(x�.��Q	 x����CA���'��.D�(҇�|���O:�n�G�oZ=�
�CD�ڧ7�(�`�����DQ�i��H�L<��~���"�F�T��LЗ#�>橙(+plt��H�}9VЙ����?��Q��T�ǃ��4��w(D�`�bBUkr��%oX� #�3�Ȁ�+>���Q*|V�\��i2B��a�:a%F
%�~U��X�=�JiC���]t�X�4�?�'ۨn��\-6\0���dTa�\H�ф�}�F��DM��w�'���z�	[�+✂q��
(:�4�O�����J�bΨ����7�Xk�
�A�"@�F�9G��yi���6k�d<%��I<7Ɛ��֊�;qQ���	��LL���)j���7e�̟$��̅hچ6�v�,��D������r-�П�CЉ�$��@��j�)f�)Z�7O�
rAƪ�ēO���0F��+�PH��M��\��,�v�I�`1��	�k��鳕��l����=�g�? "��"�A97FҨ��O�lh�@�x���%�1O��q��;��=�|�xdk��q�vM��G��7㦘�s���F��I<=��y���|�;n�ִ���W�R'�1�3"ڻ�Px��6��h*A�\	I&������D>>I�qn��Ɲ��	dR}@
Z�aC�|X%�2;���$��j��ٓ�$����;t�5�& ��/&8Y���R
�'_��D'˥u�8��'�[-d��Y�L<ѣϔ6X�>)�N>�~*� Q.�
L���b���ʧ%�i�<��CT�P �s�
�Kj݋b+Թy=qO�M�5�<�3}roF� Fꍣ!dO�x*�Q��R�ybK��P�F7y�L�3�"�/�y���^�p�����kt����AW8�y����8ۖ�!ŌX;aMZX�G�&�y��2}�����3����ƌ��y�� n����0�5��$�a)�yRF4Rr��B��˾-H����y���t'ް93�K�=�L�p���y
S���0��"%�4���F-�y��@, C
��Y"lR� d �-�yR��.YSL�����,P�hRAmM �yB�,=�0��#�M� ��%pāٔ�y2�M24%n��k�I��]4�M)�yH�g�}a��X8�� �$���I�r�����(pF�E� �(c��8�I�9O!�D0��HJ���[Z`$c�H� `2��Ob,C��!b01�1Of��g@$8MP���gA�ȫ��')b�t��A��;v��i<�����xU�t�aR@�(�Р��bުn����e����Ox�r�^�|���;J|�"�ٴ%1y�G�n�x�#l�A�<��H�+��=�V��qn�ReMQEy�`�����G�W��S�O����a+U!M�D���ĳ#��e�ǓU�<} 2e>͎��O�gt�P�lݞjF����I�<͘(�GH
�� ~�)��NQ�3�	6~�h��@�S�~\rdHI�hv�;�ဴhPM����oѭr��K|2�m� \�����2N'��@�'�.Kx����S����"9NV}�a���/u �H�f�M���r�i�b'	1c20p�OL^e����+s.��O�Ll��0�v����b�r��c5�OT] ��&n�7�>��y��Έ=��;BF��t�$�Ӡi*�<��<���'v[��� �>᥎΃z|��ƻ%.��#�u�'��!��ʶ���Ђ�9�v�����"?�1z'�¨;tzDZ��_I���8ⓟ���C>���GB�o�h��U�	�6.��S�g�����$��/\&���Ś6^�hQ���K�d�
�&r<�:1��I����.��N�6z��h�'�
9��g[j�'��Y��J�a~~�y�K��^�]3��� �|IF�V5�0��U�P���6�:��uZ��y7o�#��D�"�N�DBZ�E!?���,�4�
�J+}J~B�]�[����#�J�>Ԍ� �f
M&�	�_�Dع5ER�n�R�!�)��܎�;��	�:S\��g�.�L�E����I��<II��@�d�z�'V;����ņ'�h�AT*Ǩq��d9u��!C��l3�ݗ-1̉`4��m�b��,�O�m���!.�b�Ѯ�F���$�	4�0��n��(1��/\H؈x�@�!-�j�!��� N��M|�Y	h���"���`i��`�''�i"�I���B��I^FF�}���_J~�]���A�t�y!���}$���D�4?<���Z�=8��'�����DZ� $،�"Lސ
@s.O�X�.K3L285�9�'u���I��O�}�,�:��I%��}�&UJ�`᧍�5g��1N�jx�Y����+)@X��F\�N3�]�5�� �Τz�R���i֟x@��8y����.;�6�]�R @�")�d˟%eAx��)�)p�챰��R��p>��ެO2�Up��^��cb%5�Fa��R�\�`�'`��)V���(��G��,��=����jR�]�P��k�>��:��Otj!�B/�h���4��#[�z�H�������:`h@�C9����ՙ?�0MY0)����E��O�(c(ʫ
��q�5���	�t�����Ʀ1��>E���"4$�K͸a��]���8]q�(RS�B B�Ĭ[F�4B�$��������.և ��,��뚭7�z��I>��6�~��� ����5�p��Q�4� �+�.m��7O+Lo�t���i�!���sp�ā>=��Å�u^�O����NK���<�H�|xb>%�,^�f4	sg�.Ahhz�'D�0����V	���l��t�*qED[��I���)�p�R��O?�I*U�vP��7Q����%~�i���� h���;ɢD���/)��P)wY��X6E�a'zAɖ�'��0�RQd����P�*��4��QTi���~:.Ł�εd��Z�h��&��d�ȓB�Y��`"+�J��D�
�50Pd�ȓd���,�?}vD��p����2��x���/u�����M�}��-D�����F�\T$�Z:sa���/9�T�a.Ĵ9ӌXwE������/fI���(;��@�D1d{���a1R�K�ñS�} t�h� �ȓ ��� "�E��M �@''H��ȓr����4Cܻj$V�j��$L�p�ȓ8��ѥ�יn��Jr���x��]��J[��5��{�2X��i�.�a�ȓ*���0n҄KM^�$��~-�Іȓ&��Cä`p�QӨ��QP����䃗��l#���G��� �� ����("E�K�vm�����k�轅�ܮK�ΎJ� � D�V�[`������
�Ké[58���H0>e�̇ȓ��!�
�%`�i���&w�ܩ��*�`���*K�@�8��# I�6�z(��V]��¥�׵z�@��GְM�N���>ނ��o��I�G�)_-$��4D��r�� ���؄�ߊ�<`�'?D�غ�	S�j�!M��8�d�9D�|	rnU�Z�x0��n���1��7D�`(��'O�}�J%,qp�4D�,��!S�w2����'�,�BQ�7D���b��B�
Ѯ�#��B�2D���Ɛ�v���CH
s�́�f,$D�0�����l떼���r�X �.D�$Z��]�'~�4Yrᏽ�z�8S�8D�,��T:��Eq��Lz�:� '#2D�`He�B8tL`]`d�
;p�xp-0D����\��� ���Nx��@��*D�X���ߙQ/& ���2}d��'�$D���d�1	�cFM��d~�}SC#D�d"�G��\h��iQ�W�\<�f�#D�l�1Nɛ�8Dh0�O3"�
$�'!D����푕m��@��C&���;�!D��)��I ��B%@�;w�5�A?D������U4�Ņ�Z2�I��<D�$c0�X /Ц��.ņ5ԞY�Q,8D�|��J_���*׫��Z�`7D�"�×''�4u&ث"t��"��2D�lcB�D���������s�3D�T�@���i�	P�N�&	�3�1D���G�H�c��Gj�PI4�A�-D��ҳ��I�,Y�g$
���[%'D��a�d	�^+��R�&y�C��6D��IL0H$~ �t����a�$4D�|��FC6Br�i�c��6X(���ti8D�����ψ�D�"m�,9S�9�3�:D���0I�ny�Ú�K4��c�9D�p�4LN�(�:����_�o��pR!C6D��;s@\�=��QEʖٶă�+D�ܙ�
Q l����O�^�cf4D�P�t�Z@;��E^�#��)6D�Dȅ�K�qW����0��x��4D�ı2�v��9�b!S��p�&3D�$*d/�$D �%-$�� �1D�L�匈hT���K��P�h,D��z��.!FL�F��5f�x�!D�� &���ǆjS �˶��<�n�  "Ob��u�Z �L���?�6	�R"OX���aZ2vn��Sn�@Ű`q�"O
�!Q[�l_�t�Ƌ�ȔP��"O�XP�_�i�%#�EW��ya�"Ol�ѫd�@-p��ϙY�0���"OB\[�O䬐խ1k�ҩ��"O�R <{ذxYt�A���U"O����/�"(Cd��a�G<I"�1CU"Od�C�I�F�H��B(Y�ƍ��'D�×m�<>� ��LS�F��Db%D�(�֫���X�82"L+k9�3E$D�4��*�*Ar(;#�K ���k�O?D�0����[To��3�b�J�#/D��_{ 8��D��<��-D�,r�KY34��ʣ#
��͙��<D�h�0�B�BO𤫖��2V�~� G;D��p^�`P�"�퍼8tQg9D�0{��;X�v�Iq�I�xѳ�7D�xB�AуP�L��U�D&} ���#6D���Ԩ۱�����c��Dh�Ӈ6D��Ӥ��eF�PX�}�&�ʗ!��)y��h
�"��!(�!nB�!��{�pR�L�M�X� .J*s�!�F�w���=4��i�C팈"!�V#:4HQ�[��T�U��4[!�D\�)����M_���e��h!�	�sX��2��ǻ#H�]�ЌN!��]��.��+
 4JQ��F�g�!���3ld8Ec֯]2V=d�ZTk�0�!�0z�8 W�ǀ(%z�E��<H�!�DO�4Z���e'����Y%IS};!��ƪ>��R�K�2k(H��Ñ#I!�@aL@ �D� �z���P!�\#����\�d��ٛw�!�J�B�8�"�O�HOޭ �k�!�$T�$�9�!�J3s60R�MU�_�!�D��:�n�a��44<AA�N�+V�!򄚟4�Ј�V�M7�ˁ�,c�!���;^P9v�<XH���4:
!�$";<��}�Eb$0$Oz�(\�	f�BD��3����/��͒�*ѬуV:BP��,V:=Ȫ��I�u��8q�l��>^��
� \
B,� �dn+�!��1�Ɖ��F>9�l��ǔ� �d��6���K�6?���H?�#��+ox�*���ݰyc@9+�!�?/�B�	2%�t��σ��C ���qBc�	g��HQʁ����`�'Ur��'���"#���y'�_5�������&$�����>��K�M��MAĄ/��!�ªR(p�E�%U�|IZ���n#��D�V��9Q!��p�Q� �S��+���yp%��,ި���<���iw�LQ������mV��?�n�e�@9_S�ICvC_:".�)��-֒_���e���0>8uC2� ��W)z�T�8��E. �|�cGd6Eh��ԍv�P��ޟd�q�'���hŮ��k��4j��MCd% �	��-Ar��q�<�Ԉ�x�}�Q�2 �Fh���M+N��I9��Z���S�[��%�^?!�DW
+���9�w�e��m(?��90�'����P��!𝃃�׺@,uyRƝ��� �F��~��	Qw��6-@&<���I#&�ъ2�85<�i�BF-v��a��U�H�*@��(O�"䎇.p��1E S�`�@j�?�k��D>�-��h"wϾ��gթt���D���4bߓ[p�Eq�*�<%�%�f(��.и%����皳m�v�P��Yr�I�?aԻi� Ĩ��Z}q����Kaj8�%:n����at��xQș�(��4%%�6;[�@������RnO�WQPi�s%g~��hq8O�[E�շ9]�,̻g���<WUru�,9�|���v���˥"لFq�De;^;�k!g�$�z�+&a��UZ ���4�?���z�*�v�
�u�|�?A���E0d�1�L��q��@~�'[�1J�%�#3�qC� �<u�'7Z�� ����ͦ(�ű2�]�@u��0p�84�L�"�Q(w���DT�K
������D�3F���y��X?Z�H���8bV�Q��ן��:�⅁g(��2�=����8_ b�"RD+X4���`���yҏ�?�>�i��)i	�9��J���Q��!�fZ���1��>t�	��k�n	@@�H�[4�C�ɭ<G0�9𩂺 �"@q�@D�����#D���	�%v����|bOh�h9!���q�l��Sm �Px����uѮ퉀M	�O`� ��#�X���[�ޜ؇��)\��h1�Sa���!xD��E�M'�����ܰ���S6t&`+L����5����X�!�d�$2��� E�E2�6�p�)�6FƉ'�}���S?l�ɧ�O�h��`
UF�����:&�
�'�5;����>��t����9���0B�0`�z��OV��@gQ#ڑ�Q@Q�~^�{6"O�{���qb �Q�σud��ʳ"O���f%�L�����<[t�R0"O�$Zb�Ԏ����0g�+W(�3�"O�M��؃]:V ���� �d ,�y���7J�"��D%�U,ҽ0�͛�y��Ȯ\k2��!B�._s��h���y���e[��J�Y��飇D�y��M
'9ؤkAi@D��(��ʫ�yR���F�d̜L�4�����yR�]>	�����8ARȊ���<�y�[�5��,{0�^<k4ʙ���I�yr'�+M9��y�Oזcj�c#ȵ�y�ON;-��ԡ���]�~ Qb�
��I3���P���	(|�� G�5c�t��Ƥ�4R�!�+HSȀ��Ww�re�X)=�r�O�R5"(?�1�1O H�p'�S
1Hw�5,�}�s�'\� g�<C,Jv	
�L�PDȮT���Sa��`؟l��#	�Xe��S��>I��)ؗ�/��%<n�!��OE� ��U�3�'(���`��U�"{����"O�d��l�Zm�!	%Ʋ�V\��C��C�(��֓>E�dD��v����eN0ލ�g�nX���ի3h�O�x����	2��� �� Q��!���&��;=���Vl�3�3X($�Ck�l)��`7�I�N`,�"�\�Ñ�JM��PF�Di�-���M܇U]�*��Ύ	O������o��u���(k�줋��Q�]���!�� 1@�↨.?q3׋e����vWD��451�;'��HT��-Z-�0�VJ��Y��i#��0D�Y![M,����Y�V���r�Xoߌ=�%���Su��!(U��'>>}���)(�ǐ<jȲ4���6���H$n��D��=�ʟZ��tM�m?�yJsh� ji��%�DI"o}����d��j�̄�SOwC-"��*Y�F˓{�p<3tY�-�j�
���ɵE�Ȕ���@$�{�F_/ܶi��̩��O
�P� ]�Fi�O@a(���`��[���Nh9�2�T���$��E��4� ��
4n���Pw�E�y�^8���$k�I�!�� �K�H��S��*׬!c�Qu�)�g,נr�N�Ѣ�ʿ6�^L8u�'�<:Rm���-@#âێ*�*)RM@#��l=�T�Ԩ�D+��O�n�ƨ�N���$�yo�8rWΒ�&\`	iB�Y�����$�"8~+��@k�C9H��!C�2uG�A���Qg�&��'>I pe�:�>����¸�v4�a�*��\�n����� �ɟ8�A�l�*3�nԑ� ��!��#�$
�#�+1���JMж�3W�^�㒌Pʕ|^��-y��3�;-P�qE�D�4M!ФmCud)UF�:,�$��4�@<�JنE�~P
c��xUj)K �1+��e�'V�I�e� ���ϸ'�~���+Q��2��˱bX��X��t�r�H�E�t,��i�ҦaإpW N�vQ �G�L��0?a�F˿9��[A'�seIk��NO�'���2��	4�?	rD��VH����V�Ze��E>D�@QÉq<�����͚h��5�6�??��a�7��K�M&}��i�*DX��D�	��T����Ub�!�D�6y}��"���1�샧M< h'�蓇�>q��'�l�eΞ�ư���
.^R*�X	��� �<`�*LO�n�xU+�?r����"O�	"�h�T�h�0IT4��k�"O4<9�n�'�ФE�:��e"O"�`�3�Ȉ�s�Խ-^r=��y��w�H])G��&�N�A���3�yr��9W`��<�����Fِ�y�U�>NP��Cڑ	`f�1���y���&L��� 
Z�{�p-X�$2�y�)�q�-@d	'q�<�!k��y��8іL��ʬj�j�� ���Py�l��`��eívFe����[�<���hYp��Q��.jpt����_�<QRC��e�"ɒ&%ϨaRD�j�#RX�<��jڲ(}Z�)�_/D0�*4��@�<�ï�+%�\|рO����-k�Vp�ȓ!^\��wa�o�`�0+¯i��y��{D�*���3r�9p5JR!	*��ȓ@��-���F0�Ha�c�:�v���b �� g��I��\�f�K=rM e�ȓ&@$�VN�;F��p"A�]�U�ȓ#|�Hr� ����P�+�\y�)�ȓ��X�#W?!���ĆC%c܅�ȓVLx��'d?���%W�4�\���%֜��%�F�}�X ��Z��: �ȓq6X豄���;��r�.�U�zQ�ȓn(@�)�|�CW��!�� ��o@��8E��/tyX��|�����\���`U��IՀ!��B�t^ZL�ȓc��Q:e���$�������C�I�p�d(���vÂ8 �ɐZ�lB�I�D����Qb��L�H��$���9 C�ɵcʴC5
2?~< ��X�M]�B�	,F3��Q͍!#L�� ^C�G��	3Ռ˶j�M���5��B�	;���0p����0�
C�i�HB�I_������[����*ߑr�C�I($!H0��"7ӄxtΜ3�C䉹w���"�O��J(X�-�~C�� p/�1
���p��5�
�qHC�ɛ����f-w~�Ń&�ǰb�&����2@��� ��OFz�ceHݍvq>��!B�t-!�d[�:tЅ�T �oz�p;��Ɣt!�����dQg�bvH!��j_�^!��/! p@
�HQ-`jx��(�q�!�K�Xo�Y�ؚmhr�[Շ�=�!�$��DŴ a�&�GV���GGÙQ�!�D��x�a�!��#S�0��7�H�/!�(\��-�-�� ۣ(J:?%!�$�x�&p30-Sz^E�ΗK~!�$������U�e��VH�G�a{��!�;y��1��# �qJ�>+"��ɉ�P��Sl# ��-�"t�����K��5R���&"��ذ㞢2��.P�uPFjد�Q�b�ߟ����=9��/��U8��%dnh<1�A	"��������b>eq�J7j7�<05���QJ*}rJ��,���=�g�I�7�!��%IZ��8�.�z��I��,M�?E��dWbF�南�^�T��f��jIt�80F$�)��M	��K䩋<6��a�I�u���҄��6��O���'o9� @�,�v���TH�]e�=o���'B{B�"��h�p֝�(丄A���\�P�!�S8/��݂R���U��)՛�?�B	8�l��!ɬ/(�;W	B:.��A1�ƫ8�����<�bh���a������Դ���� D$l��c��6x�=p��O%*qǞ������'G� �Ò'�)����d&U��x�<�N�d�L�':2����O�"��i!N�Ь �����̬�ڴC�<i*�)]�4ҧȟ� ���a��O��a���}D�`w�ٝLD��'�J���s�p�B����w���r�'� �b��0h*H�P�`Y�`f��`�'+�lI�*Z�k��p�lZ$�qC�'�!�	:8�a�J��,��'>&刕*�3:X!s�ώ�%`(i�'�N�R�'E�D���8�ե�h�!�'��!K��W\*J�x�c��| ��'�0���W�����A|J�`[�'J<ꃏ�4��!�&,ɍt{(x��'�����gL�j�t�Pa�>MZ���'
���E�0K���gHח;�@��	�'9>[$�!�z,��hߏ0d�@	�'�28���'aK.�k ��Tu�9
�'!�h��Rk�0`0ϝ=E���	�'�\�:P�*�<�����l)�\��'D���ց�Mk��0�R�1˰x��'�|hb�o5��� � v�Ј��'�~�{'�q �@�cK1D���	�'��S�hA�-�"E���3>Ǽ���'�j�r�"���\�4�ې4m$y;�'��(�� I3z~����h̜{bN	��'�^1��@���>� ��ȏoM�,��'͢�� 	]������C��m���'��ĚQ�ӷD�LШ��'���'_<Y����A�p��A+C/@��'��l�7Dޞ�\�Sѣ^7/ҭ��']t�O�$M�|ʑ̄!�b���'�V�Z'�4u��q`%��rTr	�'�4��?LN�uY���^8�
�'k:�	&����uc׮�r��(	�'d��t�]
S8@3wF��5�n8h�'���tK�=f���Ӿ&�`���'6J��&��C�Б{����*��[�'~Ő�i�<���Ҕ�ܼӸ�Z�'+�٫`�ih�ys��:V�ȓ}��;W��L��E�#�E>�T���m�|8a���
�>�(����챇ȓ.����u)�E�Z<�rLZ2V)���Jm$�˧�	?�|y �Էz���ȓ<n6�Q�&�q��x r��6���ȓ
��X��DeS�]���T0!�����&� O_������+�ܥ��]�4@���6N.t�P��%zl��@�Hp��	 Lb�sd�E�w� ��(`�hBW��X�p%�b�إPx�U�ȓd���[ЁՄO��MSŅ�f ���8�\�����J�[pC�: �х�3�j5Q@�0jj�z1/]�k_&t�ȓfK��h�)I�|�
���.[�xЄȓ(ZF�2��KrмR"��6���~����h�{i�z�L��Ψ�ȓV{<���(,ty�q �ȓT`b��\���#`n�=Z��U��e�B\q�� �Z�ⱦ�5h+���ȓ{�Ʊ���f;�@�� 
��ȓc0$m�[Z<^�[�M�h�@��8��k���10�v)�w�� m�X�ȓ_���O�4��4GԒC��ȓ�z��PI<Q�t���p�ȓ*�m�鏲o���B���K�Pu�ȓIݼ��cl��Oe&aQ�Pr���ȓ0\�� @�Јdf�0�VΒ\xԆȓq)>)� �V<j�L)��(�5?h8��S�? �9�T�j�L�6�\t�:"O�	hޖ#��$95�9�Qq"O��(ek��3��@qmGf���"OL,B`C��l��$j�-��l��|1!"O"�!�(F�(/��xЁ�aۄ}��"O����DJ�THF�G1��]`"OԐjf�Y7:6j��g�g�и�"O`}���#��kUǈ,�\�#�"O�h�KܹD-������9~��T�"O��1R$�!_K ��"1��"O&=+L����d{bVb�,	�"O���완!'�y�#��%-(Juj�"OV�8�� O�x�H�@1W�|s%"O�x�%�&���I4��-E(R�d"Oj�8f.�(�VM�Y���3"O��X�L�1V�ք2�	ul.�"O�� 0�X�\�}RP'�����N�!�dA�~�1�I�c�|��u�E�X�!��4'P�9�ʜ�J�{�E_*Y!�D�������-��hjB.!���/�t�Brk�R �9'���FN!�$����áF���l�,۬a�!�Q9��U[d!C#�V�Q�=�!�DO�zC���FX�"2����D &B�!�DX�:�rl1�� ".(Z'iU�*�!��ӷ^/��K��3"
� �7r�!��{�� ���$ �����p�!�D��o�=��Ef')�f��O!�N
J�jTҷ��(ƀ1���&d3!�d]�
�%�w��((�sfeݼ]�!�DШ(�2�v�4	�!8F���"�!�đ9e�@���/bɺ�h@��!�$���P$P�g�f�*a�F�?5b!�ҡ.8pԺ�l�R����p��gF!�D�+�zٸ���:&��d `A-+!���EI�u7DN#��i�O",!�$� Rl� K�|w���
Y�K!���3����ǼcH�w��2�!��J��s楉,~oD�G)��f�!��*ArnXSpc�5~^��e\d!���="�����ޖ
�h� &I-oG!��ƚQ�}�$@��d�$� �P��ȓH�NM�rH= �
�F�ĂQ'�A��{8����m:=\���b� �tć�D9��4�G����=Ay�d��P����OE�51� RN'H �ȓ>�^��p+�'Y�!� ��"j�9�ȓ㺭�`,��b4���P�I�ح��=��I�NDa�yä��	HX=���42$_6#��@�� ��(�ȓQ��ċϖD�
4H!O۸Q�2��\!0�ɅO|��3A�ϝ!w��ȓ�Ɛ2��#鞜;g�E�2��0�ȓe>�UcuHA]���sҗ'�DЅȓ7ꔜ��	�dI�1���͐�lD�ȓwc2�����-){��D�<�X<�ȓ9��S1��V	���6L�VZ�	��,�����!XH��"/�:�6ȅȓ~]T����B�0cj� ����Nk�8��KP�2�V!k�ʚ3^���ȓS��9��M1$6b@�b��H}�H��o.^�8�I,]��s�&�����ȓ_��ӈ_�`��rV��P�t��+`P�ۦi�%d$��r��W�A'�Q��S�? ���N��6`��C��9]O��[�"O��: %��,�?Zq	V"O*uB)�#cy`P�ci���ӗ"OJ�ҷ��+���c��8���"O�v//R6��'Ƚ�� �"Ob���D]	Ն�!'L�^vLI#"OJ��%E�2+@1.�+����y*7����ŏ%���y�͘��y�#[2i)7K��R4r�*�(ɚ�y�v�(Q!V�^	?h�3�gƛ�yZ��	�BA13��rC���)
�'���d�8X�
��g�B�4�H�j	�'H`ěT�A�N�,@�7���,��'��|2p�C���H`��( �)��'�`�{��~f�A�ϸ O�y�'yT�k(����0P�f������'���q�U�6T0�@�{=�,A�'PL ���>hX��v�������'��T�Є�Z���;��C2QxHq
�'�-��i���}"��ǈ~!P0	�'F������Bl��#�?rԵ��'.����#r�E'2s�a(
�'�^���n�?"����$%$0S�'��%��E^����B	��'���C�Z���UO^���c	�'B~�)j�V:`{��P;�x��'l���W�!RPkO6G���'����(�<q��� ��QHL��'�&�b�%\�x�*�it�x	�'2R X�J@'�h0AB�:{�h��'����ga��s���x���#yM±��'��02���qc�	X���?T�'(<ЁgØ$�x�@��n��#�'i�����-�!��J�5D�X�Qbϗc��Q��2W�pa�4D���׃̓���g"��P��e�0D�)W/V�H��1��O6j�[@d/D��A'M���lb(O%a��i���/D��'T�q��yH����i�-D������t�쀑 �'i���6�7D�T����y��+1aZ\ИSr 5D���a�So4q��WD����*4D�H�d�X�Z�<��%,T(��	�dG$D����#	��X�0��.,�`#$D��B%h�P��L�$ʷ�!D���9_�Z�Pd��<Tu�m2�� D��k��.D~A�Bn�8�c9D�Q��� ���s�Ю`5�ZA�*D�x1F�>"�Y[Q`�	-8d��";D� �$�ͺYC*�蔧��ỳ.D��z�ȁ$fhD�A�c|�F�7D�\�������勝Y���3��5D�A0�D�9�"(+@�E(hf��`C�3D�@Z��Z"?�d����?afYY��-D�$��d�.I����4:�Har��,D��8��V첀�`��u��p�w�?D�Ȉ�Q�T����nJ� �wI3D����O���z�� ;���Ң�$D��9���[s�ÕOT"<�l��#c6D�T���Z�U��
�E��N.���7D�,¤��
"sl@�`�S�S��*:D�(B���7�Zhh¥,/���@/9D��� f4aJ�ӕa�z�ڑiB�6D�`륦ռ�6��m^�3U�9є3D�� ZX�A$Z�TA�!Ş"�^��"Obu��`�+3n���	�=/�|�*�"O�)����&��4��fR�\Pm�"OL�aF�[_�(5�@ ��V�\�"O���3�߷-���R"�E�b����"O�D�    ��   �  c  
  a  U+  �6  �B  �M  �Y  Je  �p  �{  ��  ��  5�  6�  ۧ  %�  ��  ��  8�  ��  �  ��  #�  w�  ��  �  R�  ��  �    � � $ 4" , [3 F:  C �I QQ �W �] �b  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z��Yb�с�5|O�"EG�;֊�R"�O�~Q:�F�'VP���Œ�'蠢DO�	J厈���4D��@Q�Ђ:�|@��Tfs���(D��`D�J�=Np�A��׭7����Q,%D��z�oV5H�r��.Q�����$D��p�L���Uk��B�����F"D����`���2����{�& �E�<D��PL��j���H�G��:f;$��S���T����t��n�����^�D��� �F��9^	�F�=[`�͆�Im�)H''��*-���t�S:E��ن�	�H���
�e�pڶ�3<K�̆�;�؄�c��v�`����֭wXވ���t~� �6XvD�e �8�HP��E��y�D�9;�px����|	J�fƈ�HO����"��aA'ݥtǽ�!:w*7�!�p��`�:�4E�*ɠ����Gu��E{���\�B��8�d
5s�.,�(�8zE!�$ǈ`VaR�킍wz�q2T�
�-!��QI�V}z�f=n�����,a~�V���J^X+ָ{�儏v(p�R��5D��)��?1� Zg#��o�2���(D�p���%HА�(��� ��Ȁ�"lO4➼�eO\;xz\���%$��1
!D�p
`f	 CHA�0���-ƵH%�<D�pZ��CX��wf �B4F<D�<��"J!���#����.�aDO-D�qU"Ո0<�i3K��$��X��0D�� @��#aǵu0�IՊ[�zl�s�Of�'�6�NQ���I�k0L�F�_3��݃�!X8Xaa}��i�d	x�Ա$o��\�j�� ��Vhm&H�(#<E��4'u��D��* a�<x��S�RU���Ms�B��D��<3�Z�V��#YRy��,�OҜh�k��Z�:i��m�N[S�'����O�4�V� �ń���/( H�"O:mKw����b�GF	ڷ"O$��$L�GE��;A��t�V"O�p�##�&6yK83�� ��ݬ�~��'�̀�=E��' �R�yB&Ӽ!s�$�DH�:�y�DކE����B�
}x�^��'J�{�A�^]~|ӄԅ<(��B'	I�yb�����1q�E�-����ȗ.|�B≎;삔t�+I'�h[���8E��B� :��)2��a�,���	�3HԮB�	�s@�@���d�j����P�B�	Z�
�"�7d|�b�KD]�B�ɝIhZ�q����*�y�JO�jC�I�ynD4�7@ɫ	�8��B->0�>��}b�f�qiA�'-P�i&�G�C�z���DI^�<�sh�E$4���(�D7�)Z`?1�]��m�|yr�S�\Ӥ�#��J>�+"
E�V��C�I7B�F�v/��q̚���2j��tE{J?�����3>k-���I���A(6D��u@I(S"���n�#^�u#S�y���>9��'��	�E�l���4�\#�4����'|��R��-Mu��;�!a*�e��'��D��EY�3�F�4���Q'��+��D �S��퇺V�N�ر�	�<y�0��+Z�yAP2ez�=Hb��##�А
��~�ў"~�Tӂ���`�[�$��iD�Rԭ��a�$��΅�U)�%a��.P�l��\�.��hǾ �8:�a_� �����B̓'@�1�F�z�BQ�M����ȓVN^��ؽ���Qp§ ���n� �EE�0��Qtn
&V��_�<�ەi�#G�L�f�I� 	�ȓ=�r!f�,`� �2�1�t��=fPH�bd�3!��,�
!H����l����JƑ@��\��OC�f�4 �� ��Q���
� ����[�����-��l@�m�!_~����$��2M�ȓ^`�ђ �8z�Qb�1n�Z���.�C���J�~4aC.$@�ȓp�D�z��

�V1�S)־�ȓM��%L��	B�� �
S"���|/���%�3-Yt��N׋]�����.�ѕ�Q�F&~���̈,M�]��t�����^�U�FӅ.��S2���i�{�J���?N䉇�����fE�,Mq�(�,D��Ѕȓ	� �� ɠ�:��Ơ��j��-�ȓjJ&]!g�B�x���blV�k��U�ȓ{R"q�N�!r$0QR�&z�}��T��a��W(x�]���"^���(�ڢFC=�8@��j�g�pQ��G�"�BG"f��lљr�4�ȓ�M�P/W>o���x5�ŕ"��
�''�#r?B��K���a���
�'\�P��mɀ)%�;���
�'�����X�v\�[4	=oH`	�'�����U(���i˺	0����'4Z��[1����p �YL����� E�����Y0�)�J�iw�!q"O�q�ʇ�gs܁�˓�*I!�"O�Y�6���I	@�R�`M�"O���# R	
R��0K�B���t"O:�!ck�a��L`Æ�'��xi��'��'&B�'�R�'r2�'��'u��W)��C�5@��J�L��'��'*��'���'�r�'���'���L�1d���XC��qՊH���'���'���':��'�"�'p��']�e���nA(\�ƪ�u��Y��'�"�'���'|R�'���'��'�����M�	`���r��k��y:E�'��'j��'���''��'��'h���@0
����V�V)qJ ��']R�'���'m��'rr�'z��'MD� �^9D��8R/�)'M���g�'4B�'�B�'|b�'"�'���'Q�����Eg�j��4@�(��4�'���'���'u��'$��'���'�ژ��-���J�_���ze�'��'���'M��'J��'��'�\];���u�eナ�'-����c�'u"�'�B�'/B�'�r�'�2�'��+I��``I ��7Ȱ5�#�'}��'��'��':b�'R�'�ʱSA��,ol`�2oH�=�����'�'�r�'Y��'zr�'�B�'�J�-9	⬱B�W&S���A��'�B�'�'K�'���w�
���O��[�G���"�|�2�:��ay��'~�)�3?A��i�BU�e���Z0d8!`%֘ Bh��������?��<A�M�	S^`aCN�#s�RI ��/�?��:u�\��4��dz>���'���5!]ZA�0��~���mS�`bc���	ly�
ff�ZF��Jo����&44,�ߴ>�*e�<I���'i����!T�(�+6��q�'�4s�n���Ox�g}���M��3W�V<O
P��dٳ2w6�a ��>
t�-�5O�牛�?�@':��|"�Ql�,°a��A���Bq� 5t0͓��$%��F˦M���7�I�(��9��������ߦP����?�X�������������glJ�
0�H\�Ũ'ʗ"h���l���^"#Exb>m���'Dx��	�Lxf��+P�N��dr�h\�$�Jt�'L�	��"~Γ��Gf��F.�9��f?i:�ϓjR��偫��$�ϦQ�?ͧL�|hh��v��$��hb�FAϓ�?i���?ib+���Ms�OB��+���L�f��:�=R�Uj�dKFUO���|z���?���?����t�'��)O�X���g ��(Ob�o�t�,�	������?}$?岁	G#��`d��]iH���KĖ���C���ݴ:������O;�$/C�Ty�����Ս@�`Ԡ�ݗ|\�h �ih�˓2�u 󊦟�&���'�]���ȈW���c��:��8�'���'�"���\���41
<��_P��n��m��Qt�!+=��������x}��p����IԦ�"Ջ�9؜sW�Lu�Ը��L&�oN~r㊍3�N���6��O�fT�E:<�$�N3�N]�����y�'�b�'��'V"�i\�j�0���I;t�:��b����O��d�즵`�gl>��I+�M�����6�3Q�\0j�.�n�:WN�$�� ڴz뛦�O�Θ��i��d�OB�w���V�`��$�[8��$��lP�`h>LH�'��'�	����t�	�]�D��P�f
!���<I��	ȟ��'�6-t#H�D�O����|���}*dt:u��'eP$`t.~~RĮ>ac�i��6-�J�)Rт	����kb�]�g��,#To�-<a/�?�MqX��xm��9�D�&6"q���39��°		9.���O
���O���ɷ<���ij���lѧ�r�˱��?��Hq!
.,�b�'�7M1�����$v�~��'-�Q����Ty�T�@����ܴ<,D8޴���H'D�U��O/�	�R�>���LD6I�бʗ�M��	Oy��'B�'}��'|bW>���h�=0�j��-j�~��o���M�kM��?����?1K~���w$�Ҥ	Ͽ5�`R�H?��<YFfoӴ�mڳ��S�''���ش�yR��7�!be+6Np��p���ybA�V�@q�����d�O��әBIL����i�������)K����O�$ca �O��m؛��?|��'��*
>?�J��>dд���ٯ��S�������ē��9k�4�?�)O���F�GuhB�f��,v~ũ�:O��D�&?h�0���LF����?�y��'��9���v���kD�)��Q��6Z�8�	����	ݟ\��J�O���<Ab�41f���i�w�����$l�I�c�<���iM�O��3BS,�����a:��3�N�&5�dxӔ m���MK�`ͅ�M;�'%�wk4��'-oj��BՏir��H�ќt�NԛH>i/O$�d�O �$�OT���O��$_�NB��!L@��t;dϲ<q �iA�M1K����'*��֟���'���e��N�Z��'c�@D�i��>Q��i��6��Oܝ&>��Sߟ�PcŅ�l,���B�zv�IR.Z�<Ϝ4�V ?y�d�z��������dV3oU�HH�`�	x�ܩ:LT��$�$�OPa{��G>�4������q�;k�Ԍ���4�d���D	�0pG)�!'`�Q�9A���X}��'���}��2�iϜw�v���.� �81G�Z,8�P7�u�h�	3�a 5֟���*�{�? ���gcD6I�HHI�I�*!�F7OD�$�O��d�O����OZ���$'�n��D�%-�(�x�M |m,�u��Oj��Ʀ�@B�MBy�'��'k�TF�U���Ր2���B�a���7��6�q��	M{(,6�}�$x�fK�0���ô"�x�&��&B!���)M�M�0T��N��h�Kj��?9��?���t�}��ÍEO�����A��q���?)-OX�n�%�<5��蟸�I�?���-$p�1���a{5��62�����D�'aҴi�D6*�S7Z^�@��Ɋg��4�CDN�;��`���Մd��y�&?�f��h(#0�m��`��?ͻ��ו�-Z@OC$|��x�&��Ɵ����8�I͟L{� p>-�	iy�p�]x�o2>�,�qT�I]����h��t�ܟ�����\�������[��a�f� ���-�b�EIXw2li�`m�Ϧmsܴ6I2D;�4��ě�&�&� ����SR�h8B�cY���Fȁ-iLz=)�4����O���O|�D�O����|ڠ�ܲ��圳M>I�sh��9�X��ݴW��e`!O��?Q��2U��?�'�?�;.	4������sw��	F��(�:aⰰi�26]ݦ����O�`�v�i���}��2Um@�EP�$�v�����,X�H�h�d�Z�c��R���۟��wC:x���,��.�qA����|��럄�I]y�x���d�O����O�p���:����-@�K^��f�O�˓�?��O��$h�lody��Ee�(Q��5��y"�����j���� G�F_����u�FM��P���'^�\��I�,�\],B��D�tg˝�?���?����?�����'\2�ޱc~���"H�#����@�+CREz�� �g��O���O���<��Cs�Jw j�y2BU	To���aT?ٴ �v�mӪ}�d����ӟ�j����Ĥ�nzd8�Յ�Npt���bJ�r�\$�'9<7�<ͧ�?���?���?yW"Q(�u�Ҋ�|��\i�m�����榡��ʃ���̟|�OB�'���CDX�A����!��)�1@X�X�4	w���~�
����	�B����T����Kw��j'�tSAaA��u�@��\�ƣ-2R��Py��{�P�1q�Q�K�;r���`,Ǖ9=�H���?i���?�$�VA�6�)(O4�o�:f���S�J"�"q�߻#�6�a$@M�:|�ɽ�M[����O`��'���i#.7m�	���fY�=��[G��#5E� q��r�t���$xćH����-?���n'֍Z�LNbi~%t��l@�D�O����O���O��+��H7�LI+bOF&<��geahj|	E�H����Or�l�j�'���'=�	�8[��*	U���h&�@ `� <�۴��$|�!Dx��R�6m"?)���:�����ag�`Dj�?��m���O�q.OT�n�Uyʟ���A�3�g2�!�B��"<Y2�i��Q���'v��'m�2Q����D!��At��<���G��̟(�I���S�D@��u��,ФE=
gIG�Z�lG)����<ͧk8��	O�	(��%�V��=hv�iѕ��q*N�������ß��)�SGy��c���1�πF+���WKR�b}��"������O� nZt��L���Ŧ1�!d�!u������C���"��?YߴI��t��4���к�����$v�˓l�,hs J�mi,�y��g�P�͓����O��d�Oj��O����|�q����`)Z�(Ҟ_U�h!!��a��䐧E���'/ғ��'�7=�8<B��M1K�P)�� E�m�ń��=!�����|�����5�Ɍ�MØ'2�LS�1��`�㚘z�Y�'���J�˟��1�|�Z����ß<qKS�t��	!F��L�:���NX�� �	ԟ���^y��{���Rf�O����O����P�?BP��%�/�X�>�I ���O���1�d�hb؝��-��M��a㎛ a���O.�Z��+(�&	@Vj�<���O���DX)�?�4�67��2�"�4/���C�/ɟ�?���?i��?Q��I�O���#X�$F��b��d˗��Ot4lڥ\�����ܟ� �4���y���x����ABJ�,
V<{5���~��i?�6m�ʦ��p �榑��?A��ޫLD��)	<
쀡�t��'
����R#$p���J>�.O����O|�d�O��$�O���BO�r���:��]�tw:�Iϼ<��i�ɲ��'�2�'t��yR$w���GF�¤������(��Fl�F�&���?����6}d��.��v	��D�	;��b��H��59(O�HH�W+�~�|�[���q��3`,��'��cC∫�ƚ�4�	����I��Siy,~�zةq��O��%l@�$d:�+N1�Q2T��O�Ql�F�5����M�Q�i�7��=�] �%ڪ$Gة �G�a�B��q��"$J5�?e&?��]91@Z�jr��
�]g((X�9O"���O��$�O����OL�?�fG߆|��+7�� YVџT���@��4<$Χ�?��iS�'��pf�0�`4�dC�1*d��.��Ʀݚٴ���NB��M{�'�b�N47�Y�����pȬ[3,ڣ��5M�T?�I>�.Op���O\���O)�GV��L�@lD�\�eJ�O*���<�i��*�'	��'�Sy��j!E��|��`�7� ���	)�M�5�i�XO���$2˔?_qR��W&�f�x��H�H��eF�o�b�'C�d�q?AN>9��t}���e�m\`	���`<A��i�l���k7%k �1�a�>IV���J=���'��7(�I���d�O��� ̝4h<!c&���BA��O��m����m�w~�N4��%����� �Z�H�SsRl�@��h �(9O�ʓ�?Y���?Q���?��򉃳t�JH+%�7"@%�q�L(�f�oZ��f�'j���ܦ�ݛX�N�SQh�1����E	ן+L=�	Ɵ�K<ͧ�?��'�>aK�4�ykT�$T(�X��%��	�����yb��ue�l������O��D�^�ʹ�RE
��r<���%hn2�$�O����Oj�C؛�hq�Iş8�ֆ�0/.t�RR�//\حhDO�'�$c�O���O|}%��Z�LL9s	BY0�Q�N
a�e�������jBwQR��<��'_nJ�I��b�
0Pj�K3�ϛN'n��A� ß<�����I��PE�T�'�0a�&��W�H��I�0f�|��'�7ٺt6�����4� ����A��I��	��U�77O����O��l��A�~ o�g~Ҥ��u���'`�	!cJ<)��	)�KN4��TIL>!-O���O����O,�d�O�!�ǋ.c<A�T�Aú�Rb��<�e�i@�X��'��'��:��C��):�q���p�4�82��B}��'6��&�󩘖b�qs�B�f_Z�:��č_�����v�z`�'%n�S��_l?�H>�*O����%[z@Q���	N�.�:`m�O`�$�O����O�ɱ<'�i��p���'�!�L3C�5�%�
C[|�W�'��6�(�	���DP����4�6�	g
U
�d� E����S���o?&�ZѳiU�D�OX���MS���tP���S��	��L�O����C��N��y���I��	����p��W��,`2�AB�ǙGO�`�E���$�OJ�m��I)\��֟�*�4��l��y�C@��aj�m!e@�R�&��V�xB�`�ʽnz>H! �=�'݈���]8� �YƍE3?�I3b�S0�ҥ�������OZ�D�O��DT"��Tif�ށ@��4�U�Rl���O�˓A��fL�d{�'��Z>�X�N�Y�9�Ck	j�!5�"?)eX��+�4Tꛖ�$�4�l�I�-�<A��2�VɁ��>}1<�A䎞�z(r7��xy��O�����[I�	Z��ހ.��[S+C�n9+��?!(OB��<���i��t��ʊ!Q��A���T�;w)���r�'k�6�;�I����즍�b�P*D��`�pX��DG��M���i�豓Ѽix�d�O^%bA�۬��dR���G�8�* [�$�=3@T��kx�T�'�B�'�B�'�r�' ��`���	I��bR�K�>� ش��A��?9����'�?aw��yעܦ(B<X�F�P4"�$�� J-���c�.&���ZM���Ӥ�	�F�3��N �G�)+��?�P(�$�OܓO�ʓ�?q���\-�q횁0P�vH�Wv�m@��?����?�-O��o�
pM*%�	��.U����j�#��)Dǆ�a� ��?�&^������!L<�Ѐ˶p��@���ϙ�V ��~~b�	�3�e�i�����	��'�W�+�|��M�b�N4��%�S���'��'�����3
�� ��H��)g|�#7��ȟ,�ٴyt��?A��i�"�|�w�.l�C����q�̍�b�YC�'26��ܦz�4�\:�4�y��'��p)f��tv��t�d�e�C>v��R�H߅�����OV��OX�d�O��\�x]�m���
����d!���P����)$w���,&?�I&c��ч!Fu�؁9"��~hn�I(O���h�"�'����lJD�>h'.� �D=r�FA�u�ԸO�6m�wyb
Қ��m�����D�>D��$-l��ى��?B�|���O��$�O*�4���C@�V�ǷS��/�p�r���<U�N�bd�Ü�y�&s���0�-OJ��c�:�lڥw0�x�fO~�\܁��P5k�BC������'0����M�J~��� ���V�R�&&+2
]R����?9��?���?!���OW��Iq��*a�NŃe���.�A�'#R�'�6�B"�)�OxnZ~�I�:oJ�(M��)K:P`�����]�I��@�i>�r�Ϧ-�'>��(e�_���J�哶M�-�#��������D\�'��i>1��ݟ��I�7�칷'	$Z5�*���40��Ο�'�R6ǇI~���O����|j��'�i��L|�9�V(K~���<!��?H>�O���J ^����ѓ72hx���>
�`	H0.Z	F��i>ћ��'/E'��0��6IK �J��L����!�ٟx�I������擖6���Iy��f�R�aU#���p�0#�&dQ�
I	@4f�$�O��l�Ɵ$�����>Is�i���F�7f�d�q���l�p8��yӦ�$�� *�6�q����]ȚA�Q�O���`ƹ�U�\:Rq���d�.�]͓����O����O����OJ�$�|:3��%P��LbD#'�2��$��DIN�ݘ��'��O����'C�$p���_2L��1��	B�a�kS
�5o�> o��M����4��	�OV4k�y���ɹ���P��#7�F9)0"Φ*��<bR��O�lI>i*O�	�O��/�P�)N6"]��zV�W<2����O����O0�LV�&�G.Q��'^��>=�8�3�M=y� }A�'޺��O4A�'�2�'�Ot� ���m�9Y"잩��cԝ��s�@-eK�lZ���'Vɜ�	���q�h�_�*��V�4P��r���ҟ��	�����4E���'ߔq����8ެ�U������1�'9�7��"?�����Oz�oZM�Ӽ�Ҡg\�}3�D
�VA"}8q���<q��?y�is��¸iH�I+ �>�  ӟ� f�U���
[�ѴK�D�gA?��<����?���?���?��hʨW1d�QD����Â�H��d�ܦ�h�ן�	��$?�	�{�Y'�+/y��T&���PX��O�}m���?I<�|:�!�1�`dD l�ޡ	&IͦFv���	���d�$(���E�8�O
ʓe�J=�U��W�<h9�O�&G���{���?q���?y��|�,O�=o�	��=�I*~���çV�P �l�wT6V���	�M��b�>����?Yտi�t�z��N�T� �ň�;�؄�E!� tϛ����cSf�����:����p�wIßWR⽐��ҍ1l4Ɋ�'��'�"�'2�'���ec��������m��@Q*�Ѐ	�<������^���d�'��6� ��_+xb��
�C�<8�<}�2n4:���&���ڴћ�O����b�i��I�V"���"斃2��]�7C�VeX͘�#�;-f��+���<����?!���?Dm£S�6��ro��F�����R��?�����$�צ̀����<����O����&j�
�(���6���Oj��'K46-��IkN<�O� ��c���*�n�{cC�9�Y���<v=� �i;���| k���$����cܤ��W�P��L�3�ޟ,��˟�����b>��' �7��
t7*�HA�g~��Qu�N:�\��e#�Ob��Ԧ��?m�>q��i���{w��/ ��Pˉ�$bEz�l~�HTm�z2�x���U� ����?��'�T�ץ�>b�ظ�0$�*��8Q�'Y�Пl�����I��p��d�$@ڶ����|a�� ��8-�7�K�A��d�O�D!�9O�nz�� [=9B��	ufް	2�RAɁ�?��4�?�O�O���Q�i�dO0_*S#�R+Ov��� �<^���1>�f���D��Ol��|��%�:x�w'�3*�j���y
����?���?�.O�m5H����I����ɇOk�
?���r�ݑ}U�����j}B�'���=�d7+�J�*r��9"����f��X��OF��j�vRQ��`�<	�':'��$�?���X7F���a�5�\��,@)�?���?�����l"!L�j�fa�a$�%�l[�ԟ��46N�����?�%�i��O��<k"����I�>h|� (Ѭ|��$��1����M�r����M��Ox�jh���&�W�05v-sC��s�e[��ȾN,�O�˓�?����?i���?��
�j\0�T�*��\��;s����DO��y���xy��'P��|ꂈ]�o)td UC�K�t���oy��'|J~�5 �"G��r�*�b\40`�4+�T��q�;���ş'в$�e�^�O��Z�f$ӃbJ `���W�js�a����?I��?���|�*O��n����'	ش#�/�]cࡑ���:�0��'�7-,�ɼ��$C������M��#]B�&T
�΁Z���5K ���4��$�.�.����UD���0�.�:��1�`H ~5�A����-e��O����O����O���-�ӰxV2�R�h]90_N���җD�f��韸��4�M[����|*��A��|��Ǯn;�8:���1a��XHtKB�	xO�im��MK�'+���4�yr�'z�`�B�ʌ�↏+R ��sG��I�('�'�ɟ���۟h���
���ŋ�=R9�׎N3B����̟��'�d7틵[n���O��d�|�ˇw��т�'s����~~�+�>���i^27�y�)���˃X�D���M43�̚�k��)?=��NV��M#�R��t���,�d���RX�U��$�Q1
�"sK����OV���O��i�<a�i3�Q���v�~Y�PJ��T�qH>{�"�'L�6�9��+����OD '�ߜg��M2�a�)-��S�b�O��mZ���oZQ~b/Χ}�"���W�	S--�tI���?O�2T0t@4 �$�<���?���?i��?�+�캥
���|I�����mE�a��Z�	ß<$?��I9�Mϻ��,�5m$l�����z{J�� �'қ�-��O����O��$�6�i:���`8�(�B-)f2�8�������&):غ�1騒O<��|���}?:�a���V)��AUc�q_�����?����?�/O` m�&#�P�������iʸ�wF�n���Ɗ&͆��?��Q�������L<a�j���m��,Y��S����-)p�U�[���|�P�O�h��krݙ'�҄)D	�qhZs��+��?��?9����zxx�¸U��;nr���`�������юH�y���M���3�?���?����4��N��Q�&<��V	p�n �1H8w��d^Ӧ8�4�?�B �<�M��'U�X	A�ơ���r���t��}�P�T�M�;��%ƙ|]��S��P����,���@��� ��� �.�.NCǃnyR�n�䨠�Ǽ<����3_�?���.��ZV�9:~�,ڲȕ63o�$�)O��m�>�MK���h�R���*
�5��EI<yP�!��fP��3����#�� ��f@�	Cy��)�^ų/�:��ƭ^M�R�'��'w�*�O�剿�M;ū�&�?9�\r��0a�EVb!�ٓ���?���?).OL��>?���MK�uPځ;'���-&�5�ė7p|@� \��M3�'���hȦ��S���������u�Cm�0Ud�ɧ������O��D�O����O��D3���T�,��@�t3@�'V:���j���I<�M#g@'��dR���Iyy�	DFN��e� �D
G���rT��A�4:��O�\	%�iU���0� �E���].%�LP�B�<Dݞ�)����?���$���<ͧ�?Q���?�2�Z���(���Ew衸!L�'�?Q���?I�h��tZ�tHB�?���?ֳ��4��-������fS���r#)��${}r�'�BJ?�4���d�� 4����o>Z	i���0&_��+@��/_�6MMyy�O�z����Z���hh�
KV�:p둿A��#��?)���?��S�'��D��y����H@bրX�m�8ڇ���]������ߴ��'��#���m0a�� �h���b�.P�6ML��dMRܦ��'g��#��T:+OXu#�l�AE�K�)�a��D��9O���?����?A��?I����i)pG��]F8�SB\3��mrFzӐaX���O@���O�����I���3lJ�xz�nB7:�ި+�� kU���4?n��.��Ɏ�o�6�k���G���.����W@&GnH4�d�d���'	~1�� �Ĭ<)��?�q�%SkX�%��L�&F�B��?���?	����$Zצ��$�\qy��';��څb�$��PC��H�L�X����a}�@q�p5m����a7�1���9�B�&V�_�|�'v���G�<Nw��D1����~2�'��"Td�"�a+�ߞ?���a�'R��'"�'��>U�ɎnK�8��EqOF���b�$��	��M+eh�(�?���l����4��i�E�8t��c�I\� 1�Z0=O^��O��n�[�T�m�<���t�"�HR��t��A��7;5ąR�#
M��R%�D.�䓈�4�~�d�O��d�O��d�vC������/!=��
��{T�q��vW��'�B���'Sޔ1B�ҏOv@9E�7 ��A�˩>���y�x��tb�<����M�`��@��i�b���*F)�]����'��%���'��I{3L06�ꉹ$��[߆�{
�f����/'��FS�b�p��Fe^�Ie.�9l�b�<�p��OJ���O�lnZ%._D-R�a�3miu���!>4*숡�\Ҧ�'������V:L~��;q,V%��E���id%�l ̓��?�� �P݌�9s��(�	2"�!�?��?�#�i6��������%���W#�"	���Rk��^e�<3s��?������l��i9�6�#?���\&􌀹�Ɏ?9���b� ES�չRO���$�T�'7�O����J7�1X1�\��RY���!�MóF��?����?-�v�ZQH�D�]�6`���P,h`�����O�)l��M�ґxʟLl׃�n�,�X +� ݖX�eĆ=���z��%����I�f?L>	4n��	�~x�f�4'�5��U<qU�iw\� �WT���R��.�^�q����b�'��7�6�	���}�j��q��%֦��F��E?�8����ڴjL�%�ش���ДL֔���O%�ɖK��Dd�w ���P�@�o���qy��',hHCW�őA{��Z�/N�ƨH6@`ӊ�� ��O����OJ�?=����!hC�����Ř"<��E.^���Kt�4�%�b>��D�Φ��>��Ö���"b�Q��K�73d�Γn��Xp1����$���''��'��DO�"A�T=��,)�Fu�5�'�r�'��X��cڴ3�FL,O�$"�e��)M(><��n��54⟤9�O@`nZ*�M����d��&V)1���8-�(�n:?\��O΍c�I8�j�;�����S�q>��ܟ�i�E�@�6��G�P�r�(D
џT���X��ş�E�D�'�.)��D� l	�184��/����f�'fh7-�!�"�2��&�4�iSte�e���q�F���$Q�<O�|mZ��Mk��)\�Ѫ۴�����(a��IW��#π'[�0mj�\�X�
(���<ͧ�?	���?���?�t葓�(I��m�(*�>9Cb�&��dO��135�<��ȟx%?�	�R舩Bl��9-
�p�L���p�O��m�3�M+���O}�T�'�4ER�
RL�0�#�/p�3��::p= �O0�F�ȝ�?� d*��<	��V%U[ذ�c':x6,�z�� �?���?	��?�'������
�,�П KtHI,N�����r(,Ui��K��y2�w��⟄�OPnZ�M;�Q�����ΌXg��H2�K�l��+2���M;�O��л�b��d�wm�@Rq�ÛGd�yP��s�x̋�'���'�r�'q��'�p郷*"r����C�
�"��0��O����Oj�nZ:i;d��'�87M&�dB�&���F�*{�Y�n�&Zv&0'�X�I�p���C��oZ�<�����H
BWܨ=KČ�~�R����'Gt���3�䓥�$�O����O����J��pK�d8�26M�5TT��O�ʓVY�&ň.`TR�'�BX>9$�$�KEj��VXXJwC8jO�I����O���~�i>q�	�}-h��/ޏ2�`�j��I��I�w��B��*3�Lyy�O���I62��'NJE ����G��y#�%�l�4pv�'�b�'k���Ot�I��M�i���@%�iQ�hk+[�Z�J{��?�6�ih�Ob��'��7�� x�tC�OR5���z0k؈q��	��m��!�ߦ��'z�IÇ��?��X���Iq�|\�UgM�e@!�wDj���'�"�']��'"�'W�+{�ra86�R��-���kR����4��Q����?����'�?���y�nJ))2a���Ue��Y�(X32
��'ETO1�8d�o`�`�)� ��zW�@=w�P��1
� &/t��v5O
��%�W>�?I�b7���<�'�?�rE��:�$���ab�HpC�ϖ�?���?���������g/Mϟ ��ݟ B�
D�8�2U�����&��e�D
a��]��I���	<��(�вg�&pzi�h-z��!͓�?� '_@�"��4��?mzF�O��d�#^#�T	��P�i1��Ir�@)	��$�O��D�O��4�'�?i�II)h@�ͪ���j�P[ ď=�?�g�i�X�R �'��w����]!�
�`2�˔ �>�{�B�+'�牖�M��i��6M��Z6-*?�熟�rVF�H�Z�qfa��كL��J�X%$�̕'��'��'[�'�h�RY�](�!`A����)6�前�M�3�'T�LB��?��'U3�ub���?a1e�7l$�e	�m4	��0�f��ZW�I �M�s�'������O�����$\m�K�鄉9���I��� ����>��	'qLl���'��x&�h�'��:����`���l�5�BL��]���I����i>e�'��6�\1C^����GŲ�KPƃ� O��aBoRJJ����e�?��^�<��ԟ��ش`Cv�3���B������N5*8h$)�I��M��O������Ĝ�4�wR�}�6��<�)�f�t��p �'2��'xR�'KR�'�,)���J�eI`�g�U6)�P��B�O��$�O �o�{�R�'ic��|�hW�J��Yp�(M1v�ۃ�tO��l��MϧCq�](�4��$ѮW�BDõ�")$��6Łm�T�j� 4�~��|�S�h��ϟ,�I`�D����<��%��	�NZ�	[y҂f���	d��O��d�O�	��T�X�GF.n�F<���XŐ��&��s�O��D�O`�&�������dʛ�[�m"�F��6�P!���U&M�=X%�æY�-O6����~�|"��R�H��/��a'
��T�_�x��b�6(��E�3a��Q����H���aM�P^����O�lm�b�_z��2�M;�o�L�ED�<s�����)ڌs���M~Ӥ,�¬d���l�MUİ?Q�'�����R-\D�a��+J�:"͇�O� �bćO�(q A�5��Z��W'thP�b��:D��ς�[�h,�PɊ*(J��g$�8;
�l�w�	9���"bE�/vR:�cȍk��(�
�%6qhiB�5!9��X��v��S��qo�=d�\$�GA49�"e� k�Y펍�FN@�l8,�3r�U��N�1�m�3x�,�j�B>-�r����4?&� ���"L)��$�n������6ዲA��a��A�>v]@1��>7<�P'�z<�=7�N�H%��B�O<��pdj�,N
$���y���ON�d��`4�'=� ;��Dk��AzF( ��^��)شNRXy������OCB�UF��l!��Zs*�eΘ�f�"7��O����O��R�l�d}�]���	B?1W�J���������ئe'�,3�l�ħ�?���?�R�Y�ک�`�R�lxzq
�B�,]��6�'jD�a�>�-O�D&���h ���ԋojfZ6�(m�4�FT��i4/��\�'��'�bU��p�H ]���D�#��ɀc�l�&��O2��?�L>!���?y2�E��8u��!`A��h��ɷC�X�<����?!�������ΧYX�I+�F��}��(aa�A��n�{yr�'��'#b�'Ĝ �%�O�TD�H)R�2�h�B�%|�z��X�P������TyBcX�EZꧫ?Dm�<$��]�a���9���	4i���'�'7��'�������
�W�X���'��X����r�Q�x���'z[��Z !�����O��$���3��S>j;D�U��m��D%�r�	۟\�	���q�?)�O֘�i�+M���q�+K��Hڴ���Ȕya�Qmɟ��I�\�ӂ���ƪ������>�$hx%�S�V�6��v�i���'�h�ß'��'��>���@3J00qMc8��I����TL���M���?Y����P�t�'��a��a
�+������7�"@YQm|��-�QE2��F���?)0
0n��}���R�ȡaG� fٛ�'tR�'�L@@�>�+O��䤟���JO�bE� �-g2�,��%:��7�Th%��������I�*���cH�5��¦
��dj޴�?i�'�5��	gy��'Hɧ5��_,�$��ɑd8L9%M��dS���O
���OJ�D�<)��A�dR$�I��
�V��Q�ֆ�"5�U���'�"�|b�'���$c�T����&`d���J{�d�u�|��'��'��2]�q��O�.ə@�_?�h��Y����O����O|�O��x��h��,Ԭ�G.�	{`Ґb�E<,�1P���	ޟ��IHy���2�J��+)S*>�>�3��צQڶ�j����e�	G�cyB ���b�~�ֻ���)� \`�:$h������ԟ �'��p��=�I�O����Br���7a�Ј�b���z���x_�p�	���'?�i��ːJU�lA�(��!ļJ8y@�v�P˓ZTQ��i`맡?�����I�ru��;�"��XXP1C�Х'�27��<���?і������4-!6�:Պ\Lx)ʤ���%n�,w�Xy1۴�?����?��'[e����&=���u��TD�S��6��L����O�����<y��$�NP:6��<��-K����X״i���'"m���O�I�O �	%�h�c-^�bt%ҧ��	�@7�O�˓<�iq���䓔?��9�������A"�byX�!�vӔ�D �I��L���P��`M���FS�f�T4¤FD�K�MC�Y��z�ܙJ��c���IRy��'��� 6�Zg�u���G��&U"��@H�(��D�O���+�I֟p�I#%����c���hTxn�%}<��FR3@).b�p�IyB�' Ƒ�Pڟ�$����	)��9���N�|�J�i���'�Ov���O���a��G6�6��	`�@�����U��Hbcj����?-OL��Ư`���'�?	��Vf�p*�Ƕ\H.]��G�WK�����O��DHH֌�B��x�e�@��񐲧��"Oʱ�$���M[����O4m @�|���?��[��;8lN=�"�W�Y�M�K�I��,�I�J2����h2�~2��Ec_�� 7�wD(���n�Ŧ��'���*��}�"Y�O���OA��C�l}Y���4v\$x�f�Ϝ_d%l�m~���?�������4F|<���ϫ1� �@ōDy�b�oڥ�VPcݴ�?)��?��'����\cNpu[BĲg²��3gՏ#H����4O�1���?����?��'�� Zb.�29�PE���Y� ��К��ǁ�MC��?��.-�x'�x�O��O��q&�P(������V���8`�i�rR��H�GHʟ<'���IX?A�M��;�f4�?W	X0��ͦ��ɪ2T��'l�'��'3�{A��kȼ�F)�J��e�$�d��L��	ğ���ϟ,�'��Z��|�҅+4��U1���7O���O�Ĳ<!����Į�.]*� bԨzL�-ڇ�P	�M������O���O\ʓ�Bj�0��)��O\�[��c���J��!P���Iß\��Hy��'��ßt�n��*
ι�r�����KD$������O��d�O��~�x�cR?��ɒ*����ׅHmH}p�#N&Ei�$��4�?!(O0��O��d�����3}�Ï&┓�(NLGV�@ ɝ�M���?�)O��r�G�S��':��Oj����M��t�r��Uw��q��>1��?��R		�����Tg��	��lڀM��j��RŬ�?�M[(O���Dꦉ����h���?aS�O�.�4CW���ФZ�`�f�/�v�'��G��y��|b��uQt���M����䬝�盶oFY�T7M�O(�D�Of��Aj}�Y�H���I�T 0ĊU�� ����M�g��<�����.��ȟ��jQ�s*����
#U���J�R���O����O��E�_f}�V�<��{?Q�꜄}��]�$ĕ�aGȁa�mQ䦑��}y2���yʟ.���O��Ĝ<�|Q; +�<p
v]��ɐ:Q���o���4k���$�<�����Ok�D6&����F�J|��1�AU�&�'�2��'6��'u��'�rS������o��F�1ke)4a���O˓�?�.O���O`������%��(P�1�&�&K����8O�ʓ�?���?+OR�(6@��|J�$�%\}��BO1�F�� ��I�'S�L�	ڟ`�ɥgrr��%K�\ѠE�3�bYn�JuP����i@r�'���'s��`�����$�����U�"��SB+Z-Zf�oZ���'�"�'����yb�'0�$��x� �@	8���4(�ܛ��'W���%�?��)�O*�$�7@�3���r�սwD�����l}��'���'�V���'��s���'S�b|���u&�'M�<o�mnLy��ΩiQ�7�Ov���O��)�|}Zw���E��#{Zͨ�OԨ7���4�?	��y��9ϓw��s���}*���b�����D�'��A������hfi�*�M���?����rX���'��DX��@�����tp��@�@��v���y�|��	�O���dʝ�~�f��$(�H@���U�E������ ��I�X��Of��?)�O�L�����A�c��?�8���4�?A+O�X��6O���� ��ݟH�r)�-5 ek����8�K��M��H��4��P��'�R\���i���#�)3������%jN.8���c�h��&Y��<���?Y���d�s�\���� ��$Sc���B��e��Jh}�V���IQy��'\"�'��p	���;_T�u�Ԁs3/�:W�D��?����?���?�*O�DR�Έ�|R�Cڼ$�NԀu�_'�P��sk@��i�'��S�l��ɟt�	M���	�y8 �zO��@D��	G�T�n���B޴�?9��?������Ҹ��O�Zc�b�{5����m*f,i5Px�ش�?a+Oj���O�D�<(�1��F3�U�߀g:x	*�o�<�M#��?(Ođ9�[G���'���O$<�a��3n�,9Z3L�<pbY��l�>���?���(�͓��$�O���'+�Y�I�>�j��rK82�7m�<Q"�M1�v�'���'���N�>�;n���ò�>S!J� R�n���x�ɕ_���	����O8�>}:��P�hʪ�Y���|�u��~Ӷ�3M���-�	ݟp���?)��O��9��({g$�5J�0Y`��"<�H��D�i?&L����=�S�h3��ӟ36\��D"�"߽�M����?���1#��{�R�\�'��O`�s'ƞ�(1���EDE�l��)�Ծi�2U��+��a��'�?���?y'f�:{�B=I7(=��d̾-����'�F����>�*O�$�<���[b���8����h�F-Y#��Q}r-��yRZ�T�I��L�	iyB �$s�$	elr����F�ŘB.I�h�>a,OF��<i���?��.���T�����+�/ `�����<!��?���?!����E�1-�xϧ7f��@@�'�T�2� 2,�o�Ny��'�Ο��ҟ�z��a��8�9	| 9���/Q�h<��b���$�O���O��0�ּ�Z?e��9�� � jՄC.0*���dA6o�"d�t�i�2W�|�I�4�ɀ_����v��K�[�pi����cL���$͎��'�BP���� �����O~��Nŋ#bݑi��"o�����u}��'���'Dhųʟ0����+��;���Ղ��H�*���M�.O44Y�EWȦ��������?	�O뎚�T��Q�ĭ�/B��j�ៀ����'��τ�yB�'���'q��=��%��-3z,����'$��F�i�ph�3f�����O������'%��;-�����=��K���6����4|��`��?�.O��?�Ipƌ ���/k��e�P�[��� 2۴�?���?	U�\8e��oy�'c��C�3x�f�A�$� ��Qd�"CR���|�(�yʟ���O����Uڨy��8Uj�{1� Q@(m۟ B �J3���<I���$�Ok,=�i�Ѧ��A��h �#�-�	~���	؟���ߟx�	Ꞔ�':�t��(�2 �@��VS�E?*s�O&���OĒO$���O�42��T�v�y�SY4�m)�g�J�L�O��d�O�Ĩ<�U��+�	�	�z8�/�t��\�KW:z���� ��a���$��y�p��Zh*B�ο\��:���U'���'r��'��]�܈�����ħ�\D�F�{�B%sPf�	"t$��i\r�|��']���yR�>1�ґ^^<��Y�J2�hXb�����I؟$�'�R �Շ(�	�O2���IR�%3�D����|��BT�*�Ĩ$�p��蟸Q�D���$���'H�J-1V��6	����2Ryliy��� j�7M�G���'��$I;?!�G@"d�� ��&J����,ɦ�I؟�u�ߟ�'���}rW����CsI�#��(�����R'��M��?�����xr�'��,����%,����#Y(��Ox��(�%6��F�'�?yPO�uKl��c�8B� i�rb��)ћ��'R�'�b�Q�J:�	����]�z �`��P��&���%�0��>���Qa��?���?� X	?\�{��'f�@��Њ	�ݛ��'O�8�D�4��˟��'8Zc��h�	X;�x���? �-��OQ�#��Ob�$�Oʓa{n�"�Y29��`�7e��Ey���Ƌ�]!�'�2�'��'�"�'+�-�W��Sq���1�~u��+ˊ�y�P���I���ICy'�XS��R�Yz@�оp"�c%n�"SӒO"�d>���O ��*!����8<����㊪/��!�r#�}����'P2�'��]���'C߉��'n���pd�α �|ס?ހ�Ҹi��|"�'����u��>�1͛b`y�.�*�����m��ş��'Q�U�f�(�)�O�ə�'��EؠQ��)�:
�=	�i;��O��������;���?sAb�1���1��MG�P�ՠm�Jʓ>7ȼ`��i8���?i�':i�I�kE��g�+Do�m��">z�6��O.�dҾ0P�/��-�S���"�_�l�"��S�P;N7
6G�kS��oZ��I͟@�S����|��	b�=2��n�R���[���N]<a��'��)�'�?�"�ׇ� D!��°�B�I�7AN���'���'���ꦦ)�4���'O8h c�d�zdA�@ѝ�ҥi�4�?�)O�e�ЈFS��۟0�	ßl �+����	S��R����Ѩ.�M�%�\���x�OkQ�P�3%�1Tt9��D�g���0��>��
<�?q��?1��?�����d�?;�8�i	/us�U8b$D�8i9�cSs�	ޟtG{��' ^l��I��:���cG <�b�8�G<���'��'�"�'���	_A��O�|��AɅ*p"�u&Ǒ+�A��O���(ړ�?Y�-б�?釣ÃYX�TC��wu��"R�I�����ꟴ���`hU$S����	ʟ��B,Q���1��3&�pK����M������?���)��m�1��q�4mMR�p�O*">�XT�3y�J6M�O��Ģ<��ڶR*�S����	�?�Ig�<Z����C_�Q�*х���M���lR�5��On���^	��7��Q��ZF�f]���i���'��`�'���'k2�O��i�q�T��hU���L�(趭S�j�H���O�<��	
51O���y෫�(^�,u��ǟ�Z`���iM| E�'u��'4��O�B�',��]��P���������
���P��4d�N�:��O�S�O��߄մuQW�2.$�������6��O���OTM`��BB�i>)�	����F"�1d�#���v���GM����'J��y2�'��'�V|2GC�<7|��W��#T���lp����ԮH�N�f�����&���P�T�}�(Q��A�>K4���,����Dr�Yv����	�����qy��_l��(Bâ	����D�ڕ�� ��g)���O���-���O���I�I3p��f4N,5#fO5j������O��D�OT�4�
a�5:�������t�hD���&�%����ē�?�N>A��?�2�L}�,����S(.x�Uf���$�O�$�O�˓H�yJ��TF&%&��4���)�:Y�	��u�\7��O �O����O樨��đ�}��@���24�e�ݔ)����' �P�X�m���'�?���u�Q�� �0$���b��nR����x��'����O�$���Ϻ@-2��ӣK.	��7��<���M�g^�6;~����ѕ�� �� 3�T~��kQ�(>�%�F�ia��'c\�ʌ��)�2h�.x�5�F3P��#�^.��h��G�7��O����O����|�H�(���e+, �8�d��q$�q�i��-���d.�S؟���AM:/w$�4G�8!����u�&�Mk��?��a���S�D�O����^6�=צ��4/\����% $c�dCU�#��۟��	���pgi1oZ��Q�_0��m�j���M+� -���Q�$�OT�Ok�$[� ���,G5!4�8���&���S1�c���I֟���ayb��/~*��$ �u�؂ G�49ָ�7�"�D�O��d<�d�O��$�- )X�ýB)�&�8��ԫ����'���'""[�h#�OP����$,��p���kS���o2��d�O�d*�D�O�җc��I+.���
z�x�D\?O28��?9���?�)O�ԘQ��\���'.���G�(��k1��>,s���E/vӾ��<����?���;p��?��'`8&H	�+A��r&L,si�Cڴ�?������ſ�\ �O>�'��dm���7��"=V�$f;kB��?����?�efD@~RU���86:p�s$Ftb4�Ii͵�J�oGy����HԨ7��O(��O����u}Zw%�,0''¬�ҥ��#@�][hEp�4�?��[�:1̓
.�s���}*�-�=K\\�C'K�:����G*����T�K��Mc���?A��j'^�L�'��iNڝQ�ˇJ�!Ȃy���hӴ@g8OR�$�<��D�'���$��1z ��+�+���Ƅe���D�Ox�d�R�h��'1�ğ��ZZ����]PN��"h��% \�>���ZS��?1���?�g�ȦJ� �b�/����Eʵf��F�'d>i��>�)O
���<�������Qh��A^,2���E�CO}������O����O���<a�%�oն���C[���H�^�H�1a]���'�RS���	�����kL���)J�:dG�Ύ�Ь�g�$�	Ɵ�IߟX�	By���4è�.?^l�s�ٿR�}��B�4I(�6��<�����O��D�O�٠�:O`�h�F�,+JH�5K��Y��&Sj}��'UB�'��I8�d�í� �d>?���Ђ�N�$�"�`���">��n�ʟ��'�'*r'Ʃ�yrP>7-Mg��xR� z�0���`+(D��fU���)T��I�@,X�#�Tu����%z��ɬf5btH�� ��TC�I g���c J.�R���_$�˗�QV�X]���u�X�E�GȂ�_J�A���N��!��V�d�T�[䇗#8pX����.�|���A�Hܠ�#@ ˲�B�I�f�<n��d*���9�|�`��B^#'I�\��Ic�b��H'�����#����8 �7E�Q�pP�Q� 0�,YB�c��
Sd��O����Oɬ;/�<��FS���\����*y(���GI�����Θ-��x�ba����O�f�'��q� -�NRQX��Z��Hұ�/+� ���4�����9�.��3J�|�0 X��4�ݴr��B ��1W����B:����a~b,��?�'�hOR�㧣�-Q�|�q��.o@�8A"O����������,X]r��<���?і'�,�Z����,Y6�ې́�{-��6Lٙas&mʒ�'�B�'���`�a������'Mn�2ӊ��W�|er���p��+����X�Hvl>`9@9ϓ,��$�e��d0q��"Q��x�V�X?V xC�	`�+�[<VP��m~�cA��-Jq��)��̟���r�'��O�%`�,ι(Tܰ�B׸X�0hA"O���sM3%B6�{3B'N�F��e}�_�tB�	����$�O����4��Ei₄0'�mz���O����1X.j�D�O�擠 ����`)7�V�s�'82�Q�j��H|�� ��ݕs|���	Ǔa��U0���DwTu���O��I�Aj��0�#Rȴ]���'%�!���?A/O��6�� 8D��r���&�4����'|OTmˤ쑖�XJ��<5�L��eO��lڗ@@�l2�F�V'����F`R �`y¯Z B���?�(��Xy��O��� ł
Mx|��",ߝ3
i���O����;� aH cX#hX��O�a��i�#_�Ԓt��*��� C����	�V!L]�BdY H�ra�Gn��?Y8���Qp\T��I;z;����>}�K��?���h� ��&BJdf�N�GK���Ь�:)�!���(<�H�+�:f����e���axR�5ғO?��ې�~�dq R�V��.���[�����<A��ˡT<�-�I����I͟�ݓn�b����(T � �3Wy����O%�I�2DL�@�)�3�$���`:��(%$�RS�|��Hq�=3}@�!q� 1E������]��剶H\���#��E�Ä8�̡��q~R���?�'�hON%�MX�G"�x��3 1��"O>LrwD�Ce0@�F���h�F<ّ���{���?�'����u��3�2苰�D�����/��~�� 2c�'���'��y���	��d�'�"J����n$Jt�@�$_��N׹4�����Ј
�H�Dy^}�Q,�w�
)�$�� �`����`X@7iÞJ�[t+T%jx�Q�ɘğd��)� ��)��E�vo�!�$�'[��$e"O}��M0I8�r��;B^�b�dD�]�,+�i�B�'�R��`�~'V���O�t�z�B�'�m��A �'��H��|r$Q�?RB�*T�T�	Ɗ�����p<1G-]D�YR��(���9���Z,xv���S�x1��[�	���bG�T�K����D��JC�I*�@k�Iy{�����$3�2C����M�"Q+� �$m͐l����,���VW���i��'�哐88��	 /���1DG�z��M��`ӟ|R�)�	ǟ<��ԍfvE�$�����|�+�A[����L�����1��>���NA�ab`�v����'I3$�Hf��s��$��ؠT���'�P1i�ɘ��O=�QT�(���#�B��U����'��@%����C��y���Ó�X��Wm���v(�x��릋��M��?��S!T�q怯�?���?��Ӽ�-�[rlV�r������+0z�
P�;O���Ӻ	������|�O�H��:d�ñDЪ%
��*�x����z���̶lƠ骋�L>�2b
�c8̝���ŠN���c�$��'���S�g�I�#4�� T4)/$Tp�A��8B�	/p*�s7��;9�X]�6B���@����"|2 O:NF�;B�Y?y�Bx��`�9�Ys'�;�?q���?��M���OH��v>1��R�O+ - N߶j�.�PĬ���C��'xGXD�q��MN��6dH�L#l*�)�X�q�]�}Рq"�ˠ9,��&݋<���(�O��8���:.���@ړP�Z-s�"O��P1�EL��b4H�Z��0�q�Ni�(}�C�ivB�'�ֈB풴	�>P���R5K�x�@�'���ոlw��'��	Z�?b�|�e�.mB���%�NQhG��p<1��O��FB!;c�?cY�9�&�ӓB�@�㉍����9�Dİ?�<����J��M!�>]�!�D:{\Pc1�ϸA�F,*���6!�!���q��M�<D�x}��O!9P��N&�I&l���4�?����)�2����"A0���Ơ�2�P�s�P2�d�O�%���O�b��g~"�UJ��qR2�ʮ���$呐��m{�"<����kLLc�{��yY��T�DF6a�'��O��O�ư@��^�p/�\A�%Ä9gTH2�y��'k�y��I�z�JQ�X
��Ց!���0<�!��c��@q��A�F�)�$"�z�8޴�?Y���?9R/��cv�I���?����?�;un)!�o�7<,�[��֓!TB�Z�y�ۈ��<	�l�r\䀐F�[!^R�b�fܓ)��9�牔1@"`:�m>�x3��[�(�0��<	��[��>�O��t'�'*�05�� ë)����"O��9����U8�i�¨_76d������(���Ӕn9��Z�)³g��MgƒM����޹8m"�	ʟ��I՟�R_w�R�' �i�L���Ѷ���C����D'@FHGL����$M�{ r�
$�V'Y�jCk��]��"�ɦa���䉦aEn��� `�:��B�T-~��Ȉ2�'���'�B[��	y�s����&C�?ynv\�'g�4�<���e���@%L"h�{k�3k���<��T� �'Uf�#V�iӺ���O���*3i�Ջ�#P6���h#E�O���Fc9�$�O$�ӻ�A���
&�pa�'
1q3i�y��h�`D `8��z
�z>5;����"�e�%�O��K4`��$R@���;�-@T�'�z�h����	Fd]��a>��L0�>����(?
� ���|�ԡ��ϒ)oYn����W���,U�@�j h��)�'ǘ'��\p�	zӎ�$�O�ʧ1a�82�"��7��Q��y�R�J>HI�����?�UL���?��y*��	0\��5���,���#Q�ܫW���'\�b���	\���B2d�c�����>1��A�S��_�<� D���4-��_�2ͬ ��X�{�!.N^�B�I��l+>Y��	<�HOf�Z��\���RC�1HR��a��Q�	ܟ��ɅA,(,���O՟ ��Ɵ�i�{Em^DJ4�R@�L�P��D����a.M�q1�$���;��L>���>;Jxp��N�U���Ş�g���PE��A�4XYEEöc] ��}&����Bҙ&$�G�C�[������g�X����)�3���	S�ap�a�F/:�q�n�!�� �m�ʮ����7d�	�ɲ��02��4�4�O*�ǧ�W�����D��� �+&A8v�ˢ��O����O2��ݺ3��?1�O��h8BEܕ^6�tpa��`=�T"��x2�ю�����R@`Kօ��`yT9�'��Z�OY.|%j�e��5�;�I���?��SDV���Cr�je���P/����ȓ3�N��`ۼ!�XMbD#07�b��<���DU��(oZٟT�I+q��(�AȤ5�aI#�$zd��Ɵ���%�ԟd�I�|ʳ�e57M*����BL�rD]qyq��*R�&�xB�
��'��ms�lX�<��R��%�����b��h�Iz�ɮ(� "S�[�d_��P�-�-?
B�	�I��fI7�fX3�舲u��C�� �M�qb�-h�x���@H�@5#�v̓;ݞl +O����|�5$�6�?�q���5P�1�P�ũ@i�%�W����?Y�g� S��ԋj]V���kEN?�O��s�E2��H�Yi8�ѧ��<?"�'��C @�,M1����`�O@�<���Z!����U�<��2�.}'�?9V�i��"}��'2�$49��� �pțE*U�1�'M����ő�}�呫;ռ�s	ÓPq��H�� $X�P�:Ec� iX΀�)��M����?��,lSa�&�?����?A�i��T��и���	��ᓠ��Jc���P&*<O0�2LC ���E�n0¨9B���,.�yR�_��Y���O�5��JO�/$1O�%�������6pȒ@�9`�*����(RrT�� V�X����'�P�i�؍{�8��'�<"=E���W{�l.��S*�5^a���p@V1u~���'�"�'�a�i�I��̧z��y��U�\�n�W�N�'m��g�@F<A3�?>����gO�M�i@����m���=���3$CR�t9P�R4�I)x�X}�A ��P��	/��8��L]:��Y�ćК��C��f���BGU)"�x#7K �bc��؈}�
L$O?46M�O������F�X�����A�(|�n���Ox4���O���j>���O�OH5��a�d��Ñ�׵o{n0���'[L[�B�?e�<c1FQ��*	�c@�
�p<�`��ٟ�&�$��X��0� 4A���r�3D�|��"\9J�P�{UNۥ!3D #e�0��ܴ%4�Q�L�'A\={�M� ��<7�@L����'*�\>�sc�џ`�4��1��@�(��f��]c�!Kş8�	�x��	
Ŋ����S�d]>�����"Y����҉�4l&}"�/Hf��P�|��4��t�j�N�d/���iԶ��ɾ���Oj���O��?�����bd��XDa�?l�1�C$�I�����I�aͰ���F	^���
���[�p���@a�'Ͼ�Ru锋@��I�%焬B>��(��{�$���OH��)�.4�J�O�D�O��4�L	����,�1s�� k6��#��4�	�QU(I
��'���&�?@I��1�L�"8� �{�ߑ))J͆�	�O�(�Z��NmaV��"U���IG~��3�?�}�I�����+�\Â�
�<qqd�/�>y��/�4;�HM�i����5e��H7�,�����D�O��<�r))�U��
�!��|蚈�4�'5���ת��as!��DkҵA���6���9���+�!�$+��DB��+�L�b��	~�!�D�?\|J��2�Th�B�ʢr�!�dJ�Iܱ�!
�����C�۳!��R	GN�$�R��6��@%��7r!��'ef�X�hj�j��K�ei!�d�q�T��oҠeV�{�˵sM!�D�K 2�B�����R%��,;!�d� A�Bd*C���W�,�+��Q�/!��J�xe��j��ǋ�\�Ze�BY!�(X��%aѓT���	�j�-�!�ܦb��t����&2`�z4$�{�!���tB�A�(�h���3����P�!��>6P��:��'9���Y� �<�!��̭;���+��[���a `�9u�!��  �+��/|	b�#��:����"O�h�Ă%LJ䫅��q�z��""O�IcT>S�hYu$����U+ "O�iS�#�����8S�T:v���"O ����:?��e� �O��8��"OLxq�K�+s�b�x#_���� c"O>��FC���ءe�W�P�\� �"OD<yū̾��83c�S I��3"Of�QdK<u��jS0l��7�3D��S�i�q�n̓w-X�t��X�n1D�� `$ݘRG�����5Ya��`Gi+D����Z}R%�4�ȕ^�ț�>D��e�ћI��0b��&Y�^��b�>D�@ E�=����V%�J�dd�ѧ'D��I��9ØL���_�-Lr�1�!;D�,ڳ��7`!ND�c+߂-�>0� �$D���,a�.�{���*�P���4D��k��C�D�씻��D��b��1D�����*u&�q!����n9�Ђ0B1D�8�c�,~�Ti�4KQ�`J�9˳l0D�h�·z�>t`��0�v�(�2D�ԣ�lıx���M�
��P�'<��.�&iR����.=e��T��kK �I����}�|�'̔kJ�� �i�@�'�w�T\�A
�(9�]��';����"C^�۱#_Z i����:3���w""�'/1�0�6E�A^r��^:0��ȓ5!0��u��>SRȹ�/�9.{\�X�X/�sU�|���'FL\�	��Wl6ɩ���/t��p�
�'t�)��˅Z�"�x�
L=��R�'W>�ڔ�ƩRha{bM͞Rr����K+$ȗ�7�p> ^�C�Ty۴S%V	����a( �A�ѷP�v�ȓm�\}�O
�P�
E���k�b�Fz�c״a�.}Ï��J�����/g��M��( �!�d�5a��`�R�ܤ#�T�����!�Z�A��ip2H�Edl����l�!�D�/.J�iTӸ_O�|ѧ�N"c}!�����aZ3u���s�IT�o!�d��$�A�(�����Ƣ�)>u!�ĿN/ұj+�%|����&:k!��	B���(_������-9P!�A"P� ٪ h�R����#jG9!�$"�YX&�=�~Ah�`�7?2l�O�ștC C���H?��P���U��uk��� q��Y:d!#�Oy� kC?�:M�b�I�����	�3��K@��: ����~�����$	�����ڇf�ҭG}bg�;�Zm� �P�]�O���íP�b%�dr�˗�}T���'/\�VH�cL�)�ҡ@�8��'R��X�NC�%JF�Gr>�3@�^�n��IX^2 �3	3D��Q��7(�y6��'z�:,���"��ɱ},��Ua@j��g���y��)� ^|B���+8bU��	�\�ZxRܘ@����b�-4�*�͒ 5h<(J䯚*)�~��ǒp��`��Dy�n4;�� ��y�&3� d�� @�L`Sc%'�y�`5kq�M��?-�r\��f���y�(F�EQ��e�P��=!���?�y"HТbi��HC�+F J�ˤ��/�y"Bʋ	�8����X�o���2U!���y�+	`@ݰkɞl��r�ߕ�yR�[_F%�č`�(���M�y2�����@RhɌD,B1��V�yr��5M@�� ��=5~pɐ�`��p<yp��t���!KR�	���jqE�
����f�6�\���)B�zBڠ��'��C�oB��w� Q�Qz���>)��C��q�f�L� �%ėB�ȓ�� J��
)���Nϼo+�|���^j�<� ��� � 1s�"�+ ������y2π
r��Ђ� )���r��	��Ɂ7,A�p���p��XҐ��/^���Ă�L����+vL6�;���&=�5�"��n�R �lۏ~Lmїi�>��"x�I3���J�4�2�s�����S��@��6�|�`4�	(e�����K�q9�A�k��`��
��^�4�*�A�'"�[S�&m,�ȩ�M�韰�u*R�u��x�i�r̒ ���J	LTb�l�0�"�$y�>�{G%��*L��'d��(�R�(pс q�D��v�١$ɒV�V��,gJ�At�4��0��/Mڼ��$H%w�,�1aJW>�,�#РŻ?Ts5Ί7���2��~���1�t�3���VX��H�� ؚq�ל!��|X"�B����1o�O�����C�����!H7j�8��>&��哇ƚ:��v��>Y &�x���Cc��{u^�g�j�����'�!s���:%�%I��W�~�*я{�R1U�p��;$���j�!Q2m��Q����2cbW�G,�}�4�C$2�u�c�G8w�fd{�
�%�8eC&�H7}Fz�3gjG�����q��7>����M�j}N��1��9��q���=0����>�8�r��~=���E�*�N��'�M��l�v4z\���(�قuȈ�N�] ǣ�'n�a}���	����!�
F�D:#bX���q��d�j]r�a��H�jeH�=��	�Ϣ�7 S2.�̚R��92��AjeT
���qo�m����J��\�XggR�7/�| @�#z�v	
��J #��0R��A9��m�p?it-��^���
&�	�,{�Xw-��F�B���z�v!��cF�+2�$Q�T�~i����O�Z��ۃ�B�y�>�HY�2Ez4{��¯H���/��$:���H�=�ņ�/x���T�C��@���4ر�I
��OȤ��T�O��0�
I�;(�娤�\�|P���r�	=#h����C�jJH���D�W�2�Y�{�����e�⌨}Ҭ�� �"J��s�J�!���G����>	��Uąy���yr��`���o��Vi��&O N=c(�?��H?9���hh۷�Awϔy�"F��Yt<|1e(|OD9�A��7q�iر�Y	z�Șk�*����*����Y(��-]$L�@����R&Z�Ia+�x���B!�R��B�tLɡ]�jȰik��
��O�\�s��7\(���E!�`���'�|�Îu���y�F��$1À")���u����2(�9FLH��iך k�#=Q�l�0H��U�I�l�$U��<O�� �ix�<����j��q���O��Q�Y�,^$T
Z���Q/��4�h��C;��	d�^u��I��6��|�D�E�>���`��J�LJ�����4�Z��c����iɴ4*��*�L;�I���;���rUO]�]m92u�,�,7�O`����;��k5̄(%�Ƹ*3L]4\�:����v������9ʤ�sQn��d�h��q@K/m�+W�ɞ[�>�����P�T����h����ė�����µ}�F���l�J`qǢ2`ȭ��$�j|����Oj!r��**�"A�¯�1A�`s��	�OQR8�K�&xԔi5m�T,��
��+�b�$F)X�c�!Z�@��}��Z̓h�QB@��;@*�  ��1(�	�n	D���"�O�!���P�� CMU[��*	�>��)mI�I��eQ�;��|�2����Υj��![6�J?C�d)�"O�T��.]/5�|��)�dm�I�R�L�'���O%m��P7�W-2�H�O�2iߒ&6d�r�5ȮpY�ܵS�,kfK6�̕����%+��\�ι~j��O? @����ǀ�05��IԎNw��A���;�io�Fq0��Q1��Gz��<�)��m�<	��q�w�]1�PM!��)X�ȑp�=���,�1O����콲�a�;K�T9�(N�����	_��Gz2�+*�D/�m?�"��;gh��jCHG&z�p@�C��iR(�q�'�1O������',����w��-��̇�tA�r�3E�2b�yr�_2`��r����b�fNEa"
%k����� ��h��	W(ڰԈ���3���|R��i����v!ƖB�|pBG�P_�̴(7��,/�bm+��4���)O��A}��AJ�	8>��aש
L�0�i�:I�3	�G8���pO���	��V� ��Qɨ<��4�n�c;6�є-ô31*h2�C��_zȷ�ծ�0=ѥM�J=���bG�,����c%[�FK��I�^��QT-Wn�Iʟ��'�l$�g�y;NA�9�Y�l�1%i� E	��}!kޱ:!1O�| %cΑz�Q�)�N�d ��R��̓A�T˄�H0袤��M�H�'��������M"�o F2�1��d۶��M��CYzx��d�5v�l�4g��0%�����	��|�'s�(9�`5j��$j� V0��N��sVQ�B�^��p>)c��� paϏ3{v}"#�Uy��i>��'��٢�����Pa�ўqҎ����-3az�`�)�h����Y�0��ᄒL8&�(���(��a��U9�<9U�=oШ���݋2L�Qp��{���E��,��e�H<c�1O�a�X#0���'j�d�H>���9CT�ӷ�-0�@%bFg���p@$`Bo�B�ܓ7LU=���=1@�������W�A���8C8Q�����t*��-(`c���a8�`@�fԌ`�lQxRA�X� -���&t�F�
b�'5
WaH�(
�d�%AS*
�֝aO>�!IC
��<	#˜�%��̀`�AS��1��&S��p=q��D�/��˨On�p��]t)���C�D(It(a��'����G�T	�)c��F/�� hUsa癘y���F�]�r���'�y��T�8�� K@��+{���Q��ۯ9̅0����17d��O>1����q�d���D�<U������LhܓN�2)��"buGj98��<	Cb	C���0!�� ����$*Fg�~]�t"R/V1nz٘���mbhH���Xbub�B���IaX���
N\2��C��
��"�I�I�����c�<��t���oB�y��8w�
P)V 5� ��G�Ɂ !��J-p߶h���6wHf4��HI5y{�y��7�f5��@Y9��� ���i����b/�%��eh��b�az���2c2�ks��)��L���1&�bY9��ۼ} ⫁���=�"棑�|�a&��y���=��
P���'��>�Q/Pp� N�� H�������xy �&�����ɾf�^� �c��U-�oy��i�E+r_:�3
�S.�����7%��D�����'�J%*D��&^�@�c������S�'b��@��ނ��Dpae�S�ć�0 MCUBÍ�D=�����1�J�'��4�z�@��h��y̧h��'re�ւ��z< ykCK-&>L��'�rd�f�6�h���@�Z�N@�#�%�mQU�(O�tآq�}rz1��I!\�^��@��4o~z�8D�^�n�t����%2ܤx�׃�w�t�� �/� ��Չ0G }�t�Оaޜ���A�Px�ϙ !����9o�x��A��dW3�ޕ1􄋣l,�8�dI ����Z�6���� M�TE�<+��Y�y"F�;H?L�s'Ó7O̺�J�Н+ⴼ����7�<x����$0ܻ��ԝxB����ܵbv��2�xa�ȇ�yRɍ�X�ȱ�V�[�I[vl���y�%��r�f�8!ȗDJ�5:���4�ybfW(L�-���7@������\��yRG��aN�`k �Qan�k��P��y�c)iL>X�gǎ>,��"�IH0�y�N�<�uZ��͚"<�W��	�yҪ��WX��3`�`Ț���y���Br�T+ËL�6ʣD���y��ݶkd��9�m^.c�$P#jG��y���L�,%y����pbc���y��-�T�&�)r	9�Dʻ�y�H:��@A� Rܰ�Ԧ���yR`"KtJ|�N�,!��D ���Py"�P4v�z\˴MԌCM����t�<qg(;M�����-�}���)��Sp�<���I	/oJ����	P����J�j�<فC��	�|�
��ẔjJ^�<�E�U|��9Z'�W�!g���"�GX�<y��G�n|c�I0A��<#unFZ�<�E4�ƀI���25}�X�f$�L�<��֔<�+��G$[pă0�	A�<����i��ԩJ�Y$Yۂ�r�<1U$�@�8�����
�.�y�<A��^g���E�Ջ?��}��'�N�<����L5�P��2_��0�jFH�<����R��
��
R�ޕ���]y�<��N�/y��Ȉ˄e��p �Xr�<i�!�3Z�d<c�a��(8%Ęj�<1�.�����f�C)��y+F�g�<�����p�3�Lu��ۤc�d�<���:M��}@�
�fC��b��d�<���F�@�&��Pxl� �X�<��d�ЭPu��c�ڌ���<��$���S�Hc�Ԩ%Ør�<�w�BR��tp¢GUTv�X5h�t�<�&��:�H��ED$R�U�3�j�<�S�/o���"$n� `]���b��f�<1S��6#��]�b��������N`�<��ܺ�6ݡDؾv�����\�<���1� JPO��e[|Ų�BIr�<I)<D|�M�r�Hv��ы,l�<�T
{L�edlԾy{�J�g�<� �#�,Po�|A�Ȟ&XިE�a"Ox���)G�%PGIׂlI�"OF�xf��'|��`0� �8;��Yk�"OԠ��	�ao��� %A�pM �"ONQ�V��Rb^��� S�ް-�"O�H�f
AwH0��$���*݉W"O��ٷ)�血���48����g"OLh�A˴z^�P���R� ~@<��"O�܀�&�.�D����R8STu��"OB�ȠJ, '*S�؜�I"O�����RY'XA�#�����"O8X�5j؋R������Wj��CU"O�m�R������ԤANn1s6"O�Ͳ2J� ��	G�õ��Bf"Oh��p�2l�T<yU`ƀd���e"O��{����z��/ȥ �-��"O"��u�N#�>���\�H �,�@"Ov��2c�=�ĥ��$LI�"OL�2"���~g�	� �V�٘�"O�8ʃ��`Bf��2/��2��%"O 0�Cy���A"N�,���"O��S�u�r��Pi�OU�˴"O:��U��wk�m ��7MB�)c�"O �R�eψp|b��g�s����"O��� Ũ~n �����V�4e2"O�qq�P�>/��A L�*i�U"Oh[��F-Nx���嘸A��ec�"O6I�a�6J�< rE�6�|�G"Od�����x羼`��K,v����"O8���l�7��0��L4�ࢄ"O�h@󋌓-�,���
���aY�"O�4�FiV$�骇c�G �hp"O6�i�+T�zU�Y¦Ȇ��ι�"O.��%��(N�*�*2H��y3"O���T)�%y*��v�8+��=p�"O��x!cC0h��3�ŋ�W��!��"O�0�q�H"$6x0��I������"O\��ċ�.�`bI�^�h"O`-�
F�5� 5�V��8��"O$�K��<I����cŒ�t0�"O�	i�̀�z��ݣr�E�@�(�"O6U�GZ�r<P�E-F���()�"O�y V��y3Ȅ1�L��q�@}�%"O�,y�mO_Wƕ�f+|��!"O���m�<�HYБ�� ��)Z�"O(تe��$PWt\B���8�0X0��'��'���h��Ö
��p��N�	^@@�'��8�A�F0�aT!�0 �����dԷk�����g��-[�?W�!�Ą1)���qEȖ%sDePeJ� �!��ӽh2��:��	7Y*|��	2�!��P	)8���X�J�
��%�9N!�O 8�>ڲɛ+m�\��AL��!�D�<2��`���_��h���D�!�D��O7j���D�,�P��2EX=�!�_�T�����C�`xR�ɸ�!��&lB̈w��4�J�ƭ�!��	�y�F䂕D�5$���0�ͻo!�E�n(�����K�����-]�6O!��.�BD�[1Et�TA���r>!��8kɒ�*���0n��Tؠ�!��%)4.T
��S#nW�t`&l��F`!򤝔:4 P���An���Л>9!�K� "���	k
�!S�-!�� 
�I%CI�
�yQB�=|*��"O�-�Ql̨*6D	�n�\^�R"O(1�3ǊC�ʁk+--���R"Ot](���+��ᑯ
6�8a�x"�'��	H���D�R@���q�
�'���FN19��P��9m�%��'���@���(8�҂�@-�İ	�'�
�@!��qM%b�  l�A�'��B���<P��*⮌�'}�b�'��BaD�j*$�@�IJ0m��=�
�'��LJ�O��{�/
_���j�',�@A@AJ΅���ۋJ[��;
�'�P�(�O�S|:��m_�FΊ���'�p&cЎ>��%�g͐I��'dzu�A�8|��Dg� a����'�v��#&�yK�_�K�.��ȓ3Q��pR�r�q+b*�-Նȓb5\h8E�!>���#��Ϥ	~����EȬ���2Z��Eb�o�LM�1�ȓt���Yg�9Fj������@��ȓӆPX�똏_qYIc�Cr'�ݤO�=�J���;q�,;�8�7�T�<qw��0zP�y��+J���y z�<q�c�W�b���'�?OB��Zv�\�<i�'�;f��	�#�T'Z[�x)5eTV�<Y��*r0̄�F���"l�r$Q�<���4<0��5lޅ#=(��aZO�<���_%f�x�e$��N�ػ �Nb�<ys�̼D��x���ۓ �y�C�S^�<�C��:zl��r���1�0˄�[�<�h^.�"��""�:ڎM(�F|�<y�MY���ۀ��K	��A�'�a�<�ҠY8�����.G	U��!����d�<�pG�R��8&�ZR��j1(�U�<1f&�?@�D�E�H���VF�R�<�w�J4��,�d��<	}(�`"$K�<�V��'%����[.SP0j�o��<I�G(z���ʥ�Ȕtt|�q��u�<!���.,�l"�!�%�_>-{�B�I�}�h=B�GѨa�R�Z�읓*U�B䉅LT����#1���්[[�B�	 q��p�Ƈ�5G�c�V��F{J?+��
4D^(*�<�D"&�!D�x���8m�m3�+U P�fT;�o�R"<���O����EU�e��IjęA1�|Q"O��Cʂ!K	z�x���&1�)��'ݛ..�O4�R�+�<���C���@��3"O0T�C&J-!x�)å�ۚq�E ��,�S��ɔ;��H�D��=%�T5����Zg!���c����ݠ$d��+eX3wd!��"a�ݣ�`��d�!4ʏ�C&!�D�=�z��D�=x�j$�4j�Oԣ=%>٘Ө�J��@�%ΑV��J�a?D�Phgɏ+1N]�Q�wF4}��!1D��0�@c�v剷�S�3�H#g0D�����6;����	>�Ȉ��*�>Q��'A�S� dպX�s��`�f��'4��{3�W�`8L P�кZ$ʰs�'���G!Ⱦ`AmCR&!P������D!�f��ĉ3�;^O�� GR����ȓ�j1���(�6ܐ -�$N~�H�<ы��	S���۔�!����X�!�!M>� e���
o���q'��fd1O~��C^<����A��jd���lJ!�� n�� ˔_O�miB�-�P�t"O4=�#k��hx<�c��8`���"O$E�%o(:¨ɡ� *�@i�"O^]I�J��O�/�&j)�"Oؙ�"k�qmj=��u�����'��	J�
풠�R�|t@ɢ��<��B�I�L��r�$�4ӆ BZ+Y"����7�Ʉm�.��I[#{�L��I�B�I�4�~%�bk�z��ۣ%��"?ٌ�)��$�4C3�D('�����!�Ą,�����"��~3���'��Kx�'_�i����'��41M�&3�F��	�24��
�'�6lC!�ǂ�6X"�D>/��
�'���a*��(�L@�c��+E�2ۓ޸'M�X���]|�H2C�F'$p~ i�'B"��ġ�pT�i��/��*��'����6|�Za�֩
�H���'��a#�\}���LM!	�n���'�ў"~
ceب �ֈ��D��KQ���a!�q�<ٗlwt��"�Hx83Wϔj�<b�W�!2��`7�ir�tK�a�g�<Q�'�"-Vmp��O�XƖ���eZ}�<���y������*Q��XF%Gx�<��� 0�( S���$7�:��5��s�<a�mB�+��a�kJ 
I��@�I�<�D��"K�=��͕CJ�xǧE�<A�h..�ŉrߛ�B�K���V�<9P���a.ap��TH\���dT�<y�H�r��Č`P�b� I�<1�-2-\}�ˋ�8Lؘ!�
G�<�
#y��dc�G���O^�<�ҍ�xvP]��e�M�,���%�W�<	�&�<b��U ���
c��@Rrk�z�<��+[�~j̃�K�-#U�����q�<�3�նj�5��N�P�v$��ny�<)��L�J,���ْ=������u�<r#Թ}�$(�7�B2�E�"Y�<Q0B4\��I�V�@�VF����.�o�<	�ڿ~��,�p�S_?~u�e��<q�7W�40�LZdFF�a!n�T�<i�F���7����RTq�u�<1���-�� ��Z#'�!�&q�<qү�9	U|$�g�J	gr!!MUi�<�Gj²�b�����T�8tNO�<!�FčG'`�2�I���]��$R�<�G,9N�h1��f�z�]��o�i�<�ΟZ�aҕ��g�n��R�h�<Q�`��Z��{j�M8�cWa�<	��	 �!�% �<�z�z�e�U�<Q@ϊF���p�c��͐ۀ$y�<ɡ�&jp.�A�!F @���7aK�<C��=�h�RA¤D��`�O�J�<���&$���	�7��mP,�F�<a�,�(Zh� �s�~�-�u��K�<�$A"kAF�0f� �,�:�S�IA�<	�O�W��U���k[�u��b	y�<r(��#`d��W,��f>�I��w�<)�� <^���K/2&7��/�yr� �̸�I��Z�����h�	�y�OT�xԫ#lZ�r��&�Ӷ�y2�M2>�V4#�T,8�(��J:�yҩ
�
�ii���2G��[A�D��yr#3.f&�#���r���I�y���j��mb�߀"��CW!�5�y
� �%�чI�W��e���K!���q"O��B��!��cQ�G�,q�"Of��b�?$���m܆��d�"OqR��S+g�Y�v�N��<�7"O6�x���"�xi�!�ī|
ɉ�"Oj݀C��7p��ʕ�*g� ��"O��
@Jβ50V5�e��TY��	 "O�< �<I����O�T�L�"O
r�V10�0}�E&I����"O$\�q��M��5cV�D+0���"O:X�d���������H�rh8%"OB	���0P;ȍAW���D��JW"OT�aM���xh�O�%�Y�a"O�riT5@ ��
w��w�nA�1"O}ǀ8!>R��#��,�4UBe"O�4:�O[v�p�J��H#dYl`�"O�e�7ɝ\�>�Sb	#���"O��ڴ,��fp��@�aP
gxQ��"O��`���	$<�E0�lJ6ɚ�"O��Ҥ��J�%Y��R�S)��2�"O1���4� ��d烟C�RE�"O�a�O�: R��(ӚQ�4�"O���L ��5?��h�c"O��[��V�Tc��s���	��i��"O.� 'oǒK�LPaȈl8�, �"O�}��:y�:�� :�0�"O�\���n�p��u�^>aa6"O���e��Y��,�M�5�܁ "O2�y�����.�[���i�"O����z�<��G�	� m�ى�"Ol����	J��C�O� i�ɚ3"OzU����1��r�+�C?`��"O��S��Gu(�35l��m1F<h""O��	�a��t�\��5d�8��r"OD �-\���B�Z
��ٱ"O�d�w���f����M��5�"OZ�$��&4l0EU'���"O�`iԁV5J/2=Cc\?x�
�"Ox�z�����.W��6��"Op]����8)4�3�O���>�s�"O��C��
��@��o.Iq`,ل"O:l:+Ng�5B�B�2�β�!��F#z� ���h�R�ȩ��	�Q�!�D��J�d�H%_�1s 1<.!�dq��y9qd��t�5�^�
)!���P��	� ���T���bm-!�:3����b�)\Q�Pm	!��Q��a��`V>H28��ˆQ�!�DM�Mt�đ4l@
�L  ��P7�!��i
 ���ܯD���� �#$7!�9o��Z¤ϸ~�~�:2���$.!�$ � �v�@��@�@��4��*!�� �N��e��Z
��3)�6	!��[�x���sk�]T�A�j��J!�D�8$�|Sv���I �$s C�
F!���C��e�*�!�z�Z"�
n9!��&<��x�`�S�S����i !�D�\I����� ޖ�Z�I:!��9/�
pIe	��T_���i�O!�d�9M���Z�cF(9�|m`�Z*!�D�7	`��� T��JP�]6!����e�7 ײS�"�<Y��C��n�f���^�>�`
ŤQ�C�I4��h��7�n0�Eŝ<��C�)� ���v��2��� �	G�P]�`"O�)Wg�&0�����%Ǆ>��,a�"O��r ���V!�Tb���ê�y�"O�e�u�́NU�	cmK�~��]��"Op�I
R=d4���-a�xAt"Ox�C��-vD�hE+%�"O� ��P���\�&��an`�"O�\Ó���8@�$K�XL�"O>!��<�b� �J7�(ux�"O
�SwB:7��M*U�Y�a�`�y"O4Y��Ag�k�AL'|u� �"O<aY��.T��d@��J75h�i�%"O,���./t��0@V:Y����"OL��g^�>>|��ӅVu7��K"O�JC���5���Yc �쑂"O�S���I�$���F�D ���"O4ͪ��R�r�%�V��]wT�#'"O�	�匄� (jթT�Μ.�`1�"OȔ8%}�1��Z�l�ڶ@�!��RA4�B0�)G4r�q"OB��`�܀e�<��%��R�"O�+@ �k�dys#���:�s�"O���񌘙 ,	����y��Ԁ�"OB�z�#�j�@ӧ�d�fx��"O���"K���<�j5(��T�`��"O�y�f��BUu
2*հdM���"O��â��(��D���)]����U"O�0�P�ոWN�]�`�[��~8"O�Z��FOx�ófHZI�%"Od�ӓ��&[�!�� Z/LIj"O:�k���:�ѐ���	<9{�"OL�+%I�<.[x����ǋ%�M�b"O�MZ��ԏbhf��e�#~��c"OнbP��ij���-2�0ZS"OpT�3���`��\:|PJ���"Oz<�Ve �><�mϡgEr�"O��j'�̑Df̠3@+�&Q*�� "O�J��Y�<�	%�w�"|Sa"O��q ��M�p��Q�
�u��#%"O8q�Խv�Τ1uhN�1��A�"O��i�*rA�@:ҦN)ar�h:�"O>=�����X�XRA�K��(�"O.S�FiR��U�j���"Oԩ�dO��[`#��:y���"Of�8v�3Id8��t<*�xA"O8��'�en �`�B73:}�"O���M��}&�A�$ߠ�h	t"OzѢ��W�V��Qj�����"O.t�q,X�����S�B�,�"O�vY|� �H$j�����4"OxE:�ϛ�Z���F���ad"Ox`k5 F�#��b5��r�p9
�"O.��1#D�X��=sf>Q�r�K�"O��k��A�2�<2��:�0�"ORUj��9:>�P�@�9S��d"OH�+$��y��y&�=>\��"O���U��bvtpQ�AY����'�B:OX\�e�Z(P�yPU��nk\���'"�T��(AKؐ��eI�~g܅���3D��b�N�?pˈ�;�낗EX����0D�P:@�'Q[6�Y�*!%h%;��,D��2An�(?8��!დ�My;7+��i��P�P�>䞝a�m�0�0�ҕ�+D��C�ϔ2D�����(>] I���(�O��)� ��K��;g���i���?d|J�3GT�F{R�'�1O��R3�wl��0]�K%"OBQ�`��$F24���6xUB(b"O��㵀��"��ԁQ���"�b�C'"Op�0ᇏTx���)ݟ5��0ئ�|B�'y~8yc�z62�1��D+,�C�'�b)�B�֧ ��qX�-#D�<es
�'���b��\|hxȇA�'I[��	ϓ�Ol�
��H�E��NK23�i"Ob,3F���i���E��t^�Ц"Oh� T��*���flZ6Z��"O����H�]¬�����2$A��:�Y�����)X()R������f`|!�B�Ib�K��0A`��� ��IG�C�	*9��݁(�J
���)��d�O�����BT~i����i���׬ΏP�!�Z1��0r宐�,�� ����\�!�߼Qۢ�1%:�Č�p�TX�!�dT�0і%�6[�`��
��r<O֔hse�[��lJãG$�z�"O(�۵�/�lQS����?���"O ��"	1!R���W�R�33>���"O� �1	��P��D2�F�I �p"O\q�Qj�q�N���d�F��P�""O�(�'�?�H��`톹S���7"O4�{�j�>f��a�R ;��b3"Ob��qL0(�8 �)3=�l�g"O*a2׉q��E�)��
�"D"O(Lx�N�6i+T��ǉ;aRL�T��3LO�����$��٢�DC�<����[�|�Iٟ��IIy�T��O?N*s�������J�T��'2�h��\�	p예4�Gxt�'WPEj$oU�NK����雙>ր��'"��G.W̤��&@7 5�'x.!�a�?c�b����W0 ļ;�'�������+x�h� LM�j��`���.OQ˵�	6LD�i�� �f!d���'��'��)�-
�k7��7/�� %�5xH��'�����L9_X�퀶A���
�'"R�R��'*� 1�2�L�db�0�
�'��\��ڲ]lmт3_��Q@�'1F@��Ez:P�Q�[_0�-O����O����_	c�8�* �T5M�IK�,Ȏ2�ўP��:0f�h9q%��Cĉ	� S:r�O�ʓ�0|b OUt�tl�sY+!{�`X�K�<Y���6+蝡E�V]m�\ؖfAI�<9&�M�IKh�w��/=�]�P$AG�<e�h�{�L��)���&F��<1�d	�r��]�ǢE>\�$���Ŗ~��b�ȠG��V-~Ȉ%�S;vᱬ*D��J0�"k�nu�̊-?�B0ð'*D����K�x� �r>��[p�&D��D��	�n�`�O�O�
��#d"D�0J T�q��y	�f��-+���l=D�tّ�YW`UӰMM�c�8�g7D��R�%�7���Qn��|?�x�6�O��DHsun�ѷ!O>m(�m���4o0�B�ɥW�(�#���D��A�,�j[�B�I�8u�dhSgԝ!(R��S'Z�>ئC�I�-f �P�ZiނZ�C�>V�C�I�&9ؠ��#��q_�q�V'!,�lC��B�%�V�L��v��e�0a��㟀F{J?��ж*>�Z�i
��5DG=�O0��$��i��l��r7��t�� ��S�? n�˴��&Cq �)Ȟƈ-i�"Ox�1�A0H�P�AI�s��iY�"O�i�ф�'UJ z�*3H���"O<͢v�:���i#y��!��"O��:��P~ڈ���A�o�ʥ�0�|2W�h��S�@��t
s��AhP{cϚ�z��B�	 O�9�3G��;Ц1Q��\7!�B䉻E X\IFG�R�.y���ع;)j�d*��r���]�(x���Q�CS*uj�,!D��R�ÔN���2caM8X�p%%D���O�=i��)&b��0ъdR �6D�p�$��;VM�S�̜']��J@7D��)d��2y����@��x��6�5D�T���$9���E*���+a3D��8��~�R�Y��
�&?�`bC�/D�lQ�H�����:h���) D� ���h@�ص,��%�"�!%=D�T�u�\<L�=�R�>"�
��9D���G�@"w��۔@;o�2��sB"D�D0%Mݑt�m���
�iE�w�?D�xZBN�$a4 ��U���g*OfM���e���3n�7N�D\`���z�O�����R /r��f�ȳb"|A�'ZLs4��e�2x�a* ��'�"H�+(y4�2�Q�RL�@��'t 3��Z����3�O�,��
�'�ܹ��f��E��2��-���'rtu����u�pK������,O:��dR�*��g��$,��hW�Qq`!���t\� b�l���fb� P!�$�v�� ��o�
3���bȬ,6!�ĝL�ɒd�j(s��;!�D��)Mօ(&#"���gH�eў��ቶ3��-�Zr�ݡAF��3����@_����I���{��J�zl�q�uI'U����O��$*�OPuBPEF@�D�s�i�~� 	��"OB�����z���7(�}��@Sb"Od��Y{n ���-L����"OH�`U�$1B�8�kڝu��O4T%�'8�Qaƈ�1*��&M<D���bΖZؑ�a,GTD�g�<D���cH��mAv���"Cz��@%�9��3�Ohܲ#�-�|=�UF�2gi
��B"O
���|S�Yb���UST��"O��В-;_� Q�c֮A�ГU"O�X"�����`!���9>2�� "Ol1���s�qA�N���ˀ,̊�?�O>!,O1��?V�B�Z*�����L�������<	U��yH0�1�)ѡ$`Z���C�<a�S�ɔ��e	N ~�v���$��<���%I�������|���q�<a7kU�S��\`�2�lt�w.�j�<e��,�T�p;W�L$�*MR�<Q���5b��s�V+�
T�ΑPy2�'�����BL�����ھ�k	�'{H��׸y'���� l҅b�'y�pAɈ83�L�*$ES!D<�
�'��Ax���6��<���ѡA���
�'9��E��h\ʭկĠ&�P�Q
�'/F�Jpc��Aj�����e�c��y��Y�~��W&��<�R%1VB���?����sS� ��jԾs|ءef�->�d�ȓnr!���<���G��D�ȓ%@�zU.��^�v����2d��̇�S�? B ړm�'�0y��:l�v���"Od@������eȉ+��Bp"O��!b*�a�8���V��}�D"O�e�g
$1G� S�Hڣ0$4��"O2]Q�Nٌ!�ޭHp
��$�K�"OT%���P�I���QU�,s�T(d"O�H�Tg�.�6!JJD&|lZ$��"OX�0b��#oӰiJ�揄KX�|�p"O�d�f�8<�D(�A-$W�9�"O*�ެ&�d��["9��w"O�RWDE6\$ܭà&ۡXW�) `"O�����Ӏ��0��d�'p|��1�'LO YcdH;O��t*�N/��2e"O���%.�S�D찆n[+k*�bQ"Ō������N�Sė�J?��re"O��a��3h����!�IK!N��2"O�Z�B M*MFiЕ-����"O�dKe���D]�ȋ� PLd@@��W>���
{�������D#�$7D��Cg��a�rZ6�A6kJ�y�U6D���4	٘B��[F͊�z���'M'�Ic�����m�줻��?����:D�����J�T�8�bd��C�Y�0a:D�$�C��Pl0�3��\_�	JbF>D�l�#Ù�s�p�G�:�<=A��<��0|��*]7J�us"�R�l���"PN~�'��Y���n���({��UY�x0�
ƣ�y"�� 2�C�g/�Sn���yR�B�v�����Ic\.���ކ�yb(�5Q��(0ħ˴r��bWH�8�y.�M�H<�g"��T�~�2�E��y�h�MA�Ib����c�f��v��?1�R��&C~rr"I�!�"���,ٲ���	� �'�Ш���B#�\
o]H@s�;Ҧ�B�%/D���&�լ��!�[��<Ɋg�-D�@S��ɄM�	#rJM3$����*D�lI1�\��`��U��I�(D�� �N��=.���L^�2��"D%D�L��A��6�@�4I��j�.�8t$!�Iʟ\D��'�lX�4��&0������������?����	A�g�dM/!�F�dc('��H�+ރP�!�����S�����xB�N�\�!���YB �)�,*�&�[Gޮ�!򤛙H����׍��J��!F313!��]����2/V�F]r�Oʅ!��]�J��̺���Y�ٳ�Nܢk�r�|]�"~�$$0w�4��/��{�b����y��>W�x���H8au�����yb+|<��AT���
R��b̓��yR��'����G$U� �l8��y���6�HB��U k1"���=�y���?V�X���wҀ��Ee_��yB��L$�-"�*>uʚ��w
��?�����t�t����Q�+���q��-_9�@�ȓ6+�M���9��R����vxȇȓ��A�m@mp�-����'Ŋ�ȓF�p�A�F\5΄��9#�@l�� ��|�����Y=4���6p�b��ȓAZ�K`�70��`��*EB�@���P��0��H� 9��i�!z�0���)]����J��|;��o:�,��fD����G�E��2�c�>O�̈́��x!R'X��@�r�O�i�(8����0u`I�z�: ;�E�4t�M��S�? �YpQ�kך!��H k(D�P�"O�i�L��-�ntBJO�P�7"OjU�&M8&� 03���*n?4�T"O����FIo����I��1( ��"O4�2'jC,.T �Rh3M/���"O:\�RaΨp?H!�Y�n��Y��'bў"~���Y+Ji �.S%(<�����[��y�n1��E��C])����"��y2DX$f��Q+��X�ZY������yr+^� ة�7l8\8\��ꄣ�yb�<U��l@rJ�X�v��,X�yrH��h?��HH�]�: �v���y�*6��л�Y�=I��6h�=�?���������8�C�_:6�R]c�lN&�85a��,D�P�"�:F� �q��{\l��A@+D� 6`�"<<*�
�j(��7D���4�F�*j�2�c�=i��A1�4D��k��x �$��8<m���-2D�����K����� �Юz�x��+D��ʴ�W�7�����n͊b˴�i��(ړ�0<�H�.6D�Jр����Jp�Kr�<s�.W�k���,�&����H�<�a��
�rѪ�/��yz5�SF�<�Nט��:�$�&,$�0�F�<�a�@+1��ј%JB	m+܅*�MC�<���Ųf����3��r���q��~�<�ȕ��q�G�=Ų=���x�<m�\NlR� 7X�r9���w�<9Fō<F���3�އ_�$A0��w�<)t�[�;�p��U�܀bX��2/�X�<�e�|.�B��^�4���Qz�<��؊���p�ŵ�Y�0�u�<)���F��)«�.A��`�U��e�<�Ӥ��oiV���˒T�zE�7nBy�<�䄋,�>tq�OF���}iӦ�z�<��ܡ}�f`���1�ZyId��`�<���$4,����v�r�a"�Z�<��(�\��ِA��  ����V�<Ia/�p+(\h���=��Q���T�<�� ��$b�����J�,�#���h�<�!�

F�xDs����80r��~�<!�	M,k��2��������Gv�<1@�Mm�.U
�&���m���Ug�<Y2L�Hw�L�&뛧�a�Ǟa�<�BlL�5x4��a�ڠͬI����h�<i!���5u��To�3ٜ����g�<�0&�Rߖ3g!�u�ѓ�I�<��)+��M0o����.;�C�I��)��l�%Nb<ْ$�(Wf�B�ɖN�L��5jJ:p�h�R�U��B�I�c�+%�Yd<�s��� �lC�ɜHܱ�a헤��i��j��B�I'g��P`0���4-�E�D
�� C�	�Z�A�U��5w��Ź0$�6C�	�aZT�֪I+[�mhp 65B�6�����P� ˠ�y��qd�C�ɻ=�4$�J9�Lqq�Հc��C䉬#@�W��4l��1Z`�-k�C��&
#xiI����7���w�F$K�B䉤2jv�I�MT��zո���$�<B�ɗK��+�>&
d%�Ձ��a
�C�:,�̌��!��FI��c��
��C�IU\���t�'8��U�P�Ň�6C�	 �d4�6$��h,� ��.]�C�)� �K�O�9a���`��Y�"O�l��Ϭ<df��0#�9�&�2"OV}{sŋ�4�B]�`H�%V��%"O�`�fԹY,��[�hϝ�� F"O����0��ehM�@i��{�"O�p���R0��ѩ'�u *!Z1"Oĥf	S�Sfk�L�9KJ�U"O��yP�B�+�R`��	52�ȃ"O��3
�#}�PӪ��5�E �"OPq�)�M��U��o˘mטy@s"O��'�UNZ�q����`�S�"O*`�TرU��(Y��2�6##"O�u�S�(!�SF��<���a�"O"�&Ǐ?�`���@ƽ8D"O �+����G�Z1�%lS�[��ؐ�"O.!rĈ��<�P�qa�C�1d�('"O�i�3�?=��adN�G�}�"O����憕SdN�zbN�[��t:e"Oj6�9$$3vF��6ps��<LO�H�秒�K�@��B�Ga���"O�Q��$
� �����gU4�+�"OL���pd5r M��1K��%R����	��p9��\���E:8B�B�2M�&�)І�g3.�h��&�B�8d�Ĺ��&[����ԂO�4)nB�I�:��eY�H�G�U"��w<B�� �r��P�Zj��ZE��w�B�	�zL�$��`
�>��D��޾�B䉼b=��G���%���ؐ`�=!:$C䉽V�<��6�	~�]��P�HC䉴I�%��П)�VT31��%GD�B�gh�]����0<�a�
�\�B�	)E����&"����f���|B�I3eB�Tb$��+�
���Q-83\B�I�"|�TGĹp0p���)@B�	:N��`����.>֕�4�O"_�C��	�r��6�ֈ!POM��B�	�X� ���0��,#" �8��B�Ƀs�аy'�Ƀ�@�̯8t�B䉩t��bf	R���X�"I{��C��)xv���Ū�?�@�ȇ�eB�C�	% �|� V���J�bd �)&��C�	��44�R�S��(H��F�]�fC�I�h^�|I�^�(
n��n�:g�*C��6j�V���@� b�ݽi
j��ȓa�Xؓ�.�(=i�͚���,��ąȓ�و&������ݶ9����)���"�M#;|�`����O���g�5[���i�A��#11�5�ȓV�p`�
�4�nUS�#[6b��X�ȓ9��3 A�aH4�u�D�=� ���B�z|��L�V��K�'?�Ąȓ�H�q��
,I4Z�r�P+{���ȓT�\0vnǙ)3�t�̇;ڤ��x�x�{`�BdT��k����+�p��ȓ	�l�Jfɋ�q L�S�z�����[��YK�
�XJB�X���9�����$�$�+V/_.v�`��"�:fHK2D�$I�fو9�thz��	������<D�\��ܻ9N�A�d���z�TW�8D�غ�ĩ$"ԌĄ»a���I1D����ǟ8jBfT:��@�%����3D����,B�BE�"!��}��P���5D���pf[�p6*�x��B�h�Ҋ/D�� .��&�B	n���"!(�6��"OZ �1O	�Wv���eo��G�Ȣ"O�%�4D��rP<(8e	ѣOҖ�h�"OLyp�[5P���N#t�ڤ�s"O����6+�~=ʡa,K�&��"O"�S%�,��h�`U�s����T"Oڭ�D&@�*�إ��7ҵr�"OR�(a�e�R0YĚ����$"O�`���C��h�#�Ɂ2�*	�"O�8:�'H���Ug٤	H*-�"O�q��)G�	�hy� �1%:� �"O����*�'?���V�L#6j��R�"Op}�$A�/W�h�Z�F[snL�"Oĸ����<}c��P��A8dC`T��"O��)��N/|�ݑ��n�ZH�'"O��3ALR&=�ȕ�pĘ�Q�hm4"O���r�Ф(i��9�c��i�`�*�"O��Ra�� ��u�P��� 0��4���O ���Ћp��2�KP�����'�0-�!�[�R���RЉ�"̲� b�È/!��Z*c^d�7��b)Ʌ.ͅH�!��,ޝ��	K	u��9@�#�36�!�dW-'�||{�E!_��UZdcD�W�!�J���������1�~�!�d��vl]�uj�������Ð���O2���0�Z�����O����T� �!��?R�8����I��@BB�uT!���#T6��3+Q�R0 컧���q�!�$�&ry~���
!.�`��H��5�!�D��<0��(A�&�ZéL��!��Ӫ*{N����wLx(Ƃ�{�!�$��j�-�Da	�e�\ =	��O����`$��pFN>G�6�7瘤u�!�$���Z+���9[����U��!�ěo�:M�a�V-$��#!H��!�$��W��1�'�@�S�d�$�!�ж[�ZMa�7L��@��#�!��ܗd��nM6R��8`v����!��N�(|��e,�(�EƜZt!�dͤe��H�mK���TD
`!�˴b�H4N� ͈ir�Ғd!򄑢3�<q����'#�"Q���.;(!�d�)��"Bj�(?4u�X�:s!�$?!�By�
Ϟ[0���럮x{!򄚖	�&���*�e�j� �
��n!�DB�n�@�E�W���H���u`!��[.~p����� I��� �T�S3!�Ė4��=k�AU���E*mR�{�!����JQi?!�q�MP�!�ݟe�F� �Y�<2����l ��!�Q;.d�!m��2��(ԫ;)�!���B��p[v��E���P�I�a�!�$�{�� D�B�tvfP�D�!�d�bL�pI�L�H&��!��S�n�1@F�+X˾q8pD
�F�!��ߥ~��9�B�{��S��͜l�!��\l
�K%��(u��h�Ə̩�!�K�B���P�e-�����H�!p!�$O�u��X&�V-[�(9#Ǯ�Y!��R�mEb2�f��|+8鴍�:=�!��G�V���r�k&�IeB��E�!�$$r)��Q��?Dd�e�7�!��J�v�N9�b��']$�5�U��I�!�0�� rThD�	(պWcP�B!�� �<��惥XS ��GŇ*(��"OR�P����bD3��8~x� �"O��X'�ܹJ^�
d��y�����"O>\�#�Y.g
�$۳�żH'v���"O�9#HJ�z�lYIA��q�"O�lUK�i�`9,	��9� C�yb��1x�ҕV��6sb�H�t
щ�y�� Ԩs�#W!iR�Ak��@�yR$a��{4�>]������
��y�d�d�)�f�Z'@�ҩ�T�� �yrj�Y�u��@�97FB�Dm_��y��Z5qL� `�֠���a6���y�㛊_`���B� FHH��ք)�yҢ�3m+�<a�@D��H��h�
�y�("t��)
�CP�4^���Ua��y��"fɼ����0��������y2�3h�E����)2H̑R�ڽ�yRk\�-`|�#gT+N�Ċ��/�yr*�Vn�:�ƙ���y�le�\�G�^|�*Ǡ�y�������[!z]�������yRBR�G(~��*��h68A����y�
tq��P*[�cS:�����y����.�����D*�rM�"�y�o�'D4ӠM�==H5
�$�y2��:���ۆK��
�Z�٪�y�	ьI:x!�G�U)q��A*v`���y�"Ь���g[�8�$L��y"N�E�:�s��6c=��4AS+�y�j�;j4x�c�`�ne�Fo��y��A/T����UJ�[9&y;�i��y��Q9$=��8U���W�JÕ]3�y2H߸�zl0�톭P�6�+����y��8-C��H	54�����jC䉅d#h ���
KB
]�񩂉?LC�I�C8����C�x��0Rm�]�FC�+=/n4ӔkC|��((��3��B�	�P[4L�G>�t����&n*�B�6]"���قl� <����Z�|C䉻d�%���ct�}�G��+HlC�	 }$8�b"�X��q9�G� LhC�I"/�� ��^���Ui�
ݍ�4C�ɯ+��1�В���i�Jۖj�C�I�*��(�!�?���C�3��B�	�A܄�I��X���. ��B�	V����L�GqN���㛂�B�ɪ����)�6uZ{0JZ�h;�C�ɵ�Rxb�� �qJl�R׀Y5ZVHC䉯�L0�0
Fj�`��@/�?t]C䉥=ʼ�N˔;�<)k��#I��B��3"�I�%,9�6{�'UB�	.M��5ۥ���'WNxT*3Z�6B�E>>�y��}�2������M,B�)S����U)	������KAO�C�I�U��J�J45N��G�,)8�B�	�<��Г3���8�@��x�BB�ɤ�P
mX�b����*-�nB�I���q�7H���FK�&�|C��.X��
>I�Ჴ��'
�\C�I� t�ic)ݣl��MQ�Ǡ��B䉎~dv��
�0>���7�ʽ|��B��%e�pI���n�&�H��	�N!xB�I�l%���@dB&X����a�2K�jB䉈N��B7@�ƶh�0�Y-zc�B�)� ���@AX�����cY�gz��A"O��q����|`�D� ���"Oڐ���:]X�#!�� pa��"Or-R"L��r����Օ��"OjP���"	��p�e�3G��J�"O4����ŢZ�X�� V�]!pekp"OT-Q6΃k��P� .S�v%ɳ"O��C ���3�:h""�V�Fk ���"O (�KN������hjA�3"O�t9���M��% �K�DU��E"O�uZ!$�$����*J�W>|q�"O�L���$h�N$�D/�"08*�Z�"O^1��H�4m.*���Ώ(v%8��"O�t��_z`;�mW� n5Ca"O��@Ӄ��+�j<��~:J��$�&��0|���A(p��ͱ��]�@e�}�<9!)T�5�M)S. ��&��f��A�<����:x�X�㰠�6e���cP�YS�<i�@D;t��lÝ߄�˅+�Y�<����oų$_�mz�D;�oAS�<	"R&f�z�㍰
ưk1 �M�<����M�*,آH+8�� �
K�<9�˟<h� � �+
�@M. �G�<��)Χ��4�%<k�!�%��E�<!rjP�Tf~�r��G��`aNZi�<іoηV����h��[��9���c�<)u��/+ �Cj������^�<�����*V����[.C�`�� �`�<�d`à1�ay����ы� Hq�<��ѽR��D�-�v�v���^Q�<с��OS��A�a�.=�q��W�<�r��1N��:C��nX��b�ƆS�<��!�0?�MyA��H���g��R�<�R)L5t�{b�W�an ��U	 N�<�g�����@��[�H���JV��_�<I�ρ3�(ٶIH+Fz����GC�<I�g[4IT,�u�٩W��8թY~�<�7+¼y�:��dBQ"J�:��B�<�s�i`|���Q�SV4�A �I|�<� ��:5�*�!R�7����A��x�<A��\D<T�4ǂ9?~:LyG%]q�<��*�9o�@�C��G0�h��g�<y6E��<�2����9��#�~�<��"�7Q�bܓ�Y�6|Q�+�N�<4B�_R�U�H�� _��"�I�<��ϟ;1=��i���H�����]�<�\�8h�2n�0�CUB�<�&�����Ɖ�yڑ�c�@~�<i�LǼUф��$';#FI�G%�b�<�Q'��z�x� ��F�rrX�:�
Z]�<�� ۗeq0���'T���^�<���K/%�b11�!Yh6�"��\�<�AV�]K J��"����1��_�<��G1��Qd��"}b��r�U�<�s�$��UR.��%�vm{�o�R�<�Fǿvf�t�J�!#H����XN�<1!�k����T��1/�]�g�Of�<y�hƟ%�lA��i@�"�vи�(VL�<�i�#�$@3c��,�F(�tD�N�<����Z<L�XǞ�O(|��c�<��ʛu]�
�䄽O�Μ�b��W�<`�OL��R��W5d���G�l�<��My�n�sEV�"<�x2�AC�<��=p0��#�0
L0T�<� �2��fW�Q��Ė|U�0I�"O$�
�J�a����uJ*Ѻ�"O�)�f"�E>��%��K9D���"O��#�V�_� ��!ێ�\ݻ�"Oj�-[�O��F�ב �p���"O�P�V(�M�Eڳ=E�J�94"Or���mC�)���7��=Hή�Ha"O`Y��E�3A�TNܲa�z�A0"OB�1�F��؋���U��:�"O���� �DtC��ƙ�B�"O��yS�}m��0�F����0;U"O�\`�[���[�M�P�B�"O����]Kߔ�@�D�ں�i!"O��3ϓU^����ү3ª�"O��"�GԔ�ce�%�a�"O޴)U���>�s�A���m�6"O�i�5+!TTq��Y`�d��!"O�����΅3#�=��C2�B�`"O^����3ʖ��6�J*�>H�t"O����Q�lH�1��܍W��I;"O�LR"C�v�z1[a	B�f�p"O,J�,V�#!�d��+���X���"O>듦 ?6M ���kU�C�����"OP��ą�2F��E�l��dՆ�P"OX��]�	��p����i�t5;Q"O��Iu�I�6�"Q(�KS���Ȋ�"ORe�4���x�H1k��Ez"O���H�7&�����#ޛZ���"O��׭Y�T�D���I�qmT�"O��6jF�"����.f氢�"Ol�e�P.�d!k�CϽ{]���"O��Ӕ�Ԑw/&X)�c�>)$�0b"OlH:q)הoR��D�S�4�rݸ%"O�5�!�I�+#�hi�֨R��H!�"O��a���-�= 6�28M��"O1��oS�P�.�"w�	�:�4�T"O
|2T`��I|�!�5J��6�+�"O$�;q�Ɩ(�����;����"O��R�N��n�؃q'��^�&tH�"O����Q��A(��Y/1��Y2"O�	i &+���߫>��ố"O\���l��M�XU8*��! �"O��)�*X�T��:]���`"ORq��l��=,0��Ŏb�z���"O@����"{�N��� W rH���"Ob9�r��^=6()�Bֹ&$	Ȓ"O4D��є$����+�
��H �"O�e��n	�K��:��3TLF� �"O�eq���=�K��̢heB�a�"O|a�3DQ�d�,9��#�� q���"O>(J��*IVĒ"Ɉ"p&8x�"O�=�EL��*�ʀ �k׼hܺD"O�5Yf�G$`N�p� A�v��l B"O����c��j/��X�/�1u�څ*&"O��qЭ/C��d�oĤv�A�p"O��y����v��5��YsJ�sb"O^@�/s���y1���<lĀ�"O�Ѹ0��&9�i���0�0\�e"O� �r�[�e�zY8s�̇����"Oa2�肨b�b���o�F(@�"Ofa���ߺ�����U>H/��a�"O��@/�y���@���66jq�S"O������V������5<�ᩃ"O��d�\9V��M��,Z)�h"O� n���Z
o�T؊ċ�/���"O(p!����)r�X.c��̐�"O�(��H�gDL1�I�%,��5�1"OL̊2� �DgԘDH�;`ą�"O�U@'��g�Y��T}�����"O`t�� =W��sqeP�[�$�h�"O^q�"��'U�0�*a�5��@P"O���5��)%cS![3,�d|B�"OfĂ�E��Ah�c���c%l)�"O}@�'M<��H�!oHO���P�"OTٲ�ϝ�I�0ٰC�Q�6D��"O�$���	�{eH$_��@!�"O�%	)�;?�p�ZR�S?lH��"O�	��	7������-I�-�f"O��H��UF��@�-M7X]�"O:y�b�@)~����C*7Ԕ �"O�q� `_"��ir��T��zɁ�"O�R�Z��t*�đ�@T&�"O&�Q!�D(0�N}C�c�u��U��"O0Q�O�6!_b@ʶ�̣	���$"O����Z �0}�G�Җv��P�"Oʌ���fU���Dgu�9X�"O8����U�MM�I��W�X���"O�|��쒶"evl�f� ��TQ#"O��CG��hs8H��%��<�0$P"O:a��gM���/�y���q"O�����G״����K4�P@�"O�}B�Z�RI!8E��R���5"O�ԲgO�	~]���(Xn����T"O��ZE�L	<
�`b�Y޵F"OH �FCߪ4�2e
dlP�C�"O��'�m��BLE�]16lV"O���cn�����5�}Ҁhu"O�e9�k�I`�
3@%P��y�"O|9�ꃏCb E�W`�4:򼵓"O`t`�IU�i$n[�tb�"Oġ�$n��=���J��Rp"O\����*��Y����p�@R�"O��
��~�2����P'���'8n���o6��@��?����'X,�!Ũ^�H��-�f�ɵ8VR�@�';t�`�y�^1c6N�.�l���'����qF��4��aV�̽0�pX�'�,�8cΞ�}c2)�V�%�f���'��h��h�Y:�������Hq�'Q�ɪ�d��{gJ��,��]���!
�'��Q���m��	j"��`�61�'�TEIR���E4X��'�W�F��'�ڠ�sB��3zIصč1K~Ց�'_��0
�/Z�vثŁ�4F��'��r!EQ&s��m�0��y��(	�'�h�hV+E�AD�]C e�*t���{�'�q�&F �D�GeB�eW���'(r��ŋ�|���S����`�j	��'�R���.H�4�b���I�U��j�'F�Ԋ��Ə)�Թp'I�LC�U��'?�tp���d[<����LÖ�8
�'���K�,L�y
q�L;r�l��	�'��l�l��FxHd��
)V]z��
�'��qH�̪Kxv�R��6b��"
�'�r1��f
pF�!kS��gf��
�'�~�Wn��w\��㮓*a�L���'$�8�����n�r��!,���'..�3KM+;���J�,�2f6���� �x�$I�@-���1CA�m�ID"O\���3���%� �:
օ`�"O ��ݿI"�i%��3	�(��"OBx)գN������NL'w�t�6"O$Z�99���J<V���"O~��B��Y�x�;Ak�T�4-�""On�/zY�f�V�r�R��G��$C!���]N��&�ǽ}w��q2��:�!�$�=,r$,�eǑ3V��H2nοx�!���m�4���Q��Qb�Z0"!��ŏ:����n���b�I!�	�!�\T���Ά�N<#k�)[ !��!i+�@����7��X0��K�% !��k��<+��A�W�������k�!��A&�uQ8�`�� hM�nG!�$d���4�
|�6�x"�I�!�ğ>-�u�S)��{�T�8*Ў9�!�$�A���ׄ˞<?<9��jW�!�D�j"$M�!(��e�,�*����!��ڝT�x�(��Bk��ǭ՞*!�d��8��%�ri^����E4!���Qǚ�{b���������;J�!�DѤE���wdٟ$�9y��Ff!�d_./��Aȁ,��M��� !�dN.zh2,(7���
A0K�:-�!��Հ|��M�gC����J���#|�!��P��x ��?�E1��0e!�ۭ�6dh�"��p�,Y�'�?N!���*wH����U�9����j3!�D�o4 ���>2���菀`�!�B�R��u�ܻ	C�Z�k�!��*f��4ab ź�
����Іd�!�d#!����Ɇ�`��̠'-�iX!��ȍ�"e;��u-�UZ@b8'!����"'M�0T�&$H��lv!���v�4�u˓|�`��B��l��Ox�=�������z�~��$
	0C���	D"O ٺ�O�t\��Z3q �!"Oؠ��ə�wEA����"\ܥ��"O���غM�J��b�X#t��"O�<cdA<4lM�gƇ&i�m
�'�����N0y�,S܄r���	�'�ĩy��Mb�9i�m�nҼZ�'��9&�ޜqH6�b*2�a��'����F�430�򂐋*@�i����6�o�	�e�H�0Ձ��j�N܉�"�(��>����,-D�L�t�~�Q�dН{�Op8�͈GNV1
7%�
M��u��O��X��R5'�ʖ�J�Q��y�n�,��'�ў�b�,'N_eY׌�m�h��C�'o2Q�&�/o
��X��9~x3�'��10H�،�u�,h9*�'�lL#&�%m" t�) Q��'��-q5��f�ry�Bi�6I}����'(֙����}�8B3O�C�e��'rҬC/;�Q˛	B>�9��[8�y�o_��`���aϬi��;)��O*�;��#}j �V�V�lZtl0/�N5��J�A�>�S�'FF�01$��2�Ԃ�A*	����/O�O?7�,�΁��[��,��W�U�����ޠ�F�ܫS7��sw'�"Ɣ�'�ўtGxrJ�O�^ܠ'��l���2�l[��y�Ի����h��\҅�ٸ'*ў������@1t�eS�7	|9p���.�S�� ъ�!<�p�kWJ�a��P"O� a��̵,�4��%�^I�� #�x�C�����Ҧ�Z;��
�g�����:$�Ȱ4ĕ/W�.DI����$.X��$�Q,\Ur��'�'o�)�s�x��NL��`�@��Z�7ݒIsA0�`bz�}bugK�a:d����G���jQ��f̓�hO1���h�hO�Z��u�3�H^�z�� �x�eB��Xe�=�~� �6��:F�M-�F�Z�'��y�K"C,�طI)+�:�2�ҙ�p<Y���
%�N�{�jQ�.�حIcE�L�p���'�J�d��iצ�
��<X
�'-nD����6��Ȋ!4����	�'��yXA'L�Őh !&�r��1	�'���p�$�~��0l�>�%%~̓�hO1�T� �o�����F9V���I"O�-�!�Cp]s���33˖�(S�Iox�p����6[�&H3��]ohѹ�o&<\���Q$�$L��O�YG|�q�"k1���Ӡ`+ ��'MZi��߫v�` ��	�<!���˛(���ɧ*Ϻ-�x�E�&)!�dM�z=��AU옃7�p!�#��g�'�ў�>���n	�N0D��ڠI��� L"D�t�$V78ܦ�`r!XN�(��!D�$k��ԏ|���>[P�0�:D�,��[+/h�M�E��7FΥR�	<LOz��J��%C�n\��˦5��Ҥ�V?�!��Q�� �̒)�Ji��*ξM�!�dؙ.�`m�F&L� ���ڡ�A1P�a~2�Ol�c��������3qx`�:2�
f�<C\�b<�(�%�2�$ �cm�m�<)��<Ȝ��2��;*�@��i�<��՟*'�Ii�b�B�I^�'��&��h��\��:���>{���b-D����E��w� !-8��y4
�i�O ��)�x��&%5�n)�Ə�|�bYq�'ғ������3���8v�|G�����-�#=i���O�,��L�G)2��d�D��4�'��OԢ}�A<%q�	��@�A�9\���ɕY��݅��a�f0H�� 48'���fڋo�C�Ʉ,c��(��8��3C�юC�I�Z>}Hf�s+�j!�R�D�.C䉴U�b1u�P�l�9׌C��C�	lL�`�
}tlzҀ@0q>�"�S�O&�!�"\�h��ke��Pq��'�qOn���i�HJ1ʵ�
�m����"O� i�)@6M�Ib0iL]�nԣA"O�!�	͘;�&�!'���S�2(bD�D �S�)B!G���g�i�����X�X��D{��v�!���:(fN0����*̪��{����>deh"�&9e5\yp��v��=E�ܴ�x���,̱L�����(c�rԆȓU��,hE��.�4x��/��DІ�(�$�1��e�(됎X*���)���;G(H�@2� �^R�8Ub#$��
���&x�"�D�Lc���C�#�~�'��)�Cۃ,�HX�R� "/�����(On���B 2��T���N,s<mH�"O���]�w��]�s�]/W#����'3!��_�7=t8AoB�>���`��H�!�D�$_��xmʠ3��y��l˿)q�}�������
�9���@�U�<�؜!�-D��a�%�|����+�n������7D������^L�(3䎁�z�Xa7D���
�R�$��kY�>GZ�;2 4D�� �BΜ7
ոu�FNJ�\�yP�"O6t
s&G�X��	Q4-X%S���P"O��[p���B��� Q���V�OH��D]2z���H�<Vre�e/	�!��ʦBo4qҷ��'����FB7{qO�����
n�:�#]�-�v(�SQ�!򤆪xIriYց��(�DXH�a����^x�������w���G�[@B�e8OPJ��dI�i�d��H�]p���\J�!��\�'����� �	��m��m�1O,�=�|⡁A�U����1��i<���'�I8��$���.ƅ;�,�ЦE�f&���#D��K��7
�y�s�a�0�F�!D��8�l�/
ր�W�K�b�&)A�	?D�Xr�
������$T�B�E����<��'�qO�2
��Q��ν:�>���Ġf���$1���  Q��q��r��i�@�R�9֬����<��OdU�'/@<��t�hPR��<��"O2�0@ I�+1�xcDHQ�:�P*a"O��!��ABtH��,**���!�'��'w�K�j�@��"���JA
�'P2ԑʙ' ����b���m 
�'a�A��E��S��s�hTBH8�
�'�0ɘed���h�'n�3��B�IX	�m�� z�:98RF��Ƥ�����	�Z����Ǖ�{����?q�E�IY�!���7g&�����D��&�����ʁl2��y��ڢ ��u�e;D��Xv�Q
_�|Z��F�QJ�y9ņ�>�I���O���$խ0�ġ�	u� �XPB@�r�!��[�n؎����O��t��#	+9v��:�O�ܨ�$H4}�4x�)ڃL0��� "O 9Q,��r*����&!S��c8��hR�9�vE��Ѻ/��K��!4�����& ,�c�"�e=~�r����x� �R�nQ�q��D��k�h���<a���$"L��1@�4+d�ȳ�ӹO�!��	4јP��B9oI�4����'�:�IR̓i���5�.Y����8d�0�ȓDIB�[�BV"+'n�H�	'V�j�IDO9k1F�,^<2i��KY�B7�4p�"Oր�6��0�R �b�S�����"Ob �M
�5��\HQL3R��U $"OH�0e��btF(��(Y: ��|�c"O��h�+�0/�Ѐ��%8Y�`]�"O�M��jƠ7�Z�S@��.��%A0"ObES�$ۖ O��БL��/�U� "O(�Kd�:R�#$L���,��s"Oʬ���C[���,]���@�"OR,P0)y5nU K�!=Խ�C"Op!S�(�Q��UA���~�#A"OdMh&fZ�$�8Ep��9��Ѻ�"O�}iѧ߽f�0� ��1N��ZD"O�a�7�Z�x���{�lM9�Y�"O<�Bu���"��|�P+X�4��1��"O�-˶���,(��#K�8"s.u�P"O��YG�D-T`J�j?*r����"OzI���ߦBwR���Hęo.���"Oxt�A��%HX�!0����Ya&��"O�r��΍0֒���@�s1�<0b"O�L�/ݶD�tY���^�@B"O�mqP`ŕ�~�	� �Lv�yP"O"Y��iʜ@�FJ�X�0�T"O  �&xY��߶�X}:�"O� ��U	�&1X`˗ǒ#M�v �"O88IS+��v>"�0�fI��,U0�"O�9"V��N��u)$Gº8�F$�V"OF 9�d�<v���@[:7�FY�"O 4*�+�1�2���ԕc_�4�"O�5 ��#?�:	��B�S*�Xq"O�%P�	�?`��(��A.�`۷"OZy)� �g�<�p��)`����!"O��J�D�.	��`A��5n[�="u"O���GU'xPV �B�W��"O�U"p��Rz8�H oRD��2�"Ol8��K
�A.��IQ�:r��A��"O��(����5S��D�t��|�"O�9)$A��0�b'I�p���{�"O0ђ�̐�M�<�l]�p�0"O��P��U�M�����+�����"O^�Ԩ�3<�hY�$(���Z�"OX�82%V��T�q�C�(���(D"O��G�5�%I�ȊY�v# "O�t�$�O�4�l��NI}��#"OFa�TO�@��DIc�+ `���"O�Z�  ��iU�b޶� f&�	\!�S�)r�� ���%�����>}!�d�2cA�T�%.�
C�B$�a�?!��Hm٦Lxp�<`�F�{���!�ד'"�PsH�Wݜ��b監Z�!�D��Ag� *  ������ �j !�$�y�tz�N8��Yo@š�1l�A��Ӹo8��(�n��y⡉9Y�y7YW�mѣ�yB�]B�L
�C��e�� �=�y"c12"h���0,,���e��y2a:7��ȹD��'9������y���m�8���-������yb&˽�jM5M�<1:��f���yb뉽^4��H]
,S.������y��7]��4��D�1^�Bh�P%�y�ET>-l,PȖÅQFI�g�G5�yro֪Z>����'I�z��ŉ�3�yr�ޣ.���l�%�� BE�E�y��.5lP�Ƈ��$�,��7�,QJ:�B�F����h��ߨ|��92�k� &�,�C�O�!�$K	F
�:lD�8����zH�ݴF���-�E�r��	$��ze`�!�`�	�f+JE�z�8r��J%�ƭ�~��Ԣ��F�(KalH��y�#����jg.�B�2��B2˸'��3�a�l�f铯6�`���oZ
]��$��bA�7��B�I�[��B �I�GD�h�!"6��څ��#ʒ k,O���Y�@��mµjI>��bd��%�&C)D�8�e��E�@q�ʧwFT�� �Y�D5 �D���hj�^�H�A��>�����¯*춱��*9�l��0+�h�r�oڻ������M'	�����z.�s�<��j�v���N���+���Kܓ{L���t��$Q���`���`�`r��1et��˦�T��!�d%+�4����&< :ʓi�]�L��� 9K�i�'er1G�,O����ƌ"�R�JЯS�����"O����H��fQ�14���P`���Q�i�9���J!��Q��I��(��Si�B��a�g@W�i���d��zp���&|�c������#"/�>i�)��O&D�,C�~��K%�Q�@�N��dj$D�� D�Ρ]Y���N�<���O�ʵeZ* �&�O?ա� �9E�����* �t�>Ա�O�h�<Q0d�#E�2l��>#><=H��l}�![�r��١�Bx���"��9���%�"����@.:�O���V+�8k>��� ���r�.W�j���O��R�8䀑�LlH<� !4���3�EIےiD�Xn�'ւ���@�#1�������(��L� � LQbhiWI�>�!��ȲHx�R1[�7<t�󓆗�;q�$��"��*���yy���'(MX�@E�+�,[@/kKX�<�j�`���DWN'(	��N?�ՠ�5!��LZ�H̰<A��44�峳�N�,5��� �HE8�܀b��$ȱ�S��%v��2��v��@�4�Y�ē�nDb��ݗ):��
!���m��EyB!���zl2�\�+8��M�,AU�آ�Y<|Xl1�"O�\1�R�[p��Cs���]R,��I,?�+��<E���)� $���4���5*��v�Ʌ�T���@c�[�Z�d���"���'�6Ųv˗�:`D���	?v]�H�e�5I3.�Bs�C���������s��m�`�ե֬U�N� ���Cf�C�	s�� �$�تښ9�� 8�C�I~��(P��}���вq�x�)܌�	�n���R�x��צ�F�ء��I�{j�B$\�غ�IV478�.U/aDN�Z�%D��Kg#G�rtP��(���9Ԧ �ɾ>��<���:z2�M3̟�v�)��.ɪ�t�^42���P*^X�H���$t~4�R�Y�bt~��6b@<��Qb�{r0�$���I��H�R��kM6�~bÒ[�Hl���[�"ʒ��l��y�e��Q����/��&tLx�ǠS<�?e�
+�n�Xg�6|6�[����?��O&vHp�瀳~z���
?��d��I�Au�͉�E�\��9�& M>���-�,��ÅT�"�x�R�|����N���� �o��4k$���>x����U��3�.'���K��P�l���E7$�`��h{��U(/8�5�t�Wyu�9�h 7}哌_I���̜����H1��^����X��؅�ahڎT�h���]�*��!��3D3b���C�m�<������Ǽn�2����.���A�B;jĻ�ꂘl�>東<^���%N�{��1°k^0F���Dކ1E�/Z�jQ"!�N�P���x#�U�l���S�@�$��8[EJ[�7�P��fOʺApQ:Q�'���(S�T�j�{�0��ʁ�H!`92M)���;庄����>�z�2ٌIY�(ДG:)��� S6�	�����H
��v��8��
i 1��O�-PW@[��6!���|�=�@]�	�����L�8U<������䦭{�z[��rg
F�7��T�� 8���ge�)��Iү�T���C��11���jZ1D��
g#�>N;�q!c��B����D�03,��J@(
���#/��a�sc�H��*M�P��6�Hza6���z ���`�O $�~�F�l}���t�S�Y2���u���p>YV+�$P㾈A���#j�
�)��x�\=i$�	;Jh�f���A��L��(�D�@������Ğ�UI�K"e���te��DM@1���J�J�4i��(O@Q&�� @GV�"�!N�F�*d��fS�<`�`î.Ghj'�w�����֖g2�o��,�u�F$4>�8A`I������#Xpxl#�����4��,n��(�U��$5?�Ͽ+�C�/����ҕD2flKAB�m�<Q�(Ʋs%��)��<0I�MK�N&�h<#W�Zp��[S�#�"H�'�HO��(7+[�z᳠(�38�2z�'��4� ��&x5��r�jȴ{�2�Hqj�4|ր�Gg\�!��d�����a}�6r
Kŗ%��d�C,hаEy�fr ���Д#��@�v��i�S I�����
a�ݪ"V�h��B䉊F�0�Y��Z�B�te�&�A�Z�֨`�h��ay4,�ik��
�h����5dA�s����P,jݸ�k�)�y��)y����'g6�؀Wꐃ4+j����ɑ1��aJ�}�p����@�q#�& t���,Ta���*B,+�OPA�$ؗk4~�8VH�#^�����C~��q��P��M�#DK�5�}�ș*gQD�1�Y +֐�T�+�hON,R�j��r�Xvh�4&5 �'W�����ݑJ����&ɜϒe��y|!��'�� �(5�$�_�B	�I"{� P*Mw�U�Qm�@�O�b�:0�!&���2I	�;�<�"w"O���/�)eڄ�;"h	=�H2�l
��~2�]�@p�X�!�R����� e�t쑁��?��J�ы.wl����@ɬ���������&)$	W蹹c(��/������6T�ܣM�
�hH���ax≚�m�T�=IP��;���Cޢ��}k���B�<�&h���t�Y��ܚ�r��J}�<ِ��e����T��:��8��+Tl�<A�k�Iy���b��!Mt����L�i�<� >DЂ�̤?=�@8����~�U"O�A��O���+��p<t1�AE�l�����Ox<rc��R�R� �҃yu�y3T"O"E���I�Ro�(+�*A��H�2�>O��	�&ϳp����B	z�z��� �U��d�E&)�{�,X�}"��ɦ�#A��Ayz�r %U�z�J�
,#D�``P�O!0q$���
 ,�$�!���G�4�`�Ϟ@b�>	Y@�I�I� �҆���Gf#���` ��i��@'ȭya��(�hA֍�x��Y�ݙB��O8�}�exz�i�F\")�d�E�Wc` x�G�TnqO�}��_ՠ����Z:Hq*ĩȯk�Ե���{<���e��&@�a{R��(TT�X`H�,��D��,�	�?Ye Č �>��8�����|Ӥ	���+ra���"F�W0�h��'fj����g}2�X
0�,��D���"��@������'2� �/G�fQD�$M�pZ���ń�/'�����!K���'Q8Lq��Zj�OVhYݥ!���Ao��W��+A%�V��E�1b=}B��PS/?�Zu`l��F�	�Ξ�6���È{B���MK3ym�EW�� t�fE��k�0����s�.	��I�e�H�P�R#62������Vn�	�.=�቗E��2`3O��u 
Q9��ƍA!�*1"O�IH�Bܙo-���"M�r�
��"O��h��4r)zU��E6��"O������P�9���P%ڭ�"Oh�adM�n�,k�KI�q3"Ot�k��2QT���U=.		P�"O�����Q�N��G�([�m8�"O:��虸Fш��ǂ�'����P"O�t�7EԾn����\"�� j�'@�����ff�Ɇe�j$��H�'*�t�1A]�l�^�)��?S����'0J���L�2��HF�e�����o�~�I<)���;g�	9 �iȘ:D�]�<�U �G<��$UlXb��XF�m] Zä8�)��\� P��aP?z0A��[	A�B�I�)�T�c�֪�0�sK�2���䍘Y>�S8,AD�Ǧ�:�����97��d1TvGζH�m`0$�;��ycf#�dp����Ťg��L�`��{�(����a�az�L?
f�O�e��g�^��"���jS�4ڠ"O�l�^�G���E
?G����DT�<@���{���'�k�f�Y2&E�$�i��յ�ycP#g�a����%&%��˞�}2�Ћ��<aUa�#S��3��5�{Pw�<y�i�)v\i��M�:K�V�p Z�<��c�VX�)�5T4���T�<vNf�A�ɰn8:qtcP�<�'nTL�Q؂	��v�Z��e$�Q�<�hΒ8F�D���	~B�XJu��W�<a��8|�0�8��w�:�BV M�<�FI�B��aB��tC�Uja�a�<���K�>��u�q*�)l��Ka��Z�<��n��a�P���)|]؜�e��M�<i���E>D<�2l�?��m�/]f�<�f��m���PT'W=9��*��k�<�" ����㦊F"28k�z�<��Ή"l(Z]Z���t��b�w�<���ɬj�J3�9ݐ=�4GH�<��j1>�=("�K�lp�KG�<9�n��H̰�O���kf$�A�<����/z�����1+e����}�<�	Y*�6�����6�5I�V�<�3	��Cp�(�Qۿ/���(�Sk�<���X�U��@�YW<��rN�~�<!�AM]wx��	ĨT
2`�R�<� ��Rqe¶��CN���@"O�0���1x &J��ڱ��"O�=X�`_�$H�+P��8�"O@iKw	D+;�4x�@
</�(YIp"O�A�C�9-�� 8!���
�+"Ob�aT@;ϐ9�s���P����"O��ʧBI+<DCU�MO$��b"O�q2�o��jH6 ۝`j�*�"O�z���7$��LcD��\	�V"O�!�!C t���⑳b$��"O&�y��#P�9���4���T"Oʄ��Q� Hs�Q&#�Ll"O�ؒb�]/P��h&1�B��"O��ɀ�j$l����A�Z�t"O"�9���/�M���F�c�$ٗ"O���0�!;I��3uJ�?]����"O���,��iX~���)8�Б"O��вj�R�(!⇇9H�3 "Oڌ�D��_�
��Vƅ��V<�7"Op�j�(I�!}�*%�B$l&�T��"O�����������l yط"O�xv- �m�ff�"'ŲW"O�$P����{F� ��Ä!�X�`"OdBv������^, r8f"O.L	��T��~�."Vv�XPS"O�X���2I�z�C7	b�|*�"OJ�X�dZ,b�:	ԍ� F�ѩ�"Ozi����^��iSmG�	���"O�ԙuj��V�t a��_&��3�"O�-��%:~�bq�T1<6f�"O�!��wY�Ͱ%'K�Zq�hK"O���A ��_���FT ��<��"O�Pj���.|R9�ৌӲ��`"O�AKv揯
����V#�VQ8a[r"Of����
�3�蹐���qW�<(�"Oڄ�F�msX����N���"O8E��O�\4R��,N����"Oj9�E�V��$�����<a�"OJ�J��}�	�0-�=˰�
f"O89�!��"3�]��T1cĜ�"O@�!��2G��H�6�\�$�:|��"O��1��ʑ<J�b�G�mf��@"O>L���DJP�5O̹\t� "O44��j՛X��1��eS�+L���"O����У2�)�r��3i����C
5:C�|����#Eȶ�b��ķH�l(0�$D�����*2�$����>~��9�RDl��trf�x:��ߓFu�u����:����۔Z�\��I,~0p��FEֵR�m�м3���rx����0��B�ɉPF�Т�努W��}��I�$��XI��y�Z�r��U�O�Z�O��Zae�S�^�C�'�P�C�1a�.is�i
~~i�S�D#?��8+���<���/�gy2$M$sn4E�D�0J�����#�5�yꄃ_�|�\�}�����Դn�J,��!40���J/lO� �"2!-��B�t�|����'�4�Ӑ�(� e"�i�E@�D�<���R�Ϗ�xthQ��'P����Uqm�4�]8dR�h�{®�6#v���`�=u��>Us�T�y�@i�$�'���	sm/D��y�.;|�� G�8����Am��̬��I� ��5�(���n`���AbĄp���0�W��dC�ɺR�p%�B�Km$�@�/P�*�6��*�D� )��=9��ȹ{�`|r����en��a�c�u��LH�f�W;�]�E��;�̐;T� 4�����4��Q�҄��"m�3&��й��S�? 1xu/4SNA�S.�
J8T2�'F��R���;�ɧ�����5(]��Hh2��21x:`�a9D�� �
�*Or]P҃ϓf<�%�G�>��k�y� �!1<O]i!��8x�ޠ�`�=�!���'c�3���DPVܠ�OW'b>43�N_�h���x�FU{�!�D�2klj� �/� a�=�Q��qM0	aD*���z�' ���&�[�yԚI�eN��c�v���*%�\��!�1,�%��[�:�P�rb�=�(� ��3N��)�������|O ��oE -��f%D���/�y�|�xD�G�z��奟����Š-0�Up�˟~X�����M���1#΅�anH3��5�ON���M�Q<���' L�HEUP3�����dM-&A��'��E�M�./���ꓨ��u1��X`��m�#�,,��b?��e�K�.Z$l2��Ϡ?���ӌ(D� �# �'�Y�L�޸Ã��< X�I⁎���2(O?�d�$^�ZH���=/h؅¯+A�!�d�ML�����3[DR�F������r��3i6�y2A�+"��L���<(M����W#��>����#u��*"�ώ&;����!��3%���y�݁<PA�JO�:�`D��y�D�}��A����To(Q5�ז�yrO�z����� e�P�e��y�I�o }�����d�+u�;�y"nI;K���*e"	��,�ٔl��Px��� ,n���;)D�Z����F�Fi⢆�Z����R�'A�"D[�e��}KD_N8�DXÓ ��9�o�"`��d����%
EU*�X��j�nc1s��*D�C�D	kT$8���-t*��5+,-B��ΟJ{pp�#IX'K��#������V���Ի1<�#׫�	=Aڕ��0>�Q��/F�(�i3J��i��]0� pp� �T*Y�Ne��_�������X����շk���g�~�hHtmG�U����F��$X�A�OtM�͌'I(����o�����p�����IJ�z,�b�a�T��RеG�<��F�ʓL*�p���)�����ʾtȅ)T#
#>YkAn��0� �ʅX�R���t���Oȴh�E�U $(a3ю����N�c=Z�⥈\H��:��8���34U���@L(����-�:�|;Nߑ�8u�2k^�K��3ǳ#��%�@,�ǟܐdm;�d kb�_�|2fNI�.��pqGˈ~�4[GUV�'_�\�cmE)%���Q^��+e��?ݪ}��"T9/�tʦ�I<Rm�S�[.ҢΦhP�qѤ#T=��3�	.Hzh�iH����@VF5˓ �DL(P��Zx� ���$Pz2H���)��,NthB�� 8��|@��C�7�dq�q�S�w�ȹ�HK�V<��D�i�����VS�� �jݠfqn�ѶHσk�~�`*Kf��=:f7��ؖHQ��(iV
\#�~R����*a-^�M>������?	m��^գ�K�$���	��O��je;GmԿY�>9s��s���j0LV6r�D˓sfȥ�c�A0X���(y�����K2N#����i��s���?��"-t�,�G�'{����f�^�}ڰ�2(�o��E�PE�4 s��R�M�A(<� ѭI�Z
�KM(hJ\Q1c�Ojy"hD/6��5A�́?�|	Xd+��W�F��~���:.7�����B�����.�Y�<�����P1K�N:b2n�䈂���b0f��U�g�v�
��JG�	�X��ԡ�� ��D��F���W���r����tm��u)*�XBh�,x�jC�	2R���c�m�#�-{'&S6�C�ɭ7�P���G:]��A����8n�C�2fĥ)v��;;jN���K!r԰B�	0,d 8 F%ܫc����6��1bZTB�	(W*�ѐ�B�P݌�7k�*d��C�I.yJ�A� �JPE���ğIcC䉐-�*X(�g@�%�6U��4��B��?��Ѣ�����R�^	��B�	%m4p�)���>c�ؑq�݁�LC��(K����!9?,�ZH��SdC�	1J��1+�1jw�\R�o���hC�	 �x���"�I��
�L�!��B�	�Z��2Gm�aF<4���=J�$B�I�c~X܃�Lz�B�b�
�W'6B�I�o=9᥎��t�K�
G���C�)� 6<iP��w|C鈷T5��i�"O���r�\7�6p8!)[=s86�Q%"O�áN�*,�T�ƏYC��"O�|+��R�RwH�QZ�C��c�"O\I	bR�&�6%���04�11"O"�b0��P��X�kǂB�]��)�)*�����O�]��j@v��Тi�!?��e��"O���Z�,�j	@�b��w��p�0O����V($���Z*�HػP%��PLjR&D�1��{bA��%bL�(3���8�i�<2�(�W��0u�Ҹ��g%D�����0f䮡`�����p� �ɗ@>90�,s��Ɂ?1^-��K"8�$�Q�N�j�!�ě�EBm��˾(S��Fb�:?��D�Յ(Z��Oz�}����X�`��r~�0u�I	O��ȓ,�f�{ЦاK�9x���d��I;j�M�tAXE�a{�lS�z�P-c�ρ���d�` ����=�`o�	
��P�,sӔ��U��U��ÕB?M�q�V"O��`�f#~}�3=�2��`�dY�0�A	�H��s0$	�bĥ�e���N�І"O>�
�HG?PN]�&b�y����C��z�P��U�$6�g?�5k�����Z����A�2x��Ke�<YINX�hbƭ��-�����<���ϧd����
�i�P��r( Z��X����*shh���>�ı�1O�!"�F��������R"Oz|� �V2Gw��1fɎ~�4� "O:\�C�O�d���5�[���`��"O>m���\�̚�(�Ă�1�9 S"Ofqha?[p4��"�{7dRR"OFMSEiӌ+��Țt��1A=��;�"O�����^3-��p�p@�+�0��F"O^���f��"q����Mѧ�y*�"O~�*Z
Ep� eW&H��"OF$ꃆ��06`�� �:_�& h�"Oʹ�ѡܳ]��8�.,[L��#"Ov��?�D�1e�<&1�q�"O C��B.�s���%_ͬ��"O�A�"n�.��i��54�V�I�"O�T��>�nܰSLGL �"O:ѓ�)P�i^Q��ɍ�9�v*�"O�`{S[�16��bF?����"O��8�J�6LH���	 �Ȁ:2"O��@�E6���g�݃/�jl��"O`Ĩ!��114������}��,h�"O���RP�*��)�!u�L�t"O�m�F̎0n<�uf�{kZ �"OvŻc�V6�\{f�����2W"O���M�>q�Y�b�ђ!�<��a"O(Xf�J9h��5�:�,3"O�5�u�	j�V)���)&:P%"O��`pfıE4dx���kϖ��&"O���dA�7���2�]0(�\�1w"O��v�h��Ѓ'#U��ҕ� "O�E��I�<{�)"U/-�TLs`"OP {���j��  `��Fp�9�"O,=�ׂϘ9�8xiW�@Bur���"O�d'��	ؖ�rP?Hij�b6"O�i�ᡃkW���2Ͷ��G"O�P	�N��N�t�q�W�I��h`"Of R��	�&z�	3��F�{�
��"O�aV�ɢ��PH� ���K�"O�E2CJW�>�xm���.Gw��"O����Fބ/���UIֲ1s\i��"O \ʔ	
^�n�CRj�j1"O�L��C"|��L��C�3Rnu�1"O� ,��i�=u�Z��B�=xZ*}H�"Ov���L��58ș�ƇoO>=�2"O��3T�Ќ5>J�#�)/%<���"O��aj��	�Ti�ǈȖN��<�"Od	b7�L,p"��ѧ�ܕtz �W"O�yђM�����c���+j�X�"O�����^&�`c��x0N�q@"O�5��B��Q< �Z&�ӅM"d�Z"O����+��\ǨtzV��/'*ijs"O��J�T�2'����^�!�xz1"O���̊�	�h�q���/P6Y�"O6aS1�Nm�&qw
ߑA\ђc"O2���:FܱahD�L0��"OMR��=k�܊6�J�j�v@�"O8M��,�p�5��E��"ɸ�"O�H���D�Ei�JG�.�be+Q"O���A�oi��e�N��`�
6"O�D��Ò��8I�C� eT	��"O�e����4��PbDl�sEnYbv"O�u�	O0Cz�|�%��'J�	(V"OH���[�m;��h�%L�Y8lЪ�"O�,!e��\����Ć/GZɹ"O�܈2��F�t�R�#;.��a�"O���!I��u�8���ßg/����"O��9� �\�L��O�)+,a "O� �p�p)H7I�m �:�"Ol2�GG�^2�Є�G���HC"O�lJ��I�8¬43���i����&�&$~���
�s~�$��(���Ӗ-&��8�]�䬐��ϱ:��i�r��c;���-O�<�O|"47O���Ov��D拪+�&|+td
>�&��AOe���')� �D�?��Ģ��Xv�k�c��)r�����ZA�u���s>	S'�D<5@����=d�nuѶK3}2iC#{ɠ��Mצ��H����Q3@�4�����B��@�O����G��T�>%?�'B$�F0f�1q�%D>?�$�b�4D��� �⌵&o���/O�?��R�A;��u��ػ^��<���/+d��`
����L&�)"ҧ`��M2Ԍ��+$ ��P-�;T�ulZ9I��$�O�����O��sӘ�6��(�VA��d���B��i�Y���(�TO�?�R��<�H�if��4j�B��J�+��I�s�$�ĕU>��QlY�G�- �G�����I��Ĕc�ā�i*�Zȹ��Nܪòh;H�x��V���5�p$��A�Z>FL��Ș���� <`���]�a��䜶n�#�H�a�+�kq�Qf"�"�4�HDK���y_�e'�(�Ak�D���çU�4�7.Ջ~�@U�擄jF�Xe 	3~�P���* m�)�' �~���Z��n�{���;
{L���ǘo��a�Y��9��OlZ��ԃ�u�x8�S��r�Y��'����d #y�{�&�
k��m �'�
q���[�Oʨ=a�� �f!j��
�'�F�j%�-�h���IQ�Q���y�'�" Z&�[?x@C�g�'z)�s�'�,���U�7�|\�L]/R�y�'y�4�"kCo6z�;�NM����'/���W����dAfE�0,��'jvP�,�0s�0qq��N�e8^H8�'�R��0}�~��g�ۼJ�p��'�: �%f�58<�a�O�T���r�'�����Ί�U�=Y�D�����'>��.�`�h�ɽ>��4Z	�'��ٙ��9��13��	8;���'�^0 �@�#����࡜8-��U*�'E�bH.)WΠ1�	�8M>��'gx�	Gn̶$V�i������Y�'�&t���͞E���dIΠ��A��'�,���ZFU:X��!̄����
�'On j$*!%4չ�N�LPҼ��� �� ��� _��*P�9{����"OP��3��Y�Z��f�U	z�� 0"OzM�4D��?8<�\T��*�"O��k6��`�MBc�ͅPJ�D�"OJq)��;=���/;p,�X�"O�!��7~hi3�n �yH�"Or�C� I����S.D�i�l��"O��Cfj�9_,ez��j�>���"O�jE��o�V�C�
K>�zS"O�ሃdȆ?��8�䘍Q��-i!"OBD���ߤP1��aj�-,~�HÓ"O޹�t�D>g����:zk�(0"O �2�Һ�&�P�oMV4|��"O�PD'ؒo�`@	�n��80�Z"O��B��Zm|x�!��#Н�"ORE�U�ћ1�ތ��J̲�6���"O"���h��k���:�L 5R���"O�A���w�A*�o=�0��"Odl�4`I}
��
��y(Z0��"O�1ˆ��`�����B	h22�z "OD�cu�ځ-��4 0aґJ<`�"OnY�D�/�V��בr
:D�`"O��X��\�	�ҁ���(p   �"O�-[`�݅a��2�J氨s"O���6��*c_��p5J�)���P"O����9�l q0jv]P�"O�5A��$JO�Iqc�!dZ���0"O�1¶Ҷbg�,��A�$\I�\ˤ"OD0�A�S��� ���]5��z�"O"ic�I�1 �Y�,�,�m�B"O���X�M��i��i�3av�4xf"O
����;@ob���G /l\ր��"O� *�d�Y��F���<��mQS"O��V$Z*��B���v@J�"O��!�Oӗr��������l3va� "O����Kb� @�ŉ�%yJ�� "O�,�PI����HՉ�EbXQ��"Oĭ�f/�6{��5s�Yd)N;�"O�|s�RI�R�P0A"��"OJ�9�&��P��4"Q�+ x3G"O�}k`�R�RU*�!�;���#Q"O�=�dC	_PT	S%;4����"O�$���١l
�%2�̿A&U��"O*d¶�Q3Ҕ�"`�>&�=IP"O�I{G�3�q��;! ��r�"Or��GHV:��B�Ǻ'��A�"O��5I8e�Z�3��~�,\�"Ol�� ���
\z���9���	�"O��!�ǹs�>�9w�H^J�Ū'"O��@ĳo#ؼ@�
^C�$��"O��b0�W;��p��w}.(�D"O@��"�ɒr��!��3_Z�M�C"O�`Y0�%[{����$o���Q@.D�p1��СM�|�a�C��b3����/D����A� Űg�B�I��{%c9D����ə!H/`��pg
$�DYa��8D�\ڳLE^
�|�tF�"E��
�*"D�d�2���7��$� )U����("D��Q�]?j!�WD"j�%x�.D���cc��h���Ui����d+��,D���gC�+y�4SA�v�[$,D� 0%ɟYApD���٭Bt2}�s/=D���5*�qy�Ī��53���*Ӂ(D�x�5��lp�MyЇ0M �ZW�8D�� ʥj���Eo.�s�%J�8<�"O<x���1"�aA�
��9��qpq"Oa�C˝�o�FD+�AR�"ܣ�"O��3�.N�Qp��� 6.$Ч"O>��lO�@���6 H��)�"O}6�Ia
��!��/�JA��"O�\�kɡkG��2ӦɴCKb�{s"O2]V���L���$UK��I "O�Ƅ�F������;e��}D"O��1�M5�*�Ǥ[m*]��"O>�h�ص?�X�9���!-x��h�"Of,I��@h����#-\L\��"O$��`�%E�@;��уpH�D�!"On,�UhZ�kC��H�ƕ�n6��"O�Hq ��;s,���E��k$�j�"O��[dC�ݠ,!�@\��r�"O�2$��eI���p�T�$��QCC"O��ҳ��*�͚wɔ�d4�<j�"O,�ZN*ea^a�����=��Q�"O�t�S�vyf��牖�{�V�C"OPPЇ��H���R/�v��"O�z���^�)�w�ǀf'��
"O�
�H*���c�b	z2��@"O�u!$��!g<���G��t��e"O��(T ^�t����o͉1��h�"O ̣��,�8$N׭&�H��t"O~��$E�-+��K��_�?�	��"O"�8�)�)8a�b7�΃p:�Q""O*�C�A�=�48�D�;B� �"Ox�J�B�2
�N����t��YC"OƐ�W?(@>\Z�ޤ�l��y�F�h�!�ԋYC:84
@�y���4?������W�MCS悫�yr	C�$��˴c����]��윸�y��'�d(���^��uz�ꇝ!�D�P��i�W��]Z~�(�	�!�$߂ �����D�##Q@��)_!�G�,U�]"t�D��l��EJ��T!�Q!���`ĩ��L�Ԥ�b.9�!�dڈ&)Hsҏ-I���;�&{�!�ː֘0r f�n&�%#�OD�!�$S$+��P��V�F|�5P�Ͽ8�!�$ƬJu��k���Q[��pD��9m�!�$�-�p] �HDZ��!��bH~P۳f�P1��8P  pg!��= 8ᓆ!�2� �R�"k!�$Z�f�%�N�g����Q��@	!�$���Ȅ�FªP�\�s&��76#!�$F�4�\[�ז����ԇS�!�$A�gL	�Iܩ/������G�{�!�ė
o&��s,h{��)b��!�d��S�F�b��`���d!�K����#jO���\�� �>y�!�Ě�O4�m�$u��hT
Ǭ$�!�H;Z�(�:�eA�-k���ܞ-�!���o���@T�oL�k� 
xq!��"Y��	�#��7����,f!�D5��q��D�H6�%�GW�N[!���5Wx�
�J1?lH�e�V!�V�'fڕ�,�=sPt��n�,�!�ǼD9,�AnR�7���g�>�!�Dڅ8-A
�Y�B��%��x�!�$�?j��I+���L�$�� �ݘfp!��ҺH>���C/z��ɕ�_k!�� ����ՆOJH�A���<OL �"OXZ�؍+�5�&T�#(���"O��z�`
�~#D�#�$�`¬�z "O�L�a��Ǣ<�g��d�ޙ
%"Oĵ�G����P�9�00��q��"O�hc6/�?1����J�Y�҅2�"Op]��/�0���#c)˶ELt�s"O8����ԉ|{b `��V�9S��Z�'�R���F��T�:Q1'L��$e(�
�'Y��z�/V!p�NT��hZ�!���'�DEbwV�4�H0��♺D�RD��'�����\�s�L���H� Dz�'��bQ,ע��1Q���x���x�'�h��(B���F�C��h0�'�6��REf���g/�k>��'��Ŋ϶D�� ���ҁw��@	�'���Ԃ	גYQ��Y/��T��'���Q�+=a��X�.W�+n��
�'Z�|sDf��s��hß.r*�	
�'�~��#ڸ57Fp��#� dR�X��'�%�&#�:27��S��_S�-��'O���n]��@j�!Ef)�"O>͋G�Dm�i��dM!p����'"OFL@�b�=B�`��f�� ~^�&"OLuHP�0���$Y�\�k�'r
����փ
�����(�	�'H�ܨ��E�#g8(Q�Mc�����'���-ـ_�Ѻc$mӪ��"O���ӥT6����D�{��("O�X��-Y�I����E�W� �H"O���a��C�4,ӃN�a��(u"O�(�@*�C'��z�L�HW�H��"O:�p�(U;nJzQ�֯�14Z�=�T"O�P����43�p:��/X����"OH�OH?CF�@9��O�VT. PS"O��s`�>U�ԣf�\�B�� �"O,�Su��=+̪�@�S��3!"OX���4p�T�Au 8Z͈�"O��aLQ�V�tYqM�=��R"OJ��K)�6Y!q��|�
1@�"O �I�P0H ,8;�Ӑ:S:M�"Oν0EN������^T�8��"O���A�'&!����i�9m`U"O�,�Ge�vH�����^�PȆ"O��Rg㗭����x�$�u"Oɱ֢�'H�4A�c�����"O"�A� �5 �*AH�ݖO���A�"O�I��͛hNx���K?���6"On]c�	   ��     K  �    +  �6  �B  N  ^Z  -f  �q  4}  e�  O�  ��  �  ׵  x�  ��  ��  !�  q�  ��  ��  ;�  ��  <�  �  : � ; � "! s' �- 4 ; �A H sR <\ b �k �t | B� �� S�  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O��jg�=Pz�Aa`�#�h��!\��̇��#=B8#���fB8%pS��H�����fȉ'�$!q!c�	^+F b�ǂ!3�v|��'��EK%�ݵXF|ԲBER�/�f�ٌ��#�
ّ���5�`��'c�6vH��C$"Ox}e��N&}A�A�3Z`X�"OJi1�Hճ,U��I�	� 4Ft��"O�D�tkI:��͠�(A�Iddi��eOuH<YS@҂+2��p�T�w޵����h��\�>y���BdlcL
�g?x<����d�<7�5�)�늁yD	�`��J�<�"]2����ܿf:����G�q�<I&��d�ɓq�:Ρ����X�<񥮀�8TΩ���y\^P3�N_�<	BdJcV�����P2.�"�J�,�v�<i��1i��#P��,+=hR ]q�<���	4M\���#���:�����o�<i���3ZJ���5Y�%ԞU��g	h�<i�-
�Z����&��U@�ɱF�DM�<����+�|�h�O��i�ʤY�h�K�<����u�
� R?
Kv ça�<���.-���4��*��ZVŀY�<��ꈍ[����Se��e:��Q�<�%��$f��F�S�r��TeXX�<��(g��K�GįDlz�iU��P�<�w(]�>c�r!�*8`9K�"O���T�W���!G�Q�R-�"OHXB�X( �i#B��)^i"O"5K!h�5��В��+B
p�Ia"O��Y�Xr�-���,�ِQ"O���j�"�U��-�~��"O&���Ǚ7�l��t,�V (�"O�a 2]`��:G���ya]�&"O2K��ƹEέ�F�� F��QS"O�%�⋖�s�J�y"nԵ'��ۣ"O�Yk��z��i�`�@�p��"ODY�̙<RE��NK�l/2!��"OJ�jv�۽;�P;"�̼#j�P"O\I�/���Y�	I����q"O�D�$j�4F  �H1e��N@b�"O� ��
�/q:��W� �!��Ժ"O깚��
=%dU�f��3���7"Oba�6� "j0]H"�sΑJ�"O촁LTf�䍐ANL�r�4 T"O�LU�]�FP���2�xX�!"Ou���]�9��]ao��)��"O
�H3 ��Y��Qo�)I����"O�u�wƓ-r��@�7c��_���"Oz9T�ȧ&u�h�IK��< D"O��!�5�6���\�f�"�"O��k�eK-fCu����:���ar"O� >��sc���5S��	�C"O���I�8-��4�nO�G���"O��X �].8pw�R�u|�#"Ob�[h>S`�b��C"4]��!"O"-���[T�]!u�v%���Ĉ�?����?!��?����?1���?����?�C��J$d�bbT*v B��?���?���?��?���?y���?ٱ@�&i��(^@i���ز�?���?9��?���?��?����?i�f�	2J�x+�QEr�5����?���?���?���?���?���?���)rev\IQo�Z��=��2�?���?y���?y��?���?���?�� A�7{��9��+X,�ᑓ�?���?y��?����?���?I���?�jȍaBN��3�N����S��?����?���?Q���?����?����?��BL�`\��ߑ�v +p.���?���?Y��?���?)��?y���?��ᖚ͜�C�\�mHP�$�?���?��?����?Q���?y��?�U΋�@�Bi@rdݭn�����A��?���?1���?���?y���?����?���<��� ���m�BE�CG��?1���?���?����?����?����?AR ��d ʽ��  T�6��'f�+�?���?����?Y���?)��?���?�֋Z.1P�u�#PR��a���?����?����?���?��dQ�6�'
RgE/\\PC񋄇6\v�{�eN"�Tʓ�?�)O1�����M����]xb�� B�av@ ��ŕ�P8%�'2�6m&�i>�I��q���S� @p�f5�T���K�����	3�Pm�[~?�ڱ�S}��[�#�d�b��-�,��`�1O.�D�<���IĆz#B-��N�:%��y�D��b�&�lZU'�c������y�ǔ���1��D	7�����J ?2�'I�Ĭ>�|B�E���M#�']
��s�R�F�>e�㣕�m���'�����6�i>q�	�9k& �`��a�����+t�J�IByғ|��w�|�kv��n�����Nd18��U&���p��O���O6�|"�Z6D��ؠ�TU�#����Ot�����G�1�t���G�J�$�(w��x� $�<{�v=j���� ����O?��6fH�ً���y\�a����Z�牱�M�&��u~��yӎ��Ӱe�p,�'e�Np����42���ҟ���� Ӣ�
����'��i��?-��"M�SD�K�D�2T��h��?3*�'�i>)��ڟ<��ٟ��	G�9c��*H6��A�F�]��P�'�\7�g4����O��D4�9O�)��L�e�=�"�Hqǀ�<����?�ش2r��T�O!�t�ϸ!.�
�A�:_�:ӎ�) ��R��By�l�3��� AC�8/�Ɵx�!dʓ2�r��M�v�"$�O(
�����?���?���|�)OFqm�)z�r��	!��s�=|�j
�NC D�J��?�M����>9��i�7��O�uʒ V��q��o��5@�iM4x7�v�l�CԦ\8E��$A.�i�	�?Mj �S���nϨ{���h�A]�n���H��d����ȟ���˟ �I���Jg�̊&\�c��NF��5JE)��?A��?��i1���^���۴��S��2��	�0"cnL�c��b�yB�i�,6-�O���eӐ������ך���b�	B�+��@b��)r".ͱ��'� Ȕ'��7��<���?q���?��M��A�}p��Q�:�.L�֪���?	������ l�ȟ��IޟH�OpA������,ѢJ�j��ON<�'In7����%���?�8�h&�,5�N$yn�`C��3�I��N�?hl�'}�֝����dy��wa~����Co��!J�@ ̀��'?b�'���O��	��M#`o�S�k �%a�AXa��j*�+-O|�oZJ�g��	�MK�/M�vK6��T��:}#�< �B�I����'.��Y��iK�$�O�-	 ��1���@�<!��8]jV�����;��=@pE����[���	ğ��	�d��ϟ�Oz`%
C��t�<�:�"V�l|J��q�8����O^��O����|�4��w�����:V�\E�6	]�OS&�z"�O�6m<���I�O��6Mb��jP�sG4�"�J�d��#���I?��X#�'N��'P�6M�<a���?q1�����PCP�����K��?1��?������F�J��O�|���|*�I�q���kH-��2dK�C��$��	���o�L�ɞW���Ԧz�\8Zӈ$���I�h�7�Ŋ(.��AB�ULy��~�͐��'�X��I�F7d]1`H�U����T�G�=�e��Ɵ �	���Ic�O�R �OOz$��jS*�3��I�:��Z�Wo�I=�M��wLz���
(a7z�:�E��@J��'T���g���U6�c����q�"x1�O��̉�l�AP���tL�&N9FE�&l
Ny�s�:˓�?��?!���?��?*�6�o�Ā���ܫMr�)Oܙn;�\e��̟<�	w�s��kT���W[�����K��� �������ĝ䦅iٴ���|r�'�?Y _�(��G�;�dܡ��D�+���Ӈ!Q��򤖺_u��k�Fy��X뛖T���r΂;`��t�M0�݉�E[����ܟ��	ϟ�|yb�k��5K���OBl�&i��/�6	�/�9'� 0t6O�Qn�f����I �M���i*��⠴IQ�$���0��,ɶ8�q�im��ݜ�`�����B��e���MA[N�� �s� m��0⡈S)~v�h��4Ox�D�O����O����O�?]�it,��M�	�E�WcT՟����l�ش�Ĉ�*O��l�E�I|��@ o��Y.f���XZ���%��[ٴ@���Om3E�i��)L|��Scg�L �0��7	;\Y��j�0L��i�ЛÂ�'���'@"�'J��'�@e���R�fR�y��#R��S��'�Q��j�4�d����?9������C$�r��#|6݉ jH�W����'���w��v�a�T�O�"^�������T�k��C$
9�U��1�@}h���oyb�w�}��'����y��Y�><4
TD�[D��	�'���'B�'�bc�<����<�'��Zj��Mz<��'�[�7AYʅ�;]^�ʓ;�6�'��'�r�䛶�ͣ��D9��/'N�`�,̯e+�6��O�p��`ӎ�H\L�xd��r,OHx�#�F��Y #�������K�צ	�'�'h��'�2�'	哵u}B��j�.T�P$	���3����4_\����?���:.��A٦��:pz��%o\�;M���7�ˑu$�q����M+�yJ~R�"�M�',h�ٕ�-`��9  ��$#*���'��FPޟ�H"V���4��d�O���ۓ¼�����&�A�h�8���O���O4˓Z��G�����'��$� Y��L�I9���C�]Vk��|Bͽ<����M�I>�7��p&�d��I�����u�x~bMS�B|2����H)R�剷�u�E�ݟ�"�'F�ԁ߳~��HsǗ (`�4�'^"�'4"�'Z�>�]�q�Q�w�5Y ���Ь��5�����M�U�
��$Q����	m�i�iA,�J�2D ��;�4q@�H��tnڐ�M���q��ܴ�y�'q����c��?u˔-W<lN%d�݃x�\q��Ԇ��	6�M�+O2���O6���O���O
�3r�U-��9���L�q��L��B�<��i&����'F2�'���y���;x��s'��g�9g�@�wz*˓�?��4�����'�?���$�"�s���SV(�N=�V4 ��.��Dѻj��;��H���B�vP�3cƠV�j-!��:��b׀���'�R�'k�O��	��M[1�
�?	�F�CX�(ŅVyH0����<ѣ�i�R�|��<����M+�SS܄+�`Ʃ~n�^ x���R	�9�M�'��,B�{������S���1�u'�w�r�8Aj\G��hs���0�
��'�r�'K"�'���'��e���#=<� �g�^�R/D���.�O����O�MoڤJA�-�'�7��O$�*܌�wJ��tOT��ˊU=��aH>	C�ijj6=�@1"��t���*2��D% H�q�k�o�d�{�`��]W*������$¦��'N�'��'̒�Ӑ`@4T���C�m���P"�'6�W�Hr�4K�m��?i����	݈)��黦D	f2kMPX��Ot)�'�p6�̦�'����?�	&�@��)��
� �L�;�NQ� ���R��#a�"��	=2�����q�\�����k�A�A�XiS��E?v�>q *��?a���?���?�|�.O��l��8x��������ѓc,���3?��iI�OLL�'�6m(	�q�4��Q�Lsf_(Z�n�|ʑm�ݦ�̓�?	���!�V���Y~2���rD�۲�M>R�0�d��6m�<����?����?Y���?�+� ѐ�K?/��p@1�fK����/�¦� %�s�L��� &?牍�M�;d��ͨ�IȌb��6k��@��i547�9�4�N���O��@�goӊ�	$��SP�Z�&�(2"�9a*��I������',���'�6��<�'�?�����4��%���B	V��?���?A���d�5j��2?�����:A�x\�8�e�%��Mj��k�>9%�iq6�)�d��6�2�H�U�6��(ՙ=;��O6�r�ƈ@�����,B_wD$�ɞ?rb޹h�t�ȴ@�ԆhcՅǨ2��'B�'`r�ȟ؀��D5x¡��\������ϟ��ݴ&e�5�'Ƥ7�7�i�u�P��^m	��M�eki��㶟�n�M[�GV\�s�4�y��'���t/��?i⠥��2��	��� /T����JRS[�I��M�*O�i�O����O:���O.b��V�G7]R'f�!i��C��<���i��A�'���'���y�K����M߮{6@}ځj��FJ0�M��fgt�F�O�I�����= ����e��#`p�A����8@*E�s��k�I�M%��$�'�0��'z47�<��2&L�\#�K7.xޜ�ũ��?��?��?�'��D�Ѧ���i���`)�&2��d����32�>f��1�4��'���'`�6�|����$	��P⑬�.6@��1`N'NuN�0/f��:�˔�I�4�~"ù���NYIe�	��S%.��yj���OF���Ob�d�O���5���vx(�E�^�~��,�bϛ�#�������I?�MӦ��}~�����Ob�YP�X(MT����B�S����UO'���ŦѪ۴�?Y�n��M[�'�b�"h�d	ԈX%M�4R�nWZX�!��Nԟh��^�<1޴��4�����O��䚂6��h��' l���kQj��kG��$�Ox�YT��J��y��'��X>u ��V2*��}���_�V�E@%?�q}��tӺ�l�p�i>���y�*�ce�� [ K0hW�:�0���o�^Q�E�*?�"���|���T�˓��[�"�9ʂ�I �qeb�*⧟?�?i��?���?�|r.Ot\l�
�;�MO~��A�s��bD�Aqy� lӨ���OdhnZ�5o`�cWl�,FD�O�"�~Y��4P���f6O|�	#\�J�(�"�վw"��$��� �-�cg�^ۜy�gA��hĴit栗'+��'�b�'�R�'h�'@�N�eT�ٵꋄp.x4q�48Yٹ���?������<7��y�
�����D@'v�Za����6�ԦXK<�'�"�' 8zy"ܴ�y�˞(*h$�Ө�r��t�6(ъ�yҢF(:�`e�� k��I�Ms-O����O��2�
�A�ЍA�(�+�K�OR���Od�d�<�d�i��0��'
b�'@BM��`5���.V���2��'!�'y�˓�?�޴r�'�Sǀ�p�^yhw"_+pY<屚'2镍wRܨ5��	W��.�u'gM���p�'��ez��:jn 9*�g�N8��z5�'[�'\r�'��>��2[���,��'�ܭQcȖ�I��	&�M�ܻ��d�ɦM�?ͻ<T�%�,E�4XN����Vg�&`�̛��k��oZ6:�\�lZs~�ݧ'�.q�S�D��G�8W�X�cꍸi�R`DU�jٴ���O���O���O���:�
��	�qNV8���
"�VʓLe�6��L>��'	���'ʄ0��Z)�!B�������<9���Mc��|J~Q��!��A��fR�H���` �
#�(��i��$�ph����~Th˓�vS�����@�8k����_K��Z�kZџ�����������Dy)p��IZ'�O�!	�ϭA�����J�t�U�F;O�n_��8��I�M+ŵi˒6�C�<�����b�ZX�4@V"IPry�akh���ΟJ�Kʸ:����Gby�
q���Q�`�R�V�5Þ�P���!0��I柤�Iȟ(�	۟��I^��XF��IX���`�ƒQ�m����?y�؛���7-���4�MI>�w�>W���S ��!y&�L�zV�'�R6M����� $čl�g~��
#�T� �8����!�Z"�t䪴��֟0�C_����4���Of���O����'0���b��.3h(A�EI�&����O<ʓ=כV
 ����'8�T>��Æ�&�)��Fؼ7֞L!V�:?��]�8�	ݦ�hJ>���?�gQ��xW�]((~�H�"�p��X��^�wKV��'f��]'2ReKyb�w����D�E��@+"��E4n��4�'���'�b�O����Mk�B�)CP6��ߊ$H>��'ϩr�Ҝ",Oj)m�_��"H�I�Ic#�\+*�T�Q� W�����8�M�T�iJkG�i��D�OBUq�"ɫ����<Q��$-	�
�5�<��RE���R����ݟ���ٟT�Iٟ<�O
F��&��N� yȀ��C!6I���cӜ|��9O���O���$Z��]�$�mޓu������UX�41A�FD=��J�"6�w��#$���r�l8����-x����$�|��+g�)K1��	K��hy�O�� H�6�-Q�9�"(��A��?���?Q)O��n���	ʟ(��#?QL���O& <I�F�q�)�?1^� �ݴ\��i;�D� �`���E1�X�:�Fį+�I1$6�q�6��_
�b>���'����<!X��A���f��!b�G�]�����П���H�Ip��y�E,B�Vb�#�H�v���D٧QW��rӐ�p���B�4�?IN>�;|�0H��E	�i��$JS�ۇP���kX�6�r�b�mڜ<ln��<���2ty`��.Hಌ�'M�0m1t�מ��	�BJ��䓙�4����O����O6��, �M�'�yuJ�sE�s��L����2���'�����'1rD�2n�7���z����`	�S����4f�f�7�4�6���:��A�.D�xqA�ƴ�X1t
 b`�����<a`��)3��� �����G��%K����N�A$�
Ae���O`�D�O��4�d˓UM�fŞ,2=2 �Z���ڭ5�&h)��	��yr�q�|�`�O�HlZ2�M��i��|�q� ..�H���χ�4��a,�/R��1O���^" a���^\$����;S]�L(`C抍SU@к3����?���?��?����O1���<*�����L�^�ej7�'��'��6픔T�b�8�֚|ҍ��"��X��Ӑ]Qܸ��OB�q��O"�m��MK�'OZAQ۴�y��'��*b��;q�8�&�c�\�!�6p~>��ɒ&�'x��ɟ���˟���3<�0����( _�؂� 6�����T�'26�(C`���Op��|��H���zh���ukr�kCm�l~�J�<���M��|�'��S���/��i�`Rtڵ:#�ɢ�.ycq'��S	<0q/OB���?���4�D�w�Zr̓1Id=@i��8z����O��D�O���	�<���i V��$A�a�x,��i�1��|�^&^K�ə�Mۏri�>��iB�3 ��+v
�!Ǐ�2/�d�� t�r	mZ#N��Qn��<��rBH]Ac�y�-O��x&��G��i� �U�>y��as4O���?��?���?������O�48���L:�MZ�&���m�h�@1�Iȟx��u�s�������JS�6� v�
�͂Q�������`ӄU$��S�?i���#yv�o�<�I�o�0����4��
�<�VNн2��dL�������OT���ET�xՁ^�<n�@'kގE-&���O��d�O�˓+8�6���B�'��l���'^��=K5�;�Of��'�6-Y¦͛O<�ਘ1gR���񎉄*�4JϤI̓�?��p��2􌙕��u3�iV>�� �1N����A4��`@2���Or���OJ��'ڧ�?I��I�	.��� �R�@���H��?!�iJr�2@Q��H�4���y'狇[3��Ek��t�)�nJ��y2j�� lګ�M�TИ�M��'T�.�(ά���ۀ �ၧm��]� ��ٳ�ᐵ�1�d�<a��?9��?����?Ѳ.�:�xi�BȴR�.��� ���Ħ��@ܟ���̟�$?��4'4P:��:[��A��	�+0�r�P�OT�n��MS5�x�O��D�O�>�J�i�
g�0�r����b�����9���P[�x��"�1i��BQ|��py®]bV0�DlұUN�)��ĝ ���'��'m�OM�I��M���J�?��L�1��Q"TeĢ;k��!҇A�<�i��O���'W�6�Lަ�Q޴<_fAS��f��5��[�5a�	�1HO��M��'2B%̧Z���S���?����4!9�leYU��9������Пt��֟��Y���6�x�mE�8����2F�1K۾�k��?��4]����q�I �MsK>�p�#L�%PrM9Z��"g!Ѱŉ'46M�Ŧu��(2pt�l�<!����1�@���H��b�����\���H$GT�$9����d�OV��Oh��GwB����11�B$�DǞ��L���O�ʓc@�栕;���'-2_>E@g%v����Fό4��(���O�p�'�*6-N��ipO<ͧ�
�А"���&�Gh�k�I���:1`Ơon��*O��C��?	p�"�D��|2�a�@lOd�<J�$4����O��D�O`��<�i����N�ʔ�qW� 
̼�q�'�<!M�I�M{��Π>с�i����Έ�V�B *��"$쬰�ha�Zm0p���l��<���tD(��&��	p+O�ӓ��t�v$�5��+���3O���?Q��?����?����iX�4�DjQ���IJ ��ei��?��Ml�,%h<�I��\�	r�s������37�͝C$���
�B�5���33��v�`Ӌ#��ɞ4u�7q�7nJ�-,p��"F�%��3�
w��b��'Nb�	my��'���
��8:]����7�]�Z������?���?I-O��m�/x%�������bTN�Y��r�N��)L7{���?iA_�$@�42�6#�=BR�@�h�*qRmB`�!n��OI`�~1آ��<i��jXp�D���?�Gd���������4����?���?���?э�	�O&0���^���Q�gS����Kg��O��o�v��d�'�6�8�iޙ�VD[w1���r?�J�n��Rߴ ����|Ӧ��եj�<��.<x�$���hc���"@��1&M� �Byq�O�䓡��O����O�$�O���T�,��ъ�c(�2��0d��uh�	*��G�!�'���$�'_�� �R�7]�Y���H�����<)���M{%�|J~����N��j^�BL�9�l!���p�ʗ:��гU� H��S���O,ʓ#�����j-i%�Ò:h��?����?9��|R,Od�nډa-64��5Nl���� ��@R�D�"��I��MC���>���i�B6���q��8��T:G6h� ��CpmZO~2D�#���ӿ<%�Og��>��� g�Ӷmo*�0���y��'("�'=��'���)�-����p���I� C�3��D�O��$Ԧ��BFvy�v�ΓO�<(�×1���B�*	�MR��:caJC�I��M��i���~���>O��ʃ:tE["��P��L0SQ�yQ䴩B�4�?!�i#���<����?����?�kSS�]��GԊr�\uZ@MT��?Y���D����(�#O�t�I��8�O��@g��$�!�B��]�v���Ov4�'�t7���*K<ͧ���J�4�n��&K>�x�����a�3Ǜ�Tk�ԁ+O>�I��?�Rg'���O0�r&E�&�[� ��5(��$�ON�d�O����<�c�i&�̈�M�2��]�%ON]=�<��"h���MÉ�O�>qҽiV�ܠ�E>N�e��I�&� �9g�m�t�lZ�^BL�oB~"�E4O�Y�S&��ɣa�J`8���~d��1�ȧqTX��Fy"�'�r�'6��'�r\>���eųzD�� I�70�|8�f��M�ń��?���?�I~�?=��w���&��Z�{ .�*��i`�zӚ�nZ-���|B���j�͊��MK�'��97ɖ!Gj�(piڪ=La�'���	rϟ��3�|BV�����ĉ��)aFЉb0�\.&
��*�ɟ �I��\��Zy����d��O��D�O����?ݺ��̈�m�v����;��2��X�����4!��'�����mx�X&��gmP���O� Z��R�.�*��:��^��?����O `!��'���ʓ]���1���Ol�d�O��d�O��}λ��p	�͍)�12�"�S�B)K��k�6
��F��I=�M����Ӽ��/K���afK�kwB����<�q�i��6mݦ���M�����?�F'� O�����e�u����;���p� �|~�-�K>�(O���O����O����O�YZq��y���5EEaX8���<�g�iR�E���'���'���R>�,A���9S%^(w3rP�P)�E�R�O�o=�Mc��x��4��/mdZE�QCZ�2���$+�'U��*��Փ?t剮l�PmK��'Q��$�|�'�t��e'G+\;�eLR-x�|X!��'b��'�����R��bݴSV���A����E/[N( j�\.k�\�"���'��'���ӛf�|��o��{Ϟ�y��^�T��lr ֟SD���HC�����?�qjƾH���������l��?pa�Ɲ?M 9��	BS��$�Ot�d�O����O���5�S�h� 3`��iz{�ƙ=��}�����ɿ�M�6!����ʦ�'�r�׈9X��"��	�is*�z#C� ��0כ�imӚ�)�t�7a��I '�z� 8��TC&��D(���^���aRcG>�?���&��<����?��?q���{��	�&�/2�%zȝ�?!����ėǦC����	ڟ8�O�m"��%'|���A��<���r�O���'װ7m����M<�'��7G\-OgJ����Z�'_0�)�șYs*����/C��u{(Oh�	߇�?���)�䓯K����,<N��D���(k����OF�D�O���i�<q�i+V�z��;��K
: j̘ӳ��>w	�I�M��K�>��i�p���Ö:m܄���D���-X�cg���nZ`�>�lZ�<��:%pҦ��ص�.OJ؆�O��i$S<#<T��0O�ʓ�?����?I���?A����<*��sF�ֻd�D��$p�j4o�=F�K�OB���O���$�Ȧ�]?1�����7C��[�FU�u���	۴����0�4�*���܈Io�,���hL�WA�#$�r�C@��(j=��I�xb�Zr�'��'���'��'���U
��H1�4� G������'�2�'�2Y���ٴYY�PΓ�?!��E�L!��ϳ<���y�Onx y���>���i� 7��o≉;{�٢D��$|�@�D7���蟬@�N�Cn�sè#?a�'Q�$�dP��?�@�&Q����\n9��0s��8�?Y���?���?���9�����R�0T20�qC��R!�\33M�OX�mZ�Ssl��'~�6�4�i��bC~��E1O�;�.Y�r�p��4,&���nӜԺ��~�l�Iğ<���m��B޹N�4m!�fE�o2
l)`�K $��&�x�'�2�'#b�'���'�V s�ҝ>W|��g�ڒ'��Q�]���4w��8͓�?q�����<iDgE�_Cn�	��E o>L �g�H�>v�I �M��i��O1�t�I��
�b^�����4�sDO
<_�1S���8h�pRL�r��Uy�ДR+��C�&�wmɁ�$u���'q��'��O�ɟ�Mk ���<1��")���q���'(��	A�I�<Yſi��O���'�ҳi� 7m�>"�=��T X��Sa��&*�&� ��o�\�I��@��xu��L-?a�'���ݱ_���#�ė�47~�07�S�<���?���?���?����؄v�-�3��>�`@�^��yR�'���v�@�J���L��4��Y'� �oZ�,�*���C��$��e�xb!g�B�n��?��������?�u�F����`�4;&h8*'e�2���p/�OM�K>1(O��O����OV��ۿ-���PC��$�f��G�O>�d�<d�iJB5��O��D�|�h،B�)Ď0�r)j�E@~RI�<���Ms4�|�'�.Ll}:w�
H��r1�_!Șm�FC�'l8,y��i�p~��O�rx�	�a/�'S��(�*�Z��U2�I�A����P�'���'�B���O���M��V7
܈��)TQ��qyC�����a+O�n�Z�W��I �M˳䚡G_8�bCt�a��7J�F�k� ݱ4 l�8�I֟$�b�����my�!�/>z���$����q+C!��y�Q����֟��	ԟ��	韼�O16�;���V.h0�q�
'M�i�t�|`Њ�O��$�Od��������W�����$_.��&��)iv�@X��M�ě|�'����j�Z�xٴ�y�b�(V�Uk c��^������y���(���I�'�IƟ�I�fN��i�薏.�N��a/Q�P��	֟��	˟��'i�7���R&^ʓ�?ѣD��f�j``���E��h0Ц��'��V���x��'�\صfV6�H�jT�B�V���Y�y2�'���0�ܱweddtU����q�@�ş��!�7Tk�!)´q� �#ҏR�?���?Y��?��)�O`�)F��2�U4!ݏ+��9���O�o�=d�$��'@�6�;�i޽���߷dþJ�C�z����"l�|B޴t���~����r�d�t��🬻��M6o*���M�b�9/ٶ�a2ؽ'x�l$�x�'�'�R�'��'*��"���.j�M��
*Z�.�#Q�ly�4Z�0����?q�����<i��ߚ�$���Ǽ�ܠ
����nN���MK�iC4O�i��(�	K0q,eb5M����`9f��V{f��Ґ)�%��$�{V���V���OZ˓)�%��՘-4֭#��P�bx�J���?!��?���|*/O^�o�`�\E���_`�Qf��ԁ`��,)y�I��M�n�<i���M#ӻika�k�t�",P��1\�P[����=��:OH���'��4���N�˓�j��_�����E�}o<1:d���bo�D��?��?���?Y����O�<�@a�P-Qʱc4m	r�4� ��'���'��6I���˓P�&�|��G�?i`�(B�S�}�ëܯa�zO�n�+�M�'0_bQy�4�y��'�~<�3���yAp,�F�D���p�'Xi�����A"�'���ȟ0�IΟ ��,��)��EĂ)�E gN��jy��ǟ$�'�J6�-^�8���O:�d�|B��Á��u�P��1N��0c"Tn~r�<)��MKa�|�'�j @K�	֩�v/ǵk�9��H$-��c�^
/�@L�,O���-�?�1�:��O�=���*���yANH!����O�$�O���<q2�i�[��I:������B4?-ȱ34�4Eo�I��M[��<��4�B��5"��L��&�A�x�A��i�B6͒�[m�6�$?�b��O�������^u�`�4&p�Q0�E�_`�d�<����?���?���?�)��9(���+H�L��6v-捋�̦}BvL�������L'?�ɀ�M�;'�Եт�HO��9���%{��r��i�6Me�)擝Aڜho��<� ��*5`�7M��c���t�4�8O�xk�HJ:�?���$�Ī<9��?Qª� 7p�ke�/��vO�?���?����d�˦�sr�ܟ�	֟ s���x;G�F#+Qqi��Kr���O��l���MKD�x�c�A V�X��Nu|L@RI��y�'_A`��7�	Q�W�d��4��Eϟ�6m�KJ]�ס�UQ���W���	����I۟�G���'Dq��ʬ��jǌ
�a�2�I��'��6͏t�˓y����4��Ha��؜MH)��gQe�&���O�6�R¦Y۴d�r���4�yB�'������?U`¢ޣ;�~aţP�0�t��dAP�vm�'��	۟��ȟ\�I ���LP���t�G�Axʨ�a��ה��'�z7M�$#j ���O^��5�9Op	{b�W�|��̹v%�=�l5$	pyr�''�&�9��O��t�O�l�qSf]=ta��"���$�	��r�ֱcR���V#��U.R�X�y�hF�_�daS4�'���т�H>9���'=r�'F�O�剩�M����?Q��ۘ�:,���S��h�U�<9ָi��On<�'7��ܦ9kߴO��]2�eI%E����R�X|�0I�M]��M��'f�&�J����J���?u�]J�P���j��`;�-C�)��}���	ʟ��	����՟��I_��ܚ�{�n�{�d�1��	TU�}p)O��d�զ��U�#: �i��'�Фs��
���s���!̰���i-����1���|�r���M��O"���D�*C��a�K�Rd��֩_y|�R��Ox��?a��?���DR�}�-L,4�t���*�xlř���?�)ORm�_�����̟��	D���Xb,д1FIDT�Խ"AL�����H}B"v�>o���S����3����g
VZu�`�BOFJ�2��зMZ`���T���A���C�oD�`	$��F��	��N2Q;"!�	ğ0�	۟�)�SHy2.|Ӵ�U⋉���P�M��)��G΂s$��d�O�	m�|�@����M��eǅ�l���'r\���@[�fu�6-���o���ퟠ@A�%#�ĮXxy���H�����}�
Bt����y�\���I��X�	埸�����OÒA�k�:E�V���Cj��9"�~�T�b���O���O��?i������,��E`�u���mт�)0Mϛ�fl�T�$��S�?����E(pn�<Ir�ׅq tCF.]-�f	���<!7 7j���D�0�����O ��u��1�J�;S:��	�+F�V���OX���O��[B�ƫ ���Iß� '� ��y���ƹvŎ ��Z��x��	��M�c�i��OH����$��0�QBZ%ei6���8O@���$����!��������O~$+�o Q�BaD�jH]ef�*!�Xr��?���?a���h�*�d�%���{�K Zn�@ #�~���i'�My2�oӊ��]8X/8�Dc&R"�d��	����8�M{r�i�7m�u��6{����=A������O68��I�*f60��cг� AH�&@Q�IsyB�'���'�B�'�N�-A*��6Cɝ3��s�L�j�� �MC�.ֳ�?q���?�I~Γt���� T<hNP�/$%�4���\����4>�&�=�4���i����S�eP�B"�	i�<���V�]^�>��d��<Qv#�y`�������Ł\�f���FR�}��`��ZS��$�O@�$�OL�4���|�f�9).���*���p�*ަX�
�j�Q/�y"m�^�R�O\l��M�Ŷim�̚B:QyTY��
N 5�1e�|��f>Ob�d�27�x��'{�pʓ�r��Sxx�@`ƾrV����E9%���̓�?i��?��?����OL�9&	H�-&]�U��f(,�S�T� ����M��B��/r�h��<��JN(+��IU�E7}�`�GV=)��'��6��ަ��?���lZ�<a�/�����e�!N���xND&Ѣ�!_8�$ލ�䓚���O����O���@�y2�EX�MM3H>��H����:wd���O����&%	����'y�S>�ka�ٱ1�=3��L��O'?�!V����4i)�6,�4�f��=xW���X�M�/C�^$ʳ"=lU`<ʡ-ѴN��ʓ�����O��H>���W��E ��\+q�,�[�͊��?����?���?�|J-O��mZl*Ip�@Q:o�u���֫kP c�Dy�b�R�� �$�E}Rnl���1��d|��ԇ3d�֡jV���MK�4	����ڴ�yb�'�R�0��?Y��Z�䛒�K'35����,A<���p
p�x�'��'�r�'���'��z��:1�'i��Rq����hQ޴U� 8����?������<a���yG�̲E@�B�>'tfa��%�9~D�6���i�L<�'�J�'tq���4�y".�n���h��^%��|��)�y�.^��i�I�<~�'��ߟ�	J����R�k�(�zQ��#{u�Iǟ�����8�',�6�J���O��䎽" �S�_��Z����5_i��"��u}�xӸ�mZ���(�E��/ϡ$XL��P�N'b�ܕ̓�?��Ł�`�J42�^�����R�waB����$1R�̖($V�z��O�^���D�OR�d�O���'ڧ�?���3(r��@(�A؎0�녶�?�b�i9x�X X�޴���y�(4y��p�aj�~ڒI��d ��y��o� n"�M;��5�M��'&bM��No���3yU<�#/�Vʴ<C$)�8K^8�W�|Y�P�	��,���L�������J@�Q���P+"h���pyRBiӒ����O��D�O:���$��n� I��VT�h�PhI��!�'��6�Ǧ=�J<�'���'12z\� ��G����I&��Y����bʘ���6:41��.�O�
L>�/O�=@aL�4E�VDD�ְBdV8���OJ�D�OB�D�O�<�Կi�F<���'"T�
��ȋB<a��*]=4��ۙ'1�6�&�I���$E���Y�4�?����5�����P #��i�2	ʍTU�T�ܴ���$N6m��'��O�>�،#@�I�g��;v�=�!�
� �H��ԟ��I���Iڟ�	M��
\�����{P��$ڒE�t	����?���Ư6�a��M;M>�����4��&�a��@6���y�Z��(�4tW��Oe�A��i�ɵ�j�b_�*����"�^�(g�,#"`�\�Ily�O-"�'�b����qh�m�@�r<�#��CO��'�剂�M�2���?1��?�)���#&�A�k��K'N�fi~�ps��0�O��lZ��M;`�xʟ�hfhܭH� 81������e%O�j����3N��]|��|j7��O�u�K>��d 5\��D�����Y:����?��?	���?�|�+O��m���:P�.��4��k�4K��+�iycr�����O�l�k�0�:�G�8�d �5/�/$�|���4q囦��.�V3Ol�$U9M<~���'{q��{��u�@�+z�IwJ��.En-����O��d�O����O���|r$b�R��
�뀱iVT��tЁ_�V��9U���rS��y�S �<	�� S�����J{�27��Ǧ��K<�'����-$����4�yb�Hn�����܁T����2��y2��Jx���.)��'~�I�4�I�yva�׎��*�I���rK�M���d�Iޟ�'�7-X"�����O��D	)IL���m[*6|�y���-R]�⟴��O�m�>�M{r�x2�L�nO*�#Q%�e^$!�+�9��$J2Mˤ5 ѠBqlҒ��98��slD�D@�n�;�O9?[�!ʕ��. �0�$�O����OX��*�'�?A!O|*$0�0��R���?A�iV� h!V�`�ߴ���y�"��oLd=�gQ7�F8Q4���~2�'���*d��i�ҍp�6�V!�)�@ �}��K�;[�����
%g�P� '���'���'���'/�'ŘM!Ž1|l��Ǝ1�P�BY�� �4�L�	��?���j+��<]䚙`�f V��ф� O��'�7m�˦�SM<�'�J�'y��K1nԳS\P����y�I��O�B�L-j/O��"���?��4���<0G��/�@T�Ձ��1�����?����?��?ͧ��d��q�(��t���5ڽ�*�#cE�m�C�h��K�4�?yL>9�R�<޴m��%~��!�V�ۖ�D��ЁÏz&��t�i��6�w�H��t�h[@�O:���']���wS��9E�'L낌�@�
J�t�'���'"��'ER�'���:FB�1���d�F��$�3e��O����On�O��'��6��Oʓd�z=���P�n�����5\��xh�x��q�n�o�?��6��㦝��?y�K��@�so�E�>Pz�a����0�g�OԙYN>-O����On�D�OЬ;��ƿMt�6Қ!
"�� ��O�d�<E�i?��e�'o��'��S�(�y�t��c�����D_rd�p��I��M�#�i�,O���R	�?;�܉����f�YP�jȠ�d�*�-��2z˓���+�O�T�O>14�ֹ1^�����3�L���K֤�?���?����?�|j*On5nڶ2X�P���.
=�=D��٨�j�@^@y2Cp�|�d4�d`}2�a�̤� `Qc!2C��!b��{�l������4a:H�*�4�yb�'�,Tj��?usTZ����F�'b�a��U�41@���
t� �'<r�'2�'D��'��S�(z��q�5*��C��!����4)U�x`���?Y����<���yl�_�8GA�:;�8�W���7��A�I<�|Z��@.�M�'����@�/ >�y�A�m��2�'�P!��C؟4�֘|�U�0��쟸#���7,?t5��@V�X�x���@ퟸ��՟���Wy��l�,��2��O��$�O�42����B�CĀ[�F�0�.������զ��4�'����s��
R�Ju{v홮<m��1�'����*gl:m*�mXq��	�?-�t�'h�E�	;Aҥdm�0X%��H��:� ������ܟ`��J�OwaR�'6��Ԡ��l�	p��#;2�d�ʕJ���<	�i:�O�Nդkl��I�J&�p��e� vq�ݦ�ܴ@2��CB$��2O��D��d�x��B�БuUIs�č�(^�Zϟ���OV˓�?����?����?��l��0�mJ�)W��{ŋ�� ��/OĤmڧ	�U�I��<�	V�s��q�Hͮ3�|!�3%	10�P�S"��'��Mܦ�۴uH���T�O����C�5�1���M�����B�lEY�^%J��2,
���'�(u'��'�l=s�lH>�����O����'�"�'����^�8	�4/P����x�����'Z*lCf��w�!���}�����_}��z�F!lZ��M�Md�f��pF�IQn@S������۴�y2�'SJ��4���?���U�T��ߥ��T�&��a��E�;鲐��r���I؟���4��⟘�Zk�3R�Ҽ�'�� �E̚��?���?!�iHXڳ\� ݴ��s,D��
�O
�8��Y���L�|��'���O͂�J��iJ�I8Ubi# "�'E䌱�`,x
� ]�,��X{�I~y��'*�'�ҡ�SՎ��v���wS �£N	�?9r�'g��6�M�ӧΩ�?���?y/�6�h@�{��y6mvK�������*�O��n��M#E�xʟ� Ne:��˱)��]Ȳ� P��JV,T&8/��@U�� ���|Z���O�|�H>�k��3��w(Ld��#�,)�,���O���OL��<��i�fQ��9A����q��0cS�K���*��ɲ�Mˊ��>a�iQ�t��b�8`��-!�*F�+�"���n�Pm��3h�El�D~�"`��1��+��%k�0�1$�Ҏ�t��,H+ ��Zy�'��'Y"�'��R>�{�'�&p��s��,
蒰���?�&�hyb�'��O}�b����F�@�E�dx@�0�Z���Qm�M��x����Ǉ@i��<O����2@F�8�]�2�ꈳP5O>-��ǋ�?�s�&���<����?!@���Z]Z N_%xb�:�Y��?a��?�������p���ޟ��Iğ����Q�|#���J7
"	�#�Q[�yu�I�Mc�i�BO�H���˼B�T���}B������8�4

�w5�Iӂ�C��u9B��ӟ�#Wc[Yx� K ͅ�k��a��F��L������ݟ�G��wk�����[-?�� Ӑ ��6G\�p�'�7�#G���O6io�F�ӼkS��#�������@M,dY4JF�<��i��7-�Ӧe:����-�'��8�R��?�x�m�VZ�֬� ��ԁc�U-T��'��I矜�	�����㟰�ɹ0ˮ1������љ��<&\���'�N6�ɇkG����O��0�9O��� �A+[Y�$��Á/DxՊ��Uk}�Na�\�n-���|j���R"��$/q�-����.d�X�a
wehP�����Y)����wO��O���H`�СEDQ�x� jUo7XlP���?����?1��|Z)O(pn��mj4���.N
�����P-���_2*��7�M���>!ƹiIB6m��5Z7�/L��K!0%�͑6Q�кi��D�O�92�fһ��a*�<9��ǿs����f�L�T���/8t���?����?���?y���O�F=�<$��TC?B?��3t�'!��'L6�^&X�h�j��F�|���fN�!0�1j5�9�b�K�2�O��oZ��M��d6eh�4�yb�'=��bȂ���Qs�j�7_-���2G�,�$H�I3��'����p��˟��	^c�c��8����m�)]4vd�Iܟ��'�7-\�'���O���|�4�����Er%e
�J�}0��WG~��>1��iu�6u�)"�)M/`���3�Ɛ2Nn^u�엩1�z��Ƃ�j9����ǟrԙ|�dX!q�h��N�9V>��ǭ��r�'3b�'����Q����4E*Z)�'+�&AD&�c�+�;n��al�"����y�?�[��*޴1��!YS �s�'��!Ό��is$6���&6�/?�#!\�	����DȊm�8*�\
&�,k����d�<i���?���?���?�.����Rf���-S�4��N��:�E��L��ş(�RG��y7�����x��S/Wh�ي� �*�Dj�Hu&���t:E�z���	c|���(z�F�s��E�&�.�;l� A�'�'�\`'�H�'���'��D1u/�*@��������I��'�B�'�_�:�4R��TZ��?)��q(�(��"b�H�"U�PwXi!���<i���MSВx�Ǹ_��t�CF6�ʅLT����^̓φ(|��f��������'	�qv*��`8:���A����OF�D�O���/ڧ�?����e<hi)��T�u�q8�ˁ�?�'�iMD���^�,��4���yJ��%5Z%z�� c #;�yRG|���n �M��E�M{�O��րE5������P�5��!>᪜ �o��G�|rU���	ȟP��ğ��I��L�QG����0#�ćIq�E��Cy� k�n���N�O�D�Oz���$���څ��L�z�t0 �� +�B��'F�7M¦�L<�|��	� d�=@�o�>��7kG/ T�G�����ެx�0��wKҒO��5�l��Q 2}*AX%l�-������?����?	��|.O�oZ�@,^)�I�Y��xH��/g�4�!7�Q(5�X牸�Mˍ"!�>��i��6m�O��"g�p�N��R.\qJ�胉�g66�>?i�#V&4#��)9�Ӗ�5@Z9 ���`�	Cx��N��y"�'���'���'���	�!�b�����?V�$L`q�t���O�$D˦��b�ryB��F�O��
Ѩ\�pn�Y ���0�`D��{��'T�6����Z��Dl^~MU;F_�Y��o�8�I!��mMt���������|�V��S៤��ʟ�0F��&ٰ�����1&z�	ş`�	Eyc|ӈ��I�O,�d�O�'%If-*���:K���%�-"�i�'f&�2���i��$��'bu��¤� ��q���O-FxJ}Vg.XW� 9�����4�.Q��vt�OD@�d"�n�~��O�o�r�KG��O��$�OR���O1�˓	���i��lt
�h��غy+\h��&�E� �fW�\cٴ��''\�Qg�vML`��KSL�!<���1�O/?w�6�֦��$�����'b� Bc.��?��1Z�d@5'�0��q@j�0|$��zQ�o���'���'?R�'�r�'��;]�p͚$�*��xц��-��t#ܴ�
�H���?������<9���yW�B�<���7�#QQ ���mu$6-M����H<�|2��Ҏ�M��'h�)���'9�J��ǥGP}��'�j�����ٟ$qt�|�]�X��˟	���.1�B�(���R��nٟ�������tyaӜ ��O�O���O��%�\�k�>��� I�@�*�P�h.�I������k�4&���� 6�2�ٵlԸ�p @3	[�����h�	���P�q��V�ӏ�⏌Ɵ��V(Y�q8T���� -�t�	"������	ҟl��ԟ�D���'혅�$�,~���)f%A(�%�OBxo�2)�Q�'�7m$�iޕcEۊ=<b�Y���96���ȧ������Y��4s�ʡq�4������ �'-��X7��\�>�C�M9xu��Q%C(��<��?���?)��?񥡚�	��uAkҽ�%� �P
��$�㦭���Dy��'�x�ӂ
^���)GN߹&.Ѕ*��W}bAm�t�o���Şv�
I��"��Ү9���J�9����+�_/0�Z*O^���_��?	 J!��<�,��ZH$fu�j �7���?)���?����?�'����=ۓ-ȟD��ˋK��Y��݊c`�Bob���4��'6,�5Û��hӪamZ�NF(�c�n?� ��qP
���m�Ϧ!�'ĝ `ɓ�?b@���w� ���.h���'�Y�w��eȟ'�r�'�b�'���'��fmX�g��9�xA��Y'q�8�I�.�O���O�n� ��͖'L$7�?�$�&����TKK�&	���3��j�%����4^x��Ox���E�iM�ɭ;;1�'HғE��%���,~�)�	ъz�"�B��Ky��'���'7b�ȫy���c��*s�B	�͌D�'Y�	8�M�4�<�?���?�.���C���'�8$��́�}�X�[đ��[�OؼoZ��M�%�xʟ���nE�51��(͇��@g@ϬJ��l���3U�R��|z�%�Of-CK>a�lΖS6\����z$�0���?����?����?�|
/Oz�o�33I�13�+FP#VN�S�rs��sy��xӘ�`#�O5l�-ot����œ�1�l�+��@����޴3s��AJ>4�F������S50����{y�Q�ɀ�r�j���yA�,Ұ�y�\�\�I៌����`�	���OZ���CnB�|�3^��U��͂�5��pM�I�|�IW�s������cvl��o��I�A� �l��:věրm�x$�b>�i�C���Γ~���#�?v�>�	 ��`�ϓZ:*�#���OI>	.O��O �PA�֔�v�h�!E3.&���tL�O��$�O���<Qֶi}؄ј'\��'J&I��A�q5P�#g�В����r}�w�*lZ��}�D��7mK;z�Q���(P \�'�`��l�qr@���dNܟ4���'��NO�i��#�
r�`�'�B�'�B�'��>��?���Qq�ͳ�nZ�:�(�	�M��G�b~2�oӖ��ݨr�и�'���&�AW�&��牳�M�V�i�6-�>9��6�%?���@.$Lr��A`� �6��$R�!����-
PL>�.O���O ���O@�d�O����	b ��%�̲8���2��<	�i�,u��'A��'���y�IN�[9��R�f�wy��+�dl��di���|�
�'�b>�z�	X`et4 �]�D �aD�F\����/?�"R<=������䓿�D�� R*�H悆Bj��Д�[R�t��O���O��4��˓V�v���y�EC�r��yђK�;'�b��n�8�y@x�z���O��lZ��M���i�v`�ͷY�� �/N�^�ꍺ"'�9�v���w�J1P������h�I�0 �\���8%��)�&3O����Od���O����O��dI�ZV�9�<��A���.UfDE���#:ҥ�K�Of���O�mZ��tA�'R&6�-�D!%o�a���$.�NxZb钄@��&���4z���O��◺i����O���&[:0�a�	�&E��l��
'~ ��+��d�V�O���?!���?��8<�,��(ɟNN�Q,�$Qs���?�`:L0B�,�
w�(�,O�����瓰j�2A[�CP
�b�T�S$*Y~�t�I��MB�i�RO����@��.�<2YP���Rd9p�kge&�@9�d5Y��˓��դ�Onq�L>!S`�C���B+�#[?��x���S<���i����@ο:��u�vF�%	���+�$����&�Mˍ�F�>i �i�^А	�>?k
�ض��	e�0��eӒ�l�.�x�n��<I��O:���c��D�x)ODi��M������T!ztv5ʠ>O\ʓ��=�,���$�k#LK14:ZI9��K�$���ɀ�qo��ʟ������y�⌓jt�H��*gV�9���ZL�6�ѦM�N<�'�b��E�d��4�yb�Y�8��$rVLR����kRFǸ�y�/�g�"y�	�&.�'���Ky�̌q�,D`ê�#� 4WǕ5�0<���i,l�� [��	�a�:���d�(+b��&��?QFQ����4yQ�fl(�$_�NV�EIu��4^����	;m�$�O�)��e�'D�.���d�<���9��D��?�a@R�6�f=4�\^��d:��Wg�<)� �1)�>ɪ� P\�n�{�-���?1ÿi���b�[��{ش���y���{0��P`O�%P��y�D��yR"c���m��M�4�[�P#;OJ�Ċ6~�^����7���8�%��s/aK5���*�|��!�D�<I����*�,�:�*��(I )6%��	=�M[)G���D�O��?)k!�:���+���'�N�#������O�6m�I�韴����x"� z�%@۰d�@5I$��y8���c�<!�d��6q����䓵��>�H�92�z�AB��a|r�w� �H���O(u�� �Q�`}�Gl�0Zk����;O�IlZm����4�MCտi�>6� B���h2̊b�Xa����
N� ��7�k���		X�Z�"��O�2L�' �t�wrl:��l���cgɏ�&��(�'A�2��/�-+01t*P��Vɇ@�����x�ش2�^ �O�6m#�d� �]�S�*i�Mi.��Ro¹'�Hm���M���q&l��4�y�'��m����"m�����%J�gH �b��:p�5�I/�'v�IE�.�1��NW�]�$S7*C�$}Exr�rӸ�X׬�<1�����T ��M �HY�"��!X"
��ra�������O 6M\D����i�<�V��%�
A<q@�)�6Jx�c5��	7�Q��<���o$���D���U�N����ܸ~�DdsA�r�x���M�˱�p�3�L�g/��Zp:
�C Q�L��4��'#����Vl�/~H��(?v2��J0�:�6M	���
5N���5�'N���I��?�J�Q����F-�~ݐ��Z��srk�̖'=�{��_��ѥ�O��'Ţy��7�G;�p��?���$Be��>@Tc7n�.*DD�b$^	V�@�m(�MK��x���f֑ �6;O�ܒ��K,[��@0��h�4O���K��?)Ӡ7��<����?aB�A�}�z�{�.G-O���C���?����?�����礪���ty��'�(њ��

���� �Q�p����f�Mw}�/j�fo��ē6?Ԍ)_��pq��N�����;?���M�1Dl�(B�X&��"A�mZ�Ll���H�D��7BM�)��DZ,SJ���'0��'���S�$��֕��@	C!^v���П���4<p`�'��6�,�i�)�����RxBu�}�����l�Hj�4/��v�d���a'}�t� 'R���|ם ?M��3�@�5L�����&]j C|�R���͟���Ο��I֟r�ɄS�ܔ��E�u9Ī�hyBai��]��8OJ�D�ON�����Cԍa@�Z.]�����
M9Aθ�'�v7MP���!O<�|*�,;�r�"�Y�"gVA�&y6`���i~B�L�n��IRB�'��	�*�� ����x" ���ϟ#�`t�I���I��\�i>y�'��6m�~1󄌌&�2�B�l
��`8� 'W�H=��U�?�`[�4��尿��4ev"Ń��G4i��2���<�U���M��OxR��ܝ������wt�x�$Nٔo'zd�#�3��1��'�B�'�']�'�(�Lڄb
Ak���m/|�y�1O����OTm���>�:қV�|2d�a�@�ځe�Z6"�� BI�Ht�O$�$i�󩎪7|7>?!��0:c��{�� ,3`$Bk_>d�l��"��O�	�J>�*O���O����O����\h�� ��L�;7��x�n�O��D�<ц�i0@�'W2�'��S�?�RoB!u�:=����$
l�:�����M׷iȄO�SG�h���1�H����1r�Y`0!�j߮�<?�'xԮ�����J�0J@���NF�:"�G"����?����?��S�'��ݦ��$�~�t!�D������Ǐ)fc��A�&�D�A}b�y�Dp�wbFj��)��I*e�ftʢGT�� �4��2�4���@��i�����SԐ�f�9,x���c�6��Yy��'��'A��'
�P>�Cc�CǮL���Z"��ܘ�@�1�M��&��?����?�O~���c��w��:'��/}ء V�T�v�����z�D�nZ���Ş.o���ڴ�y��ƴN�pAH�+U�R���6B���y�	T�Z���mb�'���؟��	�rUĜR���"-�V���}\v�����,��럐�'�(6m¶^�Z�$�O���R>M؜���(T|~��P�ԥ�:�X��OܼmZ��M�A�x"�="d#j��i��d �hU?����:u�P�d��*rΤ��h	���~�&�-5����R"&5"F�J"*"���O��$�O��D3ڧ�?qc�>-`H|z�o	�[���;0m�
�?	�i7 4�A[�x�ܴ���y�n	4}�Ҽ#�+��X�\2�d@��yҥm�xtl�M�����M��O� yt�ʁ�J��֣0c��X��B�tX|�� :n��O\ʓ�?q��?a��?��I4i!3,E�^R���C��[@�-O�lڦh4&x�	�	n�s��s��>3֐j���?j6��v	����X���47Љ��OCF�"g�8,���;e��!g�DPs N�w�&���_����`:12�Co�IFybh�ZA\�ۥ	D=%p*h������'�B�''�O�I��M{�<�A`Ժʌ�Z�N�C�82�i��<a��iI�Ox(�'��6͈��(�4-���81M �	�%��ܤm�DZ�, �M��Ol����/�j����w�-���3��C+���a��<	��?Y���?i��?���� T	\:b�M�KW�	��X��y��'�"Fz�Bl�!�����4��1HZ4�$&3\3��s�#_�� I��x� g�<�oz>%���զ��'e��a���'�l�,� df�%���eRX�	�`��'T�)�s�H��J�(�xq򰢁2?���� �!�j%�&�X+W�񟀗OP�������T�br Y o����L}Kx� po���S���^�"$2`H �[��d
DgS�&=�=8am߄i���[��3|�b^|�䈸�������P��8B�ɕ�M��f��3� �*Cj�|�0Y���U7_�f)+O`o�v�z���'�M� ����	F���]�pb��U�Ϧu�ݴu����4��$�DF(�+�'rbDʓOb�0�I�0�0T�v,ڑ�z�Γ���OV���O���O���|�Q�=f�^h�ɍ����7�B�:��D�O���&�9O>�nz��3��?B��RqטrH4������?	�4�yb^����PXŁ���	�_y6ċ�k��^4p}����d���I�hq����'1*,$�������'Q�ES�%�`�R��$�:60����'L�'U�V��9�4������?)��8�Q�G�>&�P��1Hi=�%/�I����O`7�s�8�'�����k���r@G�*�q�O�ӵ��3��TТ�Ɏ2�?���On8����|���E%�M��� �O����O����Oޢ}��j��I��f��T	f�M�z~l���GP�6E *��		�MK��w)�ht,����8R
������'�J6��Ԧ����t� hoZr~�
�� ��ӃF��1 ��3{����8z��+��|T���P�I՟P�	����g.	�EID��7����U��ny�{� �'�Ot��O�����F
h���"G�E� ��ȉ�<Ҏ��'�7���!��H����P�?��U�5�6���Ǉ�%u��仢��
ǣ�-v��-d@ԣ�N����[�GQ"t×(څO|A+�V-趥�����[�"�$Q�a!�Ӆ`Gr�Y�JۥCG*!�Q/>���5���C�l�4%�9(�r-�2��h�cj���T�T&f�B�ѓ+K 2�.��m��I�@qRf/8��0P��h�Ը;$� k�z���Iң֢��e��Ԑ[�U�|�m*!��7$AnA� �c<��jtL߹,�r��Qc��'h$p���X�H�ܑ1F̔�2&΁�ƈ�,�R���`u�d9�#c�c�@�ҡ��/^��D�خD赎�6"����q�6�G�\"E�(v����5��^}��'v�|��'w�J^�$��!Q�Z1��S�h@L��%ài�6M�O��d�O6��O��`kC�O�������c� ./�̩�3� �0L5�'	k����>�d�O��H�RV���x ��]�Ȼɉ����%��MK���?9���?y��	$�?���?�����ͷDrr�!vl�#0�R疭6�'G��'���8f����������c��)G��8W��Сp�Z�X��f�'�c��:*��'��I�?������0��y����eR��4�67��O��D�[i���f��I͖+8@�f�<|�����8z����N�cr�'�	�?���џh�'p�Y�b6�u����e�,Tk�{�ˆ�B�n��y����O�=��T	�Ԙ���A�r2��J!�˦e��[y�_�)���Zy��'��D�U����SHD�}:�5ae�ͼb�*��<y��?��'�?���?QE,�Oꂝ���@+�ԋ�2;���'?$a�R��q����'�ē�?�I��+k�@�f-E:t1�'��.�^�H�O����O2��<ɦ"�\�H��B��FpR�*c��$ ؉�cX� �'�2�|B�'���ݪ,Y@ Vh��֠0ǁ�&�|��':��'��	~���K�O .U·�4jT��Hrb��b�x��4���O��O����Oz�9#����p��+$U4�ЄR�2�j�B�>)���?����^J]�O$�	�-BY1`K�>���� c�ws�6��O�O����O���>�I�@��ȡ՟$�
1-�@� 7��Oz�d�<)��ZT�����H�I�?��v�l���J�/�ưH׋߱�ē�?i���N���Bܟ�8�G��0���U� �2��i���
t
�L�޴�?���?��m��i���w�C(Ɉ�+G2h���J�z�,�D�ORd�,5�	nܧ X�@�$�9#`�hƠC0Tۮ oZfd\Zٴ�?���?���/(�	Gy6GJZ`��?VQtu�Ҧ+�T7M�e��$>�$)���h���e��lTB£cR8A��ʝ�M����?q�<��]��[�h�'���O�R�ς�m$��qC��saf�`��i��'K(b@L/���O����OV���Rg���b��B76�4u�$�TצE�ɸ�|q�OF��?�O>��+�R�cm(=���l�&Z���':`����'��IƟ0�	� �'�H���9 ����0��,x��Jq�ī�x�����Ob�O����O�p)UFͮR^e[F�"C�%��΃=_ВO��d�O��$�<�'�N�I�bڭ`�(ÖYtA�E�x��\���Ig�Iӟ��I1����4LX{����� �C���r��O����O0��<Aɏv��\{sdX�m��ܸ��Ǣ8m�Y��-ǂ�MC����?I�}A�Xq�{r [��"|�ũ����"�� �M���?y+O��R���K����s���M�xjq��a޲E��qÊ=��<���L��?1I~z�O�z��bE��*��D�p�L��޴���6;*�oڐ��i�O��x~��5��}pS��.%�v�����M�)O��`Ť�Oܠ&>�&?7�[1. ��8Ō�%y@�x[i�<nZ76zx޴�?q���?���v̉���@�}\� A!OZM��q)G�t 7�ҷd`��$�O,˓���<	��$S�1H���N��J$ȒD@2����i`��'���q�PO�	�O~�ɕ���Di���H��։cF���4�?I*O��p�J�}��'5�'!`�����#ϩX��x��^�v��7��OJ\P�L\�i>��IY�i݉ rG�h�r���Eʎ5���9�#�>3@��?M>i���$�O�i����2�i�e5�t�dj�-1�ʓ�?����'^��'e:5��N6Hdx0���Y;V�i4�GHf�x�y��'H�IʟLHƃ�X� �8�&Υ*5������hйi=r�'�O����O���CF�;ϛ�
�5	�N���������?.O.�D�^�r�'�?	X�ډjɂ$�����)R���nk��?i�d�:T���q�I�w��ժW�	�Vy�h��ұ��6�O*��?�E���i�OZ�D��klC�=K&8�%��wcN��aJ:7�'�R[���.6�Ӻ3'`�p1���� wx)�L}��'�I���'��'���O��i��Aw/���uy�7�0d~���D�<� Jz���'L ��a�Yj�|� c�	HL$�mڹ���	�	�<�S}yʟ��iqD[ 0�Ƭ�CΗ�H����\}J��O1�h�dP (�:	zr��=�T��b	��l�꟔��ӟLQ�dٛ���|���~�F��2��A�`M�>=�6�j���.�M[����$�S6(���y��'Y��'�ʄ��+0 IX#/�:+�4pf�vӰ���?j4h$��ڟd$��݈Z`|��	�x�lq��F�x�F����$�O����O��e�()wJ�X��	�O��&� �ےk����'L��'�'M�	)*��5s�@�	b-��P�B�XJ��d�Z��0�'"�'��P�0�������d�ƕCa.�#��,;� ���
�byr�'���|b_��2����9�%���lyF	<7ص*T�����$�OV�d�O>ʓ�,�Ж�A�5�Ι�$H�Ex���P�L�u�$6m�O�O ˓RV�в���(h�d*P���#@n��sǉ`$6��O��$�<���L@I�Ou"��5F-����0{g�۹d�&�QHR����O�˓}`��B����'���욿g���mݕ/:b�AGU�����O��HC�O.���O���⟶�Ӻ3u$�Y��&�=J�P\�)G���'Y��-u��y��Gӊ	�u�4�W?v^��;PL��Mg[!�?���?����
/O���	O�D�"�%bk�E(p�S3ga,|�ݴZyܝA���N�S�OW_��xJ���$uԅ��I�:|T7��Ob���O�����<�O��p�&!B4��+܈����f#(`���Hg'֝&>�	؟���$DLڸ�ЍC�N���#�#:���ܴ�?y���	dщ����'��QZA�O i����p�0Y��$�eL�j}b�]#QRT�������	Qyb��!z2$PE�V��B�ÀS�nY"I#�$�O��$2��<���9� 03�FΗHF`��B]�B��?Y)O����O�D�<i��+��	A�AF��C�H0 ��@�J֩*��I� ��J�	by"�hy��H`�Z�I#���)�����N8듅?����?q(O�ѹ#e��d�'�Z( �Ŗ�g�"�����cV�hV�e�p�Ĺ<���?���~�d\ϓ�?1�'���c�l��Lg�*:�XU�ߴ�?����֔i�^U�OZ��'�t�R�a� ��I4���Ef�����?y���yҊ�m��^��'"N�T�C��q�ܸ4
Ncu��l�_y��3Q�d6��O����O���DL}Zw�[!�� ���H�&(i�ش�?i�dK~H͓�?.OB�>ʂ���)����HB�M�Ԩ` a��08$e��������I�?�ʯO|�P�^���GĎ\�|0d �B�y9P�i�
�a�'��'��z����dQ���S�Ūbi���֊#���o����I�ԫ6D�����<����~BL�~<`����T:n���g_1�M���?���x�~5�S��'�r�'}�E�3�?�>��!�� �H��j��dS70���'����$�'�Zc�,1�O	�_�2]�b�[PK<t��O�`�e;O����O����OH�$�<��·RY2���g�,B�a�o�IF�x�U�D�'��T�@�I�����-4Ad8H�b��t�9�<�I�4�Iܟ��'|J��u�x>qh@a#p)�NT.���.v�8ʓ�?�)O:��O���U���
jx���(͘}�r����;rՔ��'���'f�\�PX&J^���i�Oz��6�H�p�<4#�Dj;����䦑�ICy"�'1R�'�^���'��7��4��N֏N�t}����F9D�m؟t��ny2D�D���?y���2�H,%�޴u'�-XUNGJ�"lu��������8§�q����ly�ݟ8!"�
�9���#��� q��2��i��	F�y�۴�?q��?!�'3q�i��#k߬� @掍	���ȓg�b���O���t3O��d�<9��$�W"���#�ɑ7�L	��k�MCCj5���'���'�����>.Ob1x��/
HUaQ���h�������R)h����џ,��B�'�?B� �Fn�֮X�i�&a���}I���'�"�'y��(5@�>�.O0����[E�Y3C�e ��
4��]�!�fӘ�D�OL�D��OM�?���ΟT�I1g�&��#�*��ϒ0P2��ش�?��.�A��Ly��'���̟�(3G(�a�ǚ����@�]�uD�`cb���?1��?I��?	*O>�b�OѵBע�bkROx�PrX��!��>�,OB�$�<���?����|Xg��%��`Ȱ �P�a�# V�<i*O0��O����<�C!ZL�i�| 섹��W�f���wJ�W�_����|y�'v��';��!�O���V%BXTE _�(�b����M���?��?�*O�����\����5��
�H`,����/�ހ�sBO��M����$�O���Of����?�q`d��j�w���`!]z�m�ş���Ay��Z8�4�'�?A���� ��k�(�-����4��28^8V�h�	䟐�	[��T���'���
�G�-KSe�&	�,܀w$Ρ`���X� �#�F�M����?A��JvT��ݪn�B�# '�}�\)�AH�d7��O���M�\��,�$7�Ӑ[t���d�*��DlF�7T7����.�nП0�	ğ��ӛ����<a��>C�� Y�%�4����h�t@�6$0�y��'@�Ia���?ae˄N�>�"�H�C��������P5�&�'Lb�'m�y1�Ŧ>!*O�D����GL�+=��Y�D
�n� �Bp�>�/O&�2����ݟ��	���]20�e1�N�#��L� l��MC��p�l�YUT���'��[���i�u��AU�RPBa����#k&�x�&�>���M�<q���?���?Y����d� zS"�q(�<U��Uȓ�ԫ>��dj%%�[}B^����^yR�'�"�'�q�� uZ0�X�gA�b7|]�E���y"U���	��TybĂ�Y��,P��5��(G��Έ�l� CE7M�<!���d�O���O<�(�:OL����:�����R�
1���Uܦ��Iܟ�������'���Q�G�~2��C�*�/XtUUC�'oI\ɱ�զ��Ijy��'���'Q�:�'�s�#��R|�T��)��O�&�i�B�'��M�α鮟6���O6���70��a�
eq�lҁ�Y,j̕�'Z��'�B�� ���<)�OҠ��� �i�m�3��&{
�*ش���BK���o������O|���}~`M�~˘�9se��4sJ�S���/�Mc���?�����<�M>َ��ۿQ��!���,7e�!� -��M����.��6�'���'��T�>�ɾQ�4�#@%�ts2���HRC��ٴ��͓����O�⌀�_k��wA�i�'�?L�l6��O,��O�R��BM��?1�'���$�)fB��LӄD�F�Aٴ��M��M�S���'���'�>!R��EN��店$:PI�ԙ��d�����<v�b)�>a�������7X�����>'��i9b�C}2͇�A�_��I���y¨��
��U�S��\p���Z��EQ�0�D�O���*�d�O���Q�/�ҁ:�EO
)��@�B�M�WpSU�O�ʓ�?����?�+OH�����|:OP!�&r�"��	� ����l�	��$�H�I���y��f�*cŚ���9�%�� ��b#b���$�O<���O�ʓ[�l x&�������y��E��~H�%,�
)��7��O��O>���O�uJ�c�O��'v$�$�5=v�1Q�&E��=�4�?9����$��4&>q�I�?��MܵZ ��(]tڸ������?!��&Ix�����䓂����
9N�X�E�G-s(�`��!ǻ�MS)O��	���Ŧ9���.�d���Q�'�� W GhBGÑ�1�}�ڴ�?��*h�����OH��"� Q�/���
�?)����42n�$��i�r�'0B�O�b��"��I%L�<4��G�&�EQa�-�M�%��?�L>����'�0�R���
u� ��h� Q<V�r�Is�����O��S�}/�d&� �I�����]՜�Q!�>tv�Ab��2aB&@ns�	;/����sy��'���5�Ԉs)3�Ё/*�l+�ğ��M;�r/�Ǖx"�'��|Zc,����.t^�1ՠ�7R�h=�O�E�3��O���?���?�.OR��ǂIx� ��H�$�`����6Z-H��>)���䓘?!�� �ڨ��d��S3�-b¢�eҵ�.�<-O|��OP�$�<��L$��3,��J��/'ԍ�uF��r1�	��xD{��'��@{�''X�"d@�W� ×�O��1�cӆ���O���O`ʓ5�6勵��d�)J��0 �ص�<$���1M�6M7ړ�?᧡L��?Q���~ªJ(vH1���(<��lʠ�M����?	+OLh�G%IB�ß��s���# 1N�
#���$�1׌=�I��l���Rǟd��ly��np�u�2<&X�S�L(�|pz��i���'����'��'z��O2��5&I߇[�Υ�@(�:d��H[��
��M���?A&�F�Ԏ��<�~Rg"O�8����Q��UD:���W�����X��M���?����J@�x�OG2096GJ�t�b�{�c�v�Dx�t&x�Jh��	>�	�?c����)�J����� '�Y#�ʰ8%z��ݴ�?	���?Y�#�?!����I�O��ɦJ��`�fʆp���G��*?ԐQ�yB'<;�*�`��O��D�`t�IA���RAP�ǅ�La�en��T�V���'t2�|Zc
��K�'�f\�Q�G�g,.�A�O.l���d�O����O"�S`�q�!M	y��m@�JTVn�� ��ē�?����?�dpaKe8_�,D�D���>�`��q��?q��?���?�o����œ �p�pg�*'ZL$�L��M[*O��d(�$�O���	U,��i����W�ˊ�����+�$�8�ЯO(���O���<�2��4�Op��E�5JH�1�@�����c!�}�H�d�O⟘�g�2�ӄ�liH���A�JT�F��(>	�7��O����O*���/˧���&��#��!0�0�BwNKZ�bQ��U��柰��t����i �~BAD�k3P�A��:����@Ц�'`*DZ�i�꧔?��i<���#ў ���ą���n�:7�O\�Ĕ�"9� �}bq��"��]	"d9'�R�Z�����c�զ)�	ʟ�	�?�J<1��r�� >���c[-0)C0 + �A��iv����ğL��D�='��r�}@�p�F���M����?q�~�,S����Or�	(O��gi�n	�!���H�b��5�9�Iҟl���d#���UzL$`��0jת8{��7�M���B�Q�q�x��'H��|Zc�z��q� ���Cq��>�A��O
����O2���OJʓ<�Љ��d��4MfͲC�įNc�`$�FN��_y��'���ߟp�	��;�I��� )��焗 -�QPEBo�@���|�I��	���'�hU�P�{>)Q�3t0�e� H&�t��+z��˓�?�)O��D�O|�DH@���I)K45y��A#��[f/U{}r�'�2�'��I?@lfȪ�F�K�%ij���Y�w|�ٳi�	^٨�m��l�'�R�'��K��yr�>y���80�vi+rj�y���T��ܦ������'�7�x��'L��Of��Sp(	�Nࠤ?e�:,����>1���?A��`��	̓�?I*O6�/���i�䍪sF�1��ÖaѾ7;<���%�V�'���'�4�>�;-�ʼ�e�ȁIӾY�#�V>Zt�1oٟ��,/�#<��d���}��Ayr*�7fJ*��U.�M�5�]�RL�V�'���'���>1,O��K�G%��uQ��A�>Y
o����St�4�'3��)�OLP2!�Z�� ��i���[ڦq���X��0���P�O˓�?��'e��Z��A��Mq!A�!?@<�2ڴ�?�*O<p�4O�ǟ,�	y���$�>�����1N��s�R�e�ɻoKPq�'�"�'�?yH>���I?H��nA(w��+3����I�fUbc�h�����	ٟ���9Q&���#
~�V` @���A�Ly2�'S��'#�'R��'G6p���w�ҼBBC�/"`�P!gJ�N�\��O<���O����<c��
MP���6 Yĭ��-�:ot|�!��&L=�f�'���'��D].<��ɭ,c�
�a�'���@�Q���?y��?���?�fFH��?a���?�
0�8� �02���i���C���'�'�P�lr"A1�$W.#�Xȣ����$ш��!��k��~"�ֽ)����%�4
�ƫ�y2�%@\&��m�{���! �X5tp�M2�e��M���w�KQV�G�#MG�{�l�j��Q�R?`X��r���DMle�k׭wdD�{�(�LvB|��CY9D̞���Q�z�i$�� p%���mܻ[<��t- �X^ܠF�[�5x�%��W�`7@�s~�`�aA#>�ʑC��Cư,�aӪ]6�$�OJ��Ov��;;6�0�؛67 �1S�̘	�Ę��fW�10R @�
�\������Oe�'Ő�ҶL�x76�+2�I;��Ҧ�U I��\ɔ�:`֠S�]�I�x=��+�|�E�%K���݉W���2⦋�W���G/!�U�Ie~b�^>�?�'�hOYPv��:)���s�㗶U��p�"Ob��V?M�(I+�!����|�����i���?�'�\5'��xה�W�C/-؜�f$��S�
��w�'�r�'Vr'p�Y�	㟜ͧi����N�~�#���~����`D���\8�V�R����ϓ&�l����ڇ'�`٪��$utt�# m���I��4
B��;
ϓn��(�����8���?�(țt(������o�'��Ol髧K� n�6YYg�
^QQ@"Oq�����Ii& Q�1˂��M}BY���������O��cegK�?D�fN�l	�7��O��D !��D�O��S֬Sb�|K�j��5�
T�OgF�8&'N�����b,6O�!���(V��u,�*l#����#>.i��C߳.��i7��>�p<���Ɵ�Ity�Yr�j�!��*�4ੵ*B#Ϙ'��{���O� �	mj�\9j	�xb	r��Px�Bǻl���嬂��xtC$8OD�B>��ڴ�?y����݌?�����gW���V��L�+�)��P&��Or��P/B�l�v@�7�~�[>��OG�l*׋^�+�:���;2�O�P����S[����L�~ŞU��ڼS�ҹa��?�ɱ'�.(�tj�퐈aN�A	(}��ۡ�?y��i�\6��O(�?90%�
&}Yd,a�T82h���p�H�'B�^��g�S���Th�OvP�鐄Z�;""��<Ɉy2�iv�6M�OV�lZ�4R��@ ѩ��ª3yD1AaT��M����?���cF6�FC��?����?���ҿ!�B!]L����V�x����N
'Dh ۶縟��׍� v�$?c�Z'׆z4����K@/�y�GչD�m�T\�s���s�̒Q[��>5 a�<ɖ��x��#ՌX�_dT��$�^��?��i�r��*���,O����5V�\iBA$	8W��i�.Z�����>y@�D9��ɒ5G\m`��c��B��q�X�m�]��h�DP� ȲB�0G��G�� )���� D��Ћ��u����f(�ZMD�>D��2tdѦd/�=k���%8V�"�7D�,�v�A1��t
&��2M|���:D�(q� K	i(���JJE�AKk9D��;EJ��N�$ܩ&����Y�c�6D�� $�WB����#��<�D���"O�i�M�
�!�`ԌE�~��"O$˃��L�ddO�mrx$"O��.CҶ��Ʈ* �����"O�1s  �&����N˨<˄��E"O�XQЌ�^)ld��k
;Pj2-;1"O䍨C��BI9��U�-N�T�D"O& "��_�9r�"�'"I�}*�"O��щϺCd
1��=v+�ѡ�"O �J�m�#Z�|���	]�vA��"O$��H�<P�P���nH>�X��"O�J���T�f�
Q�e����"OH�!b��kj�lZ�
���@r"O�-�q`�3�L�
��a�h�i�"O����]c�>�; �T�X~z%+�"O
I�G@���@��@�s�%��"OF]�0��=�(���A�"`[d1�"O�Z�GL�?�(��`�:n^2P�"OP�p�̓.hNt)���
��ґ�"O�ْ�5�u�MP���"�"O<(J&)�6N��Y�V��yS�"O|m(�"�'o�*�Ɔ���"O|EC���+�f5�Re&k�}CA"O<�i�>/Vt!�qi҈N�^�y"OR�Qd.��Hb��kt�<�dղ�"O.C�I�\���:���,�<9kS"O�4Y!G�.y%�Ī���-sBdؤ"O\�p�ۂ/�Q@�n�3Wp|�A"O�)��#r��! �ѫ"�f4� "O�=�R"�w����KƝl�\��"OP��Nٛdv`��Ȣ��#�"O��7��פ���F&$�J(kA"O�����#&��A�"�����c"O�A@��r��B���̌�R�"O�Y�%�5R2��넏C�<��"O�0a�_9G����G�#|<��\��s�j2�S�OU��+���H0̴��Ȑ�zR,���'�D ���F�/:�W*(-]>�I>Q�**�0=�գ%���kC�V8;�A�!��M����U��Un���ŉ�
TȽ�����n8��&u�u���Ca� ��v���u�ER��i>s�'�>׶<�p���y�6��� 9D���v�C�g���O�A�>!����<�Go>���(�xIT(�<W�
Y�R���y�$"O j�jӷ?B�R��E)r�n��2�|B�D+v�az���/W4j�S'�V�lh7�{����9�n�bc*�0���\�j�L�A�<Q�"5X���#��.Q�	Y7���'�pub6�S,u$.=���޴%�hI�N3�C�ɱ��@*�Fɠ"4<	�A̘
v<�!�����i=Q�p��F�K�%n�0�7f��x�!���pf�Q+I�,�f ��PXq�'�v � �'S�Y��(�x��&į�~I��'[�0����`y��,�.i�b@�ˎ�y2�"L�ű�l�rvl\�F�G�y����2^������,� f ��y�,[�x��q䝰ZL������y��t�~����C!? �A@Ȓ�y�H�(�B�k���\r�g�H��y�e�$N��	4��� ��H���y"Y�D�y�%Q
hݢ��Ѕ[!�y�+E�<l*=c�e|��A��R�y&/wU�t�AÝV}��'�R!��'�txjL<��T0�.�fY�W�O+.7��{WJ 	����S"O� ��qG�*$:E��i��\�tԁ1@���!�0���(���)^�6�yr�Z H�����h�DB䉱T�<,��F2V�0�O�}85�'d�'+����!���R7C�&X��Ub�4=<��C�;|Ofh�C�>եJ��M����UZ| u-PU�$�1��a}R�J'<'b!��i��\�j$a#���')|��L<e&������� �|ՠ)�J(Y	`"O�̱����u^|��.��R��Eo���' ��P3��H���]5��u@ӂ��c���hQ-\�"��C�I]6�iE�<F;��h���$�打R<������6ZX����Z�'񾠻冈�i}!�$O#R)� �@�7��-B��$~X!��[=��t;�V�yL�(�A*�!�$�(K}:="�%N@f	�e�N[�!��$s\�}������|℅�/�!�$ܽP�\s�JE��U����T�!�D���t�6��%�s���X�!򄊫U� ��V��c0J!�D -i�to��V��a�O�<<!�dO�e�5k�i��,��l'��6!�ϗD�:ibpE.2�<5!�e�72#!�P�;�`���20�B1�J����y��P 1O�a����RJF;E��)��"O ����k�x`�IO���z��>� ���X��x��$��y����ӳDLd����yr���qB��Q#��G�NP���0gxQY�<�r�����'?� c�Ο#�Z "��|�J]Q�� �O�!`���Z��A�Մ;�l�%"�:��3̓- �Lڵ�'и"A�=�aې�/9�"�{��� i�n�s�öd��bE��|:P�B�B����59�Փ��x�<�{/�Q+��7�����uyB�X&\��Q��3��B̮~���`��3"��(�.!W�&��UmN��!�D�k�3���(	���u�(K ���V#L<�n��~z^�Z�e;��ON�c�O֨)���1D�z�x�oז^D$�QOV�*�̇%-(�:�h��`rJ�e��V �Ԏ��J6�	 �D�y���8ŨO�)xH�7kIzQh��Pb1h�;��'�<XT�[�XE"�G��M���P�X<BH�'R�<�x�Sᗴ�?�E#�B��l�V_8�2KY�_a��b�o)?�Ei��twRɢ��ǢM
��F��}�f	Kq+-�d�J>i�dI �LG�HxZ`*H�y¤@(ּ̉���?��1Ҥ�̚z����g�Ӭ����7�-�N���4�iR���'<�!��,��X��T2[LD����u<� �[\p�A*�P+���`�X2	VRL��	ߎxd����W�K�$�d�i~(�����G�	����
`NI�S��X�ax�C�035 qCuF��n>���+��,��K��ِJ�yA�fޤt{��;u�/$�Ař?4RjdA�@J�����-4?Ʉ@��j��p �)B� �(9�NZ���O��9��b�m.���c 6e܄8�'Wf<�� m��prF�"G��(ui�YH��	��)Yb�P#req��'R��Xr�M�[8t�P��9��- M�'C��i�a*��~�d��r^:EI��s#L ��,�G^�J`�P�,ыz��zҮ��T�!tK�����΢���/9`2p8�{�.TѨ=(�ȭ�����ݶOR�tK���-�@�b⃏,�!�$�wo&�+�
u�jЩu��%��'�z����ERs�n��~҃O�_50�z���Qn9��p�4�F���5��I�~� ��3��,���ELi7��	���Z�A��J�/.���I�9~@"|
����?�Al�9n*�!�W&Q�7��C��Q�c1�4��"'NV�_�J�b�F��)ݸ1 �cG;"d��A��f���	:�ʐD{kH�>>A�w9����*�0=������A��Ò��m��[����R��cL�sì�<X_�����i��8��ɴ+/�M���R�2b Y�*\=8�O X�"Lx�M��jj��r�E9q����o��ih-�@m;�8y�  ��{�!�D��τkEx-�6���d��\Q�K߂Δ<+�x,�2���$�|K4?�OҮ�˙w���(��&F0��E��D��	�'���Tݒ(�@��&�ݤ8WTH�0�dB�k��x�D��h�E��Tm�'�T\�,]0F����a$9o�p��ۓ<��� �% �|��2� ��a�l�'u̦�bT _'<��!P)�;&IFxP�d�
��t�ī�{X���'�N�vr̈s%��'D�So/��)rT�ٗ�4z���3'ƅ�s�FO\��C��� Mc�eg�V�؇�`H<QSF�??�@�`$��-R�`1U��=u�����+��P�&�6UޓO駻y���.�Vز�oA�7�&��怽�y�o��
N��`��[�	Z��F[|&)%���NK6���L�*v���ɕ�5��d=��p�)n��D��F�|-���,�1 �cA#|IzY�4��+[D����Ȍy��3E����
��AO XH�͚HM_x��s��dY8���8�l���H8Y��#�'k#K��1�
��<���}�T\�/�,K�u��"@>g%F�a�'c�hǈ�jxB��`��c0�*1��6h��/�J�> ;kـR��)���E�#нp�8W�>�l�r1"O4=Jd��=�҅�wa�RuBUFÃt�&�KK�tj������i�4a��t�תX�L����ҏҧ-N�tf0�O�u� ܀NpZ�i]N��[��?<��{� M�t�@cˑE����	(\O��ʲ�J"Z��������1@�� L@d�T-X�L@Z.r��M<h|B�BF�#"��a #A��N]�ȓ4���b�J�W�����؜h|J���lF��{�b�!k��̋¯ľtv����94�-�"��$2햰#A�e��?�"��#8`�?mB��YP��2��0'������͔%^хE�
S)�q�9���'!#�O�� �
7�4�j����
�^��1�A���b��E��̬}��|��H�����0��	������9�x��X�0: )lOD
�KT�ì�w�T�J� �sp�'�TU���+�DD�1TT���[>Xe�D�9?T%��)+�Q�A)�Zg�;P�[1jU�@��I��5�.OD�8���h�P��խL�_UܽCcP�@��͎.�J��b�*V<;��'ҧs��#�H�	!�5�U���*4�?�pV�b�?�.%��0Z��X�4:y{"�ڟ	�~VG��,S:]
�<�U�ߤ��g�*�2x�d��:*���I^�d����+����'��>���#�7��H�ܮu�ޠ��C]u1�l�t���G��'�(7a{�*��}�19g�ؗW�쌳��D��y�i�w��#<!��O�/��Y�!�t�L�m�{���ST�
s�8�jSM�PټB�	�?���,��C64�:s�jM����׭<w��qf�S�|4L{�c]�b"��:��\T,C�	�i��@ ����6͘�bZ���6^f0��CFY�)��<c	]�Br�	�B�����U Y�<�v��-�!1r�L�<Szeʀ	]V�<I4�p��@�A�U3Ut�D��J�<!���  ���!Z.��|�T��A�<9�kA9g�J�s��(2@=ʣ��z�<)��?a�pX9 ��*U��!B[�<�v�A�<8��ZSG�.�ʘ����V�<�bE�#T�j���O�806L0���^R�<����`C�ţ�
�5�̠ä�B�<)�"��k�P�9�E��-�mpF@�<���X�N��� &ׄ�@(��Xb�<	�*&c���e&xP� �G�<� O[]+L�Bf V 8��3U��Z�<9���!������O��t�aZ~�<!�*�7h�4�g��dǲ��NA�<	Pi�j	LCe�YQ�%�H�@�<ArER�0t�ܡ�!@�.�m��z�<������nx�i�>�jTq��\t�<�R�2eC*�{�/�R=��X��n�<�'��WLy��=+
�1r "T��	BKɫe{�)���f�P{`�;D���F�fR��Ef9#��@�S�&D�����ۼ^��tqD��4V1A�2D��q�D]�Pyd˵$�+�B�:D�+D���!�@:��0��HT�0�H(D�P�c��P�N�*�Η�C��Qw�2D��J�#��rtQ�b�+OD�<a�:D�@2�D�C��#��G���B�,:D�@y#`��t>mh�gN�|���*ǎ9D�Ԩ6��!�4��JM���`�f9D�� �5�����QZ/݄DZ���"Opt�#�35��	w.ɔT-H r"O(�"$��	lL�$�[#H50$"O�	��W
7u@�3�kD�@�T"O2���"FS� ���@�dXQE"O !oU�D�'�Ⱦs��X* "OT�:Ff���ȉd����"O8T9@�� �ġa�"���"O����&��}���@�S�s�Z�s�"O1����.�q��E�F)J�"O&e��	�Z
�Q[£Ǐ?��1"Or����=$H�#����F�`%�t"OBeS��ӫ��8V�	�C�n�"O(Qh�1�~aS�+�$d�x���"Of	ɕ�̺h�dH��%f��"O�@ȁ����֨��CW+�L�"O�aG(T7n �K��àl��B "O��a -��8��q//r�V"O�l�c垞!zR�3�M�aՐ�"O�!� C��k�(�A�Q�&D�D"O��^ �j���^Yڰ�"O�!'B����Ȅ-S�K��A"O"�aaXU:���m��>��e"OD�bC��
���I��;_��"O�kg�
5&DP�I�8i�"O��J�f� "E:S������Y0"O��A�	�RW,�맩�1-�`�"O�`�FX2o�����gS�)��!�G"O�x�t�J1q��"��X�d���'��%��+�R�`QI���0�'x�"�ڥ4O�1,Ҿ>
ZE��'�.eZ�j&WnJ�9��/>�J���'yHl�#�L9b����Ŕ;<z��+�'�N��.VS�^��G�#9�V�I
�'�~���h7m��|q́�>�,�1�'��w�Qei�I���%1v����'-T���n;FKX<P�Z�R�Z�'# 10S(_*j�kWeW4NL���'.H�F�!h�pegn�?l`��'G
���I�m�F[Fl�*'��#�'Wb�%�߇S�T�dH
�i�"E:	�'kZ@rw�%��@D�C�s#����'���УO\�.�lx�Β9p��$��'d���.��	(x�`�G�=�
Ւ�'�\LQA��l��4"D�/:4�8��'^�@i'�N�/��%"��܇5�
@�'������Xb
})#N�3,��q�'R�bI�1XHi��]�.>�Ɉ�'��h�FH��?0���\�����'s~tQF�
&wiB	��m�$P�������*��)*m�o]*��p�P&.�!�D[�c����o�+G|�2#�5.�!���dHl��j��\��a�k̑IK!��&ytֵE�S�_�a�TDT$�!�DA��9��އ9k޹�q"�?&!��#�J�$��:HUX��b��V!�DL<�.������/�����i!��f��{7��@�de#'��5K�!��2D7�}�EC�&<�Z���E��~�!��<H��en�7��m�U�m!�ď&e�Qq�B�<T#�X��
�e!��HJ���F;zr�x�cP��!�$U5'�1� Jjo��ҩĭ)@!�$?[E�8��g��y�����N͝F!!�� 4�ʖ�
>m1
�x�J�,� �I�"O���j��J� �3�G�>�D�§"O�iҗ�X����G
1�`����Iu���	��&
�����W��ECb�V'!�d���Zx��dC�R����g(�!�d�
�4\s��M�4���fN/L�!�$بs�`�,�6�@Ec4�P�]�!�d��O��h& X�G��E���8/�!���ʪ0(0,��r���J��Ҥ�!�����'�
�V�z1`i�!5�!��s.����O%Y�F@���U�	�!�߻��x��ށz͜Yxa�R1k�!���B��h��ޯ,X���9k!�	4r��3G.�5j��	��!2{!���a��8c*��:YR q�
"Fl!��o>XT�T :��!+��W ^!� ,r쵚@�N�@��1dˏ_!��@&�`��n��1(ZA��h�=6X!�V aw(qc�,ԅ3q'��!�Ps��S���T���oZ	�!�d�Z�f'��!��aSU@�[�!�$�2>�P0�0�/N��A1ae!��O�E��B4̘,i� ^7(:����"O6������O�ب!�Yi,�$��"OL�!hG�k�n�yŨ̬w�D�:�"O���a�W�*HE��҄%"O Q{ӌى\�,$C�M9~�>ŘV"OrQ;W��*H~|��q�.-�-H"O"�1�&7O�PjU��%�6L�"O�Hy�%՟z��4	Rˊpڦ��"O�I�v�ڬA�&9��J^���"Ox�6��o�~e�b������F"O�9� b��F$0�U�2��\��"O4X"%E�lԮ�3.Ǝ�2�i�"O8ŋ��NG���GB4���"Ov�J'f�qnD�F����I�"O�z��´��`R=6����"O��0�;�|P9�[)",X��0"Om����tm��Ԭ�;��U+v"O�% "�˅��m�	��l�"OHM�懌(��j��FG�bF!��y!���w�l��7�=�a|��|�#yUD9�B�?q��-�`H�y"�бad�  k�,3�|]9ceˮ�y�ś%�p� ���(U��(�A%�y2��M�V� Aj��k��Uң���y�Ʈ��!%' i~��뒋6�y2�]nAi����c�N��b�U��yR��Y ��T̀?/��Xy��
+�y��M)&8�X��O4s�̈�y� �*;[|�0�U�n`bwo��yB�O�AȾ����T�
3Hy��+3�y2e_&i��8z`m\�{��)c���yb.�8]��Me��f�2�
SG���yR�\<}6�@��?6�y ��%�y��3����)��t  B��yBA�b�j�Cu*�4�S��N��y���[p�9�&��fP[�N���y�ǘ����(�a�H��:!��yr�Ɨv��� �;=8�}���V;�y��3��� �i�#,���˥+݁�ybA'=X��5@�=�8���G��yrj�	l&��&L+}s�y���yrui��w8��*V(���p?q�O� ���Z"kY��Y��дY��9�"OV�ڦ�͛?|Պ�C�
* ��"O.I���J�V�%C�#�>\��A�"O���k�,"�x� �$
X�+W"O�\�Ǣ\�3��tC���*ɜ}3a"OJ�;f��XJ���2D�ih��Q"OXq��f���p�A!r��Y�"O
T����"�N��$E�5a���"OT��P���z:(�I��QU�h��1"O8�`$��=i��\4u���"OL���艥L������^ ,�a;�"O>��p�L�\g�i����@�)�"O�	�g��Q�X�36�h�!p�"O� #^�ZG��3 y�b��"O����(Q!�`M`q�E�ش�`"O�$�'!�A���"�!~�y�"O��Xv˝Tb�`�p!�P��9#2"O�I�� �:>�,�!�	h��x��"O|H�*?B�p��b V�2�"O�Qs��!���V��!��Y "OQ�2��'�쭁 ��,_�� g"O��`�ǅ�0����A��&дx3Q"OĤ$�ׂ?�Lz�LQ�*����a"Ob� ��x��Tp���X;���"O<AY'�T3hX�dx$���f1�P3�"O�M�OM#��� �'��+ hi�&"O��!�FYF��;�E�.5ٖ"OT� �C�-����&W\��"O�CEj��T��j!/��@�D�3"O<qb��#LŦ�"�nC�v`��"O�h��^�N��B�]��� s"O�z�$�&GS&�Y�KށE��2�"OR 2󋈾`��d럊,}3�"Ov}�0K� En�x���{�xyYA"O��IwE�=D�,="�����E�!"O��iS�s%�� ��^,z�(�"O�3 h 0i�Д7cO���e�"O�ع@C)#0TŪUG��p��!"OP�٠�ы�HJ`F7n���;�"O��� ܛ$��$�T�Hx��!�"O�ݻ�C
,{��I��.�"i��m+�"O.)�t�s��(1G�?X�2��"O$��ɒhI��r�K �8� �p"O*lhe�͊Z��eH�o�
@�9��"O<��N9L���j6ُ@+&$�&"Oz�pl��n�Њ%�¹}6��"OX�2���Y ֌
siѰf����S"O�$
�Aڒ{��|0`"���"Oā�P\8j�	��ሏ�h0�d"O\�������n��$�s3"O�����D��\Y��NI��s"O¥��E���:��_�%���"OXDY�%�(:��-soO 9�T*4"O�5cK�H�Ҍ ����(�m3"O�嘕��?�^�tOګCfH5��"Oh���IC
W�1��@"d��"O�p5�T�/	l�:Ө�� �"O�Xf I}�<4	�g�O�2Yrd"O���DaB���z����C���!U"O�B�!'&�c��$z|1(B"O�l ���	ca�)r̊���T"O�I#W��9W�R�ӄ텃����"OF�1�l�T�n�%�����"Oj`IE���̼�X�BԨYz��"O� ������3z`�H�qcC	���"O.�aw�ʡ(�+���_� ��"O��FBL_��QP+ɰG��a��"O
 	�B?�ĐuiD�c�XI�"O4l�6�@�.Mx]X@/�=VI�@"O8�x2�P�F��!QM��Y� 5�"O�(���A���땟%̌Ej"O�0��<�9��,��ȯ�yD˄�`���MD�Y�h��I�#�y��I�E�~X�#�T��prД�y2��|q���T�4u9�t !�D��y�-L)Y&���e�7��m��W �y���Hk�uB^{���$	 �y�X:c`Бh�A-		6=q�F%�y�h�m՘<�R���-��l
d��y�"I��BU��9}\��*C��7�y�J���tEJ�(t�D#�I!�y�Nn��@ '�'rO:4�r
���y�3`
�L��Ϊf$s2
��yb��*;,��J �`"(B�i[��y�KA�J���V�b�����I�;�yrlҖ(�x|��ȋ9X봴����y2*6K|:���BM�?����,��yr��"{~(ەl=m�\�r*��y"+�,2 6� ���%c��QAG�y��A�:d�9��_�f!Ӂ����y«A ,(���*ǺP�ȴ:�a��y�CH;/��ق�Ԭ(`q��j��y�ǝ���Xw��#�XH[�����y��ϛar�����{ؼ���F��Py��Kԉ�W)դk�H��[�<i3�ч3�� e�J���E��S�<�eo�) �n	���L�T�@a?T�4�G�O"��8��)A��A��#!D�<�u�Z�疝pʅAФ�#!D��H&)FK�P��P V��"*D�*2���\U�$9PiΑiX�Cj)D����րd��� �o#7��Bֆ(D��(�6q����
�_��IQ�8D��B�� �f5 c>v�����i3D�h(�Rl�TP�ڪ	�8L�R$D�Hsg+&��$�e��1 ah�
G"D�`�����;�%�R 
Su�%k��?D��c#��6�����L�y��>D��swI ITZ�Mިa���i��&D��rŃ��Lp�Ы/A�5�`ш��$D�zD��K�Ⱥ�(�=:ƈ�;e -D�,��o�3, �H5��C~Z1��9D�(��h�%3�޵���<�4Qx��2D���rm�6����'kY;>i�/D���#�.&�HjS�-	Z���(D���SE_�X��dI�f V$�m�+4D�h`!�ߍ%�����2T+�ءF�3D�D�($�%�+ɺ?X�̸p5D��	���
�����Z-|��rU*3D�$��#��'�<%��D�.�D���n0D�$ke�ȽR�Fp�0��G����k.D���E�PTX �G���b����6�-D��A 	�?K0\ �(J�ts����c,D��	݊r���8��U?S)�m+b)D���B�^�:>��Ժ��	2�'D�����/5���k�0?cz�kF%D��T
T�<DM�VMʒjA8�3��8D��Ça�o~��1��A:�L�q�:D�� Z�� �_�i=ԁ�"!|T�Y�"O\	��?"�z25"]�fE
m�3"O�0p�&E�A}�1P��Ύ+�01"O�*R�M}0�j�!\�}� ��"OTdf�5AP@mR�ÈW�D=:�"O ����4�d�K%�<� b"O�`��Kґ!�$e���T$��x��"O��3*��H�h�A�	�H��Q�3"O��"��^-n���YOF-+�"O�,�bBW�N`񠮆�wK܈��"O6HksB��D���G�nCH�6"O���,�:<���l�*1U"O��v�K��J1�&�H��\��"O�ГaB3����I�%f6I�t"O�)0K�V(@�!���m�x01�"O�5;��R?�q�07��1�"OH��5N�'`V���;fj�,X
�'�� x��Bm��,9E؉+���
�'\h`�G�9Q^Y��c�3 � ��'�`��$D|U��(�C�J�'�<9�E�':F��+g�,��`�'�pؒF��-U�+�%�"#t0<��'#$QS��[&[�.)F�k�t�k�'8�E�U�U�tƊK�y���'&|��m�aI���X't�B���'v"$b�搭}~�Xv��v��	�']�ĻBn�	�¡�U���bVؑ��'::��AS�, jI%T&D�r�',ƭ�V��l-�Xu�N
PO����'Ր��#Ͼ�3b³O��<z	�'��m!�j9�
d��˳?�8�	�'^��[g�F�oF4l(wgҜv�~݆ȓp�P5C�%xB��#1���A��l��zh
]pl��lJF-���X��Ň�C�&�@AZ+�����.ɖk��B剤�n�F��4NSr=��m�.p�C�ɕy.��� gK�C,p����gP�C��!gjt�`A�&|heE��lC�I<<9���n�;�>�7�_�d�B䉓iP9xw�!��P0SG]d�B�	�+P�}�%�U�R�,�b��B�	�pԥ7,�96�\��V�e�B�+k��a�2���ep ������NB�I�U�.���P<Ҵ�H�f��+�$B�	����]�S��Uzd	�c6B�� 7��xc��^B�~�"Ƀ�cG�C���@��ym0�!G"_܂C䉇!~��oTv�Uf�ZH�C�I$C�J�;���@J���D�١5O�B�	�Ilp�g�2���e-�#;/
C�	�#��h���"*)���.�8�B䉭L��9���"_3`�ċR��B�	)��#�'ڬ%q2��Sa�)��B䉷�Ԉᷫ�*{��tHJQ+��B�	b�m�W��8��4�	ۯb�C�I.F9h�h���9��q�D��N��C��>x��$� -��*A�q�	�#s��C�I��(}[ī�]���T$�![(rC�	�(f,��|����/��wdB�I�t��ڡ(s��2Ӗ{��C�I,V�����8��Xp�O�J��C�	�^d�)U�#��"�� ]���0?фo�-פ���M���a�s��t�<���҈G�|�҅ܓ�0`�"�p�<� ��I$�ߚyw�4�D�&"22:�"O�%��ՠؐh�b
]�0"O��)���w�^�)f�\� Ӥ�8T"O��T�	�^T�9��"��{f�	�O���e�	#�였��ޠSf ���'�
��gS=X�(��`ьJ7�{�'7Ĝ�ӧ�(���i*+B)��'�4���9�x��)�$"�9	�'���3�۔H��!N_/	��p�	�'<&,ۓ�� �b�f%R��5��'^�U�aã.EbP�G3BXTq{�'E�T�JA1@�9 ���6��q�'�ΔȁHԭS Q�#�n[�'7dI���^hxs���P	�'�.�r� ɁXHT�+H��(L�h�'$�qYƬۢp�"�z��%���@�<�QG�	��<����j��Ԡ"�c�<��!$|��0�
�z�f�p7�]�<y��R�S�� 4��N�<���d\�<ËU�V`�#D@4Md nY�<Y��D���!��l{�] ��HX�<F�בt�����51�X�dQ�<���6x�M�uH)l�d��7��x�<�%J��>����ċ�;3�C
l�<���Y4z��Dn
�K���bD�Q��y"���%�z=��J��ɘM3t���y2%�:8��B o�s�UXI̐�yr�aBE��ā��4X�.��y�d�p��Y>�Y��W"F�=�ȓ&{� G�/dC�0S�lK)&�f���e�2��_��n��7m�
�p��,b�,٧N��f:�� NW�bX\��	ϟ�����C�}R�n��i���rrB_{��O��=�}��cw�p��Kp����!^|�<Y��0d�D�!��6H����I w�<��͕$�ڝږEK�G�By0p�[�<��N(f�>R�N#O��S��]~�<ٕ�ՐO�A+pKC�b�\�cWR�<!0�I�M�:��1���|�R͡a%��T��\����+?��I!)��Y�¥B�i��$�Ŭ�N�'a���94�˴&��w��8ǌ/�yBѽ'o<����A,ı*�,�9�y"%�O��(#��:ݺȁ�*�y2KN*\�~���%�*���p��yb���\���&���ġ*@'��x1x3>�9�늕	T,�҄�R[�0��*n��e�c"M�%��C������d5�S�O���05O��c����4M�7"O�����;}�4�0��6s���sF"O�� �#�?.H诏B0d
���U�<� �4$4Ѩ��7�Xr�,Gj�<)��Bl�*�!����D��`\p���hO�'ca\E�f�:n),1�ƩɸS��ؖ'o��'/��$+��a�.%���v(�:��zR��A�<�'�:A�@�9e�[#@�y���A�<1�b�<&lj�
#7���i�<��B��1�Nh���R
��%�d�<��O�� �B�Ύ�|0ش�%a�<�� �P��©��"�\�ro�^�'�?)YC�ŪTJ�<Qw�H,c�
hz��,�d�O���<�����k����J?i�1Qj9"��1;�D%D�0롂U�v��(��Y�e&�`�"D�t�aG�<4��h1j�w$Q�
<D�`Yh[�RDIQ��
!H���m%D�� @�����g�V�3t�Q>.� �"O4�:�oN�[D�I*!�XC���b��|��'�t���l@&1:�kIe���1�'����%��3K�2H�nFX��J
�'��9���S�n웅g�K�"�{�'T�H9�ƠK�d��%F��6��}A�'�Fј��>zƬh;U�9.���"�'D�<�rB��?SDT��G���Ti!
�'M��s�͏?������6ظpH�'5�k4��h��(��.ۋpA�P		�'O萲����ڪ�2�@�<i$��'t���E����2Cۚ1ܭ
�'"�����0 9TXA�+"����'R���sfЬrܱK'U���`i�'	2@�Pϝ=�B"a_!D�ȡ��'5�-����N+�̬f
�}�	�'��37�*x&��#�^4	��в	�'
|��f5X�"�xCX�z��'.�	���:Z���b��Cjt���'M4!I&cäu�DyҌ�=5���	�'cq(�*�0��P��у/�T���'jD�� �p���j:*G���'e4����:H�\��t��7%��`�/O�=q���z����H�}�ȺN�w�h0{�/D�8�B��izr5���KK\\��N-|O�c���D���+!vXٔ��=c%d��*D�h��k��j��B��3s&����)D��X�`�'!:0("�����Q)&D�SħS�S[��[4�N��!Yҏ6D���D�;<a� ��E�|#�=���OT�=����,7��'f�*P�:��th�Ȗ�L��l�*!���p���F�_.�0Q�!��!��5n�mbfK	��Hyr
��o�!�d F� �£�@$l�0�kb*V8Jk!��S�F�J������\�1p���ZZ!�Ƕ[���"�M�7s�b�@�ʊ8Z!���2�6�;kJ�V�ڴ��O��i���'�
uY��ɝhϠ��W��9����'z!�Ğ�W,�B�ˏ$/x����8!��0va"�J�ԇ]p8��+B�H!���.��U���>2��a���|5!�$ێ� ���_mҦ����O�!�� %�:�k��>�D�sr!�ב?���Jr�7�(��K!mM��P:!����7X�����^�WP��0?���׿d+@���A|
��6�Ay"�)�'E���R4+�	q%L��ES�:C��`��:�C&?�V��遌xc`T�ȓRsT� H!x͘���l�Z��D��IIZ�:G��jC�����F�DrN���e��=�5A�C�u��.K/�����.	Yש�3��0�%��:��(�'�ў�Fx�&c��ҡ�
�����K��yR�1���A@�<3B��v&���y���g����-
��Zf�
��y�-N�[l�;'/֛nG�)��'��y�`�F:N; A�<�p(+��-�yR��,70�j�W�;g��(�.ɿ�y���;U�ȍ���(. ɤ���y�>A��Ƀ��4�&���g��y"%�)I��37nH�1%��+��#�yR�¾�R@�5�W9S����'���y2S�0�ؕ��X$E����"���y��[�h<\U�$aX9>�x1K��y
� ��	�mW�Ex�Az X�
rZ��B�|�'az����`D㊛O܍���@��y�_�0�b6�$|��I҆���hOq�
(	Ƭ�%/T��O����=�"O@ݛ�'6�H�p��Lp~��"O�E{t�]�_��tҕ��-B](�r�"O2ap!Â-V�K3�VN$�+""O��X7A�lӀ��YB�-���|b�'���#5J���O�9����6͐��!�CoI fFw�`@�Q�߼ y��I��(�L�Q�/�(D���p"�y�"Op����_ ���JˑEW8̐�"O\Dk�iU�qz0<a&I8r���*�"O5�Ί�P@����ҁb���'�:����{�&�ZG�2]�B)C�'�2���N�Ԝ�f��7V����/O��=E�䀪�f\��MU.1F�P����?���?��<�š�&EvL\�p�F&'j�{i�Z�<A���iX<��FOА)��I��K�<�Ӛ34�J��V�fPb���E�<�D��$-\��D��xU��"�Ln���?��o\XGJm\�pV��1N��5��ئ�C�mצW��X��,+�PA�ȓW��	�茳3�% VD�Gt���ȓOT�!��*B�JaL���VNm^؄ȓ)'�P�sB�r�H����KѺ��K}T�Z(���Eg��~�21��Ӓ'*�<�x�J�+[%O�2t���O�=E���/U8L#��7D���'�өQ5�'ў�>}8p
�=l�!Э[b:H4�L7D�x���KB�Z8T-E,hFLs66D��DJQE<b�ȠJ�C�Zh��2D�`��e[&�p�d�U�^�)�,3D��!B�.tY���F��$A,D�p
�呠n���i��Yʨ��$��O|�O����O��=yd�P$O�B��4L^"��}h#���?i���'p��`��ǲ�̜�`�L"]�ȓe�n��#�,hkn4diE;1��ȅȓs�D�qp���L�.�{��S6���ȓ�|\�ĤٝZ�x\suK�1{ؑ��9�.�A�g;�<u�G�ǖW1>��P<��'��"֖}k2쐎n_>�ȓ�������B�Q�"�(�H��'*�':�\"��O�1�&����hR�'��Y�t^�0�4�#���"�
�'�P�0N��_(�٣�N��y��Az�i��t���F!!�y�Gb��å��
w���K���y��H:\Y�)R��'p_��TbL1�ynH�t;e�Y�dlL��!f���y"
P��YeÖ,XZ`�Å��y��!
�h�x1��Wդ�3B*ׯ�y�	W1�s� '^�^0�1E��y�@
tH�DلbU�XO<`Q�+�yb`���lp�G�D�U�`�����y"�ʭ%H��[�K�29G�9��F�7�y�l�f�N=�E�]?,�	q���y��'c\�8j��B�bF�S!=�y҈
fi�x���tI.(á�R�yr�˨@C�9u�<j��Z�"V�y�A].����2FJ�`�@1���yb셍c��P:�(��-6��HK��yr+�1�R�`����$*~�"L��y��D!2�]a!+�$0LHM"QJ�y
� ��I֏
��3G\� ~h�0��'��3)J�9���P��8�e��g��B��%k<(�14���壌7"�C�I���ۀ"A�a�
��d��7g�B�I�wj�J�<MµJ1,�7@�B�;�*�y��(@�U	D�)c�C䉵D�@��h`�!�ʈk���H��	�j�2����Bw�B�T�J� ��B�I�'�����bv�9x7K�,���ȓaF$��B��<r�S&��t��8���pQ�F�D�����'�ń�	;��+b�8g!�ӫ7/*U�ʓ*�‡G�F�8�ird�<D�jB�ɑ*R� � W�&+8�0��1�VB�	)o�U�!)]3K���	1GđQ�����O�a0��ׯ$ʆ)W'��X6 D��%/�*B���aL�;'Ф�;D�,I��Ʃy��"�F\o���b�i$D�a�N� s�����3W\ Z�K'D�(Zq��+R�` �B�6"#X��� D��%�3/"<�p7-��S��	)D��"�a��W�@1/I	����%�O��D�O���F�1/d���T�G6`n~���&!D�����$=Ob�hA��99�n���,?D�\˓B�M�� Q)��m$X4�w9D�,Q���T��]���V^F0�D�!D���o�`�v\�ec3r��*6� D� 	a#`���� Q)Y5p�`�D4D��P���"N����iХ9X���?�O��d�Z��	Y��^l�|+@(����C�	g��\�!_�0l.i���?P�C�ɤ��H�4��\���%��v��C�	�~�h��5,Y�A�ؘ�bB�+_�^B�ɑ�y�
��M~���j�*G	*B��$>�FMa2a��M�t�B6�*$*B�7L���O�U�&����
W����z�`;�!�(�h5k���+J��	�$=��K���T�'b�QV:qM���Ê�{5ja�u"OT=��݄>�Z4y�@�$t�:�"O����4gp"��n�E�H�"O<�*@�֨�ȑ	5M/.�6(��"OL� H�h�8��%�˃�ע$H!�$�T���7m��R�*H!�I��d�!�s���	�E,q��˦EL�N��Oz�=�+O4�jU�(�| +���80K�hs�@�OrC�		���P� ٣6kbБ�FǛb�.C�7@^6Lr!/�_�Z|�����C���̘���S�S�p�1G�Ήv�B�	�O�Lzi@:2*�8Y��L6HC�so>E����?�p�Ŋw�*C�ɥ�̔Q�G��l��T3A��=�H>����J9""��ۅ`�Z���8������$�Op��'gǚWB]q�u��C"O8�k ��g(M�sI�!j�|@�"O�I���Z�zU��)�Iy�@"Oƹ�BO�����лd
>��'Բ�s���:��L����v�1R
�'�0��Ņ�\FeP��\�h ����*��p�΄�N'2�a �@�z��'w!�d�DZ.�( I�q�9��]6W�!���9�����ƘV<��	C}!� �ᤅ[����S�^�Y���]m!�DS�L�zd��܎H���aţ o!�ʳ`�b=���'`4޸XPb�t^!�� F�J�l�]6���VO^2��9��IH>y��6L����D�Z���bv-:D�����r�ԭ��>c�ĩ�Q#;D�@3fðzD�h��K�Ab1*:D��� N�}��"�疓b좥�e�+|O��<?�4�/!(�'� ����'i�i�<a�J5�h�f"_�Nn�|�<I�ϋ"dڅ*R͟1�D��a'v�<Id�(S`��)E.��v�.}@R*�J���hO�-��̘��Ņ��YD(� ��ȓvH\m
���w�r;��QRч�Ej��y�i��֝:Ao�;Lr�1���v~b���n���G�NH@�1W��1�y��Z7f��Tb�?w>�`&.��yrO>s+j��昤8a4݋e�;�yR ��	�nX�F�ڠ[�����?���0|"�$֣z�tQh�" �@��5`�I�<Y�l���x�Z`JA�(:�M���Q�<ђ�29*F�[`eڜP��x#Du�<q�J \�\�yA OH��IS�z�<�#���D0.�HU��3A���f�u�<E�Ń>�	��%4��rA�^����?9���O��2S�8"��Y�H��y�J!�DL�@! D�|}̘�rmU}8!�$RSG�Yd�r
x<��L��x�!򤀉f!01� Eי#M�r��<(�!�D/�dH2MD&=��lS���Rv!�Q�2����J�*
,"�FО1S!�-}>�`K���u&
�Ge!��Iy�ԉ�� �M�BdΟ6!�d��zU��wD�ٔ��:�!�_I����ŕ���h� ٶX[!�$�+�p�	��Att0��
�8^!򄜚R�(=�Q��xT8��f���!�d�F��)�cO/-�� ��Zk�!��úq�>@a�	�	[�`:��*m����#?(��G��="��D��\f�B�ɉj�v�Z��[�sVD�T�,�B�ɟ\&}��.ٔT��Ce[V��$Åa�M!��)�¨�!fĀ:(�'vў�>y+�&Q&eF`k�ɚ�`�R8y�a#D��5D�Xb��T+��u���qN.D���C
Ō6�Z):F��&~�����L+D��+�]��D"�RYpƁ1�.D�����N�8o���ǐ�G>Hr��+D��H���5Zz,Z�jN�~wE��3D������s$e��J�@��q %��9�S�'A�荛aa\2R!8l�5H�2�̵��~8��(�(T��X]:R	�6B�ȓ�h�uʉ��n�(���*$fŇ�S��p׭�N�������7�ɇȓ.�⁹7�G�!�D�
��(��`��c��İg�F�.�t��˷Mg���ȓ;*i$����԰�C5'#'���IS�Sܧ=|��J�g�.����l��ȓU���0���+k�D�4��TqBh�ȓ	F��+/�<p���4"4~5�ȓ%�ؐ�g,�;^�$H҄%M%�����;1"���Z������T$\��h�ȓ;�Ȩ��KX��X�▥״st������Cɸz�@��!E��q29&��$�@��m�O�,;%��2�TAy��ջX_,��'0�1ѕ�C���3-9ϐm��'S`�i��S������!<ޖ�B
��� ����A�|����bT�
�3"O��A�ӤI>~���V�O�%�"O*X���3M���Q�^�Y4q�"O���6.��"rؔ�Cb]i�l��u��m�'���9g	߯@ޤ��C�����0��"OYx옲v��(X������q "O��Z�AA�h% -��쎜G�V ��"O��k�?,(��C�ۜl|�z�"OHa򧤃�t숍+���zV��"O���"�$�p(��+
/EH�Y�d"O�	9�i565�8�aɳvA:�@���S�'u�D�I�܉g��3 \���LoRO�`�ec�urqɔ���:S"O���4�����I��]�p�	q"O�A:P�ل�F%��I_�k���2�'�ў�I�<&�T��J�y��l��M�ul�-{`�Og�<	����(�� ����"^X�<Qo˿w��� 5a�!g�Q�<��i��}��Bh�c�\*6AhB�	�K�x}0Ī�)����P�%XBB�I�/��7GB�X���Uh_�3 |B�I��m�2-ۈz`H��Aʎg�0��d�<�O��e�D���Ub��"Ӫ�q"OB�˶*?� �['����i�"O�r#Q蜄�1�_�9���"O�"C�L8��`�8���y"OZ5*t��
�h3��?ﲔ�C"O x��K/΄I䀀>Z:��9"O2Up ���x|r�+K'rf� �E�|R�'.b�'��O���<J��湊6�*����B�4P�	�'�:x���1wO�p��ʊ!ON��C	�'*�"3��n���[�OF�K��p	�'�pD�)>�<E�CP�(L��'ָTx���$���*M��d�r�'("`M&qb���g��nL�'le�A�ʅ0e�؇�ܞx��S��?Y����OJ�S�'��x��!�4A�^xa�!��E)��	�'ڲ���쓊5t]�S�C�EI�'Vf��Ej	#}Lh�n��?V�@B�'�̝��ؼ��a�*=�2H@�'@��i��χ#���%���5�$���'�T��ԍ�w��M�+K�3��"Ov�Q%*  �xP�7B>Vn�H��D&�S�I�=�֌����5o��h�ԩ3�!���!Op(�Mx%.�&ɋ�B�!�dHR |�G 
6$����Y?3�!�$�7f݆a���U���"H�^!򤝖o�h�2'��[����i.cA!�u�mi��JN��\��
cC!�$�O���QW�wh�pZ�@Ɲt5ўX���e��<	t˒�D�h��'K_>�|B�I�,#hH�7�Ù,��U"��DB�I�Rw8�#�|r�_)O:4B�	J�0�;BbJ)�P�v ���2B�I*��u��C#�)�\>(�4C�I�{V���	W�r����L#9,C�I9H���V$�K��(I��O�d|6�?щ�IS+: z��O?D��H&f�j�!�D��5k���(��eƕ"�!�E�H8p`A���aŠJ�H9�C�;y��׭��_ ��
�BC�%aG�#�-G�f���#��-�fC�ɦ"�H<���[�� TC�I6o�p�UG�
�D��w�I�T�?��� ��W%B:A h�3��ݱyL�YAD"O�1�č,�V������3D��"OЅ`��ЕM�F-��@M=!����"Opl�C��ڲw>�!���7D�k�B9g���+��b��7D����gGK�[��l��P��7D�L�Df�(�J�٥�H�@E�x�v3D�tKפ��:�SB�k�t�"	6D�<db��A��݉Uk����(��g!D��b�K���|aJ�q�r���"D��Yj��GL�%A��B�!D����=jv��a'���l�`�S�2D����]<}�⸂�dƤFJ�g�-D��cPGC =� �0���.cd \��9D���C��9�����Y9���c �8D�`���+W���&B_���ɲi5D���P���ZyI�
ԇ{��1!�@>�Ȉ�n����VWz<܂s����u�0"Ox�?Cv-��Q�L��Q���y)˘��	0�
�	����gN�#�y�HV-;�r庥��Ut�e[��O�y"j��N��W���i�y�W!-�yB��`��Ly@FU!S�q�'��y�	�\"��EL>~�ά�6b�9��'���O
��D#Ҙb��8'���BP����yRjjcuyq��&fld�qЊ��yBh�>T�<����]f�!�d����y"���v8�9ӎA�Z)���g΢�y�.�UH9cS6{8�LK�F7�yb�Sd( ���y����Dm��yr[��pe���m~�Dh�&����?)���dL܄M��J�h߼[��K���?Y�'����U�)`�ɹ���.��-*�'0B�@�fAg�C��
���'nf ��V���1AdÇ �t��'ֲ�s�4g��	�3�C%O��Q��'2D	0DŖW 40A#����Y��'ͨ���Y	M!ތ��ˏS���+H>����?açQg�	��A���fȨ���E�L���I~"d�)9�\)c�%ʁ_J:m�C�D��y���'L�:���=Y�`i��$���yҧҸk �� s
��`d�!H&C���y�C��v�R�H�`���`���y��. !,���I��/�8qеJ���yboϣh�zA+�-�D4�u� ��d ��|b�y��L*�1���\�}1�yb�;)^M��`^]l(�x�����yB�I�X�S���bM��+=�y��� ��X7�f��TQ&���y���a�$P%g۫g��x2v#P��y��r�i#$Ğp�[FJqI�ȓɔT2��C�y�f��O�D����}�$d��)Ȧn�5
 �>�
��9�ecK�%oYp���J�8aC,|�ȓv��bs � I��]�d��"4��ȓqe�%����8wT8Q!�"B=FeP�ȓ���"��Y2R	!��t�]�ȓ@
��F�RKF���%R�m�h�ȓwD��{�^'8�� [V%��6r-��Y �y�ʴ��#rE {f��ȓ���e���A�4��Տ��̄�I�֩ڵ 5��9Bd�\�0��	�ȓNӂك��:V?�hZ�ϕ�DT��[�|��#Q*�i�MǘQ�*���S�? ��"�'D�@���BL�X�a"O�����6zW�Ȫ��޼D�N���"O6���ε%�u��kQ��N�!�"O�Qi ƕ5@�� �EQ$+��ٙ�"O���ÍH&qA(�U'�B�`pq�"O&9�$��w6c��F+��'"Old�%e "�9Q�qS"Op���g����$� �5�"O a��H���3�T�P$bq"OB���M�R��M
GZ�|�b `�"O��	�����,As�D�I5�"O���N+��#T�_�e��<��"Ov�{F�2"l6�;B)C�k�*m�T"O޴Ƞ�J�>ȕ@B*��D��#s"O��CP]:� 	��(�I�HI�"ON`!�ߊS��*���=�H��R"O��ŏ�;z��I$@��XӺ�
"O������/ +���0�$����"O�%���T7y�����fRfn~4��"O>�ʠEO��
�BƳC! a"O�8#'QbN9�jܡ!Ŵ��"O&�t����V��ɳ�"O:3�b=9��(��.B(vy�Ԫ��	ϟt�'�1��tF�q���c��BQjPHCt"Oĸ�'�/l��EDH���"O�QsS�
 ��eÃY�D���"O�P��2z��usT��B�j�"O��� ��E7@���3� 5��"O\���
$Gc�xb�Ԧ�
�P"OT�q��$��0� ]�
��ȵ�'���+�Տe2����	��1d�%9��$�O���B���IP�$S���$4W B�I�tW�1�'6�j�'F�
B�"B9'�
���7�[�O7�C�I�R��ĉg�/T~�%A�AFxXC�I�9��dZUf�'��1�����>��C�ɹ*����t�\�=10����Q�zB�	WR��ضM�N%"�i���#H�B��Dl�l������YWϠe[~�K3�'D�pQ���p9���L=}NL	f%:<O�"<q ����'�=g��MR�� [�<�B&��{��q!b�_���r�j�U�<��nY
��0CAM���@���y��V	,������4��T�"3�?����h����%��B�R/_�b�j&$�?4�}����a,��#�\��d�N"���C/D�$j�*�?�} �o
.�m8��2D�k�`�^�̨+YD��)Ƅ#D�h���֜ua4�Z��pI��;D��F�0x.^m����YY�U�d�8D���/_mj8&�	%��q��<YH>Q���O$��D�b (�'�An|����'R�I :���I"O�aG�m2EA�2EC�ɺ@x��������v� 2�?a����#;�H}Qg&$�i����I�!�䞨w��*'�<y�,L�Ҋ�q!�D�t��$�fc�9��ثA@�y4!��0��n�u��<���Μf�"�'/�'+�>���l�����W2r�\��@O�t�0B��Eh��5��I�)���:�*B�	�K��b� � 9�"${r.
�btz��8�I��G{2@ѓ.D��G�h�(�ZW�B:!�D�VG�,�G��$���� �-!�d��Q�����,xpnH3Chȅ�!�� �e��L�FҤ	�+�� Ja"O`�@��C�$���r���}�$i0#"O�qya��MR24k삠�(���'z��'N�ɱp�b����H߇T�#��',axb-��W�}�D�]�V�x���Z��y�����e;���P,d��g�ǭ�y���z^d��� ٿOZ����	D��y�lQ�!��b�K��5�j�a4��!�y2��[9�3�W��PTsc�+�y�Ѿ�s'�Q
�Ε�!����2�O���bQ�t�f�0��<(��Sc"O�C�i�!�h `Uм`�>�4"O��X�f�=�
$�0���	r�!HE"O���J�v�4rd�kLԺ%"O2�9��?�"͓"��Se�T�"Oxe'ǋ^�n���S/XyA�"OJi��&��T�f�t
��K"l@�X�D��	�8��B����x���qs�A�4�C�h|��� g���x�Ã�$C䉼qI�P����喍��CƶG|�B���YcGIP
�fq�5A��B�	"h���Em_�3�(�Z/�)�C�Y-���f��:8 c��-�vC�	2�(݂f*X5/�Ӆ��n�2B�ɎZ�h!c�:Mb�$+b�2"B�I ���+��ݾ��ISu�d�B�I�{IZ$1�&o]��{����C�%9���V�F��e�`"� \�zC�|�X Ggj�N5��۫+�PC�ɒP��C&��5�2M��Y��B�I���Y*�Ʌ�欣�?A�<B䉆c[x�e-���s6�¤	<B��6����G����C�E��tJC�	�#Gi'jbx�KEᐐ!e.C��	)V�XFX�Q��i�Ȑ�`,C��^�h@q�I!;�¬#W!ٴ}�C�I�>Nl	�`�4����LH��yb��#�.=A�$%{r�,��Cގ�y2���v��*m�>���ز�yr��WZ�A�b��3��(�0O�9�y�ŏ1-8j܊QȀ�Ɛ�5�א�yr%�T���K�h�՘d�Ϝ�y"�G�H� ���`+2�z�M�'�y�#��P[���F������"D����,PK4��q�qU�y��	�0(��h�-�&lxQ�N;�yRd�	#�9!�F.1RDp��5�y�II����j�n�'�e�p�˙�y�\�i�q�Ug֯z��X`�A��y�
�3{�iq�H�<	v�QcN���y��O��z)#>Tx]�rL�6�yB�Ha��݁5
�N����
��ybl~�8|�䌝�?C��	ՀE1�y�T�X\FՋc�PE�4�d����y���\G�@yu�?DL]����y�Jt��� ��.1�������ybnZ ]C�l;�Ӫ�΅:�.9�y��ΠQ��yw)�}�&���yraܙ%����c5���F��0�y"�ʌv�B�Kq����^i��ۍ�y�LQ����+Z�W�j=#�n+�y�B'OP"���m� WP�p5H-�y�B�q���E�pTX0��y"΋:Yj�D�Pl�(<����*��y
� �lz���/䀢�ŉ�T*"O�12�C&o�`��`c� w��YBT"O�4R�T�Z��uxw�ތth��&"O�x��]=Ib����֐����e�<����	5�a�e���Y(����y�<9��)+6�xa0%��k
J���c�l�<�F"(h��5� ���x5v���$i�<�@d��H��ܑF'�"�#։�M�<�[+0�4PBခƀpsEƖH�<�P`Ls�����ʢ�l�{ �D�<A��G)�%�AB��F��"�A�<Ѡ-C8U@y�q�ɾO�r !hM{�<���1��pa&Ȁ�1Й굋m�<�v�O*GV�;q��0r�
 ��M�<��?t0-����K��m�+W�<q��.- d��hȩ9��@��B�<!�A�>3���KA��jn��zpk��<�`�a5���W�ݧ"~�ҦD�|�<�Z$~:.���s&YBծ|�<Q��4�xe-N�
�|͢eLC�<�a@2�u�$ꍀg�,TzwB}�<��oB�:��Qi%-k�pb�Ey�<��U5!�d���S�{��i�C|�<��B� b9��Ν�At��F�^�<�4�@2V\��"Ӝa!Lh� g�E�<Ih2����G=�!6��D�<�5�R�A8��{���<N���PP��B�<��EB�A�7aҴY�^U�<�%�(%@��Hs.A63�>�H5�CP�<��>8'�� ��&t{ �H�L�<��a�NkH��h�"u�>�s��OE�<�Q��'vb���l�"	2ܓ��e�<)�� �?q���(A�րYa�[�<�`l��(ؾ5\4\Bth�Y�<1��K���RB�T�>�+���A�<�E��v��Qa.S5h�@H���]@�<I���1岬k�n5!
�|b4��~�<A5k�>nE�e��R1f��(:�~�<��-m�����F��-l�c�%u�<d@���r�C��TB�r��l�<q	�-oR:�A�酿c����@�e�<q�)�xFJ4R�� ��������`�<9Ԉ���	`P��F&��ֈ�E�<!#��$Q＄�c)��<� �h	@�<�rD��&#����;Ș���a�<q�A�L60PS⍞8��1��M�T�<�.�	�9 B/�;�ݫ�)�i�<��B�1�� � ��%"�+d�J�<�'c����2 �P,E��Y� ��]�<�V��(�e9 �ϼY��r�<���݃U攠#�KK�\��b���w�<qv��3^�\a�T��>�v� c��<)2O[�{�
abFďtr2��`Lt�<I��T/D�|��F�D�
�@�&�Y�<���"���H!k��U"�遅W�<�T�L ���ll��EלYlA�ȓ%ff�0�ߡ#��uq&�ʢh{�����(it��y�ެ:�ܵQ���ȓho慡"�"��� ��/?�����N�d�X���"����!�\���I����ւK��mK"�#VX�ȓPR����.��{��k��٠R�5�ȓ%���J��$%R��
�L�`�ȓW^(p�ѿel�ч���xP��S�? �@�iWrE���Ҝ1���`"O���O�4�xqC��L�HX"OV�����\x̹#Q�ܧ3�E��"O���f�#Z,�Р%�'�>�0q"OFB"/�5^�d�h�F�!z��E�""O����A8Jt�X��%�)|���x�"Oz����vZ,jQ�������"O����$J�2< ���V��"O�C"j�@�vQ���J0\a`"Oz�q��5}��!q��BA4Dc"O�0�(����i�ЍN�2F�s�"O�X�El���5fJ�'<�0"O
�8��H�^r�y�B�s)��'"O.�P�惙_���z�а��W"O���L(>p �B�%�|Ը�"O҄��/˘u2El1�䤀�"O �:�D+jԬ���d�� @�"O6I	�Ș]t\��$�łe�����"O��؄�Ѐb⦠K�CF;����"Oz�3D�D�)������"�x��t"O|��g���j�.�CU!T�`�"O�L)aAԸq��)�B_��(h"Oh`s��	*ot�09�O���Q��"OȀ8����1�fDa[�E�l�n"D�0��矄&��L:2A�`n�ͨ��8D�x��
Q�)��e��E䪕�D�5D�	Q�� �p�;p��	���x5O D�B�a;(�(�c�I$}JX�u�#D���E�(|D�c���C;2l�!D��ʗ��;9=d�@lA-P8P��>D� S�H۴_:�:�+��Uv���B-;D�Ȑ�N��L,�&��><��dm-T�����:$h�r�,O#2�dp4"OR�X�UF+ @���[�*B�Q؀"Oʴ����%gj��,A>���*O*aࢃ�ot�<[CG1n�%i
�'NJ��EOw�颓��\j�d
�'qb�{�������G��
�'�N�H�ʞ���X�BI:���Q�'�����i[�9��膋ƫV�Ex�'����!���s���2��#I h9	�'�:`HsbHɀ(	 nԕ?:����'*"�b���:s�h��º;vQJ�'`��X�,��2q�I�%ۈ��'�}�F+��C@\�k�@Z5#<�x�'�����mA��-�g�K�J�<x�'�2����������g˙L�Z�'��A �=\+D�Pf&�&	�Zx@�'������Gt\9v�	�|����'n1K eh~ĸ%1r	:�"�'�n�h� ϛn��H���k�4��''���tC_ 6���p� ܾgI�DS�'��as�C=:زlP�@	L\��
�'}椋Q-]��v@!�e��L�}�'(d@�.��t�ҡ!�d��K��}�'�BU��O�QmX����A�1	(ِ�'���Y���]�$��]��'�V�Ӯ�v�h� ��^4��e\���<����*H��� ���L���i�&G��}���������@��A��I+^ك�7D�HCD�\9kT�T&иul"I�i3}R�)��9v�LIq� �qWH��f��c�؄�I\�����q�ӥE�F�����a?)��P1��1�D
iC�W]�<� ��E�?W��R'��\0�!t�'>ў4�n3Wтl��N$5 ���!D�<��E�=z�t���b��I��"D��j�&B��ܨA�%%fN�x�G>�OP˓���1��_i���!��Q."(�'>R�'�x�(���*R����P���;���y�>�`�3$ -�D��?�y"퉲Dr��ᗉ	�(y�@��.���OD#~s��	#*�ؑ��,"�����D�<��eV#F�Q4g��f�+ph�}�<af�U fB�<۵�C"]�n�EX� �O>��Q�
o�Q�whۗ��݈[���� S�2e�����HP��I2���5���<�;�(�2u�$�I�e�`��&�-q85���:D�$"a��[\�E�a	�6@�8�9"�"D���@[�5��1��Y�\�ڡ��H D���gNY^����?�~T���3D�ԨQƁ#`����ޱ@�L|���0D���*W)H��)��
ۗ# ` �7
,D���ƙ.
�zE ��\��'+)D�\s�n�1g���t�V�
��*�"'D�����C� �l3C*�2 �:ykP�$��hO�S]�:�k1e�\-�8�ƊP�kb������`��J��\v�6� A-C|C"�n�ş(�?E��4q����7/�)a�����?�LFz��~�b�;mQ�Di�D�<H�
ف6�[?!P�O:��dOC��n�Ix��[E(5P��r��1O\��?���JA��P�%br��⤗pH<I$LV2?,(	�mB>� !J>.��	h��,��+����x��.&�S�A6LO�⟬z&�D�K���pL�Ȝ�S�N�>)�>ъ��wn�q� ���2[Q~���[j��&%^Ni�!�@���s��p�>�ۓ�����+��s��9K���,[�B�I'R�6�!4���{�\Q ���6Y�C�	?/����bED���$��eɘ�DUz���I$�I�n��E���4(�$��"^3�bB�I,$��I��ȞZ�K'��ŰS���4�L	Qr,@.��c�Ƚ8;f8��N?I���ϙU���� E�a��-�&�)���<)�d��NْC�L�I�.L� �d�''@8Fy�Q���F4�D$�7"�6����bO>��xB�. ]��ᇌ�S%��VA�$D��o�P��h��q����T
�+4D
=b� ��'�qO�"�O>�"�'��fȅ�t"O�Pc�	ͬ|׌ԁd�)~d���&�>ъ��)�	<����s#�'.��{���fF!�D�A5��5�Ȁuwe�592���)���`vn�*T`JD�L�~�p0/9D��`��_H��;��ؙ|�@���!x� �?1�ט'Z�S4K�:���@&�Z��ML2#���m�H&��ib�́53Xg��h#��!�v�8	1H�S�O����SnS%,��rO0uf.��'k<C�Ϲ��P� U,q�ZTA�'����Ȅ�V�Jm#�B�<��1�'�s��6�P)��A�
#|uy�'�����	 0uL
q�-o�{�����&eT-Oc4x�f	r ��#��y2荿~_nT�#%[oD���&����<�OR�Ђ�*I�����m�3.8D�(��	D���	K�1[��'�+�6ذvCN\$!�����+�C���� �0bA�1�k��ħ��I�"xRa`ff�;_�썀3'��Ɠ5*r�j� fPfru��Vٖ��	�<�5�)�~�H?��S�? h�ℏǣ\ŠMC7�C���S�'��̧>iCH�h��$�T�R� ћ�l�[y�'�Jy���'��5*膤XJ`�CU@�)b|����D#��?��ɷ1�rϒ`�$��S@�; )�U��!8���s�Ж*a\X���y��C� I�#N�E��ܐRLL���M�g�Z5���?NIt�Y�!Ewar�O�q�g���̦��Q��j���'ԛ���{���U`ި Y�yA�g�,sK�B�I"1��tS�&�)a�z8 ����G���<E��B2	 @L��ѱ`EN�T��y2�>x��sLŖ_��I`�lÌ��'�$܅�I<#�n}�fi�'	L%��e�5|ߐC�-)�H|ˇ���`�`���^%A�NC��uV�}'��9iE�� �Z�RC䉃B�ja��۝'��*v#�
yvC��3k�^tz�T+D��x2�LK���⟬E{J?����o�B�+k��^�(���:D�� d�!"�jLAS�R�J�X�{Q#7D�������J*`t ���t�v�	�A6D���U���x�TykR*�oF�tm(D�04E~�U����9XM�%D��@�e��Fpd3�eݣ{��l���"D�T��E#p��� �'r����,�$��1z�%�$��}0�Y�A�=H���p?!��܄mD��[�F%Rݓ�
y�<AA ��`� ��2k_R`��I�<9I��h�݃��	�@��(*���o�<�g 'i��xjgk�
{\z��Jk�<����(>��SSÔ��ZÔ@�<	Ď̂qp�أLN��X��c����?����:%T�a;��E�}}��3�O�X�<a�B�'6�L��gG<l����`̓ט'�0�|�JH�f�PdIp懸F��]9�/IY<��85�a�Q�p܀3cPD���'�ў"|*��-,AD��KF�΍0E��v��D{��� o������:�KebK���'���$�&
I\x��BMD�9�&O�GR!�4���2�*G*>�	i�M��!o!��ڶI7l��%�+g�RD��ƛ5���gy��'� �ca!���\��BL�4�
�'��d�`�ͪ�t|Yʈ)t�p�b��$<�S��b���&��Htb8 �jɛ�y"��]�@����%,�q���mZ�Q�Q�"~n�$2. I��ژ!�4���H�P��B�I*�v�jA�Z�rrE/��.�B�!�T��N��&��YS��h���	v؟�k�%�;9B�]��-��kM��#5D���1w��үO�=9�'�J�<��.�
"�9��K^j	.��#ꓢ蟂�3�@�$v����$9�(;�"O�l؅���.%.(z�OD�+�aЇ"ORT��oÞS;�uZP��fQ�"O� �[�v�`��P�Åh�au"Ox�Z�)ǈ{��K�%*�@}J"O���P��	4�H*����^`A�"O��GLΟAJa�s	; �h�"O�ț'30PTH%ŏy�nppE"O �qf �z,Ȅ��m_�N� �;�"O`\#�#X\4(P�ވ(b���"OR���������wϞ-T��"O�P�T�*8��i���8�<���"O�1Ɂ�7k�vd�qDH#h6bUc�"O�T�q,V���-�Y�
� �"O� �Q����4X�HJt��"3r0���"O0�pqBD�D2E�sѱII\�
�"O�L GlL�Y��M����RJ7"O��`�śH��Г�+�:^$��"O����Z�0�٠�, �2�"O��s���d� 0���(�n��"OmS�Z�&z:Uб��\~�\R�"OL���ώ�k�6	�ݳjl8��"O`�x5Ș'd��"dH�N��s�"O� K�G��d�"�� �k�V\@�"Oh��AN^��y8)^-1�<i��"O�A�a
�$��
"G��\�\H�"O�Y�W���]L	���U��P�"O�Q�EW|�P���!8,Y±"Ol:s��2_��d��I�%}���"O�Hb%*�>����e,z�x��"O�օ�Aײ�� ["l��p�"O�<���7Lr�m�`�,	�"�`�"O�	A	������Ώ�ʆ��`"Ot����DZf��\1���"O���uk�m�F���<d�p��4"O�E{�%F�Y�e��.C�f�(Ɂ"O H�#R�_u�d���ƉC�V`3�"O
���A'+���Y3$^H0��"O���gJ. ����~��Y�"O�L�"e�X��Q��F�-5bΔH�"Ozm��)VT�bd�3�W�Z	�p�"O ��Aǋ��4X�m��E�  *!"O�ya�/5$�p��6%��i����"O�=�`H�6ލ��ж�`�"O�I!`��5yC0$���Z�2���"O��b�S�)F=��I����9�"Ozi����S�ڕ*0j��A��Ը7"O� R¯ײU0��ɧI�E��tV"O��	001@�0���"2�X�"O>���Y�+�2� ��=g�T�"O�]���T6~l䱁�ѕ*{~(��"O� DȢ3fA Ӎ��`��!�"O4���D<Hf�a̙{�rܙ�"O8I�!͈�c�f���i��t�$)I�"O���c��_�����G�2p��"O&�s�B$_��=A��:X�ƕ0�"O�l�1"A�RXÀKL�[��|qu"O�4��I 4E2z��'I�����"Ot9Xc�T�s�,�y��6$�*���"O����/I�z�Icg��$���0""O���Ǚ�3 ���Gm!3*5D��;��l#��3W��v2��t�Nm�<�"M�A�"�QQ"PM����c�w�<��J"f��e�Ň�"4��x2�	Y�<�`C�8�J��U�E8�| "�c�V�<I��R�qf��IG?Pxyn_P�<�ևp�Lڦ�;?�B@[��N�<Yw.&bǘ��G��81'�L� j�R�<1�eD�GcX��%I0M)x�����A�<1((�~�S蛲�Z���&C�<9�$DOǠ*5aγ+�~a�''{�<鐏ߗa5nА��)�H��g��J�<Y�H�|,Lp$`�{�2�Q��\n�<u̖�3yl��т��T�1�G�<!��DNl�i�R��\|�<Ac�2|C�E%�	�ڨIIwL�}�<a�i �E��r�]�	i�U��";T�����Ԟ�&�q0k%c�ˤ�u��I1,B�qO?� t�9�aH:�d('��
޶��P"O�q�H�;l֌@��lJ�Q��X �Q�\#B%3+BY��Ʉg<p9@�գh�Q���P��N��$!@ȁ��,��!A��"7�s�Ԋ0���u
�'�mq�)_�y���k�͇8<�J�+���_�u�����Խ��OvĔ�K	"����s��3�����'O������9���F�� "U,���4:��B����lӧ�����UDX�z�	u�D����p<qQj]'��'#Mi$iJ�7�f�h5��\=X�OީI�ㄨ/����
ϓg�Dj�˂D�i�ᇏ�z�'�����CO�S��c��r��h�������n���x�"�=n��7H@h<��	L�q�����Y.�( !�B�W̓�<,q�b��ؘx�k�*��IN���۴H!�Qr�dH�hݤd����D<���x����ϨEMv�"w���Y�����iO�:$�:t��/��I^��M�p+ҭ���rƯ'�xy:ed������}�qO���/VU\�!���C.���c_�����4 R��'"e:�ΈO���AM��~ (�Ofe)PfÛ鸧�	ڎ|9[p�S�RO��`�*�2Mӄ�9��ʄBoRT �'&j��� O�������'j��0D�P㡎 N����5
Qt*P��p�g}�O�fI@�ƅQ-r�8cC�Lp�˓	�R��!fB�D+"�\"��$�۸D�� �R��RJ�ϓN���kĨ-�)�'$��YS �
Z�4l�J�qM���Oa�b�U��D{��;�c����#�����p�O$�3R��,�0=����T�upR�Դ!�����O&g�yiP�x�B$�;�q��N�L3������#_Z���-a����$�Ԋ�Px�@\��` �H� �X���n��<��i� �(!Ҝ|��@��8�=�S$FFykD�$���KEI�7����-+��7���2��_�ZT�Q!��5�L�#�N�.��)�θ�!�����S�O�Z�"rQ�`p�8Q���-In"�
I��YҬ
]��t�eB�k�OZ�]�W�C�p��܂�m˝Bd{L���u%9��8Ǔ2B��H5��E�
��SM�K=�lx�dڋV���5GT<٨2��l(�g}BaLn.�J�	��80�$ՁH^���됯%^���ɯ$	N1���s�0��4g��X�G`���t�䓻�ē�Mki֑K�6��D��z}���5{�B�+_2\��a����L2�p��	�e�h�Do�(��DO"S�@��%l�|����!e��O�1Mo�\¦��(5!v�	A"Ц�~RF�7`9\�Y���	���c�4q �W���S�ȁ�g~�O��C��	e|�	f�}YK�;&����&!a�:yh��	+D�a�D�I:I�e�IOw�����I�y��h�Hp2�S��ɪ��};�옮�P 2�)L?s�c�\�{q(�'23��Qt*�7{ڀc�����N�P!��C�+�8L�h]����(�)�F�"a�:��t,Vu���1Ï#y[L�S��M�N��,��쎳9��%Թ&Uƈ���H�<���q�!|QX�3�N�����|0��38�@fF�)RK��H��'	�``r�Z1 �(1���`͚���B�,�%S��S�v�Tc�L�/>(��%�� x���eʐȂC���TmD���x�A� �J(u��'���O�BEƎ�X �$��r�E3!�X���0�%�M
xs��ڑE��m��o�>!p@ۂNў�tl���$�n�,�����$�.Y�h��<���ޑ~�|I2�"PH�2��Kƥ(���O�q�!ݝ@N���/_ *�>���Oil��1� ;�a~���!��!��;����U��;_s��A��0�F�5�>=8�[?%��Ϟ8����O.�X��"MT�A�hD�[N�p�C�'�*�hr旇A�:��raĹl��X�pe(Tk.H��v��2�E�=�P�5���+]�E��k�Q�2�[�|yaxboZ�kZ<@Ҧ�v ޟ]�6�Q>?�B����@>Z�YV+Z��yRJޡRm&i$ğ;��e0p��1��$Ȉ>tZ=�P@�
f�R�k$
Md�O2\4���]s���9����r�� �'(�Q�%���]�������a��lyע�']� �㵨���1�Jȗ��g�O�<�aᏠ����'ʨ2����I g�:��Ab�V� �Щe0mXQ	̖�p�ɕU=�� �SF؞hR�M�Z."�Q��׿kNɻG�;�ش����F�t�f�~��yBYw6��t��9bJ�`����7���+�'�h�؀��B!8e �.�*�Y��'ٸm
DB��b`��Z�f���;ҧ'*Q(���Q�H��e�e��N���bÂH�� �?-\���O� )3$�رd�(3͠s�j���D��f)QԊܓL���'�N�:��}2�?8�Z�!V  2sh+2oG���kp��+B�<y��4!�,`��TH����7���� �x�}0AK�}ў�)AB�15H�� ��u�\��˃�'�� 4ږ#�"�"��'׽�<+QL�cH<9��� _>}B�x�2}�l���E�%.�����d�v��E�U(U#�;��Q�R��c���=�!M<+L���'�b�[քD؞$����AH�iZ�iC�E�� ".yX�h�����_�V*��'Dh��.[~�P� � �
H�������w|�����"�Rap�"�ZuH#J/D�܊F N4.϶I�Ն��i���Õċ�n�dۢ�[Xf���/��^O��҆��6��	>����S>Y�x ��� M՞�y��I��hO�%�ďV��R�$�7#l��BbX�L�z�h��.]HQ�&M0YI"�#҃Zd�<ɂ%D�k�0�'ʰ#}���rb昪� �r&>��CG&]��D){\%a��T2`@�5 �-qh�`�q%1��$�'탕{���m=Q���������@ݽn��j�'˴@�$��O�y�
�7 ��2���K��AȔa_71��T���΃��Ƀ?meZU��� Y�u���bMV�����-\U�T0� NIa~B��&�	+R�ɼ4�6�1�&��Y�����C������A"lY��05�pɽ6�4�I�h�OE0u�4gX-~����8v����$�Mw����MQ0o7���Pg�~�s�Y&K�ɠA�Y+co"�S�+�?e�� $Ҕ��O?���|Ν�����,�R��1��-<��Č/��q9�"�Xd�Q�#%��� C�!�, �%ʀ�A�v%h����}9��чnp��$�E�i�e�fm���R��-*�epA��4cCg���fA�L|Γ)n٪©�EBy��G��Yeq�3b�a*�m"�O@q��g-d�`�r�|r�`���+?F���R�Ȇ�M����n�?9�lN�3�^�{�	_\������_�r":}�
�֙��G�OF|�v`�*u�d���ʲ��4���{�(j `�8�8�1���p>��D�*޽�$iT�%��񃦚�'�@=	�GC�t�2M
��I"b��?�� ���Hs��!�n'N��4�b"Oj�YD�� �`2�
�R �!�'vD�H���$7��P.� Hz�yd�����Â�V'Ҝ��[?��\�ȓ$�p�F)�2W�tm���ָ�v�4j��)[�ֵ�~�S!̗a���I0h@\7���y�@��ƚ64�8�F��q�S�'j��D�䌛�Tͮ@+���h���"bJ����Q��J5q�T����,�0>��3Ŏ��F���f��L ,e�`#�kV�p�Np��ƙ�?a�p�W�.�� �O�t}[�dY�@�A��5=t��Rߓ(Dq�3��>����� :���0H�I��f����j�ቢv����*�,f20���j�O��X!`��.���c�@G�օ���;8�%���ɀx*��@a�Լ5���g�M	#� t��b��N�� ~�ؐ �^>�Gx%U������o��Xs GWF	j��.�Ic�O�a@T�U�n �3�ϳ?�@9SGH�R�\X�@8B��(ӓH�s8�P����3A"yҢ�V�Dn��d��OL�	c��&��8�H�C��On�XT��9���&8���t�M��|CH3]!a|��C��l���jJ:f�{5��,&�؉��E� �G�`�!g�����#-�^H��yB��$�>;V�ٟ?����S@0X��MC�b$�0�>�wt�n��`	�Q�7��S}�y��#��LhuO���%��7U
�0Ђ��oe,��׭���ft[�-� (@��Ų'������k<���I/%��IF���.���o�$$��g�=@�]�Df�6&C�	�s����Ce��XX�MJF�E�0|�,���Q8�ЬKv�^�O���5�ѕ�jQ�Ю�0V:l0
�'� u�W�߈r���GL���|�a����� qG�<��'�gy2��[x�{����ju!jq��y��J�b��y0M3:��P�\�h���	��O�\#�#lO��A!�ԱX�z��Ƭ�<���'$�)��gξ!����i-ҽ:P���
�L��b�.*�����'���P�b�{���җ��,/�ő�{B(֖��T�GDċ��>]IGh�/Ip:��%Dq|��w�-D���$A� D�1r�K�8�pH���N�Q@ Z��l���DɩIG�M�r�H�i@:03�P��!������j]:�Q:ǧ�6b��
)!�����'3�X���޳f���뀈Þc���b�'�P�aG%G%3�Se�!	]М��'��A�A�j�5�Tm�rؖI#�'w� ��s`�Sd��#cj�'l�@�0�����A��0E#
�'�(FY%G��=+2�
�|���Q
�'�`�I���}M`�J�M�z�1)&D�� b`��ȉ(p�V����ߎ�h42�"O �����n�qo�H��y`@"O�DB�fǧ�T�)�.WA�Xis"O ���U��Jݓ��
~DI�"O^��:��лC�08���"ONb���10�r��5n���ab"O��y��!g�nd����z�
q"O<�)��X��L�W�G"r����"OT��g>#1&�{W�Fd�1�"O�I��nE�i�������=�A`�"O���@�W����3\���Qs"O��Bc�1n��0��
x�2�"Op�d�Y'/�p��N�*>�����"Od+��c#ߡCϨ�q�j]!�](4�`��pF��2� =���W]!��'Q�ȣkC-{��H�"D�!��M�,
|| ��O>�e���7�!�d��-�d�$HԛB!b�צX��!���^CJ��u+U4
�-�t�.Q�!�P7JD������a�ٌ^�!�d�r�I1�ح&���r�� 0)�!�$S�6ư��P�
(`��ip!�ޡ!�ټE~�!���	~ö��EG�`]!�䙺HwB�;%�M��ơ҈&k'!�dтV�b<h'$6y���� k!��ޯ��Yb��%s�M�K\�	�!��
.C�B�k�(��01B2�D9!��X�&-��!�������,�=?.!�D�>>��xᤈ$~����+P�t
!��>�k��X�S$ԂT̗�!�$	�"��\y`��s0J-���8$!���A�pH+1·$)�d	Q�X �!�M�0,���EnA�5a��MV�!�$��F$�I@Jj��CVfLz�!�Ā7�^E8F�|i�1��Le!�$R�#t��C�"����ac���q�!��JqZ����:�%�M#�!�DN��J��s��+s�f�s�,$~p!�䃂8���0r�q��5iJ�`f!��}���s3k9D0��8ǊT�!���F����vK)>�rt��&�!�D��<��<a� O��0	�LBT�!��2I�yg�<5��yh d�.|�!�E�JO�Uh��� i�V�[�!�D�n�"pCp�6qdV��q�b�!�
8� ��.�C���'(d�!�DR>Mcp��dk@�[:2$��g*�!򤅘Q�dMHC�z��0�+Q=:{��������$͙�Fr�Y��	���A0-2���8u�1H�V�&�P��u�!S֭ـ8M���ʀ`�@���QP����v$�􂇸{�����\��D�R6�A��,�(��ȓ>�@R8 |%�T��Q�$q��cg�M�4��� ;�)� CR���Ɇ�锡`�H�"�4W�[|X��"J�Z`A�0+%�R�i[+����ȓYi� �	@��ԎL�<�,��ȓ^Ԑ횇�͠�5��@G7Ype���ԝ�VjR��qk�!E�"nЅ�U����,R:x�2�ô�Ɔ"Q�M��4��-�U!�$.EV��O(����pI�F�Ͼ�(A�(I-���ȓ��Pa&)�$Y�!䄊*e�FH��S�? �E�*���i��էP���{�"O�r�b^�I���s���=T�4�;�"O���CS�����e��}�n�q�"O@�7؆���j�P�jhAz4O�e�1�L-Ƹ�������A��zy���V>P::!"Od;�V�+�6%�&-S*A����^������5N�T ��ɓ85B����� �f���E
���2 0@rƨk�zM*4�1L-��H�$���'��9�"���=��m� 7H�0��D��h�EA���O�4�Z�n7b���#"ƓyֈD��'( ��MM�8�X��,]Pn�xشbж�I�ǖ�?g�ӧ����dۆV�����2��YQ���y"$��Y�,�Z��A5a��s����d�#U�5[���
��<1VnG9�����A,�
�r�vX�xE�U<j���Ṅ29����E^jtEԇ�!Z�񄔚b�<��.o��c�*L�,���l!5
L2kv���	3t��Q����A���rS�L�V�!�$�)��xP/S5D��R�O�wɛF�W �U����@��s� ��P$�?�>��HɀG�,8D"O⍚7�T��͊�g^�V�t��W���l�&;�����'�f��᫁8cS@(��L��!7�H�	�Adp���V�u8�1Q��]�A�>-H� %:L`PQ3�>$���a!�$������ɝ,+�,����f�Yb�x�ɏl�q"�S�)��:��ɘ��A�tT,__^��DE�3�ɫPi�(����^���[����R Iy7�d�+����{�����(�蔊��Ȉu�~ŠQ�"M$����1C �G�B8���I<jZ���$E�X��R Q�!�$�dr<��@R�B��Ö́"⦩;!�GsyB�?1���}&�,�$h�!1mL4�T*�vz��V"9�`:D� �R�3��X4��� ���ZȄ�h��9V\�M��ɠ�H��� �
	8��A�Mƒ��$T�\�@@J�`�`2�
_J�
3$�	G�i�̈́H�q�' I��	T�S�O<�Rv�	Ad̬�PP�=�
��I��q���.w�%�u�G�O��{�C����&�
7Rj�qN<4�k����p��1j��F�()\�z@(��-�LQ�꟢d�剡*T���E��I?�.�N�[���왁BW�r4�9�#��� y��>�O�Qp@�Q�f�hA�ߏl5�[���� �D �.�W�O6m95Dxɧ�[@��I�
��t��)��q�p�c��ҷx4�r7�'�p�@�ě$m�ld�.0�-�"и�aFؘQRF��QK° ��9��(l��)U���&�	oR� s,�hⓅy������V�V3c�FZ �OT#C��X"��A�IU)�10nx��!ł��M�� �#z��H�<�4���
�5��y���A�  b2���'f� C~���q�B�6%�(O�	CR'����i�4d��<�kH~���<Ĉxp�\ g*�l5��Bm����ʂ��-H��/�O<H�b�P,C,����H%iN��K�&+��"AdB�9M�L�FĞ� �<@���.I8��	�oF��wZ�Ċv	XL�L�����wxQ�0_�����֗����W%��R_,Mx	�*cvUA��Z�z_tm)Ӈa����'�N��ҋ�(-��O�~]�W�_	2�aфG�R݆����|/Ќ$��+pP]K�fK��u��q� �@�E�C�. �d��9� �O�%��'��$>c��Xrc�6ˠ4(�A�\�9���<�F�P�
8�K�g՘#��0�-��Ij��g�I�`�u���y��`��P |���AQMV_��T�5�.J�@���j��r�h��GP]y\���O�3���4���O�D�Ҡ���p��~
��#�� %Ǻ9Y���ob���	{���Գ,�)IP�Q�dQ��F<"�B)۱Xr�X�)kqO.�N|rD���Ua0��+!�*���:O<�S%�=@����D��.n��lZ�%�,�y���8A2�OB�6��C�8R9���s�8<9/�w�0�'��yhRD޼"�Q2���E�>����1H����&s�ԉs�O4D����˜�N�t$�m�s�P���>��u���#��L��~R	O (���C�D�t&��q�g��y�)U1\&�'\�m��u�7��?ё���*}�]�&�<lO"��B��0.;&����but ��'�x9j��*W*�lZ�z�1#��;h�6��P �m|�B䉈}X6	1� )��ƯڔpBV�P�B����x"�S�Z�l35b����qb��C�)� N	q�V'.�~�QqJ�7{�.5VȔ�"ba�"�'��s��c&a��<��E(ϒ�G�\ ���$D�x��.��$�ӏ�7j"�ٶ��p��dI���q#.<O��z�EM�$+4hg������'j8���~�8��Hҵ`���L�G[��O���R�1&�&�2W�F�V�ЈO����d�#�(�"��Dc^0n���80�ذ
���� ����@c�.��
ۓn�p�v���*"���q	|�i�6O�A��eȔ�x	<}J|�@�$m��z���3��݈�Qg4�R��nB!�� �@p�`���?`����[5��*|����-a�` �e�N�~�'�f� ���GE�	?k����2ֈ���ٌnKV��:���	�Jv��)S�+Լ��1�ȜU��IA�>y���O��:�m�Ê�
��� ��AE��:Y��
��3Q"q�(p��aǬ(�|�I�J�O��r��ObQFkN1Pxh�ӓ�xA�e��K���@DHŠ�`a̓[C䌂ꋏG�Pҧ����~��E���\RV����a1�� �L `�L�0"Oj��+�l��)N�\�M�%�>yӏ��3 �t�p�ί_Nf���B#}Q?Ys�MT�W=dl(�E	8������"D� �f�/�����%A:�,B���zd�؂���J�Zҧ���ǺY��$9���P�uP�.
<�y�B� >��`��n��_>�p����~bFt���aǓf��K��=~Ozh3� ��	��t�R�;�O�����c��������Q���YE��'��EQ!m�<�3o�R�P8�m��X��I1P�/<�ri;�'�21����T�'��P�x����3)�
�J! W[>'�a~�m��H�@�+w��O��\X����H���0�"J�C��E���n\<��I�|�$��q��.45.!�"���w��=9����
�rB�+�I��H��F���to�W� ��F^D8�(3����y��
+��h8r�^2E�
��ף��?�Bʊ�&=�c�y5>Pq!K
�h�����Z7��!��p��M ��%D���vB��}�,ъ� �6d@��DF�:n+�P�G�R,K�X#�D�@a:�'�O����ݳ6m��X�;x~l�U�'|fѕ� (?�v\R!$ěh,�D����U�
�q>*�(�b�7&�S�aKH��Wȇ�R:(��J�hG{����%�QL������ӆ/��	�_&lP����b+^��h���!����^(��<sD\����6h��l*��s��D5z��AӶ͑���>-�#a���RR��n>�S"�Z�<q�g�V�X���W;]�XHkСtz�[U�U,a�v��5Hŵ�O����dMjzH���G!V" a O-�O� ��'i���8�XL "a���x���12 i�	E��p>����-hj���0�2U.�:Q�W�'ZВ�f�ϟ48s�ҮT�ӅJ�F9Ж��A7�I�gΎ�HvB�	���04
�uj�� ^5��{��A
�}E�d��<f��m�F�p�j� 7��
�y2 ?�0�����?e��!� �I��a�Sk
���>�p�d�`�W�NBt@��i�b�∇�q��l�����UaA�U��	g̎��>5ـk�a{r$R�>8$��'Ĥ}r�r��W��p=q��Y�HD�զא�M�VCD��	��s'F0��
f�<I -B��f��
f�Yx��N�2�"��2�F�Fr}����<"����J1sa���_r�!�$D=EY$�"���(�ҳ���V�+T��-G��'ft@F�,O$,��
.rb Iu�3'���#"O`���mZ�A���VlW�v��	�3�)޲U{�/�n�|��ɗG�|c�KY�,L8�XӅ[/l���dM5�\�v�$[7��U8-ƬXͦ�z�j��5wjB�	�[� ���ZNZ=�R��w�*�@9�@�@�Z E�W�O"T�si��{�������@��% �'�\�.4:��)�b��hP�5��j��^�xP�s�>a��>qB�}�H��CbO�x���E�m�<q�Ԁv�lD���7;�2�)C��x���.��}���)L�d�� �\�,�BL)���W�NC�IE7)�vk�i�*��㇨O~>C�ID��������T���i��G.(kC�)� ��JS�W)�PQK�Y�"O\yEC 2�<����@�[B"OZě�f��OT(NO�;��l(�"O�R����v�8�㵣��D�B��"O�x�@� M�B*����bD@��"O�� .�A	�!��{���!�*OlТ"�\<w��}Z���h�����'0�%�D�	G�D�04cBd! T2�'�DYp��
/F�d�+PȢ�)�'}p�;�o�6`#�|Cm�]���P�'������L�=i2�""�6�F9	�'�ɪ�"�YɄ�p,s�z��'|-X�
://�ѱ��Ĝ>cpez�'����I�5�����I��*S�4��'��1"A�,T
���1�G%]j�8�'X�)e�1����𭅇^_֝q�'hR�����<�`!��W�DM��'e����Cp�\�{�R�LU4��';t�j䫅�!�`�t�����'���9 e�K����ƛU8�'?�����شW�~p�UI!w�d;�'z8e��c��|��e��/;^t���'����e[�.H�e�SF�:ި	��'kJ��Q B�z��񭒄 ��,�'̒�4b�D�t����z��	�'K`m��Ϟ�V%��hG6"�<�'��q��� \�n���l�S����'�
��M&>��%���]�Ț
�'f#�ԧ&i8��"V�p����	�')<|+�#��b�@AL<$r"���7BB�*B��zO���F�9q[�X�ȓ,{��+��_�is��F�-m� ��bYJ���"Y7@Pj@ lG���ȓh��)	ʃo�ݓ��ttx}���̱�q�ͅE�IK�����ȓ]� �r��-~�d�w�Θ1V:���m�D�+Ui��.L���f�C�R��ȓk����eT�/ޖ�k� �4�:��ȓ!(ȂD��O�N�A�_#A�*���_���$�O�֬	�HR�(M��+:���'�0*���;eń����aN��B�7+7"���(L�?"n%�@J���ا�O��2�]7�v̛���c����'逼A�C�,-&ɧ��L���(u�)��
��r9�<)��>;����%�Pe9G'���X�((Ů���z\�S��-l�5 �R툜�O,܄ᓴxޢX#�"H#�0tzO�+\�DL���u��W�^��}rN|�K�)Hm&\�A)Y	t�j]T�A�	�t�hY	D�R��M0���M�K(�9[@��H�,;�f�.
�`�� ��@b F��6�tX���R
��W�G�R8ap��0�����p$xШ�œ6H�	 	{>�9�FM�^�����M�){��\���H#h� ���ݖ���M��<E�D�J��:U��
�$̞�)��
5�pq�좄B��OFT��Ӊ)3�HP��L6jR0�A�1j�Ƙ�"#τU��ʓ.Ū}�'G�ά�D���țg���7'ytΌZy2O�!~{ܘ S��4_?�1��@��%��y<0��#ƘO���OzdPG#&�)�SU(�i��m�r vă��Igw��o"����G'L'����T�:j�X)�^�!�d�<�PL�"A-�hKf�P��!���N�>����Z��0U'ݿ4l!�dޓu	VyfD+�4 pƟ�%h!��޺!����n C���P:R!���@���IaO�M0�����+8R!�D�653�M`�%�$~-p�`��~;!�$řu����o�� - p{�N+!�B�=C���n�|�������#"+!�� �`
)NM��M��H�%�Na�"Op9���U��}��[$`x��6"O.�3eAؗ>K�%Ju���zG�� "O��	؞����e�4n;�q"O$���Y
U��r�� ,��Yh�"O
�{��H���Q�M��V�"OH�r�/ '$��ɴi�6Y@�v"O�<锠� sPb=���o����"ON�c��$Sx�-�A"Q9���qa"O����Ċ�4��(Q O�y?���"Oz� %e�";��Ѳ�78 Q�"O�L�oa�̀i=�L#6b$\�!���0�6���H�(�y �]M�!�d��u��;$/A!F PD�<+�!�d��~�+��� 	����Dw@!�X�;Z墳��IPu��Ǚ�%!�D��Bܠ� �*�n��sl�A!�D Ft��kݐkB�A�&˂��!�d\�4\X2l�.`��3C�<s�!��+f��u��#�~�(��D�!�d^=Ƽ3f���B���#�^�/�!�dα��+���sâuq�I+�!�$��`z,����[�^��=Y!��)�!�����2+0�Ь��^�7S!�ďL͢iR����܁NI!�$�I��m,b���Ҩ�=	=!�Đ�k`P� �o�X�Ah�#M!�D�9(�����\�Xy��@X�M!��[�M "����\$4l�U�􅖒*1!�$G ��	��OȯBk��P�;$!�$ʷF\��*�K��#fqx��=!�d�Q�4c��.{Z�%afn�=$!��g�z�cq�E��|���͆�2!�D�4U�0yIUH=�H)�uc=r�!�d�0e�P���n�">�ҍ�hP;F�!��P�h�%F�G����eh\�Gq��$ʷW�茒����M�`O�6�y� N�?��$Ӈ�3D��!�ehO��yR��k<V4IRDǣ":�3u���y��B�,y+@�Ps
�P���!�g��VB�T���c�}!�d�1>�,���D�Y�� �Eˮ@!��Čt�I��	!�d���%�;!�䈐V���3IF�$|$��#Ε!�P�s�l��gY�*f9K ��7!�$�:���q�N�~��r�-�K�!�
K�MB�FR3q�N)�e,xd!��	cܸ�S`�2Z��(ru�οc!�DY.��x*c@�5!� �Y�,C0)K!��B<F%���"�ʙ�U���JE!�\�,��p��"9��4C���:y5!��ư�U��M_��D��a���Py 48"0hQ�LZ�~m`�T�yҨ�/u��I���OFx����yboD�?�F���H�&=�v�;PI��y"�E�I�l���"G:�LQ�����y2�H����Z5�?9���؅ �3�yb9
�8�)&DӬHL�a�C���y��ήW��M3� A�<��mM>�y�ўD�P�Ь45f<a1�]��y+0"���$�	�3mt9���8�y�'�n�!�9_+l耵�8�y$ڎ�xp:*
M� �ڤN��yb�PV?��kD� C�ڠ��	��y
� �q�&�8,T-qpl� R{����"O8q2�I�Z{�l��n��ɫ�"O`�hI��@�,�2艛w�"��"O��Rq��^
�t��D�Kk (`�"O�0�fd|(�)�I̢F���"On�Cщ�.���r�=fy�h�"O~H��h��b5$߄[e��i�"On�e ��I\�-��(	�,�F"O��r�%-RT�!��~D�q҄"O~�2�f_�?A����G҈Z�7"O.d�Ή'�\I�p�ϦN�A �"O�i����-��"�H��)LH��e"Ol-aw�P6_	�Yh�F *~Sr]��"O" �V�Z�p��T2 &9`�"On��삛t�����D�MuLMBq"O�`)𪅬]Q���/��L_�A "OT�X���Ze8�W�@�w�XX�"Oa!�gG�L�@9�� Y�(!�"O���*ʈr��C��L*�F��p"O�q������Ү����d"O�Y���n9jí�`Y�"O��J�C�*(��!�":ڎ��E"O`����R� ��p/ɐH�&��"O
��2��F¢�U��;�Ҕ�f"O�L*�
��g0��M�M���"O�����#c����c��b�5"O�� R	���&0����!����"O��:r�;p���1Q왉z�d�Q�"O���0�Ɠ.v��I�#��;U"O��3g�?�VA:"��.3����4"O\�UC��5-��cV�Z�ƨ�"O�S�✎U��P�مo�0��"OX)��'�86j0�"���9�d��"O���/])S���P�@��r$��"O�Hr�(�@����m�?KL�!"Ozq[6n���@Aw*��)и�!"OZV�Y�Z�� �B����"O:� ǋȡQR�Y ��X��"O��q��J�O0�@y�d���Y<�yR�v� �Td��{�Vy�5���y�F�3<��`ȎF������yB�u9���s��8�ir�g�0�y����?�M�͖4�ʩ 4G���y2"��YĒ�:�(O&)����T�ט�y�˥p��CB����~u�f`�9�y2��[��D��+ O��y��;�ybH��Ux&�S��n�x4���y�L���j�����0����(��yR'��Q�]ѣ�đ~yp1��gא�yb�Q"7��"鎤	�
Qx3����y���g��9�!"H .���Ac�y�"%>��q���1ɒpɡ�� �y2G�4;�%�dK݌(��k�:�y"@O=$<*ŋ%L�4�e,���yr�6	<��	���+0�8�#��;�yrMՈ,�u]/#��X-B9�y"%L�yv���Ch_�d٤͟�y��L7o8R`�!Cбe�z�4k���y,�N�|� ��>e�x�yC.�yr���c������g�I�C/\��yb�ǡN�rM�4'�R���5��(�y��N�����FFE��i�d���y�M@�
$	��d��Cv�E�T6�yR��(Xp��]*?h����+�y
� �˃*�&�e��(Q	Y��h "O�}�B��<{Ҫ�*�'	7�p�Z5"O"��o�1~���� HkʬC"O�]��ݝ\�"M{S�R�t]�� "Ot����j?xM�ʕ.3A|Q��"O��&j�"K��©[�K9�x��"O&EH��P?S��4H�B�&�^]�W"O,��m�5Pr"�
3AQ�\�F`!6"O�$�ƩsӠ��Ǡħ]f��	'"O|��T/3FƁ�C@�1&c���"O�a��ͧA	�ȶ&E����"Oj���H�(}�b��BRR�؂�"O����j6>z����Q.�v886"OĥE�9[����Z������"OB�!P�C�\�t̓����"�[g"O��
7�U�@⮨bP�L;l� +�"O9���ݳO����1�߄im,�u"O�����qڸr��
0l`�@�"O���`�ۚo^��J-ɛ �H���"O�|{��/����Vk��J���[V"O����僮�pA+�lh ��"O� ��菈GԸ��dʁ��F3�"O96�7RN�Z�	�E��|��"OFD�s�ιXݘ����H6�dP�"O�A�(��Jg|�JB��'늬{d"O5��	`����%���p`S�"O6ͺ�O73����l�}�B�X�"O$t��#�* �Q���!w���C"O&) �al@b G)u�P$z�"Ob��$,��N��Z�nS�\�D-t"Od�ć$!b��R�K4���"OL�����,M�"-
�h����"Op���Jߘ\7�k��ɴYZ@��"O@5Y�)�b�B [��*�j��"O��ʂ�ޞ[��pU�y�`:B"O�s�'�'��� �����@�"O<��t�\�0��\˕+L�
� �@�"Oj\*Wo��r��#@�?H�"O�5���`v>������`M���&"Oؘ��mǱS�$i�OD	Fn�v"O��ҮJ�2(5�.�)-"�Xe"O�ԑ��RA�JPx$��.��&"Ojar���q"C"��`0��b�"Ou�sF%���n�"5C��p"O��K���PzQ[Ƿ�N<x�
h�<y��.b�Z�y�,۶���S#�c�<R�O$R@DЀaM�ܰK���K�<��Ɔ�R��9:r�K�^�C�.�l�<��`��B>Y���M�6iTh�I�i�<䉖<@X�k�oPL�H�8��e�<�΅;_>&){筛�_x�`�K�d�<����E�ҐH�̈́89jUh6�
Y�<��S�&?�T@R.U����Cn�S�<	I��H��0! P�4�����e�<�-�0٣����ܳ���J�<�-�5>'0<���5xV���,m�<�B�]C���b-E�l�|ԓbC�<�D���ؚ�^V���HW�<1! �u$f����I&XB�#r��U�<���V$ @  �P   b
  I  �  c   '  �.  .5  q;  �A  H  MN  �T  �Z  4a  xg  �m  �s  ?z  @�   `� u�	����Zv)C�'ll\�0"Ez+⟈m�	�|��:F���DA$������%\�U�b(\�f��d	E/P8cꔐ�gH3]��%Ib~xݮ;�p|��'q��Yh��A�Ժ@����R��a��3|-�M	S2�@�S�X8?SjtS��ղ"�0��� �-����$H�z۴�Gc��Up@�KBT�R�B�K��Ԓ[�H}��[K�t���+T�в�4T}���?���?Y��'@&��k
�"��
�jvy������I�MS�I�����O��0�*韆���O�]#��Im��iB$����Z$�S�O\���Oz���O,���OT����'��Da�hq�Vc\]�i���(x��>�O��� !R���XV9�℀2,�듨O��.�|�Xї?Q"@�2*cv��'��1� a��O�$�Ob���O��$�O*�İ|b�wG��hǩӧ��d��C���R�E���Ks�d�l��M�����v���@6G(:�����"�^}c.¯;v,qy��W?�\�Fz���w���}��E��H�"�KG�+(�ǅR5#T�9J�B4hܮ}xS�B2�MkD�i�V7����)��U�m%�B�T��9�%��&� �h����o�"�l�UG���!� y�1��U	]��d
	Q��8�4J<��eb�pUÎ�v� ��w�ߗvO`����9�hT��
�v�`m�MC��i|���:s��{e%^���iG�
���^:��jAAU�bY`a+G [|b�᥅���X7-��q��4v����FX���Q`Y9@j,���K��x���d�F6tH�P��#��&��x�B�`�$T�	m�D�1E����$�GP^P��#��4J}h�GLn���5���<�Ia� ��ش��)l���\����j��g����'���ߟ���?��@�_�H�<`�@%�lZ/:��K���G�y��N8 x�ቒ|�`�s�4���R���hH7*Q!8�zi��o�5)���[d/2O�Iv�'�l�<1�%�h���!f^
��'��ߟ������?�|��'��|�a!��&� ��7��6�y�N��6�-WdJP��j
d�����h_���7�*�	I���?Y��3S�����c!���	�.D��-[�'v^���W(k�}�`߫mJ� ��'o���a �f�h�eˁs`���
�'p��[�[�}���B�MffX�
�'b~�����0'��9;�fC[]��b�'�ƈ��aH�g� -��N�FiZ@���3�x�Dx��	S�|⅂���(��/ m�C�	�/��=zgU!2�5	���	+@C�	*8uBZB�`����7kGtZB�I�Nz`iiq̓�ކ�S�̆6gLJB��2l�zP��/;An��Ɂ�&GlB��'l
fQ��+!9�K�O��(���{���	1f|�����"�c7n�cNB�I�T+�)2�卜��������C�I�w�hB���+��PӁ��-�C�"C4B��7�)��tk�-ʏ>߲C�	�Hq�a�����x�/[�����Cg�Xm������w��XaCjZ>d���eʟpC���џ��4)P˟�����\����\��mm��	�D���w�0�Ӈg+F��pah��.7�}�	�����ׂO8p��Ȃ��Nv�C!gS>h %�ƒ$�>�#&�M��I��O��������  MR�	����4b�{�AӼ�Vp�'6���ӼqO�aC��/j�E��-\7l-6b�@�'�>�s޴*T����JA�	����'iЃR)@���i��'�R�!��^�O:��k!c┡A~���눶c]:��� !D���#�w%�<�bF���d�f $D�X����A��Ȗ�C62��S�E4D�L��ė6:�Ԩ�d@/??4B3�0D�ȺR�S�:\���&w���#�2D�X2�A�9v�1《�>��a����'��{g��?�������}y"��|<�H{� 
�x0���$D�����4�e���lZ*6�H�j�� *�	�OҒ��$��2��Lp���7U�QZ���z�td"�o�[��`�6�n�0���Otl�uL�,����`Ԛb�ɠ�kg�h��'����Ș�?q��?!WA��%�Lɑ�[�o\z�)p����<�U��׾���87�	;Ѥ��T�#��	��M�A�i�ɧ��O����D಴a]� �.=kaN�9(����O��������uy��d�$����R*w��D�s-R1 �
9�򁁇9�.Q1��B�����K����	�b\&Y����*6�V��V�M�	E
��g�LuGv���l�Zb4P��Å0ej}�4�˻^x��b�,��X
��'��R�'��)gJٰe�`��\��0	�'̚!�%��}y��٬ifh�M>Q�i
�Z��aJވ��' UQ3A��l;@��B
�5]����Iqy��'���'��l�S�V `6k�%Z�N�� 8h�K��^������!�z<YU�'�R$3$�.p3>(��e��u{��A�G�Te"r�C:����5MC��0<ї*ٟ�	b~����e���b�%�(\Z�*�ƒ��䓩0>)!�C�{�&��E�� H��S������x�6yPUm��P���hdjC�&'���Ay�!���6�%���|�����쨖�*�n=k���&>Ċ���?!R�.R0����G>*�4H������K�aI,|����(�]�#���KFO�Uq�,�G�L W@�D�d�H(5��`b�⏺$�d�A&�z9�'/��K��?Y��Ik��@�կ{>|�ɕ��A*��r�*D�H�DΜ�xǤ��` Mgu��q�,����>�A��̱]����'LA�b1���ڦ���Ɵ\��>2� ���c۟��I����IѼ�#�9$M��� �PwZ����XN̓T{�!��I�-gD����J��lɑ'^C&b�p�RD?LO ��3*B<���Y �Ź?�ɶ�2�$Ÿ?����V#[Jh 2��,6py2�mN�DR!�ğlb��D�,��X �&AY�ɯ�HO�:�Źu�R���mHl�t�a��.ĤL����������Py���4ЪP��5����PH�z�B� *�pqAR�^�
�(&�� Jaz,7E��$*�H9oV�$�B/_�u�` ��N��a�t����	�0=y�ǜ�L�|u��ݐN�@5b��ܴ/����I��M�*O���O|�d�O��:�Gؤ[������"��b�CH�C�	V�����	�
u-�(U+M&V���O1oڟX�'OZh�Ӥ{���$�O ���,ᤈ��џAF� �B��O��D�e*���O
���<���P�f�C≹b���iG�֠c1�x���`]bŇ��+t�̝�3�U���z�R,m<"<��ͨ)U01��&?�Q�)O�!hL��c	�qO�E��'�R �<ѡo��pH�d�V����H֟D��ן�?E�t�� 8 �z�G�\�X�;��T�?��!���,I�t!�D��Ē
~�bEZ0y�6M�O��d��$7�L�'R�'|�䂝y��M�4D�@�
]ƈ��A2�B�' p��À�
���O�|����x&r"�&�r�2�����^�|T��fC�:��Hzw�u/����\�f5d���Og�����
�S�$)�P%�/ȦU��O�MR��'F�7��٦i��k�O>֝�3�8�5!��!B��J>����0=�L7S��Q���:J�MQ�L�W�'#�"=)V(ήD�,�哞5FY�P<P���B�����(�B��O��d�O��D�LI��4�V��(��r��5���񧉁�P�1�܊7 c>c�hP���Z�3�^t�r1�/U��zm��9��
t�Lc>c����\�T_�<�O�f�� ��O��I� ��䟘G{R�Z6Op>�p���r|v���C)�!�J9Yr���T�rp�z䊑$c��ɉ�HO��my2����T�u�]�#R��*6���Ւ��E���ԟ�	iy��DKȭ,�`��O?��ka'!����Ǉ�ZP����%G����M�`9��c4�X �$P+F��
3�P��d�$V,D����O�b����c�����`d��J\�@QM3 <��'uў�Exª½k��0"0}�=8G�_��y��7kd^Dqw�
�q�h��!	�����X�A�l��')b��k�!Q#0�<�f��~�����I%��3��DW(�5ƌK_$��RQ%	� p٫�ē�BI�ȓ{;���G%��_��{��҆R�8��ȓ[E�-�A#_�U6|��a�L����ȓH�"c��-��2���2c�I2q��~�ŏ��&:Fp�AI�+5J �S`�r�<�Vn/`��B!�;T�1q�U�<yf"^�@�>���ՠ�H��v��y�<!&aη"��Y+��N�k(~� �hLA�<������6����� <EԄ� -v�<y��
w)6M�BL\y{�y�*���\�`�,�S�O(���r���3�O��L�@�"O~$�5,�;;d5��ÛN.��Ҧ"O(]���9�~���ˏ�S#��1"OR5J�c�2{.EKf� b�4�b"O����J��LX��u�U<A�ޅ�T"O�L#�,J5Y�0&��"�f�Y�X����/'�O�����Z�!WI�|��Ru"O� R�"��͘Y�DTq��H�!�`��"O�$��J��:�^eh���\k<���"Opd�V�0h��)R��VI��"O�y{�h�)^�PD�Se�
���D�'An�R�'e�1� E4TV��2�K?U��5{�'�ҝC�dZ(�`T��/�S�rd�':����F�*�6�hE�ƊJ;n��
�'n����L-?�丢�C2J5Z	
�'|�t"6�*�>q+��-ELri
�'S�@@C�9Pt9P7%��c��d+]�Q?�#%��B����3�$9 �� *�!�d�$���!�o���r�I*�=�!�D�$,q�'�B�e�\ɠ6h�	J�!�dKb�=�Rˉ�>���ؒ&���!�d�5]��� *�U����̉)(�!�d��;ؠ�BE'@ZxqR����m��nҥ�O?Q �F,*���Cm@,h'*`��&�i�<y��Yf�4��UȄ+l�PxFf�<�D
�0T)�7�Ƒ���f�_�<��+��:l"�p��4�	��-�s�<хKT�Hq�l����'�m�e�n�<4G�6 �N���ʅ0�n�*r�Ty�		��p>9���)	r���R�x���ɱ��{�<閃�=����e�ρYW4����o�<�O�j��K֧� �
2��`�<ѧN�r5$�I� V�.CR\��QV�<i�F�k����ރc��h�uNx��#�뷟���
.��HA.��-:JDB�,#D�,�dJ�	�F%a�Q�pj@Kю D�@�.,�TP� ��#�0��1D����%V�9�M(��ēG���H',D��c�ŋ/�)PIC�H�Ѱ#)D����BQ�e�FA)���!�R�QF�%�h^�XG����()��H�B�:t率�y��6o38�����I��m�(U��y"�WP��=�Qf
CgF0c�DƤ�yO	#X~��#���p`X@cS/�y�*�* �r��2iq�b���y�&M]�av/űT�&Q@b���?)#�o����4i�A�F�-�I#��� 9��9��4D�xC����������s�z�3�,6D�T(���7(�t�i�جQ�g3D��B�ց��p��K
u6�Qq&i1D� 8c@K�x���eF>@ lI)�;D��;/�H�Xqr�Ŭ.Q���<��*b8�\�jM5m#�,a䫖� 1����3D�ȣ�Yd�\�f�?�:@k<D�`q���w�V=8�� &!��=�-D��XlR�J� ��!IZ
^ �22�)D�;E�&+�5�..b�0��!)�O(�	�Oĵ�ކVaΈ�7��2du�	d"O�ѐ�N��(:���Uc��k�"Ozl#r���h��f2b��b"O�����+�"C�B�:y\���"OBa��瘉"i�mؗ 5>|�p"OfZ��9|�8`zUA�v(��
��f}h�~:��[O����х'�$�X׎Dt�<ɒ�
p�p1�!O+U���KMX�<1�F�P��� ����Q�*�R�<� �bcX�0]%(��a2�Y�<�"�V�-��4�T�� K���vK Y�<�I�bCte��́�e�xyDA	؟����(�S�OH:�[4�]�	NU�pF0�
i�#"OZxY��S΀ R�ʤ9�J�["O� (գDIOQ*�$Y��\�`�<P!�"O$���虅)[�D@�g��2��"O�Hq6�Nحх發m��X�G"O:�j�D��t=�����0� %R����=�OXؠ�њ:�
�A��^Q�U
V"O(��ӅǯZ�z��
�Q��� "OV
Rn�d�ހ㑞Z�D�[�"O��cňș.���Ɂ R���M �"ODm:�iޓi��9'!�4!�J�˖�'t�0�'U4TZ5�CI�����ߧAX�-B�'���J�EJs$��MR�"F���'�F,郺J2	�G���J�)�'�hh�Ϟ6mb�����X��ҥ��'��&����R�˂
{�d��'��|�$H��q�F5ˆ����ߜR�Q?a�#FU	C����CbY<��5�=D�P���@�^z��E/& D"�X��(D�psC�G�V^��� �e�ţ�$D�81�KW~�<HKqe^1e����'7D�S��+6�z�� ����94H)D�0�� +<���SD����R���O�L9�)�Xta��n��K�"�q`�k�!9�'��⁬��h3�]Ao�iʙQ�'�T�vH�]�u�/
�)�=S�'�~B�8���#fP8yK�'���ke��l��|(��T�u	�A��'b&`�3Ǩ|��x��j��,O���'А�ꄌ��J䚔�p-�v� �'z�k��e�)JWh�)(
P���'�(���(k�D������5y��)�'��!j��8-?<U�5��F��'��ʓ��$tb�)! kO�R���mh�A��<�M�!R<6�ɣ0.��n��ȓy��!d�1�����D�<k�A��<�D��D�J�造%�"�*�ȓ"�j �r�A<d�d��"NxV⁅ȓ/?�0J�ś+� e�U�d!��KeNdpSBP:	X�=�A
VPp� E{r+�&쨟�t�L�*� \��� ]D<���"Or=(���g��|�A��3�0 "O��aa�F>��p���0&�=ɱ"OH呰lW�a��m@���-"�@��"O�h���%q�"]�s/RaV!�dA'v�=�4�L2���FǑI-2��O?1P�J�	`�Ձ%�?��C&l�<��g*Q`�yԤ7�x[R�]�<�P!_)`��!,�6@�n���k�U�<��Øe�򐻴��43�BY�4�j�<��H�S�H�C�14J�%�b
Mg�<��/֥)�a"�̰g��L�Q_y�kV��p>1@&J%��xÐl�O�z�ek�r�<YG%ë��H� ��*t�B̠�Gn�<�6�
;3�����  9DDYr�^�<)c�����үC�I�δP�*U�<����67�ȥ�CK�0dz��P��{x�$8�H����1�)Z�(�b��׭x��5�3�;D��16㔿\��Q���
�`�%��"8D� ��蛅F^̤���?����6D�hp!�9Y� 0֬��s��(gm6D���ŀ{E �R� ���'a3D�|#��XI<��y w�|���	>ړ �F�Tn�_���P�΀�f%p���y�e]<y�O��f�����y��\�Z�Z\0 �S+da*�1�K�-�y
� � A�Τ|t��Q�3��!"O�$q7�K�?����-Y�h`��"O�:�I�/Z.\���|����'a�Y���Bl>!` O���l �-�j]��'i �31cA�1���BSH�8;�XM��'gf=��$Q�3Jl�	G�-B����'.�����^������J=7p�hx�' ���6���H�y���.���c�'�0Ep�ჶs|���/��P���.O0�W�'�&�Jʕ5�M�1!�%?����
�'^�Hk�Ds�&�����7�J�i
�'�b��7K�X3��Z�!�'�E�	�'�0����  ��`�i?6�V�	�'�>���.����II�x'�x��I�f0�;V�ժR����E��v�܌��R�t��#L�5����G�dX�ō4D���Qo�)������IȢ!��-D�Ti��];5Dք
��G��8��t�,D���j߰�PQ.�\l�1�)D���Sdp݌�+r�í�@�&�e��F�ģ��bn��	�ND�
�4�80��"�y��O��T����~	�,��y��̃ :�2'���h|	�sB_<�yb*�$O�&2�dS�]�����C���y2O�e�!��P8�|cscڞ�y2�Bf��,P�)�{�b���֍�?�f}�����m+tT�U4��W��DnUX�L5D�(��r|�{��և ��`�3D�ȡ ���aW,������3D��)��U����0m�o�TZ�1D�41"�[�.�@�/ӵM4U:�)34��؃犡"!��z��J{���`hֈ=~Z�)��O(�	c������v?Y�O����JOK �� A�a��`�`+��(��ȓX���r�� hl���0�@؇�ZX2]�V�:Z��{�A
Y1��ȓ#^`�B̕�a����D蚌.� ц�Y�l5s��T�@������O�d��YZD̊�	C��)�Ȑ�Y� X�?iĤ�{����C�� ���"<r���bY-[��B�*h/j�	ݜ�zYS�he@�B�	�ߚ��e�F�(>�]� �8�rB��+3k� ��B:<fD�P�f;UXRB�	���VM�6v�����es0B�	�=��9�!M�\��x���'`�]"��IA��~2C�(1�Y @Q2H��g���y�k��,�� ��m�7�
����ך�y��B�p(*82F�7/p0a�ǁ��yR	�@����' .�@���dӛ�y��G�B���/�5O�h�٠�y2bW�?j���e�Βs�������?T�d�� ��%�)L zӠ�.]Re��=D�(�Do�F= Y�Ѧ�4b�L1;Ղ:D�8yc�[X�� �ľ�rY{W	3D���� ��S�,���H
G����i<D��hq���I<T�t�L>M�����8|O4(Ӓ>!���J�����>���J�m�<�r�: *P) �N=b��<C�i�i�<I�"_xV� kv�I�I�T{���h�<�]�� J0-�&��DjKa�<94�2/�1�U�KKR|�y`�VC�<����&k��`KU�<<j$5f�C�[\81ExJ?	zcB:Z���+ܢgݖ�y��!D�\��HK�G���U#[p��Q�"D� Y0*ٱ&��trTO�#Z�����5D�� �9A���	־ ;�j&�9��"O^�wFڢiL�� i�6_,�R"O��$�Dpp�L R��d��Qg��OR�}�^DN4��NO+6XUYo�nL��`� |{�E��4	0YrG�L8�r���zC�<P���Р����D
h)��|�k��H$�``��Ȅ�t��! ��1шp(F��N�8��ȓ'���
�{!X��0�H���Ɏ~U���ո:S�(�E� +z�k�/m�!�V93���S�� -DVu�AN��w�!�DM)N��j�G��W.�(�ClʍIz!��6I��P��-�q�P��
:h!�D���,�Ҵ�g��(�)Z&Xџh�jT��M[���?��O�tE��i�p�+VȔa�pe���/������?��u���Y�������;Z��I�>5���]���O2�0 �ӗq�&}ؖ���Ia������<�,�z]�����Orl�y�n!�� U`���j�'��5�d*�;��ԉa�:~ 5���I�&ˬ����
���D�P��%���?������|�����܏�fК,Ќ,dN�Y�L�qlџ�����E����Մ�..�<m��J i�OvAВx��I�\�
0*� ��µ�ڷ5U�	�~��7���|Γ(�2�vR�d��%�3\�eX��� ��$\�	H��-��OlS爖�M�z��� =7r���O��NL?���9O�ْ��Q�ќ�{d_H�8SS!ҬyG���F�l��O�U�O��Gӕ[d�q֫[�Z��J��~4��O<���S�z�D��wJ�>]��9�bťo���ɪz���'��'�f52L��۴Z$xq �
p����h΋%�z��'!�����ȟ	�O�9,��9:��G�n���G{?��v�T>�ɇ}��xl�i��j3V�U
��\�t���F����d@�sJt���O&�"��ɖ k���Y�A�7��P�ju���d?���L@~ʟ�DÅ#��H�YW6ip,�$ϼ�SB�W:(�"�RC؟t�4$�|���ړo����o1D�H� �. ?J@� ���(�h�X��q��D�O��?i����|��|:r��"��K�52vƜ�6�Xm���%������O����4���1��\�����aJ�E��Or�4�)���Z���B�(�Q�\�K&�&B����u�؟V�J����C�I�d�咱��0��h��B�PZ�B�&'�ܱ�X�@)�-�q��B�"0�J����V�� 6��<_u
C�ɻo<!Y1���*΄h(�)hrB�	�i�Y�gش �UK@���H�C��:�����_��H�``�m;�B䉆08-G�̔M\�bG�э�6C�	-t���w$)��1�G��'l(C䉅O��$y��X/'���"
�4C�I�>� r��* p�{ �L��⟜9 ���%*l�c�dR�ܹƁ؜	$6��bCD9(k�M�1��5���n%�D�sڡ��Y��ҝu�x܁�d@	3X�˲��d�m8�
�R]>��׻Gj��.��r9(�]�[����"�0�:��WBR�q��&I��hX�� �̤A^ܡyJ>�ê��Ӥ���H�5�T�Al�V�<��	�$La(L����I-�)��MP�<�V#�:	څ�vGN�B؂<����N�<� ��l�,���͆Z���%�L�<	� �d����u� �#&حj'�]�<q�e 3exe' [|�P� ��\�<Y��
�X�ڰvgEuŌ@j ��N�<A�E��L���! <:q�U��RQ�<�"�� Vd}�@�8U�<���@�J�<�N�B���!)�1uF��fH�o�<	�+�35M�Kq��-3*�����m�<�P�Sd:f%��L$(�XhpD�g�<�n>b�l]���D�Igb�m�<� �p�7�� ��d�ᦝu\�}��"O���A,LC~ !0刘pA �k@"OM1��R'�)Xc�HAP@�"OH�K���+X���"�H��ӈ-A"Ox�р�Q�Hh���Q���@&"OB��WS�眨�$$WV��-B�"O���S�*����艮I�>���"O��`�E�&�RmJ���k���ʆ"O���֣�9R��͂��ú-+����"O��i���
 j��w���P�d��"OШ�T��0i�<}i�!��&��0�"OX�tS&#�)��݊E�Vp�"O�ѻ�"F�|���8�@ê�Z�"OZ-T����K���N6�!�$�H�TX#�OS�?�h`'�ΩO�!�Ѳ]�i@�YN�����+�!��I�����W�V�pd�82!���
!���&OJm�P|��NO!�$[q���[��C�H�٧$޼U!���U�(���V�x�P)ႛ)o�!�$�~&�,(��)jo�lxg�Ҭy!��>xb`qAŉ��#v �J�' 'g�!�dE(3�� ��H.5c����Q:6�!�����Z���Q�ti#7�>!��^<7�d���������!* !�S�N0ɂH!{Rrhp�)^�A!�,1��K�aS�86D�����nX!�^�x���;a3Z�ꐊRQ!���R�ƈb�܊J��A3&��� !�d�7?����Apa���N��"Or(����#t�(A��7��ܹ�"O��5d�>�
��ekՃR%�("O�{�#N�+��ܳ�	ճ��Q"O��U��7w=�T�b~�>�1	�'�i��H��ZAT�Ȝ��8��'P�et.P����#NT��>���'UH�Z\C�v][������'�j�r ��RI�њ�͙���^�y2L6�cV4^"�8� T�y�,I�H�(�8�a)&o�|A�l	��y�͈�)��H*���o9 �+pmX!�yRFx�`<�`�	�j��T�W�?�yb�X� �Bt���f6lhqw�C��yBN��9�H�ň�T�� �J�<�yb [.8K�hg��RL$�Kњ�y2�گt���U�J�Z ���+M��y��eY7kK`�h��5�	�y�F��$Qa$��<�rQ��u>!�D��	|h� �ӯ3o��JǨ�$+!�$"9�
]�o�,�R �Ǘ�!!�$ȜqC���j�0���p �[�!�$�l��YQ�dDz��aDEQ?!�!�Y*N�;�k� Vj�F��M�!򄖧��ɇ�%i�i:W���\�!��g��� ��V�+����Vv5!򄅰2�楠��*#���f�52!�D\�O�&5�4�
V%Tq�+ӿ !�_��r��DL�^���HN�6�!�$��N���0ڣ:�$ha�fӀB!��P�f]
��J,V�����N�!��y�~�(�+ޫJ��0�#�9�!��C5=5�$����	���1!�(!�d�1	Ae�U��`E[S���}�!���{a�P��̻vnBP��M�5{v!�� >}�$�Ϟ�&�KPfC�QYL,�R"O4�!����a�4J0�M�hU�;"O4Z.�:M)�T�ë
�Y8�%�"OX��L�PX��x@�ȼ<�,��6"O,
rHA[�`�� ֨P��� "O|M�2jV/�@j�K>����"O|E���aeVq8r�hvb�r�"On1�ޘ��`�b�J�:����v(/D��b N]/V|dKc�
�4�Τz֧.D�l�&�L�l�.x�+9
1���g.D��@�M�;V-���>r�EBG�+D��s��-W_P )@�jŚ�9T*D���fK��б�si]�i�\Ej��&D��3RNE�KRL��nZ;J6*1� )D���Ԝ�Ҡ�b�L�q7��@�%D�`�޵ �d�G)ߡT��c�#D���d��>4a�MG�&d�1@A!D��t�_�l����O�FG8t	`�2D���#a/lY�p9Si�9qw�څ/D�ೂcȄy:�p����򒉡��?D�h��T pi�+��%�vu���=D��㕄Z�G����̇�r�d���9D���s��)~@ZQIV�Ǻ���<D�l4)�	<�dă�d��#!�s��$D�*6b�{y:�e��>���X�$D��##ᙬZ0tPFeP�^J|��/D��	WnƦ!ζLZ��y�� ��.D��Q6�$"��@Fh�o���!!D� ن�L�����鑊f�H0>D�0#�M�@@�!L��ԙ��6D���D,~�54$u{v��1D�DzE�	T���9"��:I�A��i"D��	��_������0S�,�8w�:D���aD��D��c�Ci�$��'�-D�y!�p�`���@Ϭ]�,�g�,D�B�a�@qL,{'(5Z5�\Ȧ.,D�����̡w��˷�ϊ ��$�)D��{�-Ŏ
{T���
mB�8��+$D��a5���Zg��Y�+�9����c"'D�D�V��/g�d�&OI D�� @W&D���� aN�Z#F�+����#D�L�� 
�B��B�<>7tB�3	 �qw�Q<D "�N!@�`B�	0>�I���ߦe�F�⦠�w
C�	!<Α��ee\�ᛲl1��B�	�+�b�3�ی^�ѻҪ#
��C�ɕd�F�8%d1F�b4���:�C�3�z��-�� ���+0��q��B䉄xr aIS��f[��6	�Z��B�I�E�FLѴjȪ���	*��;Rm&D�K%陆y����'׉t|DjR�)D� "���$VJU�H=LZX��)D��b�.AS�d��ԇz�ؗ�&D�tyT�	�"A�4Ԕu�`�J�`#D��	%/�5�L������	q:�{��,D�<��"ݺTOVUK���&b�R�s�d.D��1�+�,!�H<���G93��J�L)D����)V�?����U��-(
r$:��:D�zf�pD�S򠁅/�`Y�f3D�h��7!��ِ��I�Bp�Ԯ2D��5!�i�Nу�%G&���"$D��[2���Y����ņ�+k�i���=D��ƠJodz��v�_�i��):��;D�� ��h��M���[�cb HI��&D�� �غ�̉%yξ���Q�5�|	�"O"�(d�ւn�|䡧���"T�%*O4 ����j呠J�,S�Pa�'���� �_̐��S�t9�l��'��Hd�Z�����+W5k�89�'x�#���m�&9H��(b�	��'��� ��P�#�8cU���is���'��R�� ���-E�h���'�1�A.tB�rS`�=aټEc�'��I�*�DIӢ�<(�}��'�	ƣ)Ypm�G'V�� D;�'��!��_�,���c�BT�-�5��'b�����;��-���?[���'���τYe��!ffe�	�'�@�X
	�\_��PҸn84��'6 d"2���"tuyB��Hp���'�8���ɀS'D�oB5T�{�'g�a�t�̽`O4MX�2��}��'r�B�)����8eS$�X"O����Mg�~H��HM�cA��p�"O��Ҫ�q�b��'KF2AC�"O�r3k�-���U&��s4<L��"OL��j�T�B��@�p]A"O�E��j 3�T�C�;C32�xP"O8p�çc�ցD��()�Љ�"OPub!
�y�,1��4 	�ʑ"O�I;u�3q�ĝ�3�
I	�"OTѦaЭLS(�b)A�&��Ƞ"O\�S���n��Jw���{��b"Or�B�Ǚ4QI"���ڪ{��8�"Ob娕��7;ʾl��m8o0ԑA"Ox�[���J��i2F	]ʙ�C"O�,�7gň��\�C�FCr��"O�Ͳ ��|�^�!75�.hxc"O�QH�O�)M��I�����p"O�墐d6�~��ģ2��X�"OLaʖF)X�hdb�O�����"OP����L*�u+���kv\i��"O�`S����k�6��rVhR@"O���'|(��)F��c<���"OD��W�L
\�t�E�M@� �"O2�0�������s�"O���e�=z(�J�bO�r��P"O ��BY�aP� ���pq��f"O\��e��y�ܵ�⫗;r���"1"O* �.�!{ƪp��T
�0<�!"O�32�ڶ�͐�l�;j�h"1"O����B�	��m��ʡ��IӦ"O��3A&]�E �U��s���c"O�)�%�=�%�%{~e@ "O��Y�ΙlB69 5O�&(�"O��@�`ȶ<��1��M5➜!�"O� d��K}���j�2����"O$������P��Bj���HA�"O|]�Bg^�dHf�	�=A���0"O��e�I1p�X�� )_k��И�"O��ӑ�+D�L��^*s�z���$��p��e��I��\��!ZV"��M>Y�)��u,,�ҏGNϘa/A!�C�I%U�b���DV;�^`*2iY�~Z^B�E*d{�D��=Gp8�
�C?JB䉩Vèl S��jQ�u�eMF�4�0B�x"�7aQ�� 4`V�d����ȓX�ưK��C3G�~}����UׂC�I�,蜝��Y�
<Ȧ)�'�DB�)� ��� <_^ݛ����Ĩ�"O"��f�tX0�q��O��tʐ"O\10&��f��<`쐲S76�g"Om�hb}�D"T�Cք�Q"O����(Q)B���b怚�L��8�"O�Br,	'0;� S�O6h��d u"O�Q3���af$���%�B���"O"�z����A�
tq�(}��4��"O�1� ��=$���s'AW�oӤ��c"OH:�V6%���rf��.��8�"O\�h��5���P���E��Y��"OL�0P�j0��u��~Mj�1�"O��E��uB�E��Jj��9He"O���QB��b���k ٢0�V%��"O���/��2x���m/&��x��"OV� ��m��D�&P=���BD"O:�"u�"H�#��!b�pa1�"O���E�ҨQxXpd��~��x��"O�h� LN 0	�.:�0Q�"OP��Rr$[4fY3|�.I�t"O�}x�O	zptˡ��w�xL��"O�A����6�J�k��T��"O�i�wj	y��bFĒ/!�
!R�"OT�nV��`̩�˃ ���"O�"��2L��T��!� ���"O��JD�w��)��HJ�\hd�"�"OFp�p��y26Lۡ�� L�\LY�"O�I`F�Qw�|zr�.K��a "O��h�4<�sE��2}�8��"O �W��z��%���0JZ�Q�"O6`ba��"<���֮��n����"O�Q�׮^849�e��̃�O��[w"O��!S�B�l��mhC��@��Y��"O^���(��_�Z��Р�A��p�"O��GN��B�H�#'�/1�Ts�"OYC7b �TZ<<��gUh�x��"O4e�� �*b0�YJF�ݻ23 Q�"OF��Q���;���P@[�0 Q�7"O�dz�H�
	�dVf��Q�]"0"O<Qy�W7X�HX pˀ��J���"Oa`��L[2�	��˃m鶌3"O�p�T�D*/Մ)�(S�S��=��"O\���E;G�b�J�e�=K\@��"O�0B% ǩ=������ȍm+��c�"O�9�ˍ���]�l���v"O�H����Q���`cc�x`�-�"O\��%��SG:\��B� {S����"O����@ֶx9�<
B�.I(��"O�q��
[�q�(#���}fN�"6"O�e����(hJt�" E�!J��"O\݋G��
[R`��'Y@�4�R"O:ݡaNL����6&ȨY����1"O����Q;S�8ݣ�5�B`"O�qr�J�A�
-�����8�(i"O�Y��'7����f�{��8�"O~��veJ$Y�R}Ӂ���r�vL�"O,��K�7֊`ڒ��b����"O�iB���:�V��ƴB��@�"O�8���CD���E��"r�� "OL��T��"�-���Mu��`"O$� �1���k¥�)?mr��&"OX���u
D��4%�6��I"Oؼc��
 ~�XZҤ��Tz��x�"O�Y�V��*�Lа�K��}aF��"O� ��s��ݷ4@�E �!�9��"O�baV_`r��%!�3��hd"O<�⣣&К�q� M��Y8"O0|a�*�q/h���iC� �t�`"O(��mH�&��:9�����C��y��[>�8#�/��7m��qC'��y�ǉ�1!�U#P��(2��h�!(�y�
��ZJ
M�PN�0�
!��C�y��S�q�US񩋀0��ċ���y�$�;trd��ڣxʵ����yRJ��`��7j�.x�%KK��y����EF�PBpXFn���y�@ r~���$��8j�-º�y�%�pH+�-$��`�_�yJЅn��J� �O8z]ۃ��y�)1Gp<�Rc\"H���C���y�o�V��B"M;T?�옇�C�yB�԰9�
!ʂ�ۛS� ��V �y�!�0`��d:b��b���6#��y$��8��q�Ę�s�>\S�NE��yrh0'������[�_��Tɤ����y��]E��<�e�Nv�E ���y���D}+!��CX1Q����y��U;-!|S�h�5xx�P#�FY��y�gX�LDXE� K�{��ct���yr�N�K��UH��Y�\7�u9� �&�y�I�*!s��`��b�ޭ�7n���y�"D�lF�s�V�E8�6C[�y��5�:�@N�7�
ث�y@��iq���Q3[J�uW�P �y�^4��Hs4�
$j��aV���y"#�y?hUPqM�r�J��.�y�C��|N)`��h�d&d��y��Ԩ
f =Jħf�%QmS��y�R"T�!�C3b��
4���yRĔy��u��b��E N
L�!�D�<w�8}z2%ܲ"��9"�'�!�d�=X�U�%`E�!�=C%�-0>!�$_���t|QQ���
%!��"���f�	i���@�H�!�Y[x����.3[6쳂&�o�!���*�-Pt��ODaZ��S�!�@��d� �#-@A��l<^�!��];OE�xz�F�@�*ȋ���8�!���q�REC.���@{U��R'!���9����.�+e�le�� �c%!�V�@]�UC�O]=_%�p��K�P!�DU�]$��a��:r� A �[���'׬)��Ñ�
���)���$�B�`�'����5�ܩ�E׉ڭW�0���'#�ձdF��@Y���
�U��c�'B@�)a�;5n�UA�!��`�ꐀ�'�܍2��\�Y����!� !�X�[�'TQ9�-|n�9�j���.��
�'!�U"B�G��6�+ৌ�I2�)�ȓp��Т���yy����߲�8���%�xHۣ�P�P�T*B���s`i�N�<1!AP9H�����F6������A�<��Ǐ�N���6b�bTP����R@�<q��͓)�X���F�Y�i�qj�X�<�u)�(h�^��3Q;kE`|·�V�<��K��&�XJ$`�ko��Ё�T�<���X�Ht��e�e�J`
CP�<ٕb?h;������P���`�Mk�<� ���ߏ������0���"O(�9f���-@Rh��n��I��@9"O�xX6o�u�����K"\��5�"O�������	�C�?j+J�ۣ"ON�C)5P��0r���%��HE"O��[�ݺd��[�@J�n'�<��"O��9.LV����G^قp"Or8i�	�-.$M�)b4IhB"O�I����j� Y�WB�[�"O�]�Q�T�tpM�g���H�t+�"O��5�&K���&��a��Pa�"O��򋃴 ���J�G��B�X�`�"O�������Z�@DG?��$��"O��'B^� t0��E��l�� sB"O���Z--ޘ��B�ċp]��a�"O֕�c��<ځ�R<�B̀�"OJ�`��?dH���߉%�ڥ��"O����ӸP��Ћ��Ҙ_�V<��"O�$Ó����S#A=9��i""O���4*=yH�)���$��K�"O���#�X�I��%ڣTHG"O��#���\�[Ӎ�:2c<@�"O61c��	�b��T�"0:�2�"O���`�V;-0i�LmGR��C"O4�����W�xd��"�e�H`I�"O��f��Cg�uI��A/ �˗"OnI�v��,!�5q�Om��,P#"O�u��s�&EB���'1z�Sw"OH�	&EO�k�������:C��C "O�@ )�I�R�Ab�fx�Y"O��HeE�3V�.��5�B�5k�X�"Ox��$G�&�8s��� ��H�"O����K��k�\�0���/�=x6"ORXB�ǁ���5G
�A'�p��"OR��@��gН�tŇo�zPK�"O��q�ԱyxIC���x��,��"OD�p���YyX}��� ��hB�"O� 2�!�BX �)X?3�0tK�"O虓�)�:qp��894�k"O��`�醅�\�q3��b
h��"OJl���5Q<8�!΂N� =��"Oθ�#��J살�ƠG�U���c"O(
`��y�XD�Շ�$��4��"O�$�g��UoƑ��'�2����"O�y���2T"���љ@�6xh�"O=!�/��!�ƌ�PoZ-�$0��"O�P����Px���V̀X�"O �ѥ��,�Ғ-�(�ĩyE"O���%!3Iz!C�cõb�V)"'"OBu�!g�Ck�P��K�b1�)�c"Oܰ*æ"c���&/�&|�xl��"O u󀣆U�9Z҈�3""^��"O��+�S�T�2Q�h��of�	��"OVX㉙�rV() W�K�V`�E2q"O2�xY���fG�5/�y�i��yB/���Hq�]68��)���Y�y��ԁ+@���脂6�<���eӫ�y��c��ݠ��� 5)2�8R���y���
\���:��	�5���y���";�����h�,1��EQĂȜ�ybNX>)���f�)�v4*�
��'{��J�
S�riI�L�c�H@L>��W/R��TsD�ck����"Y}�<1A��/Oo����6��A@�<1�E�P�F����9v$��p�G�<� &eA	]´�!�K�`�H-��"O��3��G�K�Ĉ�I,S�Dp�"On�2"B�7A����:/��\��"Oִ�V×1C�"��7�@�x1"Orhch��F��TR��N+1��`e"O�l�BI�WͲTz��=��Թb"O��*���G>��
+��'3�2"O�weUh�,a�*ɅΈD"O�u`˃ er>�8�KT�FT�s"O�p���]�+(juP���[>����"O6M#�e�a�u�#J)3�	�&"O���#�6(?���͜�3Bn�H�"O�eH5��7@�e���B�AQ����"O�I�W��\�j��3�9=�@aV"O0��5��P��A�ԢU�}(�0"O�ty�(N(u�L�2Ca�2xj��!"O"D����v&����B�5{�*�ٵ"O��	�0��Ex�aT�x�z� �"O��	����?�vB��6M�:�	�"O� #R��\ȼeq�$s �`�"O�0{�k�b�����2g��q"O���%*̚�d��bh�<��Ԫ3"O`�s�k�s� ���C�*�A�"Oܜ
� YTm"�P6�"�ԨKp"O�<�@L#U��A᥁V�f Ae"Ox��򌕡ڎMڱFM�'��$X�"O\\�%e�	�40�C�Y�$�t"O��P�NI"	�ݱ�aX(1s �)&"O�\R#���a��l�/��QT,�!#"O���6`Q�h�y�e��w���Ys"O�+6��o�@�e'P;/Ŋ8c�"O�q8�Cc�Z�YQFŹB�&���"O���E�؈X
}k�j�,|�v"O��c��׮~^T�� �(�s�"OU�B΀63�Rp��S�2ٜ�h�"O�-U�5H�[�� 1�H��y&�@�h�т۟����>�y�L�,	� ���*�j;�*��y�M�
��U£��r8�����#�y��>W�.(�@"���`$����y�DC���a ��5/_����%�y������a	�+a�*��"�yҫ�T[h4�� ·0��3�W��yr��B�qc��U:���Vݢ�y��&m��E�$ϖ4�&� ��-�y�F�Zba�"�O!!*�U��j��y�
C�/��9��ӳ
ȕ�S�1�y��@?�� Pp땰w>Խ	 ア�y2�Ν&�Ā��Α~�0)G�M�y��@";��T�3
�%���% �?�y2��&lp�Y�#����Ԍ�y�Y� jN�X��KsdM���	�y¡1f@PE!�k��D�$���y"�'ⵚQ��1f]lY$l��y)���Z`�#\'v������3�y�a��hL*�Ǯ@�h�z�i�	�y�Ɔ-v$t�a����4B4�y��j1��(5I��T���èW��y�䔷O�E�'�Μ_�`YP
�6�yr ��35���dB�Y���TE��yR� �
%��9f\�]E�����N��y�Q�*rԙ� ��G��@�
�1�yR�B�[`�`���е.�m�WF�'�yi�L�4�3��݇$a�8
p,���y
� ��8w	J&<�{�dC #��!��"O�c�e�j=�X��C���P�"Of�3A�R0a�D�$醙�><��"O�	���w�����	�Gz�U�!"O��z�F�� �ʂ���n��"Ot4��-&k�9��㉇S�4a�"OV�B0�2%P�}�AA�,�b��"O��p��)��z�o�28���à"O�+f%2�zJC/X�V�x��"O��1�T�iZ�L0��y96��"O��襀��7�<d�`"��t�3�"O �T"�>�`Yб��+�,L�"O���B��-ގ�YwE(r3H� �"O�dqP�R�kn-���ڌFE��Ӆ"O�9�� �3�	0��OK���"O���eS_�&�����Bz�)%"OX��sVu�NM�$CL��e"OPl��-!cjƼ�A��I?��  "O٣�셷[P�H��̲<>�}R�"O�dk1��#����J�>O� ��g"O��0��L�X��:��@�l��g"O�0a�;#.j1�7��f
��t"OH�d�X&?�~TR��BIJ$R"O0��&��R��ɐw�\�L�l"�"OV��m�jڕ�
�_��K�"O���aC�r�t`8T�Q�M�He�2"O	{�BկT*հ�]�N�~���"O�1�֦��s��b�@�E��DQ"O\�Yt%�8F�"��/a��"O(�µƏaڤ����0D�$*�"OTܛ"k�B�}�"@/W��cq"O����iͭ[Ad��p!'!�E�q"O�ִᷮ�9�K�6Е�"O ����Q9L� �%m\�Q��0��"O�̱���*^�> ��Ɔ)�� "O�}�"ɒ�'���j�L�P����"O&�����t��D��[�j�"O���g̷0��cJ�H`�u�s"O�9j䋎 j�v��W#I�+�^�C�"OƝؕ�ՙ��(���E%�ꭙ"O���˲Z�: 9��5f*HI"�"O<�
�j�	6����
�mkH���"OB�����0��	��튜}O���"O��w�Ar6�8���S0
M4x�4"O�I��Wm�\ѲJ�ve�բ�"O�����
Dh�a��ݨH���:"O�!	��]7m� 8$�� �hH�"O�X�0)��.�,XԄϛ��%C�"O�e{b��x�%���-Z��X��"OD��&��gʖ��g�5F�����"O�(�ʻg~$[Obh�@�"O�,v�V�^{Ա{1A�T��� �"Od!�!�G# &HЂ�ݢa��Pr�"O���f�2z5��� mJ�?�V��'"O�,�s���"�`����W��O;��$&�S�O��)�5�G5`6>��6�ܕ"'2���'.fp��X:p´�Ue
D��'H����B�0�\
��O�3݌a��'�VU[C`JIt*�	95a��q�'�$q���<�4�E�X��a��'�@Ѻ��<8���nP�	��u��'@�ɳ"傩++
�Ȅ�Lw��t�'Z!C�,S�&������4mh�Q��'�YRv�E-�L��bNؔi���"��� &I�b�,Y��I��C��}����"O�`�q$��;�8իV텼Y�ttB�"O
Tra �*��Ĭ�4o�@s"O��a�IS#Kf��5kK����BE"O���[x:��E�&�X�"O����#R'0��s��@�D~\e"�"O$��$˚��@I˰HǕRn��E"O��[�ܬjr�V���us��B�"O"�Qާ2*��ugɸfg�@�"Oؕa�? 4���0&ǆ5 �$"O0=�c�%���!p/���y�"O�m�#F8X��<����;B|�%�f"O����H�|8pCǂ;;۠�8`"O
��D��}+�����N�N���"O��Q�C?L���5�ٔ^�F�!@"O�}�LW�,|%��l��b���Z�"O�a�(��o����p����"OlC�\��I�	��
�����"O�:��P(��lk���- ��H�"O~-�eE5y���7i��`c�<��"O���pE�9b���s҈�@Į6"OL�b�^>$��,�bH�	b�R���"O.-���:]�Pؕ�<-��E�0"O�}#k�O�\p���
 bJ���"O��9�ˍw�x�����[,)A�"Oʁhҏ
�9Z��A��C�y��"O�TSp	�90�Fɹ�a�]�ĉ3A"O~4!!Ĕ;'�V�B#�M�p$�p�u"O|����I�p8���w,SQ"O����ݫN��e�%��_:hr$"O�8���ۈxS (�%Z���"O�`��b���(1Z@XL�� "O$h��'sI;��F!ax0�ʱ�ŭ�y���;~�aJnɅc�9A���y2&�� �.󷄇_�N����>�y��F�'/b����ɱ�\X ��y�垮F��\�%� �'>y[�V'�y�O.��{�J@�d�Y�y� �4X��ҠH�M��9��0�y"���*n��S�>��HjEa\�yRJ�5I
\J ��= ��($
9�y2jРH������ڃ*O64���	�yR�ˀG?��ش�͢�t}�Eꈃ�y�. �:u&X��(�
u�� ��y��˂H�� K@DN	D�&)ѓŗ;�ybM�6~�F<�f��P��Q0��M��y���!(� �1�
F�b)�*�y2��?�J��j�P<ޝ�Ζ��y2�Ӯ[�>��V�_%xq"PG��y��4nRx�!��|��}�Q��y��E�<��w@�!�|]��AK�yª�;h�˵��c�b%)v�O��yr�FJ���s�̃]���#F��?�y2�?O��mP���.U�(����yR"��+P"�GG���!Eǎ�y� �e�|�5�Ufp��N��y�,�]�Fx��$�OӚ$����y"K�C�����#D;j3����y�G7P�խ:	����꒬�y"Ɇ�]".u�F͟v�P%pD���y���.����Q�&�d�����y�b�=*��r�i�u{2�5h[&�y��HLXr�Z5Q*8��'I��y"E�M���I���+2o�Y'C�y
� 
�� �Y$99*�G]*k��e"O��9�c�&��c�Z4`EU3�"O����k^���s��OA0�R�"O�f)�"`&}���'3.I��"O��pb�Lj�ld ���t��6"O��j�ED=<݊�e��y�i"O*}J2��7?v����
�!h$i "O�Y���5��ݛP��j|"؂�"O�x����kV��yBƘ6<� yr�"O`H�'([�us� ��̓/_���"Of$��ۻ=���`�[
{VvK1"O�%�5�K5����/Z�T0�"O���#��N6�<�aИ��d"�"O>`�E`J�k�H�@@ޫl���"O	G��{�.��m�aM�E"O�0YS�ΧY¾{1��)��1�"O���Ҫ%v6u�+Ƭ7�Ji�"O�h1r�߁s��A[�J�/T�JU@""Oک�Se�qx�5JX*�~��"O�}��j�?T� l��)^��L �"O��aсŏFW��ǩN)%���a�"OX���FP1MMάJuH��9^���"O61�tb\�h̑K �;�X�"Oy��!+t�ƹr���)j&l��0"O�31��$D̶Իw�$.&���"OF�9��P	wb��� �v�$�Y�"O�Y8�I�u�Ԋ怨[�X,��"OR�[bx��Ud�i3��U�<yd&A�a��!�ԩ�N l+�/�U�<)wA��h��țj�	c7(�	s�y�<��e_,',�����Syb�1lK}�<1u
Ҍu���*p�o���EN�<��d�,��m��+Q��XL�e�QU�<QP��-4$.�S�͉Td�}Y̅N�<IA��%`e��	�kԂS�,�a3!o�<Ɂ��17 =���B56O�9�/R�<AVD�ef���'3t�X����M�<a�+�>����)��x�<�
���E�<�0�B�=U��&��%���g��C�<��Ð�6P!
B�<C����.�}�<�cƜ0z��=K�Dk1���l�z�<��
S?�Z�nY�h�����]�<�5�t����K9l̨�B
]�<�Pm�
P������GNn,���Os�<�F�ױF�T�K��� <%�Bg�<�Sa��#���;AܑK�A�&ky�<a���.H�A�Шғp$�)��Sr�<����7�����J�XHᅄ�p�<��OZ"��1�ף�q>1U.B�<YR�	:@>�T1r-��*��1₪�{�<���AcY�PG��Ԙ��i�]�<��E8co����ȓ:4n��c\�<ysM)h�q�P��R�zxq��o�<�Tꑹq��u����|��G�h�<��D�*n6C�e�%B&�)���j�<Yg*��1?bXp�ߞ6�8��Pf�<�e���N�Ό��Ulr��j�$FN�<Yr*[�;��ℭ�a��=��DD�<�t�ͩB.��fFS��0���PB�<�Rn�=Rt�ՂaI�3Ex��)dmA|�<A�G�%����MU	*v�E��Tt�<AćP8yÔq�"(�q�d�{��V�<e�߼HX�ɠ��?�8ñ�S�<9�I��M�8@Be�Q']����W�<� ����@������^|�!��"OX��R-�\�e���.w�P��"OL�1�+���Bb��s�0�$u�<���j���&�Z�REs�<��![d;�����#M��Pjeǂq�<�QH��W�	� �Y�*��$�S�\B�<�щ9n�͓�ϋ=�D��%�R�<a��S%;�2M���Z�r@XQ�<��gR8�v���Ɠ����g�e�<iq���X�T) �e��Q�͑^�<�s�� ~����#C�d]qv
�v�<p$T*x�>�aC��"< �F�j�<qC��+MWf��$��[�r�����d�<!�B��	(@8b`%��XB	�b�<y!+@AXHs��)Gg�p�fPb�<�]�T�z�g�:x������C*�B��u�.�#gBЋ<����W��B�ɷq͘`0��7ǚ�3҆ʼF�B�	�Nx����%eD����Ԑ]m�B�	'K
�5R�b��-,��y�n��M��B�I�m�ڤ���Ι�,��M)QIVC�I�d�(=���[!t�)IS���C�	��D��i�G[lBR�52]�C�	,Li�����X�h���="6�C�IZp��sL<'���j7�Ө"�C�ɵؒ�k�R5ifȑ@S@�P�~C䉣r�����}��y�g��!H�bC䉊0Ga� c��jfK�OkC�	;0�J�ZW�Mb����ttC�	w�8���EV�e����0I)��B�	h#�1fD�'M�x��$�k�B�I�#el1S���kq��k�W>3 �C䉐_�v�;��ˇd@K�?P�B䉆@��4���YTΕ��Kl�C�	�.�Кn�~J�D����<˰C�	�9C����΁|� Arف��B�_C�Q��.��\l�H��/�.��B�I��=Q J6j�Sê�lZ�B��!FyhЉV/���PD�#��4m�bB�!A��)�ի��*���A�`����'�,hH���\��`��� �`��
�'ojx�"�և�d�ʰ �qG�@i�'�Ҡ���׬!�^-P'Uk���	�'-Bd@�o��T0��率MR^(��'nH,�U	-gZ�X)ˢ���'�@X�ds��Y��CŒ�c�'β�A�TY�8���+��6�y�i�a"�]ہ,�+�Er��J��yRB���pR&
Ĭ �t� �a��y2C2������ל�D����>�y��V"�z5c�d���c��T��y�A�
"L ��M9H�Ś%+��yR�(nD���n��Ĭ>�y��[P�3�!�?X��2�̚�y�N�F������h�b���aJ��y&��=��T�eдr�*!P(�(�y�ѻt�$z�cЅdL���$*���y����\j�3���^M:��.L��y�Ó<)�Q"�ƎZy�D�¤F?�y���;[�Bb��W* ��Z(�y�,�`�t���ĺJ��ܹ%ɫ�yR��s���u�LHe&�5�y�J�=4|����B�:m.4�=�y��*ŉ_�^��iq#�2�y
� N���#W�&�Z�l��OA��RR"O�]#po�Ex�I'�T�I7��;"O�-��'r8kr�W5����"O�M!��Ҹ~�jr։�v�^��"O
h	����4Dpq:��=yv���"OX(3���,�J]r/Z%L]z�Q "O&81V<Q'r�Fo�>[8b�:�"OZ�9E��n=�={f���8��"O.�
0h�I:�������X�"OH�Q��$@H�|!rg]�i��!9�"OD�J%Z ��q���Xm��W"Of�s1�޲DrM�-�?<�-�"O`� �G�;90�AON 8@�8�3"O<���^9j�۲ ޽@<:y""O�h�C��U2ܜ��٨q�Ȭ��"O�`��74.x���]8�`�"OzMdC
GZ���d�ۥZ��
@"Of�q!	��0�<[�ޖ1�dز"Ol����բip��8�ʴ�%"O�����9v�2qa1�8w$���"O�!ٕ���~�NPs';i:�"O������w��L(Sl�Og
�B"O(c��"�f 1p��:_�hʵ"O*�0#"X6-N$��U�C]�hB�"O$R���qPQQ�eD`���!�"O�����|�t�	VƋ�w��A
�"O��QD��A�rYP�ϙ?v��"OZR��E1@����Z��v��"Oؤ"Q�D��� ��I3c���"O��q�,�!
b�� ��$���"Ofl�S`��p��C�я;��I3�"O摺M�<e�@"C�8T�pJB*O����䖲����ƅق <���'���΄����P����ui�'8X��G�J^�m�Wf�D����'���apC�&Ode�t�D6"O���O� Y��`3Ah, 3i �"O�� �ӝDn0𩓾B^XБ"O6m��� d��U/N	-f���%"O�@rn�=+`��P$<6T�z�"O���ED+3PP�҅�`"���"O`�d��6_&� Ӳ�/@��"O�����^�w���#hQ5t��}��"Od8�թD1eJ�9��8m�Xe
�"O��� ��5��!�T�ӀT�U"O0H�s�L��rB*.F�vr�"O�-���ܽAmDU�Ԩ�0z�I��"Oadj��)gS*&x��"O��s��:kv�s���zT��v"O���b�[�@ h�Ď�UB�pV"OB!�����&%��yr��)pj�	�"O����
E>e�"m�AE%s^���"O��bFL�?����.�
]-�ı�"O0E[vbӉ|�P����ѹ,7~�C"OZ9U�+=�d���T��p�ȓ?�]1R�Ю|�`��'�/)`�Ԅȓj�"�9��"	�Hx"��F�n�l0��3_��i�/N_�bYR Pyޑ�����2&��@5t��$��sD����;��x�Ee��Ab�TbIHH��K�ڱE]�9�9�-ԨJ�q��w���B��܏M�| �L�D�� �HK!Ƅc�D�#�����*K���`'V������ĎІ�S�? � �t�bLx��S:��a"O�m�`aVA�}86�M1�ܪ2"O����!`���@���"m0����"OX��Pg/KY�eA�)U{&��"Od-�%ܰ|��i��,r�ȴ�I�J�KV)e���	�9���@�G�# E3��RU1qO����9/!~M17�k�(c�=Z(4��P�k>��
<k�8��CE옔@"�-e��y�,S�"��燏�")���#A�i0pM�0��|�:h�b@��J�5'Z�6=4�PL>'Z�Y�4^y��'��	�� �Ss�-
��D	~d��0��iL�O,F���A�Xبӭ�9`��aR��Cp�󉶩M�R�i��GXx�>�{���\ ��kG#�<�~���$��� �'��i>�C�4�ē< �d�6@Q�E40+����C*���@�]j̕�O���Ɋ��ݓIX��}Z����{��EUcp�q��VS�`YA!�b��-���A�#hfY���Ѵ(Dё��4�r�dU6�����ЛNI��-d�&�ɦr�A�O9l���M��و��㒪]$�ujVI�&]��;1�^�~��'���'~n�1g�8��(SU%�!ĞM؈���[۴����]w�����2$�D8��\�l*����<a��Q(va�v�'4���ďyDdP�b,��"����_�N;,�W��:��\Y fŐ~6��O��O\P2e�X�Q^�����׏��܈Eh	%C�J��
>_,��q/
���i���|�wH&���K������)7`yceN����M��LB�����?Y�ʹ~�'"2�'����	�L�,R�⋇L���S�E6�yB�����˵�>�0�t�Y�>nڿ�MSO>�'��,OL��t�z�q�K�30���4*��xh���G�OF�D�Ob��� z��$�O���H6x��.$���7�V�b��A�(����"�E�I��ʂ��)9�����I�/�X%�A�A�}����G���kP0aKX�S�(�1�(Op���K:'�lCƍ�%&��E'�K���O6�=���튘)2@=���@!8��a+�4�?Q+OJAm~��BP��%�����\�}|�<p�՚2!�=F�{���6o���*]�N�D��]�۴���֜X�"@o՟�'>-q�D'R���	��P�/��ğ��S��;�
���6����ǮȠ(�X,x'��Fg�G���1� � �� )*ҧ ����0�ʻ�M3�n�-:oJI/XI�b�^1tbX�jB�ڥB"��B���&��J��O��n��M�����)�+!R�ݪq��Ghʙ�C�ڞ)�b=۴��'��"}�ISO:`p�GO���d��@O: ������Φ19ܴ�M�G®b�a"�픒j&Qb�b�g?y��гc����'`rT>��6kC؟d��ǦͲӈҎ~�$4��SF?�5��nҬ3��Uє��x]�7%W�b����N��D���������'�5�a�T�Ia�Z�rj�%���L��Ms� 	(�W���4�\<8�!��I�����{0J�|�1/����E�#G e���(I�n�m�61t|���OvynZ럤�����6HA�N��<�cs�18��
��~��'�ў0�>Ѳ>d�1BI5z��@0��s�'IN6-Ҧ�	��M+�-�i�Zw�*C�^5y�X��%iB5[q-3��5lO$LZ& �  ��     {  �  3  W+  d7  WC  KO  [  �g  �r  6~  ��  Q�  ��  b�  �  h�  ¸  �  I�  ��  ��  7�  ��  ��  g�  �  ��   �  C � � � s m' �6 �D L �Z fi �p  w d} 2�  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^r�Bэ]lr"����Υc���!� �u�e|���ȓ_�}�㧟���\a�R�i��p��>�
H�?Дk ��t�Tلȓ*��5�&5y�d q%G�=QG>ĄȓGq�E@ÀVV�p`!��[�H�h���s�`HqH�Y�T}���ńi��=	�G$D��@1ib���eG�6�,�r�o�0��I�&��p�W� =O�AH�� ,P����D֪���8"s���G
�oºap� *}�C�IYW@	Pd]b��10#_� ��C�)� R"0)R�o"\�"e���v�X��"O��� ��)" u�g��w01��D|���On"�q�Z"f����m�,v�M��'�n9Z�HVYڢШw��)�8���'EИ�Ei�
G��Q�L��Z���'}�ݹ��f�i�6�F(]枅�ݴ�PxBjTWNX�Q꒘L�L�yV���=9���P}r�'[:��ƌ&)�D��h�X�� �'#I&�;#*��iYd�&ъ��Mh�OaV�������W���hc�!
�'�0��L�Hz1G��o2&R,Od�=E���N�T|v�8��?q����bI,�y� �+v�.m֦dVA���8�y�k\�0)��Jf�^�4��2���y��M��dX����Ua�uz��y��]�h=&O^ӎ	�n�/��O:�	�M1�8i"��OE,��*= ���F�B�@R��qfz؃���l�<}��A���}V�̵C��E1R��>Pe8�˱�f�<$�ץ:�f�f,R<�-�5�c�<GnX�w0&�CP��|�%C7-�\�<�lH�E�>��ߴ5nݺRi�_�<���<t����6(bf�2Ԭ�u�<b@A�'cp�*ŉ5IY	S�JRp�<af*V�o0�|�����m� �2G#\m�<�W�%�je����+\�ޑ��+��<Q ��g5�$�����|��G�Nx�<�3�Z����w'��/�(qˠ��}�<�6�F3n䬴����z��+�n�c�<���V�{^��uIPn�6I���^�<!��T�bh���Тs���"[�<q��>w�I�e�l{mH@@V�<����B�f��qT`��GP�<q"��:C,bT�! GI��b�MI�<)��U*5� �PB���'���A� MG�<��DF> U���K ^E�$j�DF�<��G��8@�M����r�~�e��m�<9 +��e� ��1 d�8F]d�<�@�ȸT`�8y�FB1�8D����[�<A�\�[��(���qD=�6/�_�<y���g,h�ʘ�峲��q�<���S}��h�BZ�\�ಁEy�<�e)ϢW����"�L�k ��eMr�<i��G����� &_����l�Y�<Aa�ڱQhI����$$t����I]�<"*̈�PBp�4]VTaUY�<� a@�~-D@�c@� �}"R�_z�<Y��נ9�Ւ�#W�|^� 6NKz�<A���$4�R!�Ҍ��a�\�<�#d >m�V��(�#�Hl�<�H\33��A;��؆���i�<i�i�1=���sJ��9����e�z�<y��|vH�i�d��P�P7	N�<��a
�`��fkB
2F�ԐW��L�<�ѦR��D�}�Nl(���B�<�E�̒zr�ዀ��(p� �M{�<��IJ��� ��o�o1�Y���p�<�#�!� ����6�9x5�m�<��l��f��/@&T|�lm�<�!�nŨ]:�)����ɤ�o�<��͹A|������>�(C`�`�<���=5~V<��)	|�)����W�<����='����C�]�������m�<q��@���v�Z<� gU�<� eI�j�x�\���X�~c����"O���a���I�ŲSK�W)L�`�"O�Q��P*.�	qT�F=��"O\	a�M�=BT����F��ؽ�"Ol��c.����2���M�N��"O� �d��Rr�LQ�ٮz�#�"O2��f ����ʣ	�1��"O��+F�(%��q��,P�(��y�"OL-J��Z�	��B�	X#�����"O<��uAf|�jG�T{
�k"O�i�!ќt���$2e��"O&�)U�+��x�A��:RΜ
�"O.��P�N�^L8��f��={w"O~D"�lإj>
̃$ȡ��Z"O�\#�� ,8&j`ò�*�L�!"O�Q@��x���qNש.͊x��"O�����t�~���M��z�Ȕ�"O޼�K��)��ae셺ib�qV"O��	D"Rd��ݛPk�2B����"O�����.`��9YqD�"E�0p�"Oa�bK;l��C�3^�^�[q"O��Z�E�:C��4��16��k�"O0Y��g�����f��7�l�4"Or�*T��O&�p`R�R��!��"O����UCeD��ѾK��Ȅ"OJy���Ԇ�4�8@ ��Z�<�g,�J��CsB?����Ϝp�<�7�FG)8�z���T����d�<��/ӿnjf	b$�/A�P�q�Bc�<aR�6:�V-��O*|�ѫä�v�<��a��H�tR#�Ǣ��!� �o�<��i	'0=�A
6c�����Bm�<YVC>T2��I3y���A6��T�<s�(!�ܛv�«xC�HL�Q�<9�B��69j��Βx2EAU��b�<��Ζ�C�dd�s�	��Ԁ��
e�<iT��Q��s�
!��!�(�b�<A%�E� ��<��G�p�$)E�`�<�aZ���c���'x�q6D�v�<!��:O�� ���MC��]a�gNl�<�Ï�,����[�17ɕB�<�e��-d���X$iB��X���|�<Yg��PW�����?}��(0!B�z�<	p�M�Y�v�C&#
�&����@�X[�<�4�6�<�����%eZ �6`T�<A1�o`MCa憖=h�-��IDM�<A���-AD��֬
xv�9�g�^�<�Q��v�h'�)Ԕ�v��V�<Q�e�H�~�耇B0\vQS�Z�<Q�^#
d�}Rff	�S�X���R�<Y�Nɟ+��$�6�A=} �yCP�y�<Q1倫,{��R��84�t��S`�r�<qUf�Y;�9���.d	�ˉn�<!�K�2.jZ	S��,=�ƽ��!�N�<�#.*G�`�'�֣mފ!�b�G�<钦M�#����F�#�&ؒ%LHF�<��,Pf:��(���E�nEL�<A�N�"w;%E��6��eh�^S�<���/C?�u��חJ�X���L�<�%
'H`lK�O�&����g�)T��c��)}�2E2�[5����C�5D�h3�1ĥPD����e�5D��:���=x(@���dB	z+�����2D�\kr�:Ǥ��a!��^�L�z��%D�� �e#P������+��[�]92�z�"OVaG�Q6m�q�?����"OBd�w��;2Tt�#k�6���"O<I[��˂c���[��ݍ�����"O� ����	��KF�
�͈����'��'9��'��'�B�'��'�0�
4��	(�T�'+��h�>��u�'[��' �'���'���'���'FY���P�?�pe"a �"M� ����'s��'��'X�'��'�"�'�<�Jvm��v|���"�m�<�s��'���'}��'m��'`��'��'�\-��7�81C LF/~L���'���'���'{2�'���'%b�'����$�BE���.zǐ�$۟��I�����ϟ�����T�������ٟ�`q�T+.Tc�7$��r'W��(��ޟd�I����ß��	ş�������(�5l�X��Eˀ6�>�x́�� ���`��ȟt�I� �Iş��	���R�MB"U)��K�`��&\Y�A�ٟ��	�H�I�<����l�I��������wKJ>�8�E$��[4,c��A��4�	� ���X�	ȟ�����@�����@&��4m;aÝ/E��CW�������0�	����I����IПl���������bz�܋EK�8��d�	ǟ���⟼�	��\�IΟ���\c7�+&tt]S��j����� �L��������<��������M����?��b0sԅ(0 ��x 6h@lO�{.�������������:Ձɒcj�P�]�dS��U'EN��N�6�4���O<
�-\RU���"��T����O����Ŵi_���|���O�c�vQj����c�Ęro���<i���1�' P�$p ԅ=����WFOT���i̳֚�y�)ʦ�+BFt��7�Up�q�a�X?\��	ȟ�͓���,}�X6�u����Ə"~w�m`��f�B�+�g�Γ7)}�����'��)�ѪQ�[��S���	��'��	E�	#�M���\̓(�p�$�ǒ<����M؅��쁊�m�>����?��'��I�F�`x��kE2�R	B�Ì����?i��� Nr	�|j���Op	#��W��)�N�(���ᄏ n��s-O2ʓ�?E��'�ФI�ND�1U:ђb��)�䥁�'�v6��sS��2�M[��O:�K4�4���)"���u�d�`�'S"�'���Z�a	�����ΧX$�D/Q2���s$�;C��°� �
!'������'�2�'S��'^fy�E��* �9��M1��B�Q� ��4P0�)�ȝ�?����)�O8�$�!=Ҷ �d�qK����&yԶ`�'26��e��4-��O6��O�JD�CT�f�%�̝�qv����R-,p�!��'��-��gWM���B��H��O�l",O��C���+���*$��c�����O����O����O�)�<Ӷi�:Qӑ�'���ɢ	�,�P��	�$\И'��6�9��8���尿�شZ����`����$C-h��c5	� ��ⅹi��䈼x��!�S@ן��e#`���0��))�ΰ� CB `1�}�UgJ����Ox�$�O��D�O���*�z^�1���Q`����!����I��8�I��M���|��q����|Ro)rI##!L~HL'V�{�O��l��M�����!۴�y�'��1Bp�%�`Ȗ��t��Gd	l@`l���l��'D�	����	ޟh�	�d����.�'T<x���k�q������'V6�X�
����O���|�c�M�nmā�f�z��y:5e�o~rϺ>9c�i��7�۟\'>���-�Ⰰ�D�&<ln��~�H�ۂkθF���#��ry�O��	��'� �+tl<,I� ��F�t.8DHS�'���'����O^�I��M;��A�Y��ň�a�6`�B�QM]�'�0���?i׾i'�O�5�'�F6��6�`xb
�3S���T$F=jn:�mZ��MÆ�۳�M3�''�e�RK����"p�	�r�qI�Nʸ%by[2�E�(��IWy��'t��'xR�'�rQ>{筂.��p�w���В I�(F9�Ms��?9��?!����0���w��TI��A^���Q5|�䉡��O6M�]��\����h�Q�h�d�ɬ-�$��B#*|�Q3�}N\�ɺZ	 ��2�'n�$���'9R�'�&�h�
�4 ���ub�]S�@�@�'�b�'Q��K�4o�x���?A�3Y�%"v*��PXqd�+v=`�rê>!@�i�7MQa�	�m��sDk���0@��c]��I��x�+N�t#*I96$^fyb�O�ر�I�x�Ҫ]2 4H���B�D���k� �3v�2�'
��'-���HZ���� �V�:�ئm���A�4|b������?���ix�O�N�/���z`
��8�=���(?m�dt��o�6�M+@���M3�'�R��$^L����B���$���G�$��%d�>J� ���|2T�����,��ٟ����dyA"I�'
Qc��2r�d9b�GyB�~�ne�Qf�O<�$�O��?q��hں��@�H�-c���"M=��%�f%{ӞX%��S�?u�S�rJ]��î9���`Iϋ@z�M ���@�<�''I!#�͟d�|S�,�!O� 0}����GpE��A۟l�IƟ���˟�iy"df�Θ� �O�Ha� 0�����>�^i4��O�0m�S�>l�	7�M{7�iJ�6��'v��2�J��#��{�(BO#�%�scl�V��ן�Hc+�� @���Zy��O<� �0�F�{��d�VM/Bs �s;O��D�OH�d�O���O��?��͒~������Y�iѺ4p"j�����ٟR޴F��i�'�?Yb�i��'��@�2�ˉ�4��5)Z�K�n,��Ѧ�sٴ��w����M�'�>-
��J5@Z�)��)��&��Hȁ��\� �|�R�L�	�H����l��%}�X,YG�ӜV*)�U�����Cy��t�`�x��O���O��'j��q0��$2�5 �ӊ+1r!�'i$�5�F�tӄ<&����?i����qڐ�C8�R:s�*KD�p��<�6��'���ʟ���'��	�l� x	�I~f��p��0`f}��ß��IΟ�i>y�iV�����'0�7-U�*���u�
%�p�4kք+p<��ɰ<�ֽi��S�d����$��8��9�E�b�J�`���M3�i�� �ƴi���9��ḱ�OT�H_Ll�p�3I�����NF�Mk��̓���O~��Or�d�O��D�|*ӀĂm�h]$,H�8׀��3β"����2��	ߟ���v��'Q�6=�N��t���K��Q��+G�\ Pg��m��<y-O�O�:���iE�B$lT��ph�&�HuF�#T��D�j��;��@gF�O��|��x=��+�J�E����%Ѿz�Lq��?݊�������%b��gy��'���{Ѭ�Q��!�Gpp>!i��$�o}�}��Uo��<�O� �()-�R9�f�ՓӺ=j$���r��*7n�exT*0�&5d�(�����)E�1֌8ae��M�����O���Iٟ�I՟,&?�*�ၧ1���imB�]/|��yy�FJ�v|J$Z��'��7�E�/.�ʓ�?	O>��Ӽ���K'����	Myk(D�<�F�inF7�Z���ʢ`
��9��?�T�7�b�	H�6�\�U+ԎJ�@3�D�O���0I>Y+O��O���O ��O��#��?(�����/V;[HPu��l�<Qs�i�,!K��'�B�'I�O����:v�H��ID�m�@P��][J�-!�V�m�.�i��?E�	�W;~*S��"yGb�{���b
.�
 �S�2~�gŌY�T �Oj�ZL>�,Of��pD� $"ޗdk����O���O��D�O�	�<�g�i�r]��'�T�z�CE�;D���-� ����'6��O��Oj��'R�i�R7�|�pa#�NƐ���>����a�����ɟtzBeX���$GNyR�O'�� �y߬Yi� 7`!J
��y��'$�'���'����;6�"��Ō6���#��L����?9�iFk�}>9�I��M3�����A� ����ѱ�@pV�"d�$� �ܴ���O|䓣�if�Ɂ54�〭��".4�2 ��s�@�sPn_��CCz�	qy��'�R�'�LW0=�@x��G��U#��A�R�'��I�M�E�ў�?q��?�)�,�4�[.�n5��"�"c�<�䙟Xj-O��DtӶy%��)��N=��h�;��Xȕ��b�X�J����t@!pK��S
���.ri�=��C��?ɥ�$}Zc��Z���	J �"ɺ�l��+�r�'�"�'���4\��+�45ߎX����Ϡ�K&
n�\&��?��B@�f��X}"�l��4�G�xЊ��m%+C��5�D¦�ش�E��4�y"�'$d�f.��?!rZ��ac�=jC�
���)_;j�0e�ܗ'���'Q��'���'A�0f#��J���>����"=^���4�������?!����'�?I���y'l�Y�Ɓ9���|�x�g�^��6������L<�'���'4�V�zش�y����V�,� 7��'z4�'Ϥ�y�ςq1T,�ɴx�'0�������Ɣ놡��iv@I��ɞ�b�����L��ޟܔ'ψ7mE���d�Ov�_�����ȨM�>�#��I���㟼ɫO��l�1�M� �x���2 �z�c1�F$;��1ul���y"�'?l䢳@�@�Q��_����Cl�LV�L�"k�c̉�šM"�&�1���`�Iܟ$��ԟ\D��w]
y3���1 
Q ]�V���r�'G:6��<��	��<)ݴ���?ͻzLV]���;nE.eq����,Y>L����hӼ,n	��5m�<�������%�j]�k�ؾ���+2���@��������O����O���O��dR�2�R�Q�Pʨ�1�C�(mp�ʓV��CFR�'�����'D�iVʂ5[v���u�P�D��b��>�$�iw7���'>I��?	9BA��W��:�"ED�B��8#��y��@xyrU'φ��ɡ��'��'JJ^	�ʞ0cB�"��=4T)��ԟ�������i>Y�'ʺ7�̹_�:�dH�'	af ?q�d�!B��Z��dRئ	$��I���D�ئ�[�4!
�� mC4�X�gE
Q��c$�ΐ\ְ�і�ih���O�ى�+���z�Φ<��'���gȁ~���P6�ڠ[߾Rs��<���?���?����?L~��'^2�����I
�2�
��u���$�����?���M���$����'oҙ|���{aX�O�=��U�+L�l6Lk}R�x�ڕm��?��[����?)u�G=a2���R��hy��gM�Q��AB��O���N>Q/O�I�O��D�OR�;6 $q쎓a �t���O��$�<AB�i��S'�'�r�'j���OS��'Mz`fG� 5�L��'R┟P���u�޴'��O~��c�;&��X1b*� Gx�@��"ar*��uj�O�iQ=
��]��?�/O8}0�A�-�0n�_!Mqꠃ�O����O���O؀��͑R����O�������U���T�Bb�<��,� �0 ���	ܟ��'y��'��6ƌJ�6��릕���}�>A"��p�Y�@���M�i5b�%�i��؟�<��)�:���O��� �a蒍M�7�!���,@"b���iU���'�r�'���'���'v�S�@lh5�eg� N��'dA'%����ܴ
�����?i���j�'�?1���?�;�\�+ă?/����Oҿ8b���c�ie�6-J��m�O���<���e�@6��l���,}�<�� ͑"����C�k�Dʲ`��H��Yy�O�R�P%��ȩs�T�%)��B�d��\���'t��'�I��Mc�a����D�O����_�I�b9c�h�2D
fx)դ*�����C��EQ޴ȉ'��Hz���i�>-��H�e:Թ�'��Өo����������?����'uh��	�S*��&Ȇn���B�c�8���ş���ҟ���m�O�Bj.л�
,���{a变���c��3���O������9�?�;�u���D�<L�5�I�9<������b�N�lZ/� Tn�W~�
��P*D�Ӷn[�)i6�3�^,i�S����@��|V�h����H�	П���Ο|2�Om[���s�=v���D�Rvy��m�|áe�O��$�Oؓ�����e���9���%��P�eU�|^!�'�,6�Ħ��K<�|�愊�MRv�FD�J� ���6/���I!� ����_���B�����O��6��a�tDM�y��]�� �U���y��?����?Y��|�-O�!o�����	�hn���!Bl����Rn�R��I��Mۊ#�>� �i��7������Ӡ[{�"갩V��V���X���%o�D~2L-b�����H��O�'���x��V!Ū���Aʁ�y��'(��'<2�'=���Cd:聁	�?g�v��U��8�$�O������6dw>�I��M�L>�R�ҽX��-���[�,$
�ұ(��'� 7- ��'w%�l�~ҥ�z�āc�G!1H� P"ҕZ����L�ߟl�|�\�<��ܟ��I����ŭ^�`c�&�� ��[���ԟ���{y�Mnӌ�"�b�O��D�O��'?1 BэC��<ɀ#ܾ!l�'� �1��f�Vx'���?��B� |oNu����l��yǩ�,�(@g�	�|�'��L�A���ݟ�'aԽ�f��.y9I�K,MJ��'Q��'R�'�*@ �O��ĲaR��_w�\X��-�s�V���/�)"�����z?C��	v���K>ͧw��7O7mى_0���eX�ú�r4�G�/�l��M��ƿ�M��'�F .��������S)b@��@D\^�Xs��ѐ��D�<i���?Y��?����?�-���b�Ł J1l(SB%�I��9���	�y�����V�	����~k�Y�	��h�i�E���O�e}���"�><�ll�aS�M�ii�6m_^}���N ��1O*�:b��
7�����`�,�b�9O.���-K"�?�F�2�d�<�'�?I��
�<s�)q�|�Ĭy�ă#�?q�i�-{��%��čڦ	��F�?�������1B�Xͫ��C�)��4"���o�	��P�'�L6mB����ڴJ��%��+���(x�xKr#�?a$�ZQta�ա6~�D�|*���O�D��B*9�����k�D�z�N���?��?I���h�~��oE�a�L�+T����GF�\lh�dڦ-�`N\۟��I&�M���ӼsM�S%�ӓ�3�@}1�'��<1�i�Z6-��!A�e�Φ���?�
Q�2|���̋G�t$SAO�@�ީp�MS;W��yN>i(O����O��$�O��D�O��aH�=#�Դ� �,[ضd��I�<QB�i�!˖�'b�'h�Ob�I<5/��a�b�%|:�e"�ΤH���4כ�Gx�p�	[�S�?��	�az搨D��&s0��g	\��/�?j�Ĩ$?	w�*g���T	����D��+�(�s�nU4���@3*�1�\�d�O��D�O$�4���	#�&cOExb�5��\�r@��^�R�!Q�҃7��n�����OR�nZ1�M��E�vA����R�����
{<��6�Ư�Mۘ'��d�������/������1}��d�D2P� hg"r�xA̓�?���?����?Q����O[�hpiT4H�(��'��"���:��'���'~�6mϥc��i�O��l�\�ڶZ�oG�>3�U��l
�\1�����Ħ%R�4�?�3g���M�'�"ă-�&�$��� b��iH�$P�.D��mo�'��i>����	�T7L�H���g�\���G�Q6��	ğ(�'At7��$�$���OT��|
�,�8[E�Iy'�&'@���d~�L�>���i�7v�D$>���+?ix����"
x��ڵT,��S�W�>0 B�0?��',8����!��r�d�1��1xܹb��y�a���?q���?Y�Ş����ڦ�PCQ�5V�)RHάG���dI�2K=���xz�4��'��Xa��k�n��=�'C�[�&e �W1P
�7-�OP\�A�y��IΟ`37����K ?)Î�+Fp���ìif	�,��<	(O��$�Ol���OJ���O��'J����j��вC��H��e�e�ie�8�`�'r��'��Osk~���@�o���)ł�j��Q�O$+��plZ�Mӟ'@�i>��韄G�ǦE̓�Ƚp���x�⥓���'2�Nu�
��	�l�O>}*K>.O�	�O��'cд&���lUl7�Y��L�O\���O��<q��ix�RF�'���'���0R*@�uw��@����Z�%��c��~��I�M��i���>1!��V�@�� y��҃�X�<��[�UP�"%(�9�'������sr�'C�*��<�Ь`�P�=�S��'��'��'�>���X�q� FW9d�aÑ���L�����MkCE�3�?I��)���4�nU��<�,��$i��Uh�l��9O@�o�3�M{���Ν�޴�yb�'���I���?QP� L��af��d9dā�,;���$�$�<ͧ�?i���?9��?��B�>J�`lZ�.�9�Q)���d���͂4��̟��	�$?����&��M�2�R q*��.�ef�Li�O�8l��M{��x��� �W�!be��*G���*�b�����@����ɩ0������'�^'���'ƀ�3��Y�Y��H$�J�Y&Nh�s�'-��'3r����V�L`ڴc���!�%c�����jh���N�}v�T[��:y����JV}"�g���m��M�E��w.�@���g
�y:�gѹ2T��Sܴ�y��'���*g)��?]� V�x��ߕYK̶�F�ӳ�J/:�
�"�{�h�I쟔�I����	柬���lC^,���WI�8u�Q3�?a��?�e�iɔ`v[�@��4��J�r��t�Ӫ!��q�BN�L߆��ĜxB#|Ӝio�?�ʡ�Qɦ}��?��l�"��x�d�[�X�m9�	I�z����O���O>9+O����O����Oδ9�c^-L �Q�d��̰�	�O��d�<��i�4���'J��'J哇l��R5�!D }G�ֶ]��R�ɞ�M�սi�R�d"�	�,1頭-	u�9�u�� qю� ؎���C�3P���bw��O|*J>���r5H)±��K��#D[0�?��?����?�|�.Oxnh[l�ie�b�0���[$V��RU�۟�I8�M����>a�in�:Ӂ�%Y�10#S�`3zeC&ofӶ�d�$tt7Mh���vܔ�1f�Oa��Ҏ@�'F�[2�q�3�C�������O���O$���O��$�|���OB�lE���P�~a���q�Ѯz�F�2H��	̟L'?��I��Mϻq�|���D�*u��=ೣ)Q����'O��>Op��?�����`Ǧ�̓>J�\�C�ƲiD����"�͓>�)c��O�,�I>y(O���O��['�F���r(r�L-z��O��d�O��ľ<װik�0�_��	�Jp�����U
����%8+�JX�?	fW��ٴv��6O��W. �"ůZ�dg��R�h�X��'��@�@X�&���ʋ����ǟ���'%�|�����}p�+O�kcH8�S�'mB�'�2�'w�>��	�DZ4P�vm6�0�`�>l�ސ�I��MCai���?���$����4�XY� ��'W���~ �u"�0O<mnZ��M���/��Yx۴����ir�' ����ș�:
�{U�]���(�u�:�d�<�'�?)���?����?�JѴ	Š�y �=u��b��5���MŦI@PWy��'K�O@b'*�,�˙�!F�)RĊiWR�̛*dӌT%�b>��D/˕��d Դ4X�e��*��sЀ��ocye�e��e���1��'��Iu:UY׊�O���CuF�ap9��ɟ��I���i>�'�b7�U-u�4�dS�H�|lA���/!�<��C�Z�G�2���ަ��?��U������i�ٴh3� CC�rO(0p���)2�E!��1�M��O^�h4E^����%5�i��(�6I%ha� �ڟA�"��b2Or��O0���O����O�������L0<>n�§���:B�{��XG	�8L�O���Q��Y���ay2�'�rU��Qa-~y���"D�q��Ph�L��M��_�l8ߴh���ONa�4�i��O�(8$�K�4��g�H�](8hڄF�9e^VX1�rV��OR��|
��?���G|h
�e֒7J\���>����/X�?�)Onړ?6���ϟ��	�?y�]/-���8Sb��L>��w��xټ��̟d�'��i<�6K���?e��K�U9|��Q��*�>4ڳc�9ʀ4���@!+>�:�#��u�i�O�U����"�
-�Q"�˅ �^Ȩ���?���?��-c��|
��?QT��.�4-
0�&�2ՅB�\���'<�'���'i�a��Ш?O�mZ�O_���pA�_������q�؅�ܴ�6��R��F����Q[��t�~b&E�	.����E�spXЖ  �<�*O��D�O:���O����O�'^�Us g�5WIw��?����D�i^T��V�X�	l��������#%�3W�2���3	Hx��be_JV���c�@��R}��ċ�*S���:O&�K�aA'C�Ĺb�lՊ7�|��F1OtR���*�?9r�7��<ͧ�?Q���?�4�C��*��X�À?�?a��?q��������� e�ڟ��I؟�9u�X�.* Pr%�>>�t)�f)�X����`��Ozam��M���'��I��Jub���7~�����j"�+oD a4�J2b�8H�M~eb�OH���n��H�ۥ�� �*ѯbn��s���?���?����h��n����M�u.dI��L5l�<��T��	����L�I �MCM>��Ӽ�E���.�~11�GuDr����<��i��6�Ѧ��� æ%��?w������i��GH�!*���$'^�A�	�( N>Y)O����O���O2��O�K�mՅ9�:�G�_�TIi�@�<�!�ip���'�r�'��Q>���wԞm�V��7�nHѯ��h�Yq�On�m��MØ'͑>�	�W�ƠA���xPL�G��dS����n:?�%�uͲ���4������ZX"�� /_�\�0Hk��2,�L�$�On���O��4���7˛��ʴb�B�߼���	eeO�=�z,��Dƻ�yyӾ��1��{}��g�T�lڝ�MC�O�<d����cN0n�豗�R�iƐ*ڴ�yR�'������?U�1[���S��q�J�Us�5�D�U�:���i��v�\�	֟���ϟH��П��`��z�]R��G�T�bQ�W)�?����?a�ih� �O���g�^�O<�QdG <���Y�JG�o��|���q��M�iT�dm��E1��2O����16G� &��@�Z2���H1I�ap,����=�?I�m6��<���?���?��Ȗ�*[V�s��@�<�QA��?	���DAӦţ�c����������O@i��6�@����{$~�I�Ot��'�z6��%zM<�'����]�a���K��L�6�4+��t��!ָ*&d$�.O��i��?��2��\�M� {�뙤K�H	�đ��n���O8���O���<!��iW`��� �Ȝ��a��k� ��KS����'5�6-2�	���d柌 ����M.-Z1�_�b[��(�LȦ�)ߴ$ T!:�4�y��''�%c�*��?)ۂP��A��_�М1��ǥd@J0�t�t�\�'���'$R�'5B�'^�L~(C��>�ē�@!
�	�4M2,8R(O�$+�	�OJ�l���I⡞������E��-=z`NݦUrٴ�yRP�b>�0ק�Ӧ��a�� �jT0gꌀ�N�>*���f��`�2��Ot�K>�*O�i�O>���C?	"*���Bf���4��O���S0V�&�˓i���'T]�D�'ERF��g�nIHd)�)&��P��۠vmY���	M~2�']���o�jt�'��iA�8#j�B����6qp�'�B"�1eXi0h�����埞�R��H����h�r4�g�q��e�P�i���D�O��$�OB��1�I��t��/Q��Nؔ~����d�-/v�p�S(^���sӸE飥�O���N���Iwy��y�D�V���'9t����)�y�lӐel���M+�D��M{�'��cǠP:��SV$��Z�b��w�l}����@�j�W�|�Z������`�I��(L�Va&U�	öJ Mt%�fyRs���(�<!����'�?��E�16�����'��i2����Jͻx���M�r�i}�d/ҧY$��#D_%&%JF咫n8�-�Q:eB���'�p�P���U�|"_� JR��)��TY%),\1h-��P�I���	ן�Sayb*�n�$�')�I(��L>aF&��T�Z�O^橊��'t�6(�I���d�O�7��O�|yE���G�X�0�ǐ.�������1�7�+?AG�
+XJ��4��5��-��I2B�3WP���"W�y"�'`�'x��'�"��
�o���St�ԥJc��d
:>��d�OT�$����c>	�I��M�N>i�ĉ�p��;s��h>��;�I�WJ�X�D�ٴQx���O���i����OJ%� ���G��Pm�18���W��8n�p�)��լ�Ozʓ�?!���?����>h�3**:�N�`KC9AX�����?)O�`mZ#�6���ȟ ��^�4�I�Eyd�g��ˢ�B�q��tyr�'N��'&��O��4�5�H�yg��M�69�1ŀq0R �"[�>��`X���ӌ#���r�	.B0�A:�"! <ԺU�F�|������I��i>A�	�^��9�'�:7m�&4G�X(��U%0:TK�ėvA.H���?�M>q����dG妥��!R,Wx�}Q���L<�1X�k���M���i ���iN�$�On�r��Ψ�ќ�4x&dڌ �����Yx�$肀l�ܔ'W��'Lb�'�b�'H��?��&���*&�Q���wlz�1�4<���p��?1���'�?Q��y׍A7��}@ ɖ�J5�L��睛&}6����I����4�R�)��حHGLӜ�IJ9ʐ)������e���6���	�R�LX0�'8�'�\�'�2�'o�A�sN���狴Mp��2���?����?)�����ڦ�8�mZ��D��ȟ�Rc��4���1IW��#"bl�ed�	��M;0�iON���>���B�j���đ�X#��@����<���NK��D �5���+O*�IW��?����O�-�@�ۈ<�*�a!�;>8�̻f��O����O����O£}�;eu|�����&EjP\�6��6\��8��0�&�C+K���'�6�&�i�Efl�&Htɨ I����ӂ�o� C�4<�֏a�l�� Ab���ԟ�b�mZ:/V��m1k�tԋc-��u�f]/��$&�x�'���'!�' r�'�\$Z� ����ju�\���Z����4OĬ���?a�����?�c,ҶY���H��� Yo� ��?*��I��M�¶i��<�	�j�����Ȁ�hHjNe@5�4{[J����L��5h:�P�W�'�%�\�'�n����i	�U8V��%Q�����'�2�'�����Y�ċ޴��t���]�d��FH�f��2@�s*e���6N�����[}b�`Ӿ�m)�A,h"2�Zp��5@��U��� +�*�l��<���$;d��"D�d�'A���h��[Pǉ�f����!��Eq�$�{����Ɵ�������I����%@&P��Ђ�Y�:%�[BB�5�?��?�³iü�O�xӪ�O�"��\<bs8�@�%.ff@0p�a���'��6-Ŧ��Z�Vhl��<�� ��1h��� `�r.�/~� �iN,*����䓏�4�p�d�Oz���n�|-�1�о#�ْchQ�qx����O�˓ƯvD�$j�r�'��X>�s���>2P�)�`�,W�`��.?�RP���ٴ*j���,�4�l���uoƍq��נe��,��D*�zH�<-��6��<��'E���d���eD>��N�-P��u�C>G�nq{���?!���?a�Ş��d]צB���<!U*�B�{��àׯT~B�'y�7M0�	���I*�i��;����ʯ�j��	��M�F�i,����i���5:���s�O輦�'E6���K�r�i�M�v.Კ'�����I���I�� ��L�4�X#*~H0HL�Q"m�1��)��7�ҔDHH���O���7���O�4oz�]� �Y�jR�.#b����5�Ms@�i���>�|�aǋ��Mۜ�� `Y��Uܸ˶&Cv�p�5Oh��s�Ⱥ�?�2�.�Ĩ<����?ABn 7Z�`Kٲ6�5��D�?i���?������Ц%{eH�ޟ�	ǟ�i�C�D��Dq�ˁ%l7F����	X�%��	�M�׼i��O��qFe�2u@-��A7D���Q�;O��$��hOn����[���S*7�F�������<�0���ִl��Pz1e�����I�(����`D��w�� ����
?d���cXIt�0��'(6��#�~��O]mZJ�Ӽ�a#ߙ;`6�G�0�Le,*���=�M��i=(7���r�|7�|���	J�6d�U�O��ۗ��X|�D�F��C��Ź�'�`�	Sy2���j������D-r�b��� !������dK�v�2�'g���̯V,4����\1��w�|�'^6�	Ҧ	����'������h���j\D��G��3DR�,б`��-�,O��s���?1��:�D�<A�J��'�d#7�M�W�@ ���q�<r�4Z�,[��+�T=0C�]�C(F�ڑl�8d~���'4���E}�iy���m��Mc�Ƅ�z�	r%�1%7h�� $o�~]�ݴ�y2�'�X�����?$^� ���u!��M3w<�*m�eN���mq�p��� ':����l&8��w��L��I������M����C�(��O��Z�ǘ9G����� iy�x��oX�,�'T7M֦I��i�>@o��<9��d���YS�׉\����` 	�B��Ϗ�# b����䓡��+���}Z�K�䟱T�\���P�^Q#<�C�i���c��'�r�'^哲D��X�R��25���8��[�n�@�uJ�I��MSѸiT��d)��T����Z$t��"��w��p�C@�T�vU��� �����!�O<�BI>i'�K���\�4�#y��q!RR<i��i�e�W�Z]���`��;��������z���'^
7M;�ɟ���Ŧ��b�";l\"�@�$i�X&�L�M��i�Z��Ҿi����O �HC���2�F�<AWGN����e��=|^\�OV�<�,O����O��$�OH���OF˧m�X��,_s7z�(�(P%�Q�W�i�hb@^����w�S��*����3��&D���I�/T�� �J�xF��kdӠ�	`}�O�T�'�f�ƺi�󄒍(���:FD�I�zP�F�]0��M�EF���
k��O@��|��
6ٹ�B�7˶Ej�!� Z	q��?���?	)O`�lZ�X� !�'��	=t�ĕ�$�AU��Z�"!	�O��'��7M��M����)G���RF�U'w~X�Rn�+0��O�u��['_ے��0������L�BcV�)�i@�4�TDA𬏩4�6���Hԟ,�Iޟ����E���'x6�Z��^�(���^�
<.ts@�'Ӓ7M�;Ov����O��n�w�Ӽ�+T�X7��`�i@���=8���<� �i�+P�?y�J���M��'������u�S�Z��Jǋ)�d<��'ܲ,���|�^���՟��I��I���o�U���I�t�Jw��GyROlӚ��k�<����'�?�a
�$ at�ᒅɎf��\H$�[�	��	�Mku�i��0�I�����a��ժt0KvĻӁ%��y��M�^4�	=�
h�S�'�h�%�d�'�(�
����w~�LQ�.��C�,���'�R�'����^���4.5ju0��]�d¥�L�2���5E*�����JʛF���z}�'yӔ�l� ��Z@�I��٬��z��øn�r�o��<��Z��t�������'���&c�Ei�j��*Z��'K��Lj����a�|��ǟh�	�4�IΟ���W�O�i ���NM�57� �cA�;����O��l�6d����z޴�?q)O�ͱ#�P�'�bU�7d�8	��x���'��7����]�� =l�<1�dst͙�i	�-�v0Y@�$���i�8!���d�䓠�4�����O���X�'�89Bm�c�yᇯW5]��D�O\ʓN̛��C@����ЖO��X9��δ.����9%�jp��O��'6b6-�ڦ�Γ��'�"�_��hq��+y�(1"�D��]1`����԰[qʵ�'�����4k1�|B���8]ڹ�C�!��i�fe0O��',��'J��$]���41O��;p�~���f�:_$͛Q���?��v���'2�'߬�I0���L'gD���ȓL�V0�1�8Z��6��O*��s*f�~�	㟤q*
!E�D�'?����.�!�@ˋ@�� g	��<�(O ���O����O�$�O�˧!�f�3J7p�����T�>��i+Rm�&�Ѣ���'B�$�O���'H`7=��!p$_4�`�'$=
N�ɐ�ܦe��4ٛ�'�>�'����$�M��4�y�R�x�r���$5�l��oӭ�yb,4qh�Iy��_�̕����'� T��A���p  �|[Hժ��'���'�\ :�W���ش`�Z<��'�?���c�e{���9���⯋=��|)���$�O�w��&vӜ�o����D7a\��Ajg�p�(��Y46����O�1�u�[�v��D������4��&��� �I
3y*�Jf��)Wf% E֟�	��4�	֟�$?���)O���-�	! �:s�	.L1x��&��5n��I'�M�'	F/�?Y��?����4��(���X �A�"���Q�II�6���ɦ	��4Zx��逓Q��0OZ�d^��P��'��p�)�!���*5m���а+�d�<�'�?A��?���?yQ
N8z$![�lY%`�L
Eo����d����������	؟�ӺO�������1T	H�d�|Y+��.�Z����X~�'���j��&>����?2�.� 8cd�B%p*� � &7h�IC6P1I��	 n�*ӆ�'�j]$��'�^ח�	4D@9�M��d��ܘ��[���	ݟ,��4V@�	Dy�zӶd����O(���.��X
4ሂs�m����O�m�ڟ�'��b�>1��ia<7MS����B�^Z(�pcE�<9-�F�')Vn��<Q���$(�r���8��'�$�k��������};dj^9C����0/t������ڟ�	�����Q3(t,��E�5IR�M�,@%p@�Ȑ���?��i��$^�x��4�?�(O�7��)rr�5��6����ڦ���O��n���M�'��9�4�y��'z�X
�h�I���R��(ԥx�ϟ&E����	-E��'��i>!�	����ɹmo�h ��O(HZ|�;�b�!q�28 	ڟ,�'��7�P47N��$�O��d����8CVr�jT�Xj,\Պ��	�d�O������|�h�n7�ħ���H�.B�V���储b���Ad;T���ds	� $?	�'DI��B��MI��RկD�Bv�p�t��+E�K���?���?Y��|R��2�2�C.OvAm��ޅ�>����ܚI�"]�c��[��(�'p�|��'{剿�MV�Q!�r�
P��2���h�*YQ��~�,��js���	������
f���./?1��6}�r�����*V(��Y!@��<�/OZ�D�O��$�O����Oʧf^�{��=&��i�O� �hw�i�Q��'R�'����Ȑl��'��w�lUBQ��$ 2m� ��%&��Iv�J�l��M�A_���?=��kE|n��<�����-k3��*v�M2�N�<i�-S�#����ߤ�䓢�4��l�� �H�?g�N�Aq焴B�����OT��B�k�ʓ[�&��3x����'����%^�a�5E�u,9x#'·SS�Q�`��Jy��~Ӧ9nڅ�M[Q��i���=|�	!f�(`���#?YB�6@5����f�'U=��ߦ�?Y7?s]Сz�
�M�B���I�"�?y��?����?N~�`Ƌ�|B�&7�$����+c�~�e� "@���,��蕯^���'�'��i>�]�Tv�-����q2Zmڦ6�.���M�f�i��7M_6#�T6M,?餍S�5d\�	M8�`8�AI�q��1@JE;2���yI>Q-O��O��d�O����Ot90W���`��7��?`�N%aG�<�4�i��PR�'���'��D��%���'K�dU4u�(Rv,�g�B��Rh�>�3�i��7�Ȧ�J|B���"�IJ WV^�8��ɤ	���C�ͳ���R`%Vi~b���f"ȱ�ɫR�'#��!90�1����$Qz�YE낶s�\���՟��ӟ��i>��'nd7�M�
�� �\�B0�\6& s!��
�馑�	x�I���Ȧ��4 O�f$�<���%,��X��(@B��&t2�(��i0��O�H�����3k�<Q����Å�R/.s5&�4����<)���?���?��?����oЂsƅS6�� <*p�c�R�'R�a��M@q<���D
����yy�����;%F�6@vX�É	k�O��l�7�M��,��#޴�y�'g�a�!!&[ϔ��g�d�4����9P0h\�	�?9�'1�	Ο����\��	D�
���"�?:���PA��#q�	П�'�d6��Z����Ot�Ĳ|b�I9H��̰%!��}��ɆD~r�>у�i�6��p�i>5��p�6I	dK�-Gb�&��g?�	g.�m�ZDp4AVay��O=���IY��'0�HbҊ� J� �핆Dp@p�'���'�����O��	�MSw��._��$]�/.JB� ЁQ�������?��i�"�|2ť<��4|fpyK��5`�m���\� "d��&�iV6�8|6M}���I�o��(#�O�� �'	9Z�灧 �Q��� �~��'|�۟�	͟`�Iϟ(�	f�4m��Cyܬ��HU'D�f�	�e���7-�����O��D:���O�,mz���F�?�H$����qN|(���8�M뷷itO1�<$��v�,��8�a���c/؄b�Љ��	�
�ZU�'��%�P�'f��'}� ����ҥ�8]���2�'���'|"V� *ش�l�+O���8-�y�dcPri+'ї:B��@�BE�>��i6M�v� Y��E�A� q��9!a"%�:�IП���E��r<��P2��py��O����I#��ԃZ�>������5@�ەK��'Y��'br�S۟x��')'�,]�b��^g��ÑD���ڴk%�H����?��i��O�Ζ03���5$F�e�D��dU<8��˦�Jܴ.����E��6O���LO���'<꘥�T��%�Q�ʴ|<��FI߷t�69argй,	zk���b��-�W�0[nMk�#��h����Kعh��|:��Ʌ}�b�p���J~L<x3�ø-�p�yd�a $�	�FǄ9��{�Q����GÕTB:԰�HE57�<�����P:�<y��?7�Vԣ��
�Dy��N~o֨�#�F:d� ��Q�A��A6�5#�t���zqR��7SHh�9� ��+'
u��)Ѡ��F��u��#S 4���@я�!���F"��?Z��B*�@���e��rI>�*0���Ț`�
V%D��TC�6]pT�w�i*��'�"�O��Uo�Y�d�	+
f8C�	�#' �o����	��#<�~ī#�%����
	8���v��}�D�M����?�����x�O^�!�P#�΁E�NC�e"w`u�,���'���y��'��Y��^�j�&��A��n�Bu�0���O���H2b�&������Sf��n]+t�*M:TX!2`j��'���1$�b���IʟL���S�Y�3�T~�4�O�!����ݴ�?ae%Ϟ������'&ɧu׌C�.�m9�AF &B��1��ѱ1O���OR�D�<�3j�]���iTΐ�f.R��$��)&�h�ҞxB�'�'��I�0�I�׀ 0�����B�Ru��?I"�}@ciQ��?���?!,O�p��P�|�p�x�>�Z��F�A&\`��[}��'vB�|�Q����>D됍b�TYу�p�,q��*S}��'@��'p�	�U,x��I|*d�H1{����so�=�����
�kH�f�'z�'��	*K:c?)مM�;[Y�Z����x���S�ad�����O4�rݚ肑����'t�\c����i� %d�<(4h�4`�K<q(ONt�c�^ҁFE39��a��	;���·Ӧ��'U���e��8�O|b�O�X�W%��
��׸P9�]p�`� mZ|y2뗄���?'?7�\�WQ
M�E�ެ.�I1�(�*;��F� )a.6m�ON���O��)E�i>�"o�aur�)�ՙbw6T�$dʳ�Mq�Ku~BY��$?�	���FK�<3nH��  ;Z�P,
� 4�M����?q�����x�O[��O��*�D�B5F��B7hlt,��V��'78i0�y��'yB�'$����Q��<��f��#�v�`��jӒ�d�<�<5$���ڟt&��ݯj}<%���W��6���EA�e���\��<����?a����!��\3�?l<=�P�IaҢ�i��O����O0�O��('z�Ad�A�,��b�TZ�Ty�C̓�?Y��?�*O��H@���|±�M�f<9��$L�� #�o}�'WB�|S�h�ã>)�d	���yc_8.uV�b��O}b�'��S�(�I&b�OF҄@�}=��	`A+,R�:e�]�j�r6��O"�t�	��v���+��"[d<�C�=s� 	��Ԅo,��'v�	��� �k�m���'�O��0�4�7\��I��/P�^I�����8�	ҟ�3%��#�b��'�R��+�,P�p�R(�=-/p1�'��%_B�"�' 2�'v�T[��]56�H��LB5�n9��ʗ�@ *��?Q�ޗ(Ab��<�~�bj�%sF� �]5R�|���]ަ5S������֟��I�?5�����'�,-X��P>2�Rd��U0&"=��o��E�@�531O>��ɐC����"h�(o8#��K��L�۴�?I��?)����4�����O���Ggl,��$Q&G¤J����*sn���yBG1���H��OX�I�X����E���h�$" �b� D��,O�D�OB��1��=A��\�ԻR��� �ʌ�d�"�?��I[���_~��'8�T�h�I��n%Y��:��0�L�]Z��)��Vy2�'Fb�'H�O.�dБ� �� i�j)��){3&���#.!�	ɟP��VyB�'`�\�!џ`�z�G)k�z�M��#jd���if�'nr���O`d�P㐿'J��B�66H>�����afx@Z�(����O4���<������*�R��Yz�OA!;���#��t���n��h�?���z?��1�Q[�I�RtA���^�o��H�ύ)^J7��OTʓ�?��i����	�O��⟄�
tK�:�Rtր�3� iі.�d��?�p+R�*ұ�<�O�~d��g��	&�"�Y!��mɨO>��b�X���O��$�O����<�;9�.����X7���DP17�p��'�bK@	}tD"�y��$%P�%YH)�L=F%J :��M�0bF	�?����?i���(O���O�-	&aX��A�4�L�z��P�J������7b�b�"|���J��I��A�ԉa�e.{PU�i�b�'h�m�+j��i>������x�p�� ��]��:f�M�*���z�	��ħ�?��~���:l�L=Hq�Z'~�ELO��MC���Pc,O0�d�O���3�	�F��eZ�G��+�`�@Հo�O Ż6�����ɟ��'B�A$v��jة+<
�[�NO�-��IrV���������]���~2�%�ҹ��#s�Z��s����M[U��E~�' �Y�4�ɋ��}��U�@�q#���L�HIVnQ"�lZʟ����?1�;F@mq��
ަ�pD�0zD��A��J.T���B�>Y���?+O����
i��'�?	"	
0uo>��fdS.��Q��=F���'�O���4p[n�Bטx"hO&.���[�v������M������O��B���|���?���L�\��ԋ)��x�(~E�9�����O�p�Ae��-�1O��=��u�R�H�_H��q��,MrV��?9����?1���?9����.O��ZI���"7��<]��!�$�&q��I���8�˙N��b�b?�B��H=P0��*��M�ZI��iuӶ�� I�O2�$�O0�d����|��M����a<yk�Љ�lI&<�(�"�i`�sրR�Ř����$�Z����^�N�V�R%��0O((nZ���Iʟ����IAy�O*�'�$�P�ly�UV�?�R4R��>o��<��ڦ�OSB�'�dU7`*0��A��X�Bx2��=��I�~΁�'r��'�DW�6���[�/cb���\5���B�"���??��?	/Or���x;��q�M��'��d:!�B�#�aR���<����?A����'��懖���#��#.T�,�q"I�[Z�Q�@�V���$�O,��<���7un���O�X{Q F8_�>�`Ҁ��H�A"ش�?)��?��2�'��-��f_��M3�h�8<M�HZgHM$)�h�
t}��'2BQ�H��
W���OY��[�s�օ�Eh�Y�<uK �|��f�'��O���~9���x
� p݃7�B�>j�b'S�n�p����i��S�p�	&	��ŗO[�	�?�#L֗[��1�L�:"y�$煀��'l4o�����y���l�A�M��c�����%wU���Ɉ|7�a�I���Iʟ�SByZw>�����/.8�TY��*[�(J�O|��cz�\#����_�>�q A�>�l}��.N,6�&IN�2��'���'2�P��S۟L�@�˿[�X�:�F3����B���M{�cE�r�7�)�'�?�u�	�x�`��'�h{����^����'�r�'��k�Z��S��D�	o?y��_�bAH��!�#jY" YG�Dh1O$�QB�d�ß ��e?�����:���ЋX�;�D���%��)�IAyxU�'���'R�M�T�!Okn4��_1T�cX��0MS�xt��?������O�l�똲`��!s�\4^zȹ·�L����?���?1�b�'�b�/˭t� -���?i�$m�&M�{L!��O6���O�ʓ�?�����4�
Y�.D9D$�8b�� �����M��?����'��B[�UUq�ܴ:�DK����p|�#FT ��'��'���ȟ�c��WN���'$�](�(�p�R�b6�)Q��$;v�y���d1�	��4s�i@[�O�9`iڬYEP����^b�\y"־iE^��ɊB��	�OZ�'��4��6�
4��(�8�.%��S�d�b� �ɪ ���'4�~:P�X�	^�Rq.��8�p:d��G}��'�$݁P�'��')��Od�i����Ё\>2e3cAS2.��C�>��R�4h��`�S�'Ov�"��Z��Jɟ�6�6�o;L"b]��Ο������qy�O�R��(�БB�!׹)CJ�b���-a��7�"��#gk�S�O�]�=n�	"s�M,kGR���$�ͪ7�O����O�����<�'�?1��~�J�8����Wl�7J��h�ŌH:TJc�<�AD���ħ�?9���~��X�8((I�@�F�re+P&�(�M��uy`.OT���O��;�ɯ_�dŋ�*8�T1�sᛑaN��L�QYPe�c~��'��'��|�rY���$q�PN׊x�Z���;��Ħ<������OT�d�O���-[Fp 3����e�h�*�;D�1O��d�O��$�<i��\����'H5\mP�]�v0\@гlد|ڛ�Y�0�IZy��'+��'��Xq�'�j��%/4l���N�/�0\�k~�����O����O`�^|��#T?��i���Po�"[��)�I�1��cЮ{�(��<���?���$�hqΓ��i�|H ��2&��
�l��6|��޴�?a����%Z?��O���'h�$�Љ!������H*X
�0�Y����������z�x"<)�OĔ���oM�'��p��e�+o��ݴ��*�to�ğ��	���S&�����]J&�� Pp|H4�Iv��+c�i�R�'�����'b�\�(�}R�%�&*���� ',Y��6i�즁�6���M���?�����[��'i6QA�[�&��YhF�_�Jn��rio��񗒟��''�\��7[���J1��7��]�E��9��mٟ8����4hu期��ĸ<a���~��W�S��L��+x� ���ϵ��D�<)T��R~�O���'��ԓ\@}j�(k��Ax��ФL�7��O�l�b�v}BT���RyR��5&�/_L��V��`U]	��G��M�Q�P ͓����O��O�ʓ�n=b)�L��j��"-_2y���3\��Iyy��'��	��l������D�<s�����2��i!��}���	Py2�'2b�'A�4H��˟Ok�5�C˞�RH��&�q@ڴ��d�Ob��?���?�!�	�<1D�dw�����,T\tu���ѵJ3��4�	͟P�	��Z&F��M���?v	?�L�)�k�8��Xh����&���'���'��ޟ�T+z>E�	B?abaO��I��	��Ͱ+��=���0�'�m�0I�~"���?���5�]�a4z�V���K� ��xtX����� ͓���Iy��'��	χ<�@�#�k�� H& m��W��� ���M��?	���R'_��]�n>�}�جJ
�HI��^ @���n�ϟ��I#e``�ɺ��9O��>���X>�e��$���@�C4�rӔ̫����=�I�����?u��Od˓M��=���Ү���s0!�,|�h#�iB�%!�'	�'���:9[�����(@#�O�e2�%n�ҟ4�I�T:�iF����<���~�C$E$y�į��r���`�Y��M�L>IP&@�<�O{�'-IQ50�؉j6g�!D�]�t�>ǌ7�O6%� ��t}�\����ky���5��P�@p!O�h��B������ ��<���?������g|���G vT�ㄨG���0�b��_}"R�@�Iuy2�'<�'``�S��2vL>���,Q�x�r��Ǐ��y��'���'^�X>牖9,�@�OEp�9TD-$�� ��?]Y�K�4��$�O�˓�?���?��L��<�s�ɉB�*��$���o��0����Tc�F�'���'q�Z�d@��ȍ��	�Ok�ΎH$ b��&�4%�1LF��'?�I�d�I��(�T�c����f?!��	H.�*�4.�YQ$�Ѧm�I̟�'l��d�~r���?��'Dp+w:mH�2���TlPST��	ן�I18�����$�?�ñ�КH/��ɔjq*hf�T˓��f�i�"�'.��O+j�Ӻ��_Nh�L����(��A�g����	՟��@{������*�3� $P!��7]��g�NWbABf�i�,\��'bӤ���O����
I�'��	.rn���Ar��a��^�%%�8�ش d%͓�䓞�O7�����Q��/	�L���1�76"6��O��D�O�yZT��D}�_�d�Iw?�^�Nً�!�;s�����'�8���k��?���?��#��5r3�)�2.G.(�	]ś��'.�SF��>a(O���<i����F�p��:Kұ
�8jE�Pn}"��y��'���'Y��'�	���ADDY�`�mb�NG>c�b�;�����<	����$�O���O�b ��+>d= 1T cO4����D�X/�d�<���?�L~�@��g��i�O��6��_R�5���Q�x��Ty��'���'�͒�'�T ��s�X#���V<���&s� �d�O����O��H��WS?��i����m��G2AJ>0L��t�o�z���<���?���9�D�̓��i�#�N��O��%eF;f���c���$�O�WT"�z�Z?)��Ο�ӭWT����ϙN}n8k��g�z�I�O����O
�$�\����O����O���'{��x�`�^9[���@c�W��
7�<Q2lNm��檰~���ћ����ƕv���k�NĈ�xT�i����O�Вp:O�O~�>�����&6:bꂨqd��F�g��);�D�¦i�	ß��I�?�I�}B�5SO���FJfV��G�Ȕ~�(7��{��8�2��8zb� ���'k���i���'�����b۸O��D�O����H��.E�:�R��wl�6M=��ߔW���%>-���L�I�d� �h�%ޚ/.Ra[����#�>�x�4�?n*��O�$&��ƴ�����*hD�閇[0J�Q4V��1v'd�̔'��'�"S���F�IT%�N�2e�,��7 6��L<q���?�/Ox���Ox���-LQ������2A8f�;�hI�W�� ZR1O��?q��?Q,OF�����|
6#;�8���6ΦyЄ]��ɟ'����ɟ�k�ì>�d!@
�P�g�Q3z&mQ��~}��'��'|�?)���qN|*�G�:\jL�ȫ��S�-�F�'r�'9R�'�L�C��+t@����.ƾx��	 �$^0D�v�'c_��f���ħ�?�'|@Z�a�&S��r��6FV���x��''��!�yr�|՟B��閒4К4 �'96����i��I5�:���4"\�ڟ��S����}wf��ר
:jL�u��T�`����'���O��'�~��&�41X0�	i�����

�M��L�&j���'���'��b!��&�i��5^�D����߰@5L 8۴j�H������O���-�6�	`�B9���A�)s�6��OD��O$z!eQS��?��'���+���#P���X�L�:-H�}�c�H
�'%2�'5��)���:��sZ^	�Ӭ�a\�6��O�tNk��`��l�i�Y��G�^�P ����4B<ҡ�<6Mi�Ĕ'(2�'_S�j�/M|P����M6b(>���n��p�XP�L<����hOT����6dLI�ͅ�]�Ȃ$��Ӟ���O��D�OR��O����|2�Ŏ��?I3EށJ~�̂��ˇ��ѫ镎sn���'�"�'��'�2�'����O:}�t"n�%�^�s�I�
� _��� �	���	�HA1�D�D�'�Nb��D�}��B`R6Er�qb�jӚ��2���O��D$D��1Q�xr�	 f��	8��G�s�>���ꐩ�M����?a/O�����s���'���O���pR��=H��u���VB��;֡w���E��B���1U�Y����_��zS,Æ".P|nZݟ<��GH�!�	��Iß\��֟$�i�y�dX�����R�Ͻ�Nȹ�fn����O��P��FH1O��&�s�FR7-���j�&@�o������iϪ���'���'�r�OhB�'�品7܎%A�+�D��&ߌt���40�&�k�S�Ox��+
J�PQOC2w|�j��C�G�f7m�O��d�Od#� l}B_>!��ɟ�(�Ǯy���3�� F��Q�֣��'NV�(p�|��'j��'�晈��N�`\�C�� $z�P
vӴ���baLʓP������$�`��+O���<�f�X~@,���`�(��D�8������(��ܟ̖'�E�cΦm"����	l8����L
388U8��']r�'V��'��'W��' x�X�jF�j�\ Z�fձ*R۔�Q�cP�iS�OL�d�O*��<�Eo�� ��	�?o�1�qD�L�|��f↻k�'��|"�'�r�ȉ���ʣ-[j����.f�����6�I�|��ܟ��'x���E�1��˖Ybj���A��M��.=�x�o��'���I�����?���?�vQ'O�@[F&��&�6��O`�ĩ<���:��O`��O�E��,\�6��V�,/"���*>��OF�d(����'H�P���=KJ�2�2Y'TnZ�\��
P`������	�(��UyZc�x�:�.�+��$!%+�`w$=��4�?���`ՊYGx��	Z� �>I����c�0���фH�BL��Eg���Ն!|OԊ�	HK�����D�<����U"ON�� "H#�Q4�\+����փxQb�OO���pNT�@] ͨ�(\�����[%�l���Ӊ.�%*�M0O�T�I�#��q�!�R�X�̱�3%M +���Z#���D�jDO$g���#J	�9������W�L�� H�2w��Uz<�v�A�B��a��ƈ�i0kV��Oh�D�O�������?џO��8�p/��ה0�2��\iT���:�b��C+B45��@ՠ*5"?�m�6c�D��5d[�[Y$�svA�)�nD�V,�RF|�)Uc�T���2Aˊ�R��(��b��Q��#5�ؽp#���Fhܼhr��Q`�[bh<�u�Q�q=��u3!	B��P��M�<��䌦
�<�04E�/Zt���eB̓%��IFy�,�)vN���?I���*4@ּq�(9R`�3[?�?�����?a�Ol��iŠ4 Ⱥ�+W?q��R�]`T�D���&�1W O��p<�K\0�:���d��I�ߴS,.]#�j�>:/"Q�`䂑?���	+�����O:ʓj~A���� ��EI��Q��]�<yߓG�,�`���L}�� S�]�u��l��|��&b���48�GK�Y���`a��yB[��BĄ��D�OR�'[�~\��O�-Q�Lրo&�� >r?� ��?yV�6o.aS�E�`vV� ����|�į��D"*u�p�ӝO�=;'��u��޼~@�z��\O�:��r�(ҧ�rp�S��2B(8�ɞ�m\���O�\p�'���ǟ��D��>+��t��֤V|��J�!#D�Њ�#ν5���!E��?��t��f OPFz�fB.X��!�D�l��W�ܛil&듎?Y��;\hKv�	,�?I��?y�Ӽ��X�k��	�'gU�({�q���ǻ|��U�5��
J���xF�<���L>���Ϧw9�GW {�|iH@j��~<�L�b�ܙJt��N�0�l,�}r��eU\�I;^�2�)*1xA F���|��R~� ��?�'�hOb5	����O�p��F ��F ""O&�Q��<hhꓥ��ٜtbǐ��+���?Y�'�л����PTa���]Q5���ڪ[j�$9�'��'���m�E��ͧCĆ1 ҈�J�,%��j8y�pXW�I��ȡ���k�$8�ϓ=� j�f��M\���M�lqU�H QV �Ǉ�����`�b�G|R����Ed�:N�(m
���"���� ���`��j�'��O@��v�H0��p`��9p��	0C"O.����F�1��m����/�n����$r}�X�,�N?��d�O�[P�̦��x�
ܡ$�� ���O��$(Y����O���2'�`<���S�4�B���'N8b��ڶOjά��'�T�0��B��@P��K��%K��O�({��!0�T�p�C������'��lP��?/O��H7o�Έ8�W5>L\V�d7|OUb�#Պ^����%D�!;I8I�aO�m�&E0��*�V�À� Nc�	fy�
:7��OR���|�&�R��?aĉ!�t���@+a�@�����?�Q��0kӰi>1O�3?9���	�2M��k P
Es��Vq�߃pex��?�!4��l�����FL�A'���)1}��?I��i�
7��O��?�Eaڽ�t��3V��m��!=�	�����I=[��xӦ&Xx[�}q�=8N���$DI�'_",��X�,��pgBN�#6��*�b�"�$�O�̛M�r����Ot���O��$��dD[���k� 3KR>�����*�	����i&��@.�-K�@�}YB��k8vB�#�y��Z�1�X�}&���g� ���V�����M��i7��$E{��,O��$Z�z�&/z�B�%9l�C�IOt������|f�  _�DW��>�HON�'����:4$��v��=y��9A�.F$/=��3ugD3��d�O��$�O6��;�?����JN\�b2dD Z��!��: �Lp�R�'f�h��CG�ƴ
`@TT*�3ƋH�iT�rG�_�Z��E�Ν`��aqGPI��b��?IO>Q��?ُR�'YDmR`c^1Q���.�0��\$���HC1G�����0-t��<y"[���'r
�`d�>1��+B��ɰ�A+=l�Uie���d�. ����?Q lE��?!������ͷ2���y��U�ʤh�� ��LS���jH�H)�H�Y2��8�����t�� G�:EF�Q�`%=�p��#U�%3�t�TcW��t-���
T�'������q��&.�>ae��$B.�0�c	� M�B� A̓�?	�|�9�gԞY X�I� ��R�B݇������ a􋐥5�z�ˤ����y��d�>�}�'�p]+�-��yV���ũY<P����'�2%�ac�>bY��Ia�1�
�'����q���y�
�>�de��'H��!�.��8Z��<'t��	�'� �ӳn\?�zY��C��"��m��'��e�&(i��:c$�*��C��� �Y�'ܡ�V��:��hD"O���e��W�l��@�JM^6��"O ����!+aBe�0�Q�	��di�"O��*w$G�4�i1�b�)�"O��zq ��K+�����TJ|���"O�p��T�e�^�6�I�yX]�"OJP�b/D���Gc�\	r���"O�MP��V��E҃Z�x����.D�<�SDI�[��I�lZ[e���h(D��Sr�4e�� %W�b�y�v/(D�\jc�у-2�Y:��զuoҐ؁f%D���w&G.o�:�zqi0[:��#*6D��Q�@ҫJ�q3�a�^lٗ�1D�H��ԆS�Ex2W(y���p �$D�Hkv*���%�Ժ01��p5D�HR�`�"?�P	���T�P~� c��&D��� ��n�����<\r0`a�&D��:�(����- ���;<�h`b��#D��g�I�O^�\ɠ��I?4�c� "D��b	��n�HY"r,�	@2���?D�HAf#�Z Ld���$!-�xDE1D���L
�I݀�v,]N� e��"0D������k�`�2⧇�S�q�O)D��0 ��=;�X�Ch9"����3&D�Hb���/�%�B��Q� %D�p8.C�9
x����!<� l�d7D�`0�
V�����5I�����'D��Ε�BM�`��fʍ�Z��o)D���r��G@rhn�)(\.��P�%�O�q�PSw�*�Q 7%ZA㒇�&l����&��S��sU�n��@h�n�-L�r;	� $~8e�ւ�z'��)F8Dx�)�(g���v"҆}��z�B^�ҍr��@�<��5�,���r��-C x�������BMI jLDI��D\p���΀�pT���H��;�D�Rp-��	A�iT���tc���M��y7 [�]�4m�v�>$
M� �ɱ�y�@�PO��B��X����`Z����
�'8��WJ�-- 6t[�O���@���!<%4��X�(�eÛ(�ZDBϽ6��q�7;�O�;a�ʞ��g�$p,�`��7�<��Se��<�a����f�9w�R={��)���/��f�<ڕoP9xr������Fx�+�E�0;2'ǒ�`�q�N�_7"q�U��C1�!Z����F�
��U /r�:+����	O�JF��gÕwӺ�
ϗL���l��5��}:��R� 8l��$	N�NV�Y�oӵ7S�sޭ�
ԚxQ�ܪ�|͋u�2D�4�3�����+�@g'���4$\9Ha���я2�T�q�&�(�B��]b�h3L=�r�'�����)�\s�aP.���OS���^q#���8��bS�\?:��8� K�g�ZQ��IRm���ˏ1��y"����Ox}IW`��zq!���Z�r��ɶ.\����شC�J�� N 1C9�Lyd��+�T)��^O�i9&����x���K�Bx����?�\��m��K���2��w�P�q�ą!Hf���?L���9��=�L9�Bm��p����y��4=�$��d�;^Kt`R�IP4�yB׆C�(pZ�M��<�Da�T�F��dMx$��d؊UNj��K�OZ(qX�A��\e�`�RW����C�O�����U
6�H���m'�OR��A*�=�@��'�=+,��*ˆ
D ��(��@�+Ȯu�Z�mS%b�PB��M �I�I��H<���).�
``��D�D�A�#<�2��8�h@��ڶ# ��1���i}B�()z" ��l(fr(�W�
<���/Ry"L1X�:b�b>�Po?U���v�
;L��Dk)Auv�Q!��?w�-���L�4&�_^n@Z��~Zc�}���D�����0�/Fb"�ˤ�;���L�"#|�'�,!�U-�w|����T�h������ē�B�sqW�Ժ�˞G}6�	�Ӽ�k,~�f����n����.�F��'\�x�%,+�l��Q�zuf!Ad�E,B,���%ơ�M�GW�`�l�Q�����i�f C��T��O6$
DM#M���j��E)�����I3�PlJ�
�,�I'R�W0�a�$�V�hR5���r�	�Q�LA�cE��0����E$���&<��er�I��"��h��$m�.��dp�A��bd�i�	-�|��Y���R$��f��|jԩS?$��{�	�,M�ONE�!�3?��	P#[2E�C�
�/���2�� 4�=�@�<���5t��8�a��y'��NE�EQ�OP9� �[���/6�(�Ԥ:<O �Y���vj(�� ����ɻ ��р�Pk����4��?��	ͬxQ�C��|b�&�-�$�aP�x2M�"az2|�JI9*'���󦏤�0>9���w�$욢E��qN<(�.��;�J�0ǡBZ�3�ԣh"����D�Ik`=z��d���ӵ`[����/W��@������z� "<P�+A�I9Q�O��N�Ha�{~��M��cD�K9F��0���Ť/X�0�`�9�䚉MW�E~b�B�z]�@�u�7����&���*ūӍ���r�ɪk��ٍ��ywC@6]@)���/[�	˄��3?D�P5�O�@�EG� �,��M׽tPu��4����;`S,��Eǝ4�Pt�2O�-jѠGc+���+�zʅ�BOZ5z5	����@`��
u�0�2��]?a4g"�T�Y�aΰ)N�D�f�'q�T��j�Iu�E�#��if�(˓a�)�BO·YR�!�U&޹J>����I�%<�� ��_\��Lɋ9>��XF�#�OL9�w�A�1`��E��5o`F�T�x�'+^�� ��	Gv�9�6���T>��u(�d�P" V! �t�d =D��iCmΚx�t8;�iׄ&TY��չvT歋CB��#vLdZ�b?����˼�c�A�� �WY�x,B�XU��H�<9��@�F���є疦.��1�g�ʿ3z�m��}���Ѝ�qLX��O&"=)�@F�5��dx���~�T�#���Z8�P5���
$��m b8�&Ə#+V�Ѩ�͓ \ P$�iR��s`�:�O��;r�K?7:�be���Eښ�� �'Z���<Oz!ň�t'@��U�$l���`"O
hbBA��Qi�'-ހW�(��I!�(#~��F�#dl�AR/,0ek"o�m�<1���R�d��E��k<�Q&	��<i�@�������	�tk�>x�0Q*��!]jqB�"O��zЌ�@�Y�kN�KBҀ
2����b+�^���J�GA��d��@CT��fh	�2�O�$��I�O�p���ؽ>��H�o_�f�&L��"OxsŢ�2g���*���:��3S$*	3���#%���?��S� $\Y8U���E�|��4D��������U6�|Z�"�	K��d�`9l���RǬ����V�I���W�dE>�"~BÊ'%�&٘�B�Kl�Qe(�|̓ C|��(�>0��QF��Ō �`,����U�qX�o��yR+>4|���'J�D��SN�(��A�aC¥�����3X>�:��
�`LG֊��%��qr�؄�TuR#���k���htH�
�* �'4�
�f��N��Y#G�B!s�iѕI�
@�B�8LO���4�˦S�Ta�<OL�`�b�)w�>=�&鐶��4�B"O�%�f�ٵk��Mɂ�G�n@���F�jP�S�Y�o?Q g��,��qGI>/�9�)#D�Pa�J������Ó!ɜLx�  b��Ѫ,?�pb B����d��pD)�78 �����F�!�$X�|�J� ���,���7Ւ���Et�^����'	v�kԏ�?;��d��JΰS:�*ӓty�e�gَ-�@5ϓP��!�NG�9h���r�
fj�d�ȓ}����p�thSl��Ҝ��<)�l�� ڌ�g�YI�OR���K���Ռ֬{��6IK�X\1O��)��3?��'�^�2H ©W&U ��Aa��w\��,�F~���6�����dq�%Z�`U-]������g�
��\�<��0�'>x�M@	9��qQBk�;"��ӓH��5͜K~B+R�p\�a#E���R��g��;�yBo��9��
%JF�Z��E�'�1�D�p|J0#OɁì�+>[�W��y��=r(Hْ1��(
\�E����{���c�yr�����I?4-j�K��Os+j�R���'i�iy�`�� 820I"oV0y�~EK��s��J
�M�*ը�M"Tz��`9P�j��hO�ĄK�b�O&-��A͑y�����U\��Q��"O$$�db�qX�|���K�p�V �R��J�t�F ���O�\�	�)͌#A����)a��x
�'Ƣhzծ�:5��@G��W�����,��Ә'�����𙟘�%�$$q0�8p!�d,�H:D�@J���y�z��Ċ�}VB�:qF�0&0��g�&�OԀ�g�A4x�H�HL3s����"O� �p�"����P�V�E
�@DR�"O��#� ����r��\��@�"O���KM�.��ܢ�(Q�*m����x��P�T]�82�c��ȟ�P`�܆5�p����
=4�1qq"O��RR��&��M
R��7T�=)�
(!��P�'g�;��$�3�$�7Rr��GIMv9�Qr�#r!��?T���5w�����k�z)���*ٰy3׹i�ўb>ݡ����GȰqjҏZ N��p�v�&,O�A�T���
9��]�\j����s���h��#D� s���#\�¹X"�(y���j!�D�U�����!� d��?����@�a����|��U�V�!�d�P:&l���T53d��E�� ;QJ%c�T~B���E6fb?OҼ1d�"�,yY�9N֡kO����N��2���Dt��"O���t�[#�a}�iҴ'������ܼ.�R�Yb��"�<i��Ի}Uh��3�Ga}���\��ҡ���A���yrZ��lr��4��I@'
��y�Ty��C��p7�!0�& �n��ȓ8-�|��b]hl��[ӭD�w�
i�ȓV����T�CAV�0a��Q���X�ȓ.�X\i#�B���U�A��(��I#Dxc�ֺ����@�ESa��~}�h�b<�ܔr@��)H%���ȓg����7���)�&!
@�L</؞Յ�]i� ���gxL�)������k_ h�1퉄/�Z�!%-�99`��J�V$��'�
4_8�ɇ̋?�LU�ȓJ�m���ԓ���9���u��ч�c��9&�U5a���C$�V̇�$�,��Uʚ�}��-��������ȓI��`aS!�,��pR�݋p����'�N�Ό�)s(ɽ).̈́�Q�8�8�*I)|�����I������B�`t����P��ıP%<���a༵�w�CDS��k�����@��ȓְ�$Nf���6��ZU�8�ȓt��,�V��:hU���Hά2�C剠;�Jx�ï�yE��gΓ[mB�I4�x4�$\�>��P(B�P:`����lL(qQ�V-(���`&B�!�B�B$<�k�ʕ�[�j����$!�$]%E@v�I�Mݽf`�Z�O��nZ!�d�k�*P�O�V��2�	o�!�$D�R��Ν�|Ru���޺8,!�w�u�S�]?�{E)w!��!�J�y�hE�R���c�J�>X!�d֠;(d����2/|��'�3�!�\*�\E8G	��N
@���i<!�Ć�"b<k�#����)�A+&A"!�dQ�t�-�!يxЁ`P	F�!�є4�%3��
)�,a[�j�#zo!�dӼh����-@0�����i�3X!��5>~��I��xzh�yq��9K!�$�&�N(�� -��칱�45.!�d��8���E  �U�J�fG�'"!�DD#n���T#¦v�� �rL˃�!�r���H �Ƣ}�����?o�!򄆺G�����X"L�H×獉|�!��O֝0veJ�9��ɲ���!�ĉ&AT�Q�Ve�ezRd�Q��!�U��V��&�
pW~�;��=	�!�d-�*Y��4X:\�c�l�U�!�dی~"E�&�&"��M�`!򤓓�<�,�Eĸ�gk��tg!�� ��P�jK%I��A�C(n�^i�!"Ozt�"l��:D��IVr�b��P"O�ig�I8Nά�òJ�#�*�y�"O|Ă".$��!�0�ؒ@r*�Ѵ"O�8b2&��`qaD��\��"O����{6�r+T�Hp"O@�hD �]�Pk���2C�h�2"Ot�0��K��Q�*`�iZ"O��D�Tq�tд)�+Y�r|:�"O��PL�B|���߃(��"O�}
e���~�B%k@�N\�Uѳ"O�C!7#�f��lC�+�t�	�"O��e��moP�"�.B�6�4"O.�qc�b���1�. |�8�"O�y���5����C )`@qA"O,�鵅��,�ź��&T�R�"O u"r蛲`q��bg��7����c"Oz�2��V��B��G�.z�"Ofeq4��Fε�eoY�#�j jc"Oz��&�$��3n��((8�`$"O�xf.
�!��Tb��
���J�"O�B� S�h9.Th�AD b�$P "O�Q��ᅿBWb�;��Y�5�"O��P�+�kИ��dB�'�� "O�!3�M�W��i�%䍵K���R"O���cG�"[��KS�{�ޱx�"O�	c�ʡ80y;��^�r�f���"O�����4+bu����{��)��"O �p�R�5�"q+Q�.�� Ҥ"O�8��n�5X]|�p�ʏ�&�ܑ3&"O��P����q<�k�o!p��;"O굑Έ1gj�3'��@��S"O��iq��e�8�d�ھ\��ٕ"O��iq.�5c�<a���X	�mx�"O�=�RH_�9!l�^AF��n���y�<=w��֦�a��L����y�E�&M^�c��(�K`-��y�ېA��i�o_#��@�����y�����r�
*�W!ґ�yR��_*aR��D=9�F՛�$Y��yB�8|�Iá!�?5q6eEoɻ�y���"!�X��IF@��`R.�y��	�@05҆GM�oV�+��ѷ�yBoȾ��<J��8>궥X��3�y�`��=A�o֐��9���y��e��H�FM
~����5����yB�ׅ?�`d��ܦ @��^��yć�x����-B7,�&���y�)C".��%)Rj� 䩉��y��P9��-���6m�a!�� �y�/D!�xR֏���vl,���;�'���"�3���
iUֵ9�'��9�Ē�}l���͟�P���!
�'���K��L����e�Gj(�	�'��P�Y_�Z���X83�^-��'�l0�C熑M��h3�	�':�~��'�Z�3+�e]� �dP�h��P
�'�t3�,��5{��AF�	�Uj�}���,�S�T+E�l_�Z$���U� "FJ!�yBBǱmMb���Ҹ=$ƇR��y�J\�+T������0�j���y2�S2p%����t)��AE	�+��$)�O��!= 5�U%k�G�P<��"O┰�FbC��X��~́�T"O� d��eǔl��e�C*K7 ��"O��2ÂU���3Ԩ��4���"O,p�ʁ_	z ��L-b,���"O�	��;�xh��EF�B� 	r"Obe�)� 4�ڥ27��R�v]�@"O
m�&dDoXƱ����x��%"O�ċ�e�,��$�Ta:X�a�2"O����@�M6�ٓ�o!Bδ�a"O���B:&�S�n=h9���"O�;7�	�2��2L��y�9i"Ot�RԣHIA���k� L����"O��`U�ӭ����Qi��:hr�pg�:�Ş��`���*A]��BAL�f�ȓGF����ϙbD�r��6)�
�&���ɭոqK���9�Ht;���[�B�	�V�H�d�lӥb%f���bK>D�|�
�:�q�aC�U>�9 �>D�D	�/K$bD��4R�Q:�yǩ=D��� �0ZڦJ1��'+@��d=��U��ħ9��@��/:�^���ǌ�IO�|�ȓ`(�0�1Ɏ�Z�.�#��Gp��ȓS�(��$< �|c�f�I7����N	�c#�#,z�Y� 3VH��%D�PqMCQ3��$ �:@��87��"GD�(�����	`���ȓk/^q %��*�J��?<����Xؠk".��v��
 OХ2��$�ȓs�݊�g'4�q"��#	
X���:�b�a7�\�",	k�
.�h=��ql�eQ7�ͤ�~���SG��х�}�f+��2�YI�Uu� ���	M�ɛ"l29` [�������ɺ��B�ə`�*2�4[:��˄#lB�I�p�R���aX6�2|�2�B�u�>B�	�#1��JUHM��
��ѣ�g�6&�DpD��I� �2'�5s�?D�t E"�6P/�AS�W����3D��yW�
/O,XQ#����A��&1D�X���
`bE3`��a
,�G�0D�؉!ȞN4�m�vl�K�+Ђ:D�(�CX+u�0��D�_߾M���6D���fh\$@�&ћ ��7ͨ�*�*D�x�W�Ֆ<��Sg��jAy�g&D���@��?]����D5PPK%
$D�p��UO���I�
;o4�RD�!D��B յVq�d���#@s ��+!D���FO��$��쓽o\���h9D��B�)�Tr�$!d��0��	�$!*D��Q�F�I7�<���C;((��3"�#D�dJ_&x�8��p�Dλ�PyRo�n0L�J�o�z�Rhd�Y�<�GS=P�Yz���[F���KV�<��,X'q|$��F�b���gm�<��
+I��e�R�Z�D�UHq�i�<٣k�:�j��r(�C��`�d����?ф@T�x��a�#��+D¬c���z�<Q孅+���S���$h��v�<���Ė��qP��A	~�,:��u�<��+^�`�2U�۹%��4��	�x�<ena8�3�1<��BKJ�<��� %6�)R"�_2G�4q�7�HE�<i	߳v>�B�d�x�����HJW�<��Y'��� �$r����
S�<i�͝�I�,�B搥"���7��K�<� v�
�ME8+*`�(ĉߕ(Ez�RT"Op0G`��#̀��F��k.�5C "Ovu��jL(/���j�F�Y�"O$�P���	���8�d�2ulE""O �P�n�?9�U���ܙ5�E�"O���e" k�,��P��7�X�A"O�)�&$�,`J�R�m�r�j"O�pPAH�n�����RhL@�"O��b���=id�#�e�:3��� "Oz`$)�&{QF��P�@���E"OJpka%ͳ%��y pÏ�h����T"O��X� ^�ìh�'c��<wL`��"Or���.�bS܋%�Q�S��4"OF�z�
T!A�LŲ���
E�B�Qc"O��FA}L�cԬp��H�P"O01�AaC6Y�Z�L�yn~��s"O̡��͟T)��	��*i��"O੊U���\	v���XO�!�"O���CXK	@Kօ�Z�Ђt"O�=p� )2�&t�k�*>,�"O�غ��&�N�J)�D$�)�v"O�Q�$��(���tG?v8���"OtL��F\�F���g5躑"O��Cc�+_ 4	� G�M&F��W]������g�.���ܭ�������2<�C�Ik�T=��+�K�ic`��L�C䉘XV.P҂Jˢs�ڄ�W�B?4nC�S�9�iدJi�HyP�B6{o�B�ɚR�$-لhW8s�J���d۵��B�ɶtR����Щ�&�r��ّ.D�B�I�]��JO�>�xQ&8e�B�� ׂ��'�W8��8��L�B�	IT<�C��#�V��EG-MhB�ɯo��8�l&�F��kE(~ C�ɗ:�%nԒc�~���hőZ�B�I�{�\�@6�T4bR&`����B䉈B�ز����@x��ݬ8��B�	�*���S���^�^L��m~B�ɨ<贅3�eāe��8�L1�:B�I*S�Mj���Y��\�5/�2$B��7>����LCZ����h�xB�	��P���Bv���!9��C�	�/��%��gJ�*��H���hP�C䉍$X��! %������U�tGDC�I�!`����"����O�CvdB�I;;�(D(d�ȎAz�;slA�{T�B�Ir\<K�$1M1p��VA�!$C�B�Ƀ�T���D;X���[1(��q�C�	�;T�!C�Q��Ƀ�LD�
�fC�I�1�Dxx�G48i�����o�C�ɹD��ؠ�>uD)���]�XC䉚`x��$��?NY$�z�
, ��B�I�V�[��0 ���� �TB�%&`����L�� YR,QU��C�I�l��k�/W)o`ʌ9�+ҭJ�B剠Nl�L:�hݼ7��I1���.!�$�&($2LA)ݤ+������ֲ+!�d1�j�����k.��T��"�!��Mr���BꀇHZH3�kߝ%�!����.r`���pT� �A�)Y!��Z�ok.�Gm_�A7X��M��$ !��>k��A�o�^m���@!!�d;"<5СƊ$�Bk�� �!���|�ɓd��1�l���D8vC!�� ��(E��DjL�{��fJ�b"O����%J�|:�	��0>*�!W"ON`�*�)@w���mQ����ѡ"O���g<$�~Mx��[';�|��"O(���(��6�MH1�S�E�	RP"O&m��
	]��# V�쬘`�"O@g�3��0�EU7x��!s�"OD�a��_:����E�M(3�4��G"O�`���ŶUPpD��  .{����"O�R�I �X�h!�>/[X�ʱ"O���ŋ�e��<��GB�����V"OD�
�J�/#.e[RfӘ)� �r"O\Y�@�;OP�kÅ�LаD��"O�ʴ�]�I��a��.#E�Dt"Of����7B2,�.	�A�Y�"O��;�م@z���
�r�B1d"Ou��i��ްAW��7v`XX�"OѱTD_	-U0�Y.ƕ,ֆ��d"O�e�����h]c���D��ݚ!"O��w�#.j�	sQ.]��P��'H
��������VD�WJ ���'�|�pf�v|ⱋv�ދJ�!�'׮�c$�h@�Õ�Ğ5�=p�'�<��S'�6mN��J����-�V�1�'�����k����S�nD.d1�'����c�#1V��(G>���"O��A��Ɔ2���q�	w٢9�"O�Y�� ��6�N܈uL\�q�R9��"Op���+��\��t���Yr�j�zR"Oj���-.m�F���7�� �"O����^�SA�t���\�.�X�"Opj��G�N*���@��P#"O4���cH1,e�yh�HF'%q6"ONq�WG�� �4��%g^!1O�=!�"O^�zW�!�ʠQ3�[�;���X�"O�l�� ��G!�K�۞y����u"O�����
O��ce+Q:�6Y��"O���0�݀1FR5RA�m� �f"O�M���W�ygv��I�,�"O�Y9��T`�9������e:�"O,�@P�A�Y�a�2�6"O�=�$�Q>a��M
��F7�4�v"O�2aP0%L\�a�Q'q���"OX�I��֜À�(e��2$e���"O~A#7'R�U�Y�pIKÈݴ�yBDȗ��Jǯ�79�ӏ�	�y"��_R���T��>2����i��yfP�BL�2C�S��})�fɟ�y-߂�b����"L{ĝ�r���y���&p����j	vT��uG�=�yb%[�|w�fME3rdXx��b���y�l��Z� ��h܏dizQ 境�y"��2Z�.A���`�=�a��>�y�C�-C+�̛GA&dlQAH��y"��+$�
l� z��OS%e8ЅȓK2f����R� �p1��p\p���;�bW� �w눉�"l((�2���bYs�돮~R��Ёju�LE��@|�݈�%?9 Z���nY0"�B��ȓ':b�����E�4#ڳ9��D��`|B�aa!���;�뇯8`h��ȓ��lY��*�d;�H��tWnl��d���Λ!n�R��͇W�d��A�8� Y g�{�o�� H݄�S�? ���hʌ7�JD;�3	�����"O���q��x�q╊�Ltx���"OnH��(ҔuU�	S����iqFA"O��:�/�A�t���H�`�T�"OT��a�+v܊ {�Eן(���A�"O~����@�IP2�c�i�:1�`�C�"O���$
�-%(U���!d`u��"OB̚�B2I2����'�
A2��"O�mѤ��|��ǠK�P�0y{T"OdAB5-����:2`̵T�&u�0"O�cC_6��,��mcH�7�yB.�&!)���ġ4p�4�Ҥ����y�  �{���K�U�i|�1��X%�y�bŊ�H����-�I�2���y�Ú�km��J� �UO�h���T/�yb��?(|b<6G	#O� ���k��y�퀉l���� C�Z_D�z��ْ�y��H~t(m��*�#H����3�V1�y��ޡq�)� ��</�h�jY��y"
�?m6\��w��&`���B+��yRQ2)�䔁gЦ�@Q���-�y�Ϝ7AB�i��e
�@�*Y:�yҊQ4/�<�"����-ۀCŔ�yB��b񲖪�3}5� i��y��|�����w�Q�H��y�@\<C�0�`�K�n�f�!c޷�yB��#a��R��2���;����yR�T�~��dЦ-�r�H�@��yBΗ�MO �Ȇ���1�~�������ybX!&����3��9�v}��!O0�y�KB�9�����?ʨ-c O��y��ٌ
4a:'㜣Iif��f �y��J2E�������*J^���H�!�y�-WFҠ���ϊ$8H�TKL��y�ɞ�xݑ!���M88��a���y�K%xn&�Q�.˛������y�b�#k��9��כ�褚�JQ�y�[m3�����@uA�ǹ�y���Xvع�Uj8�^y�W��&�y��Ǉ!�D �	E�3F���R��y�J�6?
ڐ���)�"���!�1�y�oV�
MX���#�H�F֦�y� ��K�qg��� �b� 3
é�y2�C�B��p*Գmr��!�X��y��jX:�q��-5B�����X�y�bàm�J���$#h40�J���yrR�7�z������,.CEHߩ�y�-�=��b�C�A��&��y�gR�Y�aFG	�b����\��y¯��$��ŉ�8<,P��Ƃ�y�o%��F�</���(g��1�yb�ȶ ��A��ޑz&8lk�G�y��+Ir����7vj��#B�yr	�0Wr�<���(o>������y¨S%K�$�;U���	��U��y�&֙w�z��C.�E��JO��y¥��v�����HEt �D���yb��L8p�I�ރ	i| :�Q5�y2�W�0R��qĀ�Q�BSMC��y�@&Z!r-�h�4�xՑ3���ybMX�Kz�8R�/F�;�rI��	;�yB@�)&�2����,k�+t���y�
��U������*���3�3�y�I� e������;0��I�����y
� 
�Ɂ�Í^�P�K�o�<%L2��"O���b��N{@�����F� ��"O��1���7?z00��|~�-*�"OD���ϗ:4��D�R�g�8�S"O�t��\2 ������eg�Q"�"O��Ǌ�+��=�����%bP���"O(�`wQ=���!��0�8��1"Op�!�č}�dH#�k��n�����"O;��/H}�ǯ�L�J�Ie"OR���)��-�M�<�P���"O�X���5�F��*��Y^�Z�"OJE��Ο�|��Mb��ʍpV��"O�a�ė+b�s�%�8���c"OH,�K�8�@�DS1Fz��A"O
m#F���PH��AJüu�
`��"O�@�l� �ؼ'	�Q�h!�v"O�� � ͝;�L	IF	��8;���u"O�1q���U�6��w\�/�<�"O��Xv��3w
TS0�Ŗ 6L��"On��%��=�FȨ#bQ����Yp"Oڈ �G�K�fu�ԂN�i�ƑP�"Ol����Z�q/xա��8�����"O�X�m�%���&*�ʌy�"O:p{5![*�:�B�\*_70h��"Oƅ;C�� ׈M����f*v��D"O��K�@'8Z5Ò�ӑ��l��"O:�s���9�zt��j��"Op k�%N!{�)pe�� ~���5"O��������~@z�	��r¡ "O&;��ӘR�������zDXh�"O����X,�Y"e�P�=*���"O2�A5L��fi8���.r�N�b�"O�lI#�%(ߦ��%�T����"On�`��ظ&�:x#`FV�)���G"O�] Ud� j|"M8Ee���"O���Re
.��C�%�l葈�"Or�%I a���G �E�U"O����E ^5SCFt]���3"Of��0,,c�x��
r.�a��"Or�0v�J�ظ��X����W"OIk҅�.gv�8%��p?��;`"OZ�C�	�&wY|Q9��#/4��)%"OJ�����. ���CJ�~#^|@�"Ot J�C	�h�숫P�^�%& `hT"Oz����b���H�S�	X��r"O���r�j�q�j�<#`�A6"Oܝ�Agɂ#?Z�S���ab�"O���Ņ�a���� �'mmD �"O��+�-��E����3 ��@fr��"OJl����2��\	��ѝ(��4*%"O�H��%�~pȓ���h j6"O*�*��0�Vв�+��v�𬹲"Ov��Ǩļ��Bshӊa��D�"O^�3ca�y�¹j�&ה{�䩰�"O"i�\*֠B�@��%�:q!��A��y�,�9��#��\$��1��f��y�,��<�~E�3#���~H ����y��ڹE�1j����~Y�5�B+��?��0eL�Dئ��dX��ͪkj�� ���x� Z�/8���G_�xJ�(�E�C��y��=C��ѣ�j�F���ħ��y���9I�2]�t�[�DG��C#D��y�)��Ҷeב
�( ��"�yr��=|�pFK��n!p)�a"#�y
� ���V:b���k%����	F�'��ߖ5�ȣ�k�Y��Pg��'WoBO���1
70~V�W`�)ՌV�<	���L�BgϼS��@��P�<���+\�RQ��Cޮ+����c^b�<9� Χt��pqua��C��(���_�<�6� /"����lI�$l�ȓ�p�<16E��(����:r�bl��n��p��]aVѸ��3���[!揲q�T`�IW<iu�)tV�yPK�7���b�Zb�<��m������El�R3%k�Ƙf�<12Ɨ�?r���a�L��1�G�m�<�Co��'��q7-��Q�`陷�k�<�1�]�昨��˂W�
(�㡃O�<�0��:� ��5�MRƬ�9p�G�<Q�!�i�<�8r��pH����@�y�<�f�_C�M��I��4l��y4)�J�<��A�)��]��ۄ���!�m�O�<)�$@�Y���Q$�m��0s�E�<a�o�'�")��Qj�}�@�l�<���i�쭹�j�0�B���f�<1e-ޞ	NH��� r\f����^�<���V<��d�i�p)�5� b�<���<A�f�q��-v("#��x�<�%�P�촠�V�Tvz�A�%}�<1�g�%D���RE�&�})��r�<IƖ� ������Y��\�Hr�<�d,�
8�$B�1@N��R��D�<с͑[q�e:�lL�7�ҥ!��BC�<	��!!ݸi8�n�JG<�I@�{�<�G�I�xH��ɅS�DP!b�b�<Q�U�N02i��I�?�tQ��D\��z���O�t�!ޡ��M����?,�Y�
�'&��Y�� n��ئK�#)ӤŃ
�'b�eA�IS0X����%`� V�L�	�'$��cK�6�� ���\��D[	�'����'��.W�L1P	���D��'Yf(��֢E~bg��(�0�
�'&z<�ĞEJ���.��ey
�'R"E&���M!��S�&fF��	�'X� g��|��p��ETS��X	�'��#�aM����B��v���'HZ�rW��2�����ޘzt��'>�8��mP���m��������'_,a��OT���th��)̶}S�'�2P����G�l�l*������0�~Y�-�WÖ�|{�acg��6� T�ȓH{���d���TȰq�֌v4t��IN��@q��22����_D9���ȓ7�d%��3	��q@�čI��܄�8��䢥�q���k�ʁ7�<0�ȓ��N�f�xk�e�?m)�h�ȓ��1qB��
'����My���E{r�O��h�ҤשH0�!y�d��	�'��iȵMx*�sW���pPֽ"	�'Bf���(�,2�2ұ�B�a$"��'�N�# C٣b�Y�nG�Z�ڈ��'@�!�c9|M
 cї)?HX3�'
 ��B�Ғ0������P�U1"�X
��O>�!hEê�c����@*"��i>�#��Z�u�ba�%�;��$O9D�dp��^�}��ݒ�U���pk�j"D��{R"�>*���A���iæ?D�x��	}p&8�?�~U��;D�� ���&?:֩��#C�p�b"O	��K̔��Y2(Qo58�"O(eR�Ȅ|d�a�^:������T�O�V�s`��x����"̠1���Hw"O����+�1{4��N�;I�ִb!"O�ř�9xː��a��	��Ih�"O"����*H�!J�O°{�8 "O\���̨:�F-�!��Wݘ�Q�"O��1q�ˁQQ~}�珖�Y����"Or%�j�=T�����Lʷy�(����A>Ap�mFg��	���U�u��)D��2g�"^~hPԁ�*M�jE��f-D���+�Sg�E��c�(}0���.D��֩��p&��ӄB�#$
����-D��z��Ь1�Y��F�c��D�4*O"M�t��DX,�y'͕"�=0��'�1O�� ���[�jM�����)�d�IS>�Xp-٩�N��B@ЋjR���B.D��aSe�U6 x ��?�4��!.D�X(5JLG��Y8&��q�^R��,D���� :x�y���ڗ4�"�+D��ᶪ߀K�N�GO��<�:"d(D�C��ˢJhj�y��Ct�� +D���PA�
e���1q�h��	$()ړ�0|����FQ両�2
�r!��N�<񄥛#��Ԡ��+G����P�]t�<!��m�&����ɨ �h�*t�<���N*]X��k���!dNQ0��s�<���"Z@�A-�(L ��PhWl�<)g��2G����ל@���Qu'�h�<�iI=Ɋ�ځo�2m_DmiRa_a�'�a�$���g��wbt�b�K_�b	.8�ȓ�� ��-�3Dl����	B|�p��C��H��-B)����!�<�J��� �d���1��G�D�.�"݅�)�H냪E�x��[���8<����ȓp��iI�n�/��ys��FbpA�ȓK�j�c&L�
B�����¬arn�D{��'�?٫%%֙��$���E�S�:}q��'D�X�oі\�
�D�6� �C'D� *�i�<}��m6EN`k����O$D�`��ő�t�E�Ŋ c���!0D��b��`��ʵmC�"��<��M��y2O�����+G+'��5����y��G"B>�أ�Z� �p��š���hON�b��ʿq��8`N>�^ �4Cן�y"��;��M��,�0�|������ya��X��oU&o.1R�G��yF��PeS��W�~di���&�y�C�*�I�q�HC��
VHZ�yҧ��4����H?��e|��S��%𧂅77�`"MD2k�f0D{�OѤɲe��k� ��	4��'1R`�� �4#�TS$c�!�z�<�Ď�z�C Gc�x��6͟r�<!3T]�Tz�ZKK�a�r$�H�<��9kTU;�(9ڊ`&��H�<qU��;;�`�"�Dr_����m�<�W)H�;��:�Xx�Shl�<9�O �SMj�����Na��]�<�f"W 
�*<Ȳ�ԗR+�k���X�<��jR�"#�|��/A-2�T%�C��<Ѧ!N%M\�z�Щ �t@0R�M�<t%ܴ
s�mj`a�9�IA���w�<� Z� ��B�H�тټ`�8 R�"O���Q�K�7n��@'o���P"O��(��B�c��6�ߪ!�(��&"OP�h���T�(۴�ΐ1Fd5��"O����ѫ(8$��d���6d�F"O��3v�^��]bg���E�3"O�dB�@�
�
�	QY��@�2"O",�V� !@|�2���^�&��"O����/.%��&�ʢ`p�i�"O��h6B �t`bux�-��W����d"Oz9)T�� ��0�d͉!��C�"Oܬ��Or�ꜣ�΂<f��m�"Oz�s��?�1��N�;E4�Aw"O|l�D%C���U��$�"�7"O
l9��J�ETxX"��~v��w"OA�耥e�]@�
�/��\�E"O8q�`	��l�GGʡ?�0 ��"O���]�
�*�Ɂ�J�򤜋"OB�*�$�Q�X�
3�0e�P���"O��#���d���w"�%ݾp�"Odق,�u��1��
Y4Z�q�"Or`�T��@|Ơ('/G#�q��"O��+Q��~M�uA��	��"OR�F*A�dר@�$S'x��)�"O"�;�O�&9@0��lTc��D�"O�ŹaeT�D���ŉ�Y�NP+�"O�h�5��rk�NU�McC"O���cG��	y��0��M+HU�U2�"O��RlF�\>�m͎*OD�9�"OP=a&%J-.��`��^�GARl"u"O؜"�LE�e��p��)ސn%r�E"O�%�dRpb��
�C,���"OJ	[p��k?,��R�J��Q��"O�q��Ӫ"�|�gF�	f���T"OZs��.&�zx�Ŏ����I�"O�	�M��(�y�B!t�H�G"Od}�1JB�H.q�ƥ�>a|h�"O�\sĞ�j��r�"P��Sr"Oa���T������?]�����9D��;���(h��9��+s�jA@-D�l%��hk�*��G'N�v#',D��SU⅊!�p����9U�4m��a(D��IU�F�A'��[V���=2"}��K'D���fBԘ[��Ś��K$��A
'D��  % �ng������5��qJ6�%D���d� �
���Cj$�1��&%D�`�!�(~L���fBƽ������"D�d��(�׈Y�6��4'�ri"�*3D����aA
z8.�xq��e�Z(� 2D�lbC�:N���qW�+U����p�+D���q,>t\&Y��$M��ɷ�%D�@����Oy�쀕��g��ڗ�$D��D�S�L� h{q�̓�hmi�d"D����w�a�O�;`�)���2D�`�E�h"�$Y6�3 "���=D��!���nˌ0� C	hTmZtf�<���?�M>����|�zt+�L�_�0 �a�=7��C�ə!��,�4��,_|��` �ϸMTC�	�Z �7ċ2,��y[��EeDC�I�="p ��ędV�QҗKΦ^�C�	�-zpچ`6$��0�˕j�C䉨V���ȷ��|�Z1;��L4u�FC�ɷ.����F��p�i�O�(P%Rʓ�?َ��)A�V��	B�J�:jP�csH"u!�� �p�g&J=D�� ��<[ܔ�A"Ol ��,K�y����g%ЍD�L�p "O�� E�Wb�е�ʰH�<Ÿ�"O���T2��c��8��+B"O�3FCo�,��%�����"O-�¯��gg�쁦"L�;����'�1ODjq�'��>]+���1�L�S噫?"N���i�<1cY�(�lI[V�(x������I^�<	�)��b��I���\P"$j�	U�<i6���V��Ӧ-����NN�<ل�Q
?��Ƈ�%~�U)�)�n�<�p��8�q�DӖT��O�l�<�$�>e��S�K�V�P%i��Jk�'�?�³,,P5�t@Q���twr�B4D�l��'P50,��st��:Y.q��=D��p�`D�B}$(3a͝lO��"(9D���Ņ�rB�y�� �0@t�,J$o8D���M��&`�)�����z��1D�l�U��7��H�ge����2D�|�t��5(ʪ��2HK�wex|��-5D���GJW�Z?��K�,3����1D���E�T�V���j[��$4D�l9A+@;��ҮZ�l
�\Zd=D��;Q(G:|(*�#Pʗ$m�<Z$-;D��:���4`�h\�#Gի K�2�.D���*ݜrID����ѩ� H:�+1ړ��<�Hu��C�|�MC�[�J`�w5D�P�6m ^��"n�,;$T���?D��Y�#г��@ţM��@PU�>D�Ⱥ���!ܦ���nħ�r��r�=D��ѥh���xXFnA�-f��u	<D��i��3j� e�GC ��0!�;D��p�J
o�����\��:�%�O����u�6�qNF��<�k19B䉰F�&����Y����P�A:V7�C䉺t���`�ʚ���A
��˓�0?��J^'< x�(@�2�Ak�<��,�*/��Da��26�B��e�<��eT���ٺL��h������~�<��!R�qS�e�sn��XD��Q�G�}y�)�''�4P���0�6`
�J �Ba�����#bɟ/eĨp���%ĺX�ȓ
�TaũsIVQ`��ة~.��ȓz >����of�}�#�_Ά��ȓ?��A�K	�L#QzA*�[j`��#��U��kN�a�z����w�R��ȓ7����Q���V�I�B�9�|��	@̓��
�\�p<�1࣊�0D����tށj��1]��#�Z�=��Ņ�W�Z(�E!����Ǆ�L`ԇ�,�=�C��	L�`T�W68���~r��� $?��T&��<��Ȅ�.��)I�&=\��(fjD�=�TQ��B~�y�PE��!���6�Ȗ'�'����y>=�͉s�萐#�R�zIQ��3��p����B����}���E"n�"\BP�&D��
E	�-��H�!A�6B��Z�m#D�����1�j<jE(L2ie�&D����AZ�4G�\8:�H�6�$D�䫲GUrA���p"�<HҰHHA�'D��a�b̽s5:`�V��b,r�ɑ�#|OP��!�ٮ!ܕa��B#�4e�|�Q�E{�O/�����}�Ja��f�~HX)��'	���pLJ�稜ʧc�4,FP���� �yC���"nF� �W:>�(1��"O�t��ڍAV]Ac�8%���	u"Ophȃ ř?@T��5 �h�c�"O���ԯS {PƜ���.���&�'��<i��N���Gnو	�va��<A�r�S�(%�;�B�	E	B��a(�iDXC�� ]��8��
�P"�pV��'�BC�	�~,�eȥ`Q�b����M� C�	N��p��b��Z� ˴��e��B�	�C>4��; �P=(s�	b�B�I+2�R�0���!�Fe�#Ǽ%����d7?�&Ć&,�aӠ!�Gc�!Xf��R�'a��힄I�*d���X7 fL0*(�y��ŷ/Yb���G���hOP��	��s*V,�f�4�ȌQ�(�t!���#:T��
��7��B��I�!��G4[_$���	��y��	���>LP!��1ؼ,!%�M��FT[��]`ў�'���|�eC*6���j��H#?e԰` I�U�<@)R�J���@K�Yv�Q�<Q�)Ln�]��c�]�`�6�MJ�<	HH?i�1��Z�=`�1��H@�<�&�'�͘��1>�I��!T���F�<N����`Cl��貑�7D����6���Q2d�8eX�$�� :���3��h��Vm6.2�|�R��)t�ڒO����K6Q��x� ��[��ڀ�(r!���2
��)H�R2�p7�{����H��6	q �I�`b�0{!�$�J��g9x���
�=O]!�DN��e�"�K�B�¡@�n�!��%��� Q.�o�F���@�S�!򤆿[�E�Ū���ʹs
j�!���i�tЛ�g۪?��l9�I?�!���w��'s��U@t(��^�џD��۟ �|2ECE����@6� �y��Q4oCc�<�v�9t�U��(���y�$�_�<�Vo��uZU3"��f����t��[�<��$�*,�ţ�G·y��i.�m��X�<�B�%Qч�/�ֱ�@��ry�)ʧ=9����\�J�D'
WƎ��b������3�n�@�������m�E��x`�i�I�����U�vC�Ɇ���%A�D��&"���FnJ�����ȓv��0�V�%!���F�Č'��]��u��sr�B?Jހ�S�֢Dq���I����<!�M$��1�Ĥv���,�Y�<�������'R�Rt�xw�	X�<1�G��U��M%�p�#wFR�'���'�1�F��gJ���)ꠌυZr6ySq"O�-�A�E�4�l !���eZ�][@"O%ZVB��4|���KJ7p�<��"OИcT��o�
�&�Īq/�ᨒ�'#�I�.��tYס���܍�0d�pm~��hO1�:�	9R�Re	ƀ�r9���`/��l�$�)�����ջR���h�ԥ"#��$(!򄒲
k��;��N�6��!�uM��[!�ο�J�k��S`�;�N�,]�!�dɛ�^ ��.�.O���V���!��Tw4��c؛u,2| ��P�!�d
�&�I��b��P�x�!�D.*p	�P�A
Aᲈ`�BT%8.:Y�Z����I�R[ę9� �4b��Yb2��z�B��3#��2��G�0���"˟�G$C�)� j���� 0<v�ӉR�aƞ���"O��q�aƭ|���0�D�~�d�Rq"O����U�/Q"��E�\�l���|�P��%�8�<� ̔n\bL�1ő�D��u�������&��L�&48Bm衤Z,$N<��ȓ}Ҍ p󥜐gt^���-�*A<���o��=�N�70ڀa$�E)HΊ@�ȓNz��z�݅~bB���̌�v΀$��)��T��8:���:��h�zx��.{�XQB)n8�Ш�dA	z��X̓)�8��]'3W���(ΦJ8L�ȓqʴ)���-��e;��A#=R���Iv $"��	�}S`��G��\�'_a~�F�' �ē���d��$�W���yr@�&	��<	��:�p�iW���y�LB�Jn\;wǭ��8��9�y�ş<|��P���˳m��]!r���yr.��2�墒LJ<i`(�ٔ�-�y�>e�Ŋ�]�ٰ����U��y��Ի)�}�B��(	���SU�:�yb+�?�I�R���,��}���P��yRd	׀��v��-�E
c���y�j�6]�� ���B<W�}�sՑ�y�@�|��8�":���)���y�;��H�%T+Gn��խܪ�y����� �$��bk���g�G��yb�P�%�,�	��<p"�U�&�yEݻPb��#�K�[K�Y�UM��y���zQ&pKJZ M���� ���yr����쐊1v�u���C�d��'H<	�*�.\��p�t�Q�m����'��*���"o�L�	�X�=�����'�p��(I��}Zү�h���s�'}ԩ[GcU0U�v0��ē�sYZ��ϓ�O�Iv�(�^��j�%u2 Q"OvhH��]�kYJ��uK��1�N���"OJ���$��`c�9�&,����`�q"O~D��F�j��\�v+]�"b 8k�"O�\��ɟ��ԑ ck��)��"OHBw�ěQ.dpC�J&N���[�"O���@C��Z���(�1��'�b�'���똼�5�>�@��S��Rm!�D�!�(53`���K|��rJ��[[!�d�R@��9SeS�&4���E�J�bQ!��245�Q��n�	,x�L�ŋ>:A�O���D�a���œ�9�NIs�ي�yo�kpd���KG6|�Я�f�6�$�<I5�����f���HV��J�l�Feɽ��m�ȓ���(��)G�5��iV J��ȓ,:��cM�BaC�ԇHe4}��H�&��e��[�U�$���|c���#�^8��
�h���M�� d�?���?����ƣ~�4���4:9n�2�\�4k!���,Unu��K(8|3��S�}Z�2Oެ@s�|���M�Ҏ��pFƍWhAcB�l�\C�	�kD����E�U��Se뇑g�:C�I$9�����@�Y���
2�h{fC�I+*S����*ip�Ѡ���FH4C�I�+c�q1���6�l-��웣L�,�4�'E?	9���/�X|(�ԲXkji{�(<D������!z@b�N��t���;D�� BLI�S���R�a�th�gA:��/�S�'R�(<`0��v)�U��ՆgB�T��M��aK�S/i�P)vd� ��D��S�? r`�MJ?06
H��!׃v�>��"Or�;7 �L�� �-�´�r���O���2�'m��q�]������/ήP;�4��L!J�А��E=8�"�' �TȄ�W�jܲ&�ærV�l
gHnA�Є�m̓U�v����gdP�! �L	Zn̰��
x&`"&��y|h���O�kM|��*�ఁ�NF!f�ʵ��f����q!q���2_L���JT�X���ȓ�<���N�+�6衑L%G
���?)���0<�s,�5+�$��ϙ��
��ě{�<���U1#�Nc%瞝�Up'/�R��`��N~BoL�:����H�;n�<j �];�yB��A� �s�5��t�B3�y�/K�zI>��F�.:Y�M���؀�y"�NSX(����pH�B ǚ�y2��&�U���q�E�e��?���p���ѕO��m�å�5�f��3B+��0|jri�V�h���G�jA�T�<�@�G<	K�s��u$ޜ�6��L�<y��_�C���"JԼv^N��c�O�<��a�O54Ѣ�a5�p|��)Nr�<�ƃO�Qa1G�+�H8���H�<1 G
	��q�*
0k� ��#N̟�E{��)J�j���"ڥ`D2����M��C䉚*�� �	������B�I.1�Yr�L�B�
���@�<�B� W��qQȴP�� Xe�ހA��B�	�%[�RRGK71������^/ ��B�ɗ!J��Qd\�M���J��dwJC䉃08D͋��Z"zAta���>8�vC����U1)J�Fo����L p
bC䉕B_���B��șp��X�kNC䉴Yn�e[lt����a��5vB�	8��#҇�� ��l:�,E<B�	���ibMG�SܮLx#�ڷ
�C�I�H~ɇM�\�)���)�NB�=\�����Y\R�����C�B�� (9ణ�*��8|&@ەg�
8�B�	,Oh���JV�*�<�r�ܡ~��C�	�)(u��gSB BD��%��C�	Z�6�;`-�5	�0��]���C�ɀ����ؽW~�P��L��7��C�	/��&n�"�X�K�g8��B�	01O�fVx`�y�7ĳ�B�I5Y�ȣ&	�C0��cO�-tb�?�����Q��J%!p,l��E��'x���"OA �Z�a�����DjD�w"O�ȡ�C�*��E��$�%Nɦ`$"O"��w�*kna��b��&�l��7"OB� v�]�9���a�|��8*r"O�a�$P�s칻��3�8}�"O������C�&s����M������a�OP��Z/��%��2seK�v��E �'l(�y6��ir���B�5\y�4x�'%���h�#PĖ���K�>*j c�'��X���@;P�3I�%��9�'� � ��çQ$���B��5[Hhb�'1:u(&�S�b��%S�e�%�\���'�z$K���q-Dy"t��$l�Y�'����(l ��P�_�B���'�N�$n' �&8m`�p�'q�mb�P%<e:����&g#\�'��t�����R� �3�eƩ/�.�p��� ��6��]� {5)N	 �.�G"O>��D�NlS��v�6I�r�Ұ"O��g��0G��0�O
�܍"Ox�t���� ZSk��
��"O��Bu�B6dց
Dd�1��d�t�<���H3:-La�)�T���%Ft�<9Ǩ5jC� c��j�.��Tk�<чc]�[؜2�,�7[Lx(�(�R�<���B�~ٚ���<��Q�M�<��E+F��  �ؐ-g�D�$�D�<���x@Sb��{��ԂtBID�<�#L��t���1gѓ::-C!}�<��Ak"y�D%Qr���{�<��0κLp���rrbq�1́y�<QF�żBV���!�>Jl�gd�\�<٤�GB@#�C�P 4#T�U�<Ie�1$����qdN�.���ҁT�<Y�H^i���^�z��UR�O�<)��}��ȧ���,�8i�N�<��E
kn)	$�܇`�0�Y7L�J�<-�i�H@��#��5�ʡ�
D�<	sJ36$	��I�j�A�<��'֐���#�o�B^�b,�g�<�sg�8OE�)֏^�L$*%�C�o�<	�A9#kj8��!aY��c�o�g�<�BMP�b��*pf�!>".d���M�<��(��U�Y�3����3��D�<Y�"P7����qdJ?��HR��i�<��(O�y�3M��q�W�K�<y��F�ɒ�/�tI@���BI�<��`�n�bK�D��!�p:`�]C�<��GI�j�挀�J
�.��42`�{�<���5�^E�"\�V���i�ɃN�<)��6O�}�VH�;4)�$I1)�a�<�-�kj����ӎ�HJs�<��DLF1�.Éh~̻!�Mp�<�g+G�Q��4:R,�]}Z<�lVh�<��BA�)�TQ�MQ����#ro�z�<A�E��T)�-"��T<1�.�r�<�&E3Md�5y����^lD�(�l�r�<�f��_�,K�AF�:X��G�l�<9f��4zM3S�׼E��% ̓b�<��Ù;��2�o߂LyT����v�<)6"K�-��r �<e��IpC"�u�<��
m�p�H�gR��!�}�<�᭞�`�p4)��_#C�E�0�v�<�C�M!C�L:�ˀ����H�r�<Y�������e@�J��扂i�<�t�AG�%�	Ҷ'��وV)�a�<��ܛ_)��pddE�e@l��&�I�<��Z��f�����+	��H��M[�<Q1W�o���
� �����W�<i��B6OM������w�Yyt�R�<1��S�L	��� ܮ)��H�GK�L�<����,6�q�`N,R�9���I�<� �	v�����ۤv���'�I�<�P�ם:���%��ecT89R�B�<iE)�  Мeʄ��$mBF*@{�<��F��" �����Vd2#��O�<!@�G����'�[�ԭ�|,!�D%j�H��D�x���؃��:n{!��C�DDx��0'��� 傱I�Dw!�$M�)�6�҃m�-@����G���g�!�D%=��% Y�r�dRw"�`�!�� ��p-=`�j����P1y��@$"O&�{!cȯ_t���e)6��h�W"O2�	C�	 ��=��S�\��	�R"O���r/��Da������wמp�"O�pJ���Z�H��Ҁ ��8�"O�A�g��eI�I�BW9e� �0"Oh:�A�)y"���dAC%QE2���"O���`MI~��Bc�/4A�RG"ON`Y��޼7ʄ�S0K/+�9�"OFmc�K�R?��V�\8.6���"O�y��L=�����̮<3�Q9�"O ����V�$66 �r�F���"Ol�(ƀ�N!T�z���;T���"Oذ!�
^5Td�*$.��%[�"O2ԫ�*ʐ"	�% g�9+iJ1��"OЍ���8-MH�4�ˤ`�B�"O�ˁ'�,�`�K5^(�0"O� 2�D[�/��p�6-,N��I�"OJ<zpF��̴B`Jʔo7�rp"O�M����-F|Ha�Gꝩc}m��"OlP
���67pL��c[��Uz�"O�8j�LA�6,�Y�r��?�R�i�"O�+��]-"���I@$ɢP�@�B�"O��ۻ&��`���;h����w"O�1�'�z����|`){�"Oz�{1���x*��W�wQ��Q"O��ʤ
�*O���(!���3$�5�"OV�b%�L� �r
W�w$��"OP�����3ҼQ ��)j$����"O����̰58E��.]�)r"O�+�m��,���Hc�Թ  �R"O	M��pٶ��G'�k\�@�w"O�8�(N�h�,8c%DG���"O�`# ?:#t};A�I3*��iT"O0�8�#L)L��AXA�>_0!z�"O$�Y5�ߘO�������u<�XA"O�2 
��Cj�D�4��1w��"O�|��o�C+���q�ܒ�B��"O8e��!��8��`�?N�l�C�"Oΰ�0��j�N�{��6:���"O���C��|�L�)�H�<&�C3"Ozu���S	5��S'� %*�"OM��ƛ�tE�  �Ɩq�<�c"O2�(� H�`�ޜ�ec �P�9j "O4cv�\�<�t��B��!��e�"O�@�1�%��A�5"S37R09R�"O����*E<��XHt��92��� "O��k��Ν7�eГ��(`�Lg"O4H�ec�,'�F�U��'mZT�e"O\	���}=�8��H�z�P��"O"$��Ȕ�t���S��, Ү�s�"O
��G��A fy��X�5�,(PD"Of�0W.ա�(�Hѐ;�� P"Ob��"��@�f��&��@�:��"O.���bHs��o
�l���"O��I ;;����=Z␛�"O\�P���j�"$0d,�i�M(�"O��!a�rV���Q"xi��"O�yrA�ǚ��� �	ܝif��Q"Oi���*.j�Xڧjי_(��ɡ"O@���<&x���f^?N h="O ��u@1���2� �qlx5��"O(��/Px5f�P�akP�|
�"O��9����[ԪPAQ�}�B���"O� �<��c�$Ȉ���W5<��]�"OzC��h�@� ��Z�3w���7"O�t�dJ�K�`�0�[!=[����"O�kc	O�NKZ-�fM�~DrEw"O�)Q,I	>�
u9��B�a�<{B"O�m�+:fڮL
�ӸfԂ��"O$�;���"�j�c�0���T"O:=q��֣Kc����I��§"O�phh�R�8�7a=[�HQ��"O�Ё�
E�D�r�O@<�A�#"O�I13JӼ��]�W�.���c"OT!�*9Ұ��"�.] C6"O��C�O��\�x-� aL�+Z�a�"O��)R��S���c��
MH=`D"O@i:@) Q�m�D@ZL��qA"O
8)�#D�|�Dl3���5oaz�"Ov�ɀ`�Bd!��.OiV���"Ot���˂Ja��Ο:QT�:�"O~��sa����sM��8T��"O�$j5�A
Ǝ\�1掵�P��2"O(� 3��!	����#�_/PWhd�"Ot�@�n�X����W=|FZE@�"O�������q��^.�AK�"Oa� �' К���.F���q"O:	�$E��|������HT*��"O|�i ��]^��j�^����V"O�H���^{�n�2ՠ�'�b|�"Ohz��5�*�R3O���Ќ�v"O�`;#@�T]��b����"O�L��x��p�P$����`A"O����
�* ���+�� ��x��"O8��㗾$t��rbD$hf�ó"OF���S��q��ӓjs�}Zf"O�s�I �E̎L�4NC4N���(d"O�p��!E"$��I�k�� 0&"O��5���i�"H8���ASv��t"O�%�Ga�@�X ��5t皡��"O��0�c	� #�ʠe�r�찛�"O���7e�KĔ��%&V�?����"O�)ؠ�Ո/H�����H�.$�"O|���,S�{`��G	M�@"O��TY�9T��C�Ґ�R!"O��
���e��\k�lRD�h3Q"O��`S�ϼ���3a�ìE�~3"O�ę���'>M´�U
c�^�#�"O��g$���rt�ƩX@�h@Ȥ"O��A�B�1�\��%2kL\Q�"O��JՄ�_��!Ӫ�="�ބ�"O�pS��1:��H�j����a5"On��!jڻj��R�h�&G�����"O��<&� �1	��o��3�%ɤ�y�),p��K��92du����y�S ���M5]��2B���y��3�t+v-D�M�������y�NGm������Ƚad�$K��bN>����#D�c�٨zI�p�E'��KG��"D��1�R>g�Z����Ϳ"���$D����c�" |F�q �J�\_�:c!"D�$3�ܻ&8���#�����!q�;D�Hە<7��xk�.
p��q�PJ:D�@� ��*����Ulw�sN6D�c�ۺp$<�THշZ�wB4D�4"鎽V�,�*�H�	B�Y�c�-D��Y�M֝B���QcN�&z�u�g 
F������ �MQ��������"�r��4"O:�2�ʁ<� �4E�I�(��V�'�ў"~bE��x�\d W"�
��)�ud���0>�O>!�˓|z)@%O-M�!kňu���'�����ա4���Y���R	8D����R&Z�l�2�L�l`¨ �`7D��ѯ�t��P�
�2'7���3�$<�S�'&RliRc"s@\h�A��v�$�����s�T;rEU3D���阦u��R��:D�Që�08� p�5�.,�ޙY�<D�T"T�}`l�9"�߭'���#;񤥟l�e前��	Ղl3���d��o�d�Qvk
9�!��sք@�K�*�z�9
�y��c�1 �)�i$g�dc��y�TB�#�w��y��	.}E`��o�"�ɃC���2C�I�A��:�N�nQPd�r��3QyZ�O �=�}����`��ؘ�KՑh�)��f�<�WA�0��$1]� qЍ�|?���'>�I�<Y����~�ņң��с��#=
ny*֤�{8�$���<���li�c��]��@����v�<1$�K� Ԁ��f���H.ɹ�%�m�'fb���)3�6)����9�5BdŞ�0;�7�0}R�>%>c�d:A-����×s �D���Z���<E���x@�A��!�"R`�8���N�EՐ���HJ z�j]|c��
�a�{��l۟@S�"�"��){T���|ZI�� �N���V~�rG/�U��Xbu��<iL]��|$Е����2�� ��c�v�YG��S�=��탒kX aʍ'��(h���)�� !4�TK� ��zz�y��\�t�����1�PI�q$V*f���t�ܾB�I9�d�÷!��X&r1�׮�/P"=��'�1Ot�M��DB�*լ�Dp2�.���t�ȓ�2`��N�x��Q͉xP��ȓ/���bO�,vL��QF�$��+�	"cե�\��7&;�2Y�ȓp��ل�$/�6�C���!#\܄ȓXbt)�&Ƒ5�ԭ@�*+���a�VղP�E�$xĥ�,�~y��	1��1&�6TB\}`d��-r����ȓR)^��`b%e��8�b�r���ȓB��0r��-(|0 ��>0�J��ȓT���� ʕ&���T>h� �$����I6\H	h��� uh���#)�C�	zkN���A�/E���G����C�	�S�b�{e����8����8$���*���'�a{bE�01���b�Q#H4|<�u��X�<	E�� �����N���l[T�<�b�S�Ҥ`�]���Y�Ԥ�M؟,�B�8@"�]�I��YPƆ
��PI�?�ӓK2�0Xe'�O�:�3RF�=1�j��ȓ�, ��
Ã���(�É�	��Ѕȓ�taH$2I�P���Ңo.��ȓ6�tP����=ڎ�  ��9�"���	�'b0��,;r����Ssq���ڴ�Px� �}��I�-^�0��)�G��yRO���:p¡�½)�����I[���'��{RŞ rCB|qg.@Y"��y�VI�  �牡,r�9`���y���#V�����m?h;$�{G�I�Of��hO mC�m��4��EP�f�J��U�b"O��;��&,��U[�C G��\"3"O>Ȓ$l'u2"\2$" ��ph��'R��C�C<���0$=$x���� P*T��'��'�d#}֧� �$:�^%P�΄��ˡIF��4�'�������$Y	�*�#����L
4�6D��T���<��t��mf�p%C2ړ�0<��A�F���'�(zZ �!*�}�<�7�B"T*�8��E��(4�)4�ߦ�H�^�4��IP��ĸ� ?����$Q�=�C䉬,Ѵ�J�-\�/3Xy΄5��b�����3�N�5Y��q ��0
��B�ə�X+��֡P��)P�*�p�.���d���A��Q�_�T/��`g8OB�O�ʓ��Y�p���+{P����=ZJ�I�ȓg���LCs^خ;�P��%�	�HO�O�����/߹vTҘ���M/{�Bei�qo��S� <�ĭE����H@(� =�ȋ "Ov�t酱;��iQM�=cy��"Ol�	1�1K*��3�T�ʠ� �'j!�dݾA�h��Q�E�y� (91�@!��Ĳ'�S�vkp����L<*xt #�C�	�j�x�Aa���s6��~���I���I�)�L<��8om�4��mΞ�Z����k�<�`�C:yV�A	\{,���p}r�)ҧZ]R`)�ݎ#@���%&Ϊ��ȓ;. 0��X|��@ץ;��ȓBl����c٪{�Y0�'�
$��iܓ��쑅�1��0��HNM����ȓN��ѵ`���ǌ�]q:��ȓH�Ȗ�ߞ%��̑�-r��	�ē�q�qC�K�|xk�脠(�hr��ii���J�����l�|* I�o�!��D�<�JXkB��"_�1�n]0s!�B5	��H��焒%B��AC��/c�	]�'Q�d�=�FL�y~$���P
T����R��P�>�ь�2���.�\2�p灉V�<��b��I���[@���҄�&�JV�<a��OsO�p�Gڕ2$�A�*�Y}S�����V)����� _޾=�$�ɬoh�B䉒+�9+���y褥ӶJ	�~�������|�w�W6"$�R(Y�+lP	�2⓵�p�2���H{��P눐Z�Bԙ�"O
X��,�)�N��Y�Y��"Oz���FM�>oa�ר�YL��"�IU�����{k&�17�^�AUH豱C�����'扛�H���!H�z�R &$����`� ^�dB�	1bz0���b��?GX�V#U�Y��B��.������L�#a2)A��M�)ZΒO>�=��y�ŋ�!.�!с�L��l�b��0?�(OX�9p�T;u4�룮��N�x"O��C��"IB�����bH�`�"O����ʏ	���%��,:��"O��b�)�+">,�2���$�|-K"O`E��T�p���6��lҐ1�"O� ����kx�����"8�2s"O.�˵'��m���'�*��"O�a���q�]� �N(>�ZY$"O�JJ�1д�n��D�e"O�Y���֙*kP�����"d"Oh=��(E�i��}�`���_���ɶ"O���6�R�h2z���B��V�6|k�"O(ʰ���eHLS�֕nO��C"O���bOƸ�T� &!\?�P'"Of=����B��d��8��p�"OR(�&*�C�0��ah֙l��"O��aE�S�z���"���.:�"O�``���:����&*
����"O� ��֥ѶE$@(��D~Ԙ��"O
9�Aj�Ef>��c��6R��4"O&|G(S~>��RDö9l���"O�HqS��}^��[�-�FP�"O*Y�1��,*��U薏��X��"O������]�ڠ�M��"i�U"O�$�#�I�V�X]�5�O{'�m�2"O�Łp��)5(�S��~��
�"O�
 o�6M�2��M�1QI��R"Ov��!]Cxe(W�J'��(�"O*�P��M�8r4�aGF#0�<�+a"O����#�*� b'	#a��k6"Or��G�!�j��唎s0�,�@"O���4Af,[!"S(O	6@��"O��j�g� !���)v�?	�Ub2"O>er��ޘL�0�CW��# d�"Oz���v6,�JLG���X�"O��B��+�譲��N)b|�R�"O� ���I�rӂy��X�H����"OrM��
�
զ��.Y�t{*��@"O)�*J)^z��pCJ8D�r"O��ٳ�OH0����.U���F�0iz�H:�>�t`Š91O|Be,�4M�b�{��(z��eۅ"O���%Z!rc<|�rm���*Z�"O�ʦ��L���#!�7?8	�B"O��q�<H[�Ɉ�#�n�Qt"OzX�D�[�o=`�{�ݔP�\�`"O�8Q��6!]��R���J���"O �jԡپ8��ܣu`��0���J�"O�ݚw��=)Z��V.�|~���"O��d�S)���@l�?(%��6"Of�J����7�̱8,ԏJl�j�"OL8@+�
[@�@�I1t�e��"O�1�ƈ/d)���.0r��5"O0<��e����@mZ�}#"O���e��#cD���I^��c�"OpT�Aȼ5?�}���x.� `R"O+��J5x�B�-I.�T �Q��K�<�%J%9j��5T�y��	���h�<�U߸ry���Uqjeia�g�<���	�e؞<�@�
4��<ᒮFE�<A�����z�nT<K�t}ؖ|�<��!**�*�;2�Y��AQP�<�e(�)s��K�lD�.d|<�E/�_�p�G�9d�a}B�L'M� ]�@��3[�n@SW�J��<�`��Z�hLKg�ʖ�y�e�22��/�I��H+Sf�<1cJ�*9f騔�V'"����Z�	�OG�q�ǉ�6cD�J5�S(��@�-�	y�搸��?7bC��cK�Y�G�2��4zp6D�L�	�$�"}�y!�Vqk$,4�3���j[2չ���Y���CC[��B�k_F� ������"̺u'n(;Ʃ�
V!>HЁOZ�o(Ĥ���cA 1`"b�
]Th0�'&ꮣ>9D҃'&���� F�.T"�N�b@ �����Z�����M̏^�uq��/D��R��I<��	J���"
����F*D�P�s��!9��i��eƀ$N	�=��O>Ҡͻi����7)!(Wh ̎bRXɆƓI޸ G��m���0V�O�>�zy:`Ex�m�
a��<�C�V%Kڴ84'Q�l���=�W@�r�$��dvאNS�a���'ry*b#��|ۀ�Y=�y��nK���(R.ӒJ�LU���y�iX�'�<9�4��%i���[�<OZ<( � {9V��Ň�"�:A3�>1���)B>i:��T� �Q�oF�v��ے��%%`H�`p �&^���*%j܋&�d#[`�#�b �I�zfP ��˒<X��>M �f��2�t@S�c]�`xl1`#�$g(�ê�7�	0�fF2�eHr��3��S�18��?�}ra��5%|�m3�-���uQ1�ڦ�H{��^���dEx��M��IŨd�P��,ģ�����;u�9!&i� �^b�@�9#��c��g�B%� �!	�➘xJY</I��'-v�gC�	7�����D���h��@�<?��E	���@!�oy(C�2��� ��"5��-A����v�;$!R%!1�X.T��Rψ�kX�K2b���'��]P�H�PAXP �k�u�\sU;A��%�E�J�|��'�s��J�
��Ո!�\�e�����3	�t�0I���ם내��@�O�\��-ӹ�<��N�;|��� k�:��g�⒨�� Yz���\�W����L)h�3+ 0<���g�
/��(�4��9�,���K�|��BnπM+jʧ)�r�YBJ�˴⁑4+fʛ��d�(���d&5S�jzu�ϓ{/�@	���M��~3剃 )*�S�ˁ2j~�Р/(��)�:4��v�ƌ��Ң�����k�1llܠ�@��.�1��	A��M�f�I9=�|�5,��n�:Esg�=l%��sc��Y�d�F�4��/Uv�QO[2J���� � M�mx��à8��9�dM��6�E�re.��#K�BN��	�o²jP�]��!?���d̜�(8�&�i��8{f��s�h6 [N]9�Z��n2(]4d�o'�!hͻf>jD��c�FJ:`�O�F�3�CL��}I*R$���,;F5�H����,Q��H��\�cD�4��jrQ���	¼;@�;��� �>$!�b⮇�oT�Ӂ��NP����*!�f8(P���D�VD��h`�L�t�=���2�kD&�E8萪O��6,"0��<��G
͊��ǆX=d��-
+O*<��X�?�R|����nx�t��LZ�J��JD��9��ɶȪi�tnX0;�BX�Q �iq�X�Q��M����Jݎ}�`ahEϑ���� �	N���ň�HR�1� /� ���	��	Z�A_26�	D�9�5����!%��'���|=�s���v/�L0��0�n,�W#@�A��	7B�')�)����z1�3$�ϐu)�@ "�S"����\�t���30���ɹ�D���$%�,Q3@*q�z�����~� a㺍K&K�1"��Q2��ܶ@�H4x��a��5sb*�&��}�mDe䰝Sk~>Y*�,ܴE�R����UP�g�L���:�$^1O:tA��}T1�tOY+M�q9�#���y^�6-	R�$1�4�%;	|�
wK_1�d0�G���KTX�3 V(u��930� y4ۄ �'=j�Z�y��U�Rش�@�L�F�L�2 �'�^3�-ۏu������xuZa�'ڶ�x��Q<B�X�R�-�%�D��h�˅
E�Dq���S�����Z 8�T�U�{�<�5?���O�@E�w����Fn�G���+AI�2�`H��>�%e_0
O~�1��A90�ICg�Ǡ]Z�	� ��P����C]7s�Z88��ʹgO�,0�de���:�"O�)��E	_m M��	��^�H@Y�o\�ZT����ѧI���5��P�������u'	'&v%q����+��<U�^�3M�Z��q��|��ytoD�'���z6�V?�R��')ٹ}���Ȩe�n����-z�����(]	��:��׽	�Dܲ��@9ES0�A�.�J�y�h�i\�8��ʇ2ጩ�5P:�
�*�-Jt���H�!�; :�ۗ��O�8F�w��S ��y�z���sx��q����Z"�$"P@� DR��6"c��ubM�B9�%L3l+"�9w��=_(��`�A^�<��47�RP1B�G l�rj�<i6@a1�$�:��x�L�pL��/vu�lA��	�n$��$�&Z�������X�vB��H�~Xҥ쏮u}�@)qNȖ�yW�
4�tx���J���cT	�F��dBX��q�#͹��3��:Xn���&dўjhԜ� �=D⚨�L�jK��&ƌ������8]e��%�lX�*�$S��sÀ2Y^��g`-��X��0�1|cXVk�����`N�,;$���c�ȍBڞ-�$��2}�Z��3�Z�:���@tM�Kڐ8˷�I�?!���pC�O������v���
�Έ
u4,�t�	+t�`	OY.4h���ǂ�H�������s��j&ϋ}:8s&+F�<$ r���{�h4 �JШf�ўĚ1B���p�F������,"��#��9���r��;H�I�3�<��#�� �S��A	!���p��:�ļR�*�B�@����1���b��0ud�4xEi�����;OKU��U����?���"/ѱwa�$`eIyݡ��C�)���s&�m����:�$D��Bæ!p���W����lyP0X �M0���+
�My�OH%Z ���
�����A�@`��@�#W̈p	^.�\D�ڑLN)B0��	��蒉AAb�9�T�� X� �Va�'A!�EDPXU��dM!o�d��@HHhD�U�'VZA��dL#kjm�'�G;��c
A�N>����WJ|�HdcM�g�
�$�H�vQ�'h�9U���C���'I;H�I����O�b�8`d�P���<��	�K�a�돔J�p�h�D!S�����*�OE�@�$\�z��U2��t��4d��O������!Б�q�GOF�\�T�y��A��#������L�8egʫuV P�rmnӂ]
��� ��`N�/_��uY'&�@��OU�\����ZٌAb��+>���%�N�x��@��,Y�?�ʃ�ߡ[%�ر�8���y�#���'h��9w1Ol=��
$��QG��}������'tրR���wcP��`ʙ_~@2'��&
�ƀ�{��Y ŗ���R�G�"H���q�H&Q%�1�C剫!p:<�d�_*ĊlE�	}��p)"�����i#�D�$��a!OX)b�T���4dF(y����m��aףM�As��!dH�|ʲxِ�Ѧx�Ā����*~��O�Y˨�,6��"=��'Bg�0�QN�Kp�"C@�os>X6A�9l���"/ۥx��JSC'Ekµ��X ,�En�1@kt@д(�Ox#��4M��)[FƅO��W�Ё����+/q�i(K��_t�6�ԺRq�1+U��5�z�`C��X�SŇ��RW�l� *
5��	A��;M)�T�V�O*���M�Ukb|���ş@��b3Nt�1ufǥO*�TD|�H��4IXX���<QDҁR��9S�p��4=D6�Ed]�B���35��2BL|��DR=UMƩT�:R�r6C�e�YB�b��>��H�f��*�kѦؤ+�y"��:�+Q�% �5�`��N��h� ��="y�Q�����9�t	M$Z��� �R'�-� �YI��\°�'(a�� ֐+�0`aC�^�H)��G;�ў��d�8(�]��D�,^����(�n�D�֫���AΔP�P+� O�`�:�+�٦͑�Bh��,U"xpc�M�-�$�a!1��MB�I�3\��袎	9?zY�E�`�<�ʎ
,�3#�&Y�Xb��Ĳ^��Ȓ.ɚ:8ty�ū��w�L�pC��>r� F��088�qG��7����1 ���y@���a�x����$E��]�@��t�4ݺ@�I�q�F�;�Q�?�a@�N�-�P��<�I�S \u�2њ �Hu�X�o��Z�!��;_�������>~�%�E��+�a|bI,k����kf\��`# Lݕ3[�A�@5\1B�9��7 ��]!�Z�wxt�#T�b�p30,�3X�qG�Ƿ߀ j,Q4��KH��!`��1���'����g_�@�h)�'��0�wa
�>��W�	V��`h޴G�>h	����[��yr����ȱa�C1z�5���]'�~����O���fk̾Un���D�Y�vt;t�|�ĆX�r|+d�>Y7�Z�z��C�z�|�#0S�zB\��ڲ�2�ed�b>u�w�ĥNԠ9C��QG"�pF�zFP�T�$y!�m%6eJ= �A�0aۓ�|�̩@�6q�� X#e�N}2æU�`�ȐD�S�>�2�MV<��@R�������݆~�li�	H%v^իQ�)+�azrkʘPZu�r��QX�� �.a���1%��5*��]Kua�	s2��ʚTRU�J߷SV���gB-`���5�Y�tL��b�e��!>ph��J��Px�l�:4�(#$�#�v5��Β<{W�5rS�
�1M�T)����>�ˇ�!3�DO'�n�7N>P�9bsaJ-,�:jM)H(4�VӺl:����(4�,��@�[3H��X�J���X�ڈM�Z��IW6}�<�/��S����8v�nI����#��hU�O�J�Kg�6��\(v�P�(7iD'S�Lx��'X����O�<���iβ�Ce�)�2��ʓ�N��$���:V��0e�"�@�[��Uc�Ȥj��W\�JA��=c�NW��3��y���d����"�5D��\⃊	.rz�v�(��lD+�&>���ra�)b�����H�6B��x��
��vb�R�N��O�ĴsV����\Y` ťq���.�L�>���C�P��=9A�ؠc6�0�>�>l�j���	*�a��0�ہHB�W��i�i�#e"�9`�B����H�M�!*ذ�/��I�,�Ódk�a�{��y�ŁY?A}P�3�ϣn�}�D�&&�P �Ճ���D��;h��4���@�n 'D�.��/	"H@�'��u�X�3��҄!T4E�p=��Obx��	�*m����-����%�%�^�:���h�,B�.�딏i6@�1HV#c�|�@�'ި	�^٬��d$�u�٤\!���n��"`�< pR�Hו*>���@(�^<�c��� �n]�q�:j� �Z�i8P��V�+:��F�*���W�W��]� B�@��������q��L']��PDʧ	�J��@�'b�@B��̾@�t�'N���D�ʛ{�T��aګqXD�䌛K`p��v����b�\i�l�1�%�Z��v)�m��& X�1C �J��bH1���]LjEZ�f���z mF�6z�e��&pc��K �nhyS�d�|���ZWk������ʍ$F�9 \!%�U�$O����ڹP�zIB#��T�\�1�I"}�UxQ�:�'��$lȞ|8dJˏkDੲ�פxw<@Ҧ�)�C�����ad�Z(��Ȇ�cMZ9�0��%S:\J�ţ?�`t{V�����9���&�V4�sȇ�gGB��LN�!V6@r�>�d���O��d�1��H�@ ��	 a�b���/����Q�C�+����F�9J H��Ua5<�����fi|�C G�H�Y�#����R 0^, do�d=2do�G$9#$n�)h��X�ǪN#l�N�P"Ѳ@����.O�q�JI�5��RU���O+b��aMB?x@���S�����B)�6лg�A�(�,��p��I$x���MC}�n  ��C�#�<0Ja Q/f;8��I[?4
�(â�b�#�	d6�%��!%�("���c26���� B��!iKD&PZ׫),)H�z��2���hTbE�t��#<�n��QPB��u��f#v���	�7;�,�cwς�06	"%BG;��I��jC:s�:8Sc��W*`����5>�6����23<
EB�8�����Ɓ�v=p7�[2u���}�L�ohMzF�F� @`��iޛv����$ @�	�b��C�1o�B�9��:	�����(7���.T`ܸ�S���
�l�2\�i�X�i�����y���D��yzf��W�n�V�30`�	�-�$blk�8Z��z�L�iY[����BG��ch� �q�|X!2�(��胉+e�uGN����%�`#�|�*����u�d9j���#5ƒO���0N��ȃaa1o�1@���	�t �WJ?�9��Yw��Ɓ��aܰe��n��D�[��ÊO�_�~�r���&�V�C�D�>� ���5U���<��OF�1_�����4�U��E^�x�V��V�'4�T� %;]��w�ĸk�ze��c�7Y�}��e���L���+��
?�d���9\�ݩ�л5�j�H�J*���E�]�)��q%���#U�8!bZ�ɱ�n�..�l���D�:m�Dx���\^Ų���-J档���Dr͠�ő�(�x��^;n�Jd �@V_V�̒V�ʇiUv�ub��р=R�4)e�ȣz�B� �'$�-���MR��I�?5I���*`�������L,�I',�4{���
��̑��݅r��I��<m����O@O$�iH��6~�OTq��D��f<�8�F&P�z\�hZDT[Gd� փ��mmE���H&gFPy����d6�ӶƑ�z^�pRF��ZF��)J12uLd���9׶�����
7��<s�g�Y�:�#_ܓz~ȩ��>SX���	\�%n �V��@dr�e��?���bbf�h�tYS�!��4\L�҃�ܭ'c�&o�6@T:#�U�:���Jҩͩ+Ӻ<j��>:��x��%d���8[�R3Lk@A��e��!��鑱E�0cb0	��F��H���1�\�B��Q�L}�t� HI�}:.��-�Pf�D��5��l��0���"�(�n�H�`93���2���eJ�Y��a���ֲq�	�j�;_��%�ܕM�p%�!�9�L��JINL\��f.6p�c�5��L�d$ �,��[�b%?���j�ONX���.�$яb.jx"�CU��(�Gj^�E��xV"%V,�a�����rdڟ>��AN*A|�ɩE<��h.$@��� r�P;�(�0���5�]2D�^�#@^p)����HOa�⃞�M�b��o�� UBə&�"�11�1H#|�q�U/��Q"�R���F>>^�0�扽HdDX��^@Y3��ٌ{��ⓢɺ�����'���X�n�zp��2%���;B�X���P{� �b/nr�ݥO� 1 �_���C'��j��XD���Θ8Y��r&�<G�z\�΀̸'<*��S��'r����@U�ORV��)-�`�G�-6a�6E��qr���RP�h��Iv�g�dO3gF� �� V%��]a�LjZ�$[6�J3,
d�X*O�aE��O2�Ð�F(��a�IC�����"O.���ɕ�&��iC"E�#:ƽY��'�X�p��	7&V ��I3>n�!��.S�r����g���n=��D�	Gx��0��� ���)C*eNވ An��jun�RC"O훳��-\��Dˑ8�"O2I�S�F�\� ��m�.	h�14"OXA��]�n��,ÂkĕF
J%S�"Oz��G)�0G��U��ʓ!��P'"OX1A#���rr����càZ�&�3�"O�D��&/�(����7��1"Oj� Ư�,2Z={҂�L�Ќ@A"O<�p�N�W��q�ҽY� 0��"O̕	Ѡ����BjY�4��3b"O<����P��4�R�sv���"O������ȡ;E��ej��aB"O��X���rb��(@.K.6�\�:q"OR��cS'\�#���Y���3�"O�����*8�W�A ~�J���"O�Y�`4i�U��c�+�R<��"OtA�@{������u~��	�"O�E�5�_�g_�Bv��	GP̍��"O�	�@ȝZ�ܑ�䙀W��LXe"O�9#�l؈	��tс:�݀�"O�[kG��R9���Ē�h�1G"Oر�!.�0-������z&VH�"O�m3���<<�T�I6j�:,0mٗ"O^ܘcԫOt\�j���
��"O8�rJ0u�Ld[�%�&}��y""O���0/��9�Z6a�K(�T8D���$ΖN��\�թ�0w�*�R1�7D����7|��(��W�o �Ғ))D��Qc��|���D���mi��8d#$D�@$⌆|v%�Cƶ�bT�%D�4����y�FT���%cqd��$=D��:�m� �ܵ��J/&�&-��?D�L-R9�V�Ҡ[�AЂ:D�{���6_�xԛ��P,����>D�(��	o���k��>�ƼJF=D�1�&�7c��� �R*�֔CEc,D� c1 ѩJp���P9m�R���m-D����*��Oq����L�@�����*D�Z��V�K��9@ D�-�P �/+D��C��Ь��3���0l�,:�-D�h���.f�!ȣ�ְz,�B��(D�<K0D�>$v�!H�<1�A�u'D��qA
ߵf`	�)['2�:��c�%D� Q	���� I2`B: S�e(#D�4��hd@ى����zy�hQ D������/p�P�Ӱo�"u:"��t�>D� ���i���B�"�J�:�p�A!D�����w��;�)��2�V��a7�=ð>i��D0}d��7N�9J�4���.�ux���.V�K�2���n��<y�ڒR8���%^?X��JAw�<����x�^Y�#Nx�I�(�p��0!������c�x����*zP�tQk��/J��aL�W`�C�I���a�&B��<��X	LN)�P�"k$���a�Ÿ�4�3�ȿ��¡ #�������N���
e�
 �`��@XB��m�?V�`��H�F&�Kń�M�r��-M.�U-� V��}�5Y�axba-h���$��
E���*��ֆ&B^��쉄
X<9!�M�C��)�':���܋��""B�1�>�s���
�yBk(!*f�I���(��V��K�'},�.�0(�fM��]!Ce�� SDX�R����I�ʸ����{ݼH���Ę����4l�)5`�ժ��49D����
H�̴��,{�qO��eNۖO=�5�6Iˀ[`�����'�~�K�����!G�6C��5ᒣ@!H^��#�a̭Y��x���G+5(��>G�Ȃ��I,}P8eq�3O����G� `D��!���v^d���>c�"���WHK�6\��Tl��4ςRnJ�x��oZBV��kV&����%Ü-8	�?�!�ŧ �� ���,�g�? @����O(p��%;����=�(�0E9N���2Qɨ���!�!0T���a����		}qؙw5�t�a�J2�P�ABD�(f�C�0 c �Hy��8���p���/B�艋�$ӆ��9�u
�O��2ĉ^�	@(7c���Fu�q	A5\�,�C��H$:���r�*&�(��� ��m�O� (妼J��& �M??q���4�a ��ڼ){�$�ܕ�����`���CvcR�A�ҸY0��*��Aϋ�e4$��i剼.���n��0i\8��O,56����k�lHR�h��ц V�I�Aܞ��a� J�Ա���>�x�)����%�P���u�ݛ�z���Θ�Kwd=�螄uܱq���yb�s��a�᜙�p���^?�[T/��S�HS�v�:�QiD�*�@1�ϊB�,)'
C��D죂a����x�(����
;�T��c��6-Y�fQ%dp�h6)_2G2(���� g���`��!�Vp@���'az�@vI߲��DI�Ek,<�v�ڊF��1�MF��ѻ��m��� !��1�`6-�9{�D�e;AHB�?e���P��y� p �4Y�n��NŎ]4��k͎*��t�EM���Bذ��X�"��b)Oz�#�׌e�h�3�Ĩ:d�䕿'�n�ٰ	�	cM��PG��=�^�sR�Ɵ�b�(�q���c��>$�l���iV�aJ��0�(�>�����Qd�H"��N�*�� [�#����'>E�@Nj�� rf�ԇX>�>!���Z�P�Pd�`�M�07ڍ�ǖ�>�J�E'��D0c�{sb�s�[!S�Vl��13Бᇇw�8��_=z4��M�i�A�@H����p�����2c>� <�cRJ�F�&9����
�;��`}R�A�i��H�GagH�A�
Ī(�HyR�#�S��H=~�T��Seԍr)��8�@�<PŜ�'�E�9T�'ǚ䛧��	?Y\�@'�X	P�CE�_?v�(�yg
/_Z��F/]K��3w�C�r\�����m���3�4K�
(���@9O��堁�d�x�b��&�4� P���Е��3(@4UP� �s�0��Z��,�B䓄)K'��"C�H�jמ	g��AI��&�'� ACR�tJ$(:s$�`�OȠ���a�!z��@#��B���S�[Hb9�')M6g�0��A	�3�����W�������ۼ�.�
ΊP�����5O]��Џ<������<1T%��@:���I�u������łX*\YZ�0p��,��HP�^4��&1�v0[�(�O���@��]&Du
#�*�ę/ZXj-p�a�.����q!�8����{��{����(@��Y�7��s^yYVc��P�y���b��ꔣ�`?�ae��z��}RMC�}8��'Vypb��]�F�Y�d�'�P$��Ob�ru�&D�yG���$ɀ�W�R��0�䛐t"̑���0&���@��	ǜ���B��ȓ�䄲�쏹_��4K@��G�&����M�謓5���$M�-�������o�y��A4MI��6����S
@�a�A���V�f��3��'�J8���O�0��hC�,ݯf�"������C�O�u���F�ӛw4�9���ۏ4��HGL�,c�:��<�*�'>��*2��z���w�A�'=D���F�ZO2�`�Oc���ĝ��QB"�Nz���x����|nα�3��> ����w��	#&�৆����<Y �έ6�n�X���04�$	�mF�<aCHV��|$#Ӳ�vT���0�z���21�<%뇽i�ġE��::΀�	P��6^<r��'�0���d�9T��es�/5U�64)�l@q'�{5�_�3�u3U�C�
d Q;Q��y[�/��W�&q4��t-�n��B�G�
u��L{�&
a~"mA���,ঃP()f�`�I?L��ݒ5��9)�� �f��thZ�]۲��W#Q-!h�P i��I��O�t`i�O<`Y2Ə	���aIt��,�QA)F�M���'#�8)��pn�m�̹`���n3�-QǤ��0����]�0�4���C[qK@���D^;o�ܑZ�I��r��r����R�vVL%����B
~:'LK�Z�<�@�ՀI`�cd��r���Ui�pZX���DC��G�+.������B�d2F�D{CQ� ���"��ˬi=����kP3� ��V�����a�,S@Ry���R�)u�	��J��'�v\�� ��S�����ᜭPH@Q�`,' X�Q��D�Qo�A��/T�~�h�
�(�<Ն�*�H��G(�)2���y��D!Sj�U��O�)�u7
L#1x�$r���v�|`FI��M���_�U��`ϝ�����	T�,�(��C�-@��ِ�*�J��J<iC��OD���C	�1����7���5���dO<?��SΟ>y �sslQ�MA���I�0����`��3��
�i��0r~x�CW*��	Cf]:��\;S��];`���k�1EaQ�KT��;��|3v.Ï}U��Z��P�M���f�$̰��.#��`aܷ��C�ޟp@l+	���6t��U�K۰ �jI��A��ʝ��MF�i�Q���v���~a�bH���޵�QM��m��%[`�	g�H��Ҍ�"��`J�MF1	�܄@�MĿ*���K&�j���f�F胢l�?!��pR�-�1�ތXfG�
<Q2`̀.��ء�i�7�Mc��%C�y`e�=(�V�W�42Tx$��[���3�� k�|�8��2|TAv�U"M?#e�٥n9f(;��U�cPR9��aipS쓶7��[wª�j�)'�	���a������уK���M�0(�4O��YP�ˁ�8�4(Q�_���E�
[�������A�شT lH�,�+3�
����>7}����G��6�*#��Z��=��o��&�^����A$�D���R/d~��͎�d��"ȵI� �B&�V#9���)E!�X��)R�dj-�3��a��b�bL���q�lA��a�0Kƒl~��l�c�فh���`f��o�*E�#H4:h�	��j�%C% �´�e9�!K��P�Ӡ�jiң�iD0l�֢� �?	�,IpBx��dBo*�̧@�(p���F��d�9l~f�;ڴ�c�C�{��P7��xL p��24:d��W�	w�����$�	��##!CB�}�2MHC��)���;0d�6.ې�XT
�(G��#�I��)� ,ݘO|̀�e�6:b0}�P.� �ƹ�!��)W�Q���
�������Jl��e��=o4}��4qCn]˲�߉��ل�Ԧ���x���7/�����I&���8��5,�[(�n	�\T����c_#H�\�r+Q�q뚌٥�K\4������(�1�N	]Y���%�L�+�i�6�SsÅ)�s� :S�uD{�!�O���HJD0A�B sA�d�!��n�VN�P�%U�-�T,5���P!G	*!z���Jp�RP�о9ReD�vV@-��k�q� ���OU�\ '`�EwȊc�D!t��+&0OD�I4��-:�Z$"����g�Lg�ԝGrؒC�D w� �k��s� ���AnM�#�ȥx�$\���٣�~bN�
�0��V�~|v�D}�6_x��������5B�� �
�Y��W9ٸ�����?X)�Qq�Q5Yr����ۊ~�����Bٔ�7턪Gu�H-�5B�Dd
�aZ#V@�RG
�0>��":O�T�W�XT����O��0�$K�'���Ł/*�4a��nӒh��τ1�0���E'/:�9p$�	���!%�-�L�هK�! �tb�'[��*�[G�'8<�0%�R)ar�uk�HW�{�Xу��S@�V��;kf�:!o�*z�vtrA
%S�谫V搬�r���wC�\�uF�V�1UL
 O����M>u� N����M��k�i�6����V�)�~%�Q@ĕC�$�R���^J�����U�JL���+V]���X^9� ��C� �����	�9��΂�~g%�Vh���'f-�f�9	���! [�o�<��GF2o�.���Kϫ����%�%/p�5I������u*�=_�M�rǜ�7^��iq�'�&��fGN�.Т�`�#�'<�z	��n~�h�ҍK#0<m�Sl�N�(���GO6-֪�@�Ó%9�b=�$쒝l��D�R��t2���*�>y�'E�P:���G�Rup���!i�|�3�U� n�p��fr	�놓8�F�IbF
G�Ta8��n�d,�CJ��!l� `��ϣ]�������V8!AY8�Hã��=
rDa�نi�Sh�k `Y��tk���ׁ��oGV����n��87���x��dĹh&lqp��
q`��O�@H])��mPe�-h�y-8�ɶN���\2*A.�!l�9W4,M�Є�Z��-�R���qC�<�
=K�+G���V)�3�^�S��0Bdl�J$!X}x���W`6�b�����Wp��0��ȭ{	@�)�k��^�n�(ՇY	&��̲��Ğ0�v��EVSy��«Ȭ} P�0Qa��m�HH��JΗ4�ȸ2ǅO���(���|�y�'��i��sd�D?gX��я�$|R�B�f��D�H�sF�T�r�)"�Įa���n�=bV���o�59��p3�V�Lg����*B�z���[�B��MZ��O"L9�vK�S`�XQ�dZ��th�$�?V�"Q[U�i�h�b��*��H�gJ]&o�r�"`�5*�ɘ�)�D�	��JE�jR�T?j�CV�� �Y�t�P'�_�}tXq��+�Xy�5ꆌs��]�w�A�0��d��v�=�ׂ�	2�<5+ ��DB��:��Y�z'*�#J�3��<	�c�l�VՓ"䀂zzX�
��V6N5�6n?,I�'�-���Ku�Ԃk�N�Ӣ� ~~B�
����j|�pu˗*yJ�)���T/L��j~�@ M܇T�*H3��|<�˕�����IXu�B5Q{���'���p�]�l���e��}��,��@ۺ
ˢ��w�W�N���� ,s��-�Ǔ^� �҃������$߰lw�yt�U,Q����éj%��`�@�D�2!%��%b��GD;��B�G�r��R���'VA���>s� �˷C��!a]�J�0���'D��d�++5����N�w�dH*`��"O[&�ʂcЊ1�6U�Ӭ��x���p5#6XL�p�7;��e��oM�'2ph��$�ɦ	�r��6bT=���=,�@4�M¡.���S�F�!%�x��.�7�"���2j@zB�>)�J,(��b�q:4b�:_t
��aժ,P"�b/ʓ.�|"H:^v�?	�$m�S������)kF��Cq�ޘI� \����ܐ�dZ?���4M�R����QɌ+nL���+�L�@��ŕ\�P��!i��!%�,��|_Zy�E���@`*O�I"01Q���"J�ԳB
�8"�䘑��f� �����=Y��b-ϛ%�S6��r(�˵�ɻ$����q{��W����&$�/0������(���ɯoA��2c�m�V�M��S��ɒ��X�6��5�&*���� R�/Z�Q���hC�p�R��H��;��4BU�3��\"GJ�9��#<��P� q)JRV ���L��^���R�q���sG@E�i�ؔ�H�3�>%A�i۾r@ ��(L��D4�0�Sr���['@��j�v9�b�m}B�
 D��t��ӎ}�k���E�EH�+RC���i#�&
���\+$��2�ڽgiP��c��Hd�"�"��G,����Ů>@�y��W.w#��
tb��bbJ���DۓBp�qZ�@y��B�(|<�����*v '�B�:��B�9:�,e��bW�pY�Hq����yiB�����D����*��5��32��.BD�\1a-j�mS`�='�\�B�D����R!�]7��O6��ŉ�N���s׍>ut����]X���T��8q�>�7G^�K81�u%�N���[��¿w~�%۴�S�\UJx��m\�m�\ ��/͗`w4y[�}�ԕ�v��"/��`!6�w�.��|a���42�@x�M		�!���ESSb�C�H:	��d��@�2o�Bh@e�>1f��󐩊�-�vhDV]~�S�I���L���B.hr q�F/c�:R�Ū�(��<A���>���g�%j��)�jC E@�
�I�ip������޴퀂iT�9N��:��	�-�Dc�m[/�^��c^*%ؒ��"��O��򉔯:K��2=�.1Y�CX�O�L���(�b2��pM��a4��T�E�|�u vc�:V��M�N�S1wx@�&)��q�`E� E�<h#��#(m���A�S��$ r��6�4��)(r�X��$M�$Hs3��D*?Ϭus�N߰DH%�c�?#^��c�۴1��=3DQ Z4^-�C��*>΢mS.��CG�5#�?&D��s�X�0�1�`�^�ZF�sa/r,��`�m��	����Մѿ#
��=y�h��h�#al�m�E���O�"..Ej���"$��c�5i�lS�&cB0z"II�2�]�v �� )"Yb�@eI�4䉚Ĥ]ہˊ�?*x�Jt�۩rt���� �qO|pQƐ_QZ�y���"B�@��sDF2i��5%իf��=�V)�$h$iz�(@3 �r�k�l��]��AӤb�ˡBѩc����^���)��A�g |ت8�f,U3J�n�g�vG����i�Z9�Ԏ�xn�l���"yФ,�F���w��Q��I��o�ܙ�B�CL��uڤ,�@�i���I(����ą���	�n�܉��|��DE�t|Ґg9|#�p���$�^\ƥr܉�b��(��yq�O;:aЃ��>���ɻ9c���"�Ra�)mQHtJ�K�0��$y��� .
��&�g�'':-��Hئ=��ETl��jшX�89`J��0�V� UF��U���k�Sy�C�c�\�2-J���LläL9{��(�@��1�N{ ��p=9���#P�� �#��0���#�L�;��iR�HH?i��ǃ3}�j5}�̣1��':`���W�8ʧr�n�SlC(����-�Ky�i�=���$>躈���c�"|���#� |8��Bs��A��
=�:�!BK���$ڮ�T�?ӧ� �U�m(b�~|[U@DnZ�ʦaY�#�ܔ
&�G7��F����ŋad��4�� B�8�e�=|!�D�d@;�IʷAu�Bd�QmR@�0��p31�g؞��	5v����H�
'Fdӷ-�O(�����y2�@�z�N�R&P�N�((�����y��A�j�<if�;
(��`��yrBč@�,�x@(�+.��Ћ�y2)�p�����X!�4�PNU7�y"oT�J�"�s�͉=:L�B�	�y�#W<y�@���	�gb:�y򥎆a4�����䈁�JN��y�ǃ$���y�U4\�@���y���2�ju[�hB.}��PՋ���y2��O��C�~��Db6o'�yb&�
��qK�v��A��^��y�'��|\��a�߂SEl���-^'�y"�L+~�:$x@nI�Xb:����P��yRl��r�R"��M����3���y�L�1��4r֡��FH�r����y�"�8~��0�Uc̟�X<� �؈�yb�5W�$���Oɧy�V���J�yBn��y��H.�c7��wL���y�A[#-�L�`��(Pr8��i۴�yrn�4G6�LT�R�Z9˷��yR*�0N9^(�t �J8��+��	�ybDH=�tF!F�x�rg���yBj���܀{�̃@V�%��#͗�y��ۂ`h�|B �
�k�8:a�P��y"��+��kt�G���dP$T��yb�N�.3n�����49��@�N��'6��8E��7v��x��G*9��9�yb��*���8A��)��k�EJ�=g(���̦� E�w��L��O���s�c��M�bIɐ(,h��!v�_���y�I�)a�%M?1�a��A�<|Ɱ�� ����К`v��0ყ��c0/��*��	N~�S����1F������R&z���>�k�YN?�"	p�N���'g�á@֕"~���Ç�'"ќ�{6����ӽi}�x*��?�˱`��?ŋ�t��ܜ+
�b�Axh���3F��ɱ� ��Fa2��� �<9k��OȾ�,X��p0AA�AxJ̹�̛��k@� P����0|R�B�S�x;��<��4PA����� �z�^Գ�`E�Ք��c��-��?=�PbW���Ah@O݂r���!���$t�Q�X��) w�Q���	��:�8��W
"�V<:gb�w���IL�P��Zļkç��� �.�O.4�
�W��]��u8�|z���0P��/O�>�`O^�p��u.�L�iha�4�I
�HOP�Ov��I��O�D��b��ږ���"OzLR�m�I!,P�π�tX���"Ot�I�`C�w�2��!�M�yF��+�"Ob�Rŕ�@�0M���	��h	S"ObqHx�N�A��5���H�"Op��a�%g����� S��"O�5p�ѐ��:�&��JP�"O:L�$\��P�^��`C[��!򤚞=�&�9)YOe�i��K�!��ֿ
���p����u�p�qG���=�!�J�c��9���C�, �3ˋ�l�!��@�"Lib�\(�%̈�O��Pj	�'l���V=e��A�匃g|��'b���͙�8~T!Gf���Z(��'�4�J��A�fB��hcN��
�'��H9 
��2��m3^aF�
�'�=J�
��̼�2CB%@�8Ȇȓ?�$�i�ٖ-���H\k��P����i��WB2�/�V�<��ȓo��\����G#�d�[=Q�<�ȓ%�l��a��D�ȼ{PF�6H����Be���I9�f`��I�2Y��h��S�? (��@�ыF?�XI�k�1L��X@"OYcvdD�B�>3�埏@���"O�%��hN2n��!B%�ئBfhz�"O��E%eA~@zuM��zM�}KV"OP��BU.e�8��m]�3HH��s"O�H�.F/�"
_�vA�iQ"Ol��]�����Q��3G�<�c�"O���G,�F}��fʔ!�N�H!"O�z�I�8O���Wϛ�&����C"O,A{��0@�X��[�I���C�"O�ٙ 9K�|�:�LM(��U�"O��q� �
��8��(`h�\0a"O�$*eaH�l´c�-Y?No�x�"O5#v�O)Z��	3fZ����R"O��X�+]I�T:��P�sC��Q�"O�9ɰ�ȃ. �d1� �c+^x��"O�-�G�S5��[��\�X��"O�5��+�.��@��� ;8{Fq�A"O����A��22 �1��0�"O��D�ΣV>�LѺ�R�'�R�<I�g��g�R@pVl�j�F��bTM�<Y��݇ctts���uv:j���I�<	��5s����Ҕ)a䑱`UC�<aR�Ɛ;�P)GI�~Hhq1�Y�<ђI��KX�4R-D���D,IY�<�v����q�W*��)b���R�<y��3g��	�fՆL�M��C�u�<yg��-��и�">b���hf.�x�<��-T/s�������+s�] cKr�<6�����4J4�F�9t웡�g�<	�k��e�zh{qm��y��Y;��{�<y���?PXd)�.�IS�#_m�<�^�(M�]0����VPyj�+Dk�<�@'�P��V���q&�d�<	��ɯT�`(2�Ǌ1e��m��Tw�<A���kA������T�n��׭_[�<)��M�J�;@`,c��Y��P�<���@6e��j�M(*Ȝj1�\Q�<ٲ-�4�H���U���̚I�<逥K!�a�g	�0r�kĂA~�<6φ�$W^ݒ'�D�؜�W��v�<�g`ڕ?c�	J�L�Q�<� bL�<٥@ֶ�t����[Sӂ��F@K�<A櫒����s/D$z��p��PF�<�&h�����q	�>vź,H$C�<�,�� �ۡ��71+��	�|�<Q1,�?�P�"��+AΦ�Z� �{�<ѐ�"<	j�,]@񣔥�;|��C�I�Z����E�?��Ǝ٤[�FB�I�2�`-cקI>�6���/Y�%��C�I�3:�3��1��yib, i�C�I HHYQ��AT��J�)�
jFjC�I�p�� t�g�Z��^�txVC�	uqj�	��'^
�Q)a0~txB�8p�����$^À�
&d!^�B�I0@��Y�a�2�V�q�Ɓ�j#�B�I�etx��f�[j��%%�B� y�hy� ��%.N��F�Y:�hB�I_x.A��k�8�I���&T��B�	�n����"<.�,X:�/Z�H��B�YJ�P�\;o
� ��#�dB�IU>N�r��"��1�-��C�ɾ�"xQfB�+8����F>�C�	.PW��1���~8��U�E)�nC�)� �b�CHS�����˓�3��<RB"OVպ�:�μ!`M R�L�"Oi��a�%��٤���&��5�p"OrQ�`ǆ"Obв&\',�J4�w"O���k���,���	D"O�����Ş;���� �(G�"���"On�{�]��M#a��Me����"O �jN��hVx��Ed��f@$1�"O��
�G!��L�|2�aE"O$	��C��h����(�h3"ON��u�0qx\0+�#B��<J"Oj�Ck�J�ġ�#�b����D"O����g��,��M�k���s"OVtCԂY4�	�4�N<h�@ "O�L��"�-Gȭ8��R��]j�"O�x���̉8	��`���k�h%�"O�չ2�V�hT�|� ��9C�<�B�"O6 W�ȏ?��"��:F�,��"O cG&��rs�ak�`\�i'�}��"O@���a��>�KrAȚ^7L���"O��8�(�$+��q��]�K0@m�"OR���P>��BP��j/h��"O�u0����"	��f/КX/B�
�"O�Ĳ�J]�8�ʱ��$�!z���"OX��c�+r�*2�Y��a��"OZ���/�p?��bJ�N��mS"O���Sn�nͻv��'SlJa"O���䘐P:�E��m��|��4"ÒP䃚6����ԘfI��"O���$E�9ª���c�uX��Q"Ov�����pD�`1$!�U�xb�"OP�"$F�]݊�Ò�NXp�-�b"O�x9b�@�P�-*�*Ғ%pp��"OP1jO��&�0H�Q�U
^`)d"OJ!��IH�^ ��i�I�&���8�"O<Ԋ�ȀEBq9��zبp�"Oj9�taײVC�T C�8o����"O& �爇��YT�W�Ak�4��"O������I�J a� m�ePA"O��U�͒o��)2� G�����"O�Y �-�"=�m#.S���y�"O��O��):�!B�Ǡ
�R�J�"O���L�8H�� "��6l��ҵ"O����ҤK7n�*�"uL6��a"OV��E�T��Es2AHxd��"OH�B���3321�$̴A<��"O؍	!	R_-b�fŋ#lΞ1H�"O�Q��		7#Rȹ��P>d��G"O2��t��uPd1j!��_��B"O\��K<p\Lu�p��-m�^��"O��(7	�W"$L� PF�D�X�"O.1��%�r>h!q���P�����"Ot�a��� #`*��R�ċr��QB&"O�D��d�&^94��4��x|��E"O�="�E޾qD>E�2
�c��	��"OA�&I>�<��	�6���Y`"O�4Sq	.L�:���� 6P�z�"OT9����9�b��rm48��T��"O&�륁��948�;1�-Rp�� �"O�U�v��eȡ����M<ДS�"O��e�+ �-��46c"O\���W�a��LQ��߰�6=k�"O��������Q���1��`�"O��r��_e���bд:u��xc"O� 1�B��@@���H�)[�\�1"O��3�����Af(8��(q"O����N0=�Xǀٮ3z�)"O\e���ƅ!+��k�A)#j\�	�'L�b!��.!����#��0�(aA	�'t�����L�:?���r�\4-3�4��'����*I��⌘�9\_�r�'sR4��	ߚ+'$�SA��b���'��Pz�C�%&���h˦, @��'�j���g��K�4T���,�:`�'h��Ły0��S��E?���J�'H�rm� Hvh���#�3�$�
�'d i��E6�,T�d�.pƙb�'���ϯ+j<�9t P��B�H�'�rd��n�9A�Uz4dG����3�'G@1I"��zFu�` E��0�*�'���&���@_ =�GF^�v@��'=D��%���T�IbLs�J��
�'p"�"��,z�Йf��ewz�`
�'V$DJ7m�"!�2�����kT�PR�'�<�� \�@ie��:^�\��'d:H�4�âs����(��3j���'��y����7\�f�UjÄm��D[�'E���Ӊ�1�V�0�S�g��'l��x$��/�U���� lm6��
�'����v�[9j��ǅ3P�:
�'F�°	�e��X�O�>tƉ�	�'|N]k%,x�!/��t4�"�K�<a��8��]C�m�����YD�<�Q	�b��P��;M�D#�@�Y�<�j�����5 �^���r��]R�<	$BJ1;J	 !�	.����WP�<�7kC�Zt��ʒ!ц|8)��q�<Y�ƙ�T݂�m\�TWd��*	o�<�G�Ի��2�Q37V9S�,�s�<�tكB��m�%�~E�ԢB�F�<�@�P��h�b��I�Ҭb'mD�<qG��\��-��k��� �d�<�p�8Y���h�M �)��ENw�<!v�QP|@HCPϸ}Ćؙ�bPq�<��JT�a�����H,H(���D�E�<9w���B���p��(	�����DB�<�&�W�N�^��呢R�N���u�<���F]�&��#� !dX�S��x�<YS���(��1*j�܁Q!C�c�!��{G>	2c$0Seq�a`T��!�$	*\� �.�)>Pi���۴�!�T�_����g8Ezp:Q��2�!���8��X9\ֽ`@�CAo!��(C����/Y`�8�2�!�,8!�$��\����D�m�*D��� N�!򤞢[P���
�&o�����/C-_�!���<,*�J⩔:���GгD~!�D�h���׳C��$�Є@2
!���dE:4
�L�=\��L�d�ټP!��T/l�"��UA��~������!����d���)���;cq�"�*_�I�!��тh���I�{Q&x�0*���!��[�l@2CZ�+����'O��7�!�d�J� �  �P   g
  F  �  ]   �&  X/  �5  �;  5B  vH  �O  pV  �\  c  Qi  �o  �u  |  ��   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl�6x{3;O�1"�'"dE�>2��EN�%�D�j4Ý_�ց�Ф@�n���#!��a�w����CG�?�JS��?e3�f�x��x���4~�ABA#��j��5��Ėj��]�s�??����ƞ��u��|@�t�'oT�ɡA�T���,w�Ɲ{� �y^VxBt��O�4��a�|Lc���I�P��П`�	ݟ@�I֟0i&ˈ�	�$UyYD����㐼m����O,L��E���	�'bkۊQ1��'�r�]d��ÃN�
V��!BP����'���' ����r�R��?љ'���n�u
����j�8�^�s�@Fu�r7O.%��U5���z��GO���	�S�Dx�O`�����>����,j��8�p�F���,k�P=O%r�'��'���'���'���ɼ��h�Hy���!�$������\��4���'jӒnZ某��4J�UD�i����T�'*��i�Ę�.Af,�q�ކkT(d��+ғ?Y�0{r�7g���	c�34R�pʃ&� �С8���#4�0�3�X8i�hl�McҸi\���O�.9X�2eĈĊvF\2!������3�0��w�h�xz6$B�]t2�s�-}�����D3aBRh�U'^���ݴKl����N�vXY�	^2
p� �T9vв��4d�l�`�v�̨n��M[�%�
X��U�fov������#��#�k	s�>���,�):��:R��<"=�0�ҟ���`���n�n�Jxq��ϑ	lLq��M԰b�v�^�F�����;�|�;0����?QQ!�	c��c"�ոS��HF���?1���.�x��!�^�p��S
ݖA�����O�DS����m�h�d�U�[���s��T���D���?1-Or�d�O����$,�� �5���أbUئ��1,�v7�1�C��,_�V	bbm����]Y$�m��M~ݎ%�I���hh���Yj� �K(�X���ûo��'�VʓpS��xb����FX�U%��<H��ȟ4��`�S�'�y�H22�0Q#-��=���91d����?�s�i$��Q��}0Zh�q�G8?�iX��z�f�R�`�����@`D�c��$F��J�G6�y��TR\q�Q�IzQf���yҤ�,[4%���C $QdM�a'�?�y��CtЅ��E�%Ja!y����yRBI�0,j��#=p������yBՏ:�8��gJ�/NR=ˠ���?Q�g�f�����h��所&Bδ�%��D2��{s	6D���i�dL�*�H�MS����2D����!b*QX� �+W����	;D�Ĉ��*S�ؘ�R��hG��з�:D�� �ȓ}� -kW�)���T�=D�����.�\�!�*@KVa`�<��i�U8���6
��/7 z�EߗR�6�{a�<D�x����Vq�1�⋐�2��Ѕ.<D��y�	H0COT�Z�!)���,9D�`�c_�n�\���ُC|�=���$D��3T�� {y��B�jB#]�v��F#"<O�t��LC���I՟h�s���C?B|���4�lx���ڟX�ɣPx0���ş(�ɁeP����Ԧ�.ϻ2W�Q?|q��%� ��H��7�0<�Qn�5OFա���%߸�4N��ȴA���2����N�Otʘ��*0����OF\n������ ��&V�ř$K�_�h�{t�:?������(����QBE��qR�!��ec(`����>Ɋ������U��>|�dʧ�F�>��)� ��M�K>	SJB^E�!��2�O�8Ͱd�@XH��:��f,���U"O�#�<@�f�����8N*"��f"O�LHӃL�["pʂ �
���"O�A�`�ў��}���A(���"O���$N"��x�㈪[�`�2�"ODɸ��/�F�k2d�7 F)�bKu�ГO��C%����d�OF��<q�	σ~���-��!�a�]�J���$�i7�6- Ei��K���|ʂ���P~�� ���/�p#��,��J�]� �`�7���"�	��$X��'zNA+ O����4r�) E�qʵ�iv��N+ l�Ie��\�	ퟘ ���.���sE���`Ѻu�fNgx��P����-:QJ�≁�l.r4�#�O���W��@�4���|��'��������1	I��ir1�Qzĉ0���O����O��d�<�|''E�d��Ȇ%]�xb��y��J�2�衰��G[>���4�B�`��y�J�o���WBA�=����λ���یKCT��`F*(��t�7�G9]txEy2�W�[](�To08s
Z���E�$U����?	��D(����ڜ/4�Eѐ/�V���ȓH%5�&��(����GB�mx��$�ش�?!)O��@��@�S�)�jAZ!	F�HSCh�/4�����<���?��Z����D���0;⍀�=
� �I��@��Cm�9��ߦ_��I;��'Z��#�	�0�v�;�ɗX�FMj�\�{e��+!�ZD���Ƈ�0<)�"����Ik~��@��Qx�iQ
� !���Ӂ�䓟0>4��a~*�[��m��|J!g�[��@���&���^�����*��0�	oy��S	��6�)�I�|���Rl�@�S:B�T�S횴Q��h���?��ؽ
�r��s�L�裭]��?E��#�2C�f=�W�_�9��59�L�����x$Mj���Z����n0ڧ-��qB�0>�6��p�a���'{m ��?���)u��H�����F��	`tp�rW�7D�s�%ѱU�lI��A�B�D8!��4�;8�>}��G�p��xE�&!)�T"�b�צ���Dy"<��d�'��'0��
� %f�!o��hD�U"���!�@�g���o�R�`&��`�g̓@�>�� ؠ&J�p��7v,%M�!?{\��"�H0�J[�g�y��J�ÉY��8jP�5�V���4�?a�EhP�����,OZ���O�ē7]_,���D��/��h3�K�w�B�It������Z�Լ��>t��˓	�����ڴ�?�/O0��ۆ
�؅�uǈ"Z������QX�w��O��d�ON���ƺ3��?Y�Op��%'ȁT��T��bU3�V�$-��xR�Śf����I�.m6@@�R ����
�'����W!��y�6���0����?�q�'��}H�g����1�`�=C��
	�'',�Z���}��4�УZ�9���K>q'�ir�'���qn�~
�"���	��ޥi�@Q���֫]�~Q����?�#��?�����ԣR9fSj����9l���)E	DE葧�@�O�2�Kv��6{Ge�J�'���w�7S��7�S�ZB�L��@ؙNּ��	Q	a2zM�tG��SaџD�6��O4�l����*�lՓ�W�dX���s'��;��'M��'��H��瞑p�r�p���,;0��Ff�'Q&���`�K�<�@�^D������S|�p!l�؟���f�T�F5zo�\!C���qT���3���)+C2�'����S�ռB�.�O�n���Ɔy�I�JÆ;�`���鐽��d�=R�0F*:H7��SI�H�����d��3�O*�!� ���%>��r@�J5Qf�h��O~��e�'��6-�ʦ]��P�O��IB{Î��0@q��l@L>���0=�G_�Aڸ0�O�_��)S�ɀw�'r�"=�T��N��\�� ֹ-�I;��>��A�����d�%�����O�d�O��NuA t��k�f��� ��w��1��rf����'Z��1I\��Ϙ'�D���^W㐉JT���
tL��)EN�6A F�'��I�Y(��Ϙ'S6�`�-�Kb�[��_�!q��i������jc��'ў0��h�/YHDDV��d�J\�<���&t��A�^�D��ex�Oy�o9�S�P�����4V�����Rz捓�Bˎ	�5��ڟ���������O:��1Eʅ3"�B�◦�_X�pA-�!9-��"3�ȦXf���g9<O"<���L�r}k��IlN�!o-Z$.u���?@�D q  8<O y�e�КN�ހZ�5.������+�'�ўFx̂�r�;��4X���=�y҈W'~�	�h� ���3e��&��A�IB��,y4��'HfRA�ŏ5nW�U�2	_�3t*Ň�y�*���2ΐ�Z͞���I�ȓ}�d���*����� ��d�BنȓdjN���A^'^�L����*?����'��<���k[4��_Byƀ�ȓt�=*�KD�=ޭYZ��\{��	Y�~���	��!��J�^A��b�N�<Y��O;�~�զ�@+~�@�RL�<�Wi^�Dʂ�C��]���� '[`�<��FʦS0��E)�d�z���]�<q�L�z��,�u��44��b�c�<���&@��dʤ%^�BL� �័���5�S�O�T%	��(�& �CeY�Lt�+�"O����%|T��$dR�R<l\	�"O���-N�$��LYe��2K6�t"OF�Ӳ�[�(�e��A���R$"O>-�����LO4�I lK�,��c�"O��J*%A.�L��i����U_�D[�,�O�8���,!$(��\9a�:]�&"O� h����0A��{��L�d$�"O0,�TnuN�m#����$/#�"O��[1�C�F��t&���).y�A"OfV�yL��:¡�v���е*�]x�l+BŨ���+lX�):��26�s�+D�0��,i� ���M�>[��5�%D��S���$:�V�H�CĹj׸�K�#D�����&(e����Ő?p��A� 5D� BVgş���Y�)=2�����(D���kB�w�"�T�̱&n���'�%ړh� 8E�4D��X��@��,�!(j��RU��yr,/y�����`Տ6��p�Ui��y��^�p)�MFA��e;8��h_��y��Y�8_��{�j�c��Q@B �yR�ԃ\ܽI��0^7����iG��y�;wn@�i��HZ�r�����?��Kd�����i�4 P�ꎉ�q��ng�	�bo0D��ɤ$� �8x�̯d��`�0D�L0W�w�Ƭ�0�H�4��S,-D�(�'�98݈��t�Z�U	��3`)D�L{Cώ4Lp-q#D�2!��3<D��+ѣ� 1�<�q Z!U��8�E�<	s(�8�0�+^;bo����#mT�ܑ��4D�$ǆͫ�,����t�~��@�2D���$�P䩛��ʮaI���C>D�q�:H��R��9��4�'F7D��V�I+�p���D>w�<�#�?�O����O�Ԃ4�#��!������H�"O2}jU����)
#A��6`��F"Op� %΄�D$��s�<	�p "O���EV��؈RC0c�$1�"O<2�!�-:����gC��h�z5"Oਙ��V�"V.�
�Q1�H�퉇G���~���ʬGU��`��vw��8�i�{�<���&2�n���K:	����Fy�<�WjA�X�8� c�RjpL�pc�y�<9"��!�������z�D���`�u�<���I�O���h$m��Vg@Ջ1��I�<��d�nT	!E��(
��[V��Пl��*�S�Od��ZSo�������X�f�LYbD"O,����x<�MH��P�
3�"OhZ��HM�t��-���B0��"O��A�O�+QpQ��+O�C�1qf"O�0��*	hI�������A"O&�0�\���P�Ч!�rq�\��0D�<�O
(a���]�p8�-��ra�4�"O@����՛.�z�0�KSX
)�"O-sP�67�,���D�7:D]�"Ob� �.�:B2 �C -_�j �̫"OH��B"c岑�e����0�'�8!�'2D�1��,F��Rg�U a����'鸘"s�Z	�v��f�\4�]:
�'�B�����')
�� r�SC��	�'2h�2 E0�!A���(4�޴��'�FYZ�͎!� ��sٕ0�j��'�DY��E4��|RÙ�/`�������.�Q?�
ġ8� ��qΓ�@@�J��9D���@;b���s�&V"+����7D�<
��܋'\�`za�KC�|��J7D�@)5���DTT�*N�F��g&4D���(L8_,ѫb�N�_6"�hI5D��ʦ���M9��u�N�+�@��O�� c�)�jBQa��$� pS⟆y05B�'E�l'!K֖�Q���
c��D���� ��p`�F�%�N��%�����B0"O���FH��vUD,�`�£R�Z���"O����)t{���U�R�{���3�"OP�Cl�$[�X�X�͌}�C[���*�O���[ �����G$}�y�"OnMJ��Hx���A��V3Iwr�#"On���#)@0�aX�pmd��"O<-Ӵ?�<��ٸ+V.�Pv"O*����%
�ҝ�"Z��}��'�2���'c�=Idg�x��ٙ��$}��j	�'�.|r*� ���@��@�~9��3
�'vd(�FO6�����(!�����']=2V`�&_wx jd�6��z�'_^D�2�1ܖL�f!�eD�
�'L�!"�%6�\��g�QNY����l�Q?ىC��T�ۂ���6�l��� D�,�/�*|Q�k�Kl���� D����.�<��`.� I��()D��"��X?|'z]�(�,��xWi'D����ß�'��,���6~�ƭH#� D�T�!�C6M٘ ����Ё��6m��I��"~� ��k.� Q"M�=��ah��>�y�iM�V���X�KK&P��=�yBi�)�J]�ƃ�DNp z����y�(��/Dų�G�$Ce~}�R��!D���d.E�(�t����&,��DH;D�D{I�=J��h��g�=9�PeCĩ�<�U��`8�з*͜b��z��+O�^,;v=D���0L5W2~�a�A�<�Ȁp�/D�$ ��N�Ri�t�޺����4.D���G��}�$������"%���"�-D�� ӣز�ؖΈ�u��07�*�OZ����O
�2�hݤ6�0q0�֯CFܨs"O��v![�;
`���-�v%��;�"O�ujp�G8��U�2�7X�m"O�y�"������/]�T�"���"O�5@��nגx���_����"O�L�(�)F��YB'k̯A�N0X5�	7A�Σ~J5G̎I~��AB*Z����@UA�<�r�2f��(��B�l(�A���@�<y�Y (��!�,0s��]�#|�<�A�'QI�t�`l��!1Z�g�_�<1�Qb��L�7m�%=��P�p_�<ـ�����0m �N�P�A�������0�S�O�Y�@Hn~R1{F�>VOB�	"Od��.}gX�م$dK(T�	�'<pqU�%3&\ŸԈF���
�'U܋4'�P�����g������'�:]`�O�;-̮��D�I۬)�'*4�Q�j��L���@�Ď
)�t,O�e�'�ЭaFlƟR����'���<�A�'�$Q�AC�f ��v��3[N8���'$���	J.tRD��F��&�`��'�/v��E°�V�L^,�@�[6�ybϕN"İ�)��9�|��p����>a�aFh?�*�XIV��RMQMC��!�Kk�<y2b��[7�����s��t9���h�<a���&:μCc��:��41�AJ�<�#��$��x&�3MH��Ip�<a����1a���O�.zO��@VFAm�<��`�:y&x��a�)J�⬸��i�'X�̣��i^=m�*�8�?������4�!�DϗCZ1�w�^85Kcc]f�!򄄸teN���ߵ&0��VIT$/!�� ����ʝY\d�
GC�#PMA�*O�y7"ژ5��(b��!^�&8#�'E��B6���W�<���!24R��,�aFx��	�Iw4���U��޸)1��\>�B�	�+�b �a5t���A&0=C��<(���A�*U03Mظ{թ�d� C��1@��(į����`$��B�	o¥��b��R��� roG+߄C��!c��K�j�;C���(�j�F�
��	W�$աcd�~3�d��8DC�I?!U`�Uƍ
2��XB&O;#?PB�ɺ[��HSm�M��]��6~�B�I%9l��yr�*��\��b��e�>C�I�W�͐2�+MGE1k�:Ya����C�&����-eK�,�%i�� ��V�Qr!�d;g������6N����@�f!�$6,֜�`���a����@���!����3@%H� ���g�Q��!�$E>ܼ��@�0
��ȣ��<0!�$�"��QjuI�>A ��p-Z"ўtsSo7�'yrм�AM��@:�;E��v�ẍ́ȓz�м����\�h�+�y����T����w�"u�0�R.O !�"��ȓjZ,���+0 #4�D3~�=��+� ���Z9��x��Oi��ą�k\Lpc����i�2Ixta����ɈIT"<E��m�Ԥ#�!=4������6jB!��> 
B��k��z�Yr��>�!�ĔO
� ��g!Θ���D��j}!�D�6P�օx���G�fɐb�8+�!��31d{�+�����j��
���v�h�)�C ��t�D&υi����)}"f�^}�	`}H���	ɒ���q�8;}���L$��B�	Ou���G�v�� hdʆd�C䉾o]@���b-* ��@ư+��C�ɰ �8�����;t�$�1�lC�^��C�	�Yy���"�&�p�W
qP�C�ɺ:<�{ֈǹ=,�)F�n
0⟴8 �>�S�I
	�r CT�]�y2��p�l�*�!�^�i�h�Y����1Q�X��[� �!��I<Z�ƌC���L�r�bN��y�!�D�>���'�L�,���	�!�I�a2�a���/XڤajA�B�!Z!�$1������i�V���Ԉt�L�x��*�g?�ǚ;�m)��O0q	P<�c�i�<��u�<ٳ���)XAP���LWd�<)Į:��BŠʌ>Q�DxD��`�<�F�"_ʮ���F+�ȳ�Z�<yS/U1V.)p����%b0���m�<YVl[s4�kק�3cp�+����p�,�O����u���a���v8��r"O�a ��[��]K6#J�_Z��P�"OV��7A��D��b�*D6B���"O�]@"�\�B	���1P'"O�`Aׯb�`Y���S�e�
51��'��x�I�4I���dh���^Hq� ö�=D��"1ME�7iF<��\]����f>D��{��Y�I?2���ܵ��]�@�/D�<k�@�=T2
b�&2hA`��0D�2Ck�.��!��#V�(aX"k3D��t��B�(�&X�$� A��/�ɟ~�"<����*,�5E��|Y�ˑsulDaU"ODa��-�'E~E�iʋIR  5"O�В�j�
Y�֭cBA�K�@�7"O� �H��ȍ[�QC���2@^���"Ot��V |D� v �4��"O���P�ނ�lA:�I���`�E��O�}�Pi���7k�]�l5*Po����ȓH?vhCѦݶ"B����b�;\sv���T�����.FDtƃD:e��Ȅ��@����4��I��J��ȓs�6�� ��%+�VQ���
���ȓm�ȰcH�*uFxH�W`˴>T�I�Dy���D�=]0���I�ysF�#k	�C�,b�h9XV��g`\�g؉,�C䉀&�	ȗ�F 7�5J�׏(�nC�	�E�D��,�6!؎��E�w�JC�ɧF�P�F��w�mztGS�e�F�?	�KO�[y�f�'�B;�n����F�}񊑂����S`�'�
iۧ�'r��'��0�U�'�1O�I?3 ��!�.I�pi��4iѝ�ԛ��(�$8���g�Ȑ�ר4ú�E|��?7��J� ^px��6L�1g��g�!�$ȯ@N0l�Մ��D%�aۤ @}�}R�<!V�	Hz��w�B}����NCy��'Ҟ|�Oҟ��� �}:61C%��6��w�?��y�>�b���,J �P J\2K�H��+��I2>O��������K��� �ᅿN�)	2k�����~�K�����|ΓPon�)�˅�BA؀���S-{U�5�W����C��S.��<�OLdă��3Nݲ�HȀ�i]�\�D�C���U?���9O�5+���5Fbjm��nZIl���2t����u�Ot��O�P�*5�H�)�8Hҥȼ�Fq���PT��O(��&�S)-C$��7L���e�L�J���I�MA~�'���'�"AL�Lyݴ6�}J�)�&Q����sAQ�x��@�'�P=�M�\p��	�=�Vpy�����DJ���%U&	�AOʘ�O�s��S	!?I&(ʄ[jL��E�ߡ`>^���hې��L�-O��p��O��$֙�H�4�x�ʟ'�˅$�B��#�
^?qr��g~ʟ�d� F���3^���.T6��l�~e�*�k؟���էj����$�+4�$�9��%D�(��$�]�2��@<`��]N~Ӛ���O�ʓ�?1����|���@�`���I�(���2bԽo����'X��~����i�OJ��"�( �@���@ZqFT��lM{������?�'��	�v���+FmG+��E����h��C�*Ja��X`/F�$��-�ĈR�p�C�I?X����#M[���p� -��B�I=g�N�
6-�~�p���lҜe
C��ʤ�r�.��|�h��A���C�	$��,�s��>OH���m	�F`�C�ɩO��� �a��3,l����oqxC��/���ǁ
:w�p �A��1c�C�	�2��+��'I���׺7��C�ɣ����J�$�����@��w-�#<�&�)� �;���ٷ#2-GX�:��	D�<$�r�a�e	/?#�er�G�B�F�����P1KqL<��Gԕ-��� �5b&h�&��ڄE��CC�R�ɰg"W�0�h@���Z�P$4��	qJ��i`	�"�T��EN�f��)q�%X�����b���������i�����ʐ���`�	4�pp{�
��THa���2�H��+��G�| �l��xJ۴~<5�@-S1O���E ܸ{����'�R!ǐk`
���� �T>e�O�PE�' @�戚�g3B�M<��#ΤDɂ�"Y�"|�7O�f`�⬋�ޖ�I�F}|=k�튀��	Dk[�)��'4�9��(R�F�qӘ�D!�Ӹ=����a�/CXP��	W�B����CX�h�G�ޑDkV S�*W2�`�pT
3O�PFyr�	������iK
��8����@Ǯp���OZ���+�.A��B��O� 9�&� Y!�յV�~X
'e8��Ô���S!�=�9k�l3�ʷ��!�d�<[t���LB;���2a]$:�!�dN%�ZE���մZ�BȒ���!�8P�(Z��Џ ��tۣ��x�!�$�3%2�DH�
 '�X�jD�ȱH{!�� ��80�tL�!Q�\�V��u��"O��M�IΩ�_� nV�k"O�r�
����A�Y�U�(��"Of�jk�?d��A��R�T��"Or�zWŕ�Y��X�#_Tr�{!"O�����dVB�B�ߓ*&��4"Oti�%/��$Wb�(��L�6���"O���4ER�)����<STdɦ"O�-z�"�6m��X��FZ�dC"O�Tȅ�͇~�4�k"hK��( �"O�� aLB�u4S!n�*�<��"OR�C!�/{{�SO>�U��"O��a��U�������ҁ�"O���4̕�I.��S�Bԋ_����"O�����!�6�C��$%Y�@�1"O>�C��D����0�;"倈�"O��!p�̻X� �cV�1S�� ��"O&��C�\�4��լ�7U���0�"O�l{�jݚgE�J���6T4"O>�`"e��v֖R�l̺ٖ0��"ONmrǈ	)a��d��[�0y��"O(����31�i:�k>tC� �#"O*��6b�6x�l���jV�t�`u"O��r�I��p-8�󲉘P��Yc"O�e�0�,fP�R��i� i��"Oޝ�/l���d�t�p�@�"O|0�B��q�NL�qB�@���"OpL�v���\�\�*���"/zMaC"OxQڐ�%i��00�!�3>�*l��"O"K&bX�~�uc�Ќ/��c�"OX��0�0[�����J`�r �f"O�8h��߱(�`�d	��83]��"O��ڲ7�Fr �G2�H#f"O��zЕbY���Nۋ�w'*D�+3��p��Q ��H�wH�1�)D��3@�C�I_�h�l�J.����'D��pC��qfT1+G���87��sbm&D�D�䍄mv�#ѯD�rL��pf�"D��z��*N�y�pj��6�x[��!D����AP-F�V$ha�?m��0h >D�dY[�p�jV��&c�j\!��.D���Љ�4#�,�K1��W0|��-D�(�A�J�`	�p��%L��*D� d��)
�t�I�UBH@H�"�4D� �T��l���S��0C�$�N&D���pL��o����#������0D���s��j��c�/ѓ�e3�L*D��v@�9[�p���!�[f�)��&D�,'D�9�,5q�.O�23|��&D��JB��8y�P�p���\�N	��9D���#��	$z Ђ�G�
����Ro6D�����_�Ři��#��CT�4�l!D��Kэ\�a.���E�w���h�)D��4�8Uq�L9��Êm!�M��#<D����CT������B���%&D�8�A��Z�xR��*f,81�g.D�D����#Vb("Շ�
t,��bC/D����	�QMQ�ወ,� �c��?D������X�Zĳ� �:(Ԭ��(D��)$���\���aK��q���j'D�0��A��n}F�@��0���&D�|�C�d: �(���4-�&�Y��"D�|ڡ&^�x�&�؂���0��05	 D�������Ra� 4�]z��?D�� ��R`�nl=�#�7V�N���"O����]�s����d@�Eþ4�`"O�y)$�^��1��N�� U8�"O^	I�`�55,�c���4{���f"O4P�Ō�f�~�3�$�.
u�S�"OXe�bJ���Z����@�;�����"O�	��.+Y����G��eQ�"O� �M�M�P���
�6�j]��"O���7�E�I�5	�%3�N��0"O<�)���	8������K)�xɁ"Ob��⏒0<��B�����E"O<UH�섉lVDm��e�9h�"ࢧ"O�XZ��.8ؽ ���&@:��"Oj�3��K��c�I�TQ;"O�ij�G�9r'�{ C�1Cm&-�t"O�]C�*%S:<1ɰ�V�$S�ɂ�"O��@f��nF��bA�eJD� "OV��ρ?}ڎ��D�߽!A��f"O�Չr"��!ӦH�D.�A��"O�E"�ɘ|y@H�`M7�(���"O.��3G�?C�J��g�ߔ(�L=c�"O,m{�Q;<lty�#K��u"Ox(k֊2u�� ���V��[4"O��"�]*?�n�X�k}�TB�"O:xBd!��8U���TQ���"%"O@�6�ԹH��Kj��U!4W"OL�k"O�g� 퉵*߻`s|��t"O��X��	BD	S�@�5)��eQ5"O�݊'�q&e�qϝ�sT%A�'0��W@��V:P�`֊�%��k�'�p��c!�;` �����
.`P�'a8<*3g�4������?f��ec�'�|�˖�R�U#v�y�%]�b�̐
�'�"P�G߇4.0����=`�n-�
�'f�hB3��v��EScΜ D�!��'��9��Sy�@���#kz��'�(�A��2�@H`��- @���'�(z�"�<B �%�B-ܝ-���p�'����0�\2Y8n%ౄ۸YxD��
�'"F���0Q8ݓ�� ���'��d��d��J�� Æ��ְ��'h&@i�
�/�@i�@�^�����'>)��ױBF�A�ާ%�ظq�'��P4d�ZZ�M RN?#��ty�'	�;ǡ�&}@��f�1 ^~�c�'�;��9N� cf�+�l\��'��uy���Kh<����|$���'H�9��C	J5.��ݬn���:�"Op�;$��[���)C�R����"O@�QNO)1��iA%Ɉ����C�"O8� GYn>D�5��zO��"O��x�� jؐy����2B2�bC"O��d��:;u8�3 �n-�pf"Od�+b�W%X����Bc1W���"O��#	�;������Y��A��"O��0����DYBH �̝3w�X�"O ��G��\42Px�ˮdZ�\Hr"O�S��42BT9��$�e;�@��"O��ꔌ+��U�b0� ��1"ON@xF
��X�p�;G��ja"O����'U�7Lb�&T�<����"O@�8��
�[ ��`k�,V��!�"Ob�5ɟ�{"9 �#�
0���E"OĈ����$f�P�ɀA�� a��"O� ���G�"
~v��!H��"��d"O���F9���G-;��(A"O.<���=>�8M(!ëk$�	�1"O0�W�D�T�"�	�.m����"O|�G쌽,%蠫��]�(s���"O�L���Q{!���@C�e@��"O����W��Qp)��@Q́R"OD��T$��r��E��(]Xq�"O@u
�h�6s�]{�B�2G8�"O��I���+v��}���jU���"O���b��KH�9ڐN�S%�x�T"O���
�S 4���,�&�1r�"O�X�A�ޖsT��2D቞���R"O�p����F� � τ`�p��"O9�&�V܈��	]�g8�2�"OdJ�Үw��8�Ɗ'��"O��#D�~O�}*dݷ\�8�B"Ox����+��52u�ě��]#"OvLfƅi��a@� a�BP"O�$0��<5T�|ðE��3���Q"O�B�(�%;��;��]���2"O`1�`��q+�	�f,����"OF���晉�dhX��66�bH�v"O��٤�0�Z4��$ڿP�XQ�"O�M��*$���V��0M	0yRQ"O��e�!�zM����	���"O>�u(ȹU���၇̾fE�0"O\\�bƙ�t0AAG�c�r��"O ]�1	ѕ@���b�X�p3Rh��"O�}3`����a��REC�"O�bT�6u�\�����B���"Ot�"��VGM���`��$���u"O��`dBY@$�P���9�9��"O����K�~W
�QR,(ע�0"O$�k�MF�I�P��%�ӿb��)�"O,��/@�!YA�f�y��AQB"O��k���^Ͱ(j��![�H�C"O4�1$��Y<-1��3L�܍#�"O>���ƙ�^�أ��Dp���R"O.�H+I�D�m�$\�J�1"O.�i���#K�z���Xm����"O�a(Q̍6���.ZW��C"Ol !���=�BS�T�N:�s�"O^@���?jf�X�%ݪ(�u�7"O�UB!��E��R�e(D��"O�	�@�v@}�#eQ�T�Ă�"O�%����z�ة�7�]9c&$%�P"Ot�VZ1~y�Si݋��zQ"O,�`�I�>�=Hg'�GHE9 "O�4�C�L-D��bئ.���@"OJa�%N��E��� �E�U��d��"O,�Ʉ� �V�,�A�J�3� u�"O 09��CE_�]����!O��c�"Olx˅?	#��o,!�"O��
�
g#�X��bi����"OH��f�5����W�[OY��e"Oި[���3�4��֏UV9�	��"O\��6�M�G�jƎ]�8��a�"O��P���c(:E�l %O ��!�"O��&L���y�e����$��R"OలC�?n���c�*G5? *��"O(���aS	#�6�30H���ebv"O����$���.����0#�\���U����m1�2p�=<OUs� (V�"(���\#�Ѩ�"O� �5�#�<W^��E�Y�0�Z�Z�"Oڅ	f�;.��Ic�����(��"O��FNX�#�6{#,���M�B"O��#P&ߝT�p���c�*}��"O>��i=w�I��L�EHB�!�"O�P�3ǏP��ȟzSDش"OB�U�L�e\~�Y�oȡK<R"Op��J!%Ţ- �՚܎��"O�����nIRE-J����F"OTD I�#	] ���M�2%ĄH�"O���dͶSȆ�;F�H�K�l���"O�p+W�)+�yz��9O��x��"O�8�Z���b�@�iy
�'C���2�2Y¬mJR, �?��2�'��pԫ�;��a���Ǎ �ʝ�'�fd�􄂓s
�%���Y�\��̠
�'9L�C	\Q���I�6Na$-��'��UB���1,a"q�P�.��'5P1C��1InJ�0@�9y�j���'��)�OG*[���%�b�'��s�Q7\�jF�ЖL�:d��'�$��J'�M��~\�y�Ks|����B�a+��gș7�y�C�3P����:0~n,p%:�y�,B1z}Ҕ���J/"��kӠ4�y�0�ێ8�,�Ҥ&VX�\���'KZ�GK\9!��(��i]��,��'F,Y��U�&j�l�w���Y��%p�'VXHy���B�+�$S����'g�0��¶ʮ0BNA��N}��'s�t0�(�ر�tD���Q��'l�Q�p�W;{���g�5{H~`H�'�D�i4	^������w�օ��'�6���5Y��`�f#V#;�0}C�'�Jk��Sg�MY&�;_�`�
�'�d��䌌16&	�`
�8����'i�@Qc�u�QB�'��*�"�i�'�,� Q!j�d��Ktp�H��'"d���S�h��A,ܧh��E��'f �d�XY�H�۰.�("����'�nV �2Wu$Ըe%T�,4z�'��]sV�+��}P�K;:� �',��W�BBF��4gK�U���'�.%�-�#�uH�	���K�'��	ն� �z��	6Nej���'�f���%�
�P���G�^��'I^X&1F�����gпH�r�'��x�p�ʥR��l����-,�0��')(���f�eI���p��".��'�F�Z�WE�2I"�(��n:XŸ�'tY;@��@T������n�8%R�'��x�D�1�.IK,x�"�.�d�<Y�h�3rr�1�d��|�"��H�<�7+��-p��YGcކ+e�zb�M]�<I��jK��u��<4{���0F�\�<i�C�!ZM:Ģ�ޝ7%Fx�!��`�<� ���}��}SX(��ox�<���:ʼ��Q"�l���-�N�<pA�4�\�ze�G�F\"�iLq�<��"^(A��;f�������S�<�%�%� �WO 2��miU��m�<Yu�e�`����A�N)��Ol�<�W�`k�aiĄ�W��©�e�<As��!��U薦�O��B��<� f� c$\0y���Gw�"��"O�b$�Z�&&p�3�?6��\!�"O����׏"�� �U*��4��r�"O�����/wqfQ`�&�4R����"OX��,WT[n��� �"�䭘�"O�!�1��6&�*%*����r���+$"O�V��!iI�I*B�Ӊh �4"Of��a�zX �ۣr�V5�"Ol�#��6�e��M <�$�r�"O�܃�f��}�88,���ah�"O���� �[���[B�N;dE���"O.�R�ơ/(԰�`O�~�z9�"O��b	��&���C������"O^Eh�+S�MX����4�z}��"OE�6�T;_B�6˲��p�"O�hA�mB4GY����c�)���w"Oll8�7{>�SţE�r���"Ol�rǍ�{蒽�$��uш�y�"Oj]���%�N���/M�R�̒�"O��
���Rj��T9_&�bw"O��P.W�Ѡ�ҞFޅjW"O�@���
f�2�˒�B���h3�"O����)��Nb(Y��O��:��'"O�Ռ�>|[����C�5�ݚf"O��Y%��15�����j��%B-k�"O�B�����<:ǪY'g2��r"Opt��ɏ�$t�7��A!���"O������N�9�㰴�"O�����O�~1�b��;�0�u"O�9��أ0,�%�ł�U�Ċ�"O.�"�,ޠ~*
�J��Y;|Q�x(�"O�UkD��>e�+D"�9A��&`G!�#9��%��J`�dD0���!�d�7{� I�+T�`7��I�T� �!�D�_ִ�Y����<̮�I��	}�!�D�@�]�7YO,���u"�!�&R8f�{�@̧- ��;��^��!�[�.��� �4\%��)2z!�dI�f�Jh �,�
8|౒�ٶW��4�R���|� ���|x�R��m��o�[�<�q�_���i햝_2�!H�<����vQn��I>E��oN�;��Sv���0�����y��
`�@��2~�> �A����R td���	 .B6���X�j�,ۅf��ӧ�Y�a}�_2Jɕ)��3��� rB�j EP	:�
O*��!�Y�+�1� )K�,�~�S3��/<��T�K�4�$`�IBv�Si��kP! �/4��Iqcܴ&�C�ɳ�v� &��$ �������F<i�`."��L �B���Z�)��<Q���<  �Q�d�3f�B�J�A�<��.�j�@S��9t�����ɠ�:�@%��.tUZ�A�Z)>9��3�@~�z�c(�V�"�%�$j�|��I
ْLP�n�7 ��\u���SjR�t�*�s�i*���Q|%a��1�lA�CeJJ9�e���'Bh�§�Y.��ѱ��i�(�:$�~"rlP�(�N!>��"t�m�<���9%���礕�j<ܰ���
p�j��U�˟?�ZH���[q��F�T�Ozİ�`�n bB�ٻgЄP@b"O�$��eъl3@)֎Q))"����[�i���2��!m��&�{X�n*�Et�ٚFG�3G�|e���EY��i�퉏l���%Em
�U�ѯ�.bE�5�L#<jn�q�I$%}� �V(Fd��P��.ű2Xx���бz�LX�7�IS���AM��TG�a��K 7G�D��Fd�NZ�b�A����
��v"O$������W���l��f��!��I�K��zA���H�8j��K�>���=ݤ�2�T/W��0����P�>B�I�K������L��}{�'Y�`{t%�pͮ>Y��˛}I�٧�ϨO� �(�h��	h'˒6uZ�Y��'kt�U�A�mX|Yjp��i��
D���u4��ق͇E���Q��Az�*i��)ȑ+4x-:1�8�uE�3���y�'?y �%I E|J5b�<�H��)D��A�@���i�S�]�T�e�Tè���PF��jmB�I<E���O�d��2�M��oK��S��;�y"�Ō!�l,1��[�%ZH�C3�����ɗ˴���nN�p<����g:� ��	(=�d�o]��Љ����|�1���Cr�1� N1�2DG(\ah<�G�Ѩ��uB��D�`��}��r�'F��C��n�t�5D��
0ܳsj!f�C�I3j�䕒��է9(���$��C�Ʌ$�\�ґ�Λ/������_`(B�	�?*�`�%�?�. �F =
B�	
Hj\����/��Z�2ep�B�5$By*�����N|�a
�Z�C��?B`��ͼf{F �5V�dB�I�[Pj���g�B\��� ՜$P�C�I:S�B��́�`@~�!�.�%��C�	�F�X��A_2V��q�*�B�	�2�m���ď|�x�"�=7�B�bz.�۶�9b�!�5!E�CT�B�	)4Ƥu�֦Z?ji8���-nC�	*~Q�9#p�@�/0@Y�iJ�.C�ɼT�������ੀ�b��$C�I��^�b�eB���L��#S�B�$s������&�R�Aˈ�'ˌB�IS��c�zs� V!ˢ4�PC�	2J��k����9nU����O2C�	
fx��"f���2u�r�]-$C�I�_IY��T�9��H��պI��C�I3waX���@A#w�(��P)R�tV�C��@�Ɛ�`+��&�h�t�E.bB�	hJ���BK�"r<�|��j���rB�	�r�Zx�Wc�#�,�R�O�QDB�	MU�zĦ��~2ZyC"�OAvB䉚O��	�%��(]
��4�@�C�	,�P��,'{����o�w��C�	}/>��v�Z�-��\�E�!}+B�IE$�A�)���C�l[�n��B��w��9G�R�]?z}{W�bw&B䉀v:��F�M7vD�'/;;�B�ɏ#��|	�*�=�����B{vC�		e��I��U�J"���� )L� C�I�f���� a�8g8�y��@��T�B䉠q�`kI�C%���D�$�B���TÆ���=�xTT�F!;�B��;|t��Q���=�p��;"��C䉃:����d������?C��C䉿 ���0��O"�3��s%�S	�'�0�s3���O6.��fbE�znٸ	�'����E.9��;wl=l����'�rA����R���C�h�4d��M!�'h±�e��h�1���Oߨ��'���a���g�^���A0H�'�-)���(ۼ�RV�@3)J�Q��'Aj�%mTZ|���p���՘E��'/�U��N�1K�DI!^8�����'��h�0X	Sz�%�톕{����ȓo;���`h�0%Ҿ�9v���Z}�ȓ ��5�TA�jCx�RE���*��ȓ$"�c�:3����g83�2��ȓl�  WD�
(��K�m��1�ȓL2%CR�:K�:�Z�b��o�R��S�? �	j@� 3%�8�����xR�d�W"O$\R�"[���j����-�@"O��! S�O٪x�A$̈́xӐ%3$	�=B�������>RL�5	1<O`XuȐWP^ �G�@��8�qD"O��A�i���m�d� C"O\�p��)���g�R�3���2�"O�A)�<�5�խ���˥"O��J��R�]z������&���;�"O4��wDҩ9�J�в��%(fr	�"O��0)K�
�x��� �{��)xW"Oj@q��C����U�0�L��Q"O���G�
��7%��IP�"O�,�0�)����Ey�X�Zc"O����$�x��,����<{�=��"O���-�X�Ti_,�W"O����*s���U����"OH8����"�$�!.�e0ph�"OFd[��I��$�̃`H
89�"O�|3wI]�l��1�1,[EH���"O`������8��t�ҥL16IR@"On���H�9ON�"e�����"O�S(�}!� �Q�^F�>��v"Oh�5ɉ�E!rl�C���@��e"O��	�i�;��S̘�X�d�B�"O��f��-aP� &���3��5j�"O@�14䅖zp\��r�O�O�>%�S"O4�+3MJ�}K!(R(P���`�"Oй0ҤM �D���Ѓ`�J��"O�YY��I�N ��ˆL���L�9R"OȜ�q��{">�K⪌�����F"O�+5l��y�"�1!��0b"O��ҡB�4�QC�Ƀp���`F"Odk(W�9����F;c���)�"O�IY#C�!s���æ[�V�����"OT�EB�����'w���"O�,3�k��a�D|ɑg��_�$ب�"O:06�M����iAb���""O栉e"^�f��L�L=OFqZ"O"5��lE.�U� L\�a��	�'"O~Q������ 
 �6�P��@"OЈ*��E+%(v�{�o'~�R�R"Otxy�C�%X|H�Fo�M����"O~<Qg�I-i��������|(�"OzeSv���y�h{B�:Xh��p�"O�URB���b|��m�\�ĢA"O���.K"A��t����V���"OzͰ�d�x'�0�GV�GG�I��"O~�eA�Y �x1�+e��"O�%c�N�H��� ���.0�X9B"O,��1MΜ{�QI�@X��E"O��P�旆�X,RW�L�h.�� �"O��Pw�1!ܔ!
��4_�Ĳ�"O@)葢_3�(	(���}|���"O��bs���OC��{BP�h��}HE"O�ӷ�AM:� v��8Y��xXS"O^��Ù�#xzS#�3V����"Oԡjg%J�;�Ɣ�Cn��hNb��#"O�<1� ��[)z�[�#�[=����"O|�j��x�S󢊾9�J�+�"O�(����%�^�� 6>�}0s"O�	b*���n�藢G.��h��"Of�g�rBp�!c��s#"Ovl�u��H�|��r�V�PZ�"Ob�����G*��Rr��1���0`"O� ��	��*8�8:��A��̺�"Oܘar(H��,)��I $��)Bf"OT )`!Q.�50��QOi��a"O4�)'�7>Rֱ{A�܉zxp�"O��  �&@�"LU\���7"O���D)
������nA��Ѣ"O�����Չ9��m�M�)9,|(�u"O���oIk�\%sː�.m�A�"O(���	�|��l���
P��:"OF�"��5��pG�V��t��"On5��9O"�J�!�>@d�"O&��� �H0���14��A�"O���ʜ�`�pE"pM+(+n,�"O��a"mޙ#n<,����(!�"Oly��(��D�$Ҡ���.����S"O.t�pi����A���Ix�8��"O��;�F^ m� ��ӣ{��l�t"O]�q�]�?����A�t����"O[��YT��0���%��>�!�d	�S^ZTb�dA�e)�AcA��3D�!��
�^I[�Kر ��H�L�#Q!� !DY�Y0��?!�>��e�],d!�êJ�d�eOܛ~�8<zAf�N!�^#8�"53��1=i��h�=!򤐁BH�0B��a�\�-�	_:!��26|�%��3R�x �U�
�5"!���BcșҴ�ԵKnQ��)X�M!���|7F��A�t1d��h���!�$sƠ8���L�d��P�ح�!��]����������t&��C�!�^Q[$1P�ϕ�9�`a�E�%�!���
A�]�O�FԂ�1�ùn�!�� IJ8���kY�}�D;0 1n�!�d��Smt�@� \�����.,�!�D����Xɵ�."S�Ar"�,*�!�$ߨXTb=��AJGn�a@C�s�!�D�����T�
���z`n��!�$ʥ3���'�Z�|��8��ѿo�!�dH[�b	p��
Hpr�a��gx!�M�N<� h��o6�\�a
J�p`!�$�8_
<Ț�씺C6
B���ca!�ē�A}�{�Q!ФZ�M���!�D��*p�93�[�b6KҰL�!��)�����U�^�8�t{\!��:P_&�b�8M�ܰaOX�U<!�ޠq|����>O���e0"!�$��ip�P�M������{!��1q~�"��YN,��
v!�$Y�[g(���*f���h��N7U!�L0|>�X!�l-hf� "0�Ȉh�!��50��y *t�� �&HQ!x!��rr$|B#c���	��(Or!�Z��8��#oۨv���ㅁB	m!���+;NuQ��K�Yb��f���M�!��:)�`�s�Ú�\K��s`G%�!�䑃PM$u1��.!�e�o�	t!�DP7\d����f���AD�'qc!�$j?z�㰍�1ٖ�f�<eT!����$�W��1(����
F��]����̒�.��v+���#�?(����"OH�aï�"��r�
�h���"O@89dk.K��\ �8i��	�"O�QW"�O8:D���yI�p��"OؼSE�ME��]��&�V�:M��"O� �8C ����T(rl�%�ؽQ�"ODr 	�r��` LٟA�2qp�"Ob��U�G���2�k�t�n`�"O<YA��?Z�a#$ŋ�t
9�"O5"��X}2]x���[WF0��"O���	w��\!���4��x�"O�D�B��:�FūW+F:Z#\<��"O^d�se��!��$i��/�d"O�TI��Ԏ6o^=��'����W"O&���/IKQ�q#E&�V�>�)�"O��Ac��*!|�L2�"+nDH�S�"O>���Z�Y���d�M]���"O��a��_ :ʴ�%�8W�I(w"O L3��!3����M^��M��"OL�V��m���'D�P�Č��"Ol	*�0R�(�L�'xٌQC�"O��ɚ�;��5�� ��,��[e"ON�zWɆ��rS��7Ny#"O41+�Ј� ���a�0O���""O��� �U�*R̐�@�Ӕ���'�R0��F�tД�⇭
y�,<S�'�@����׺E�������h`k�'N��	�"3��$X�X&z �p	�'�r4I2❆!	�)�WI` QK�'C��2�n?j��M�v�������'Q��r�	��0�B�!L%�`a��'��ti���	~�J$� [�9[�': !i"�ю\ɣ�֒]Ǫ9�'�H�;�P	�&\!C-�`�<1�'d6 #3h�K��-��\?SL� ��'�̨S���|��i�. �Gf���	�'���	��G�I��`S��S�&�	�'^�I��l�9�DL�a�V�4`�'��)�F�a��i�D�;Hi� Z�'���H�"\>K��������'�H����=�ڐq���
A*y��'zd��$��;0����F��@ĲlQ�'�Z�	�g7~�p9AL�2:b$�
�'GҀ����N���� K�7�ҭ9
�'[����&	ʡ�F,B7���
�'6� u��(q�(�ɑK�)�F�	�'��$K�5A�E��f;,��"�'�.]�QÍ[�|��. x�'�<ӡ�E�Q*��aJ�
?r	��'o�h��B�<v"`�F)	S:B ��';DpI�iV�v���R����'��}����:/��	���21d�J
�'�䅉�FJ,�  A�+��AV6E�
�'�	����n)�,Y����Q�q�	�'�НЮ̙9�ʀCRjL��!�	�'�&a��Q�Iښ�B�?̮(��'Sj�J�Խu��4��oٙ4@!�'
�ݳ#ֈN[��z���3���'".%`$�$@�|8RgM�?~2vI��'���3D]�W$�F�ּH�'L6`��$4`�A��,ݡG��8�'f�8��A�V�0�?9�fy�'d�=��ǎ;�Ԍ�VhA).ƈ�0�'�u�!��\q��A6��&2�2\�
�'W��'�ֵl�``��-0���	�' FD�Si��x1
��Z"%��=��'�t��*|�@���9`�X��'�D��P
 ]G�X��,�z��'�=ae�Sqz�hao�<|�N4C���  �hRaچ_Hڴ�4a�S��-�$"O�P(�H��*�4h�Z�D�ك"O� Ɯ�tT�l P�~]J�Q�"O�L�ӌ�9�HP`���9\L��1"O��x��ۆ�z9�&,�f��-��"Od��3�*��U�#l�T���d"Of]��$$6�T����q�S�"O��y��ωT� ���F�@�"O^�`��7�%k��9M��mqb"Od]���3 ��
 �Q��r"O�!����'>���K��S<�����"O�p�ǅ_�8���R�ބ^sR(8C*O"��0`f��R%���H�T��'Z�
�I
�}/�h1ր�,s�]*�'�(QJag�FV�$�D�??�Ȋ�'��I��T�t���4k'���i�'v:���.�ҭCR��Q�T�K�'.�M��ѭ	�5Z�#1xs�T�'9���l��w������B&-�(��'H��#�iÆ�r!A�U�����'$X��B����Z�S�iHK.4-��'C�)�I�@wBU��I��~h��'�|qXW�0�=�V@�3�@�
�'�>��5�	_M.)Z�f�'xĮ H�'�̜K�N��pBf���ޒh�T��'�ڡ��J3�ڦd�,{&A��'��Tb�W[ѼTi� T�p����'�rMpT��!c��qbU���e�.�R�'g(�y�d
�h"h����J$� 3�'P�yG���t�08T�S�@d �k�'��`�K��X눜c���;�h��'�@};��Od(J�`�ߢǔ��'=�l��n�2����Ń�4���(�'qn4 �N�enXlKL�0N�œ
�':8���(5D����X.(�Ub
�'����1��(YZn����(hA�
�'�x$xwo�;X9�)����&�4 [�'/�t��M�/2+P�����/cT�Q�'N*��7 ٯ�`a!aٴu��EZ�'�~ਕ�ڵM�>M
A	�g�P�9�'G��ڃ$�-L����w!�eB�1�'��p�	B� A���H
H�A��'D�DVS�8\�S�
�98"L�	�'���b�^�/:D�O];7��	�'1N��L��Pb��Î>.�.�
�'h��V���1�f�)�љ�'���åM̈ft��E1!1����'�x#2��+UO�9a�HND|�X�'��I��"͒�R�i��?;w�4�
�'�0|23�m��SDf�7�$y
�'4�X�$�R>TDʱX�)��e�'�=J�(�$c:�YZ�"�%j�\r�'R8H#6HU0<�x�vً-i`���'7����)d�>�@�[��J���'�&�{wg�l���*� �>I��'���ґC��C ��ʥ ߷$�U��'O�Jt�W�#��e����E�T���'��M��$�$F�1�㔱<cJP�	�'�n�k�`Z>I3�ʕ-Y��
�'�|)Aw�ژ}�H%�e\�,�e��'	��������~�R�N<;ڸC�'�t�!H�R7�ɁC��7#��8�'��kc&ʇ�\zs %9��)�'��Q��%Z�� I`H�\.��	��� )�Un��o<��)7g����("OzM�E�Y�jF��!�|��J!"O�����H�&��Y0���?�~M9'"O����;+�@��QW����X�'��qA��JY�����O$v��	�'��!%ѥZ ��[G`	P�k	�'����(Ɩ���1M[�7���'l��kw�F�uv�ԭ�*��A��'��֋�	G{j�z�*۷9?�-�'���3Ѐ�� s�ޜ{vZؠ�'2��¢!G���狒n��}H�':�`�ЇQ���Sg'�/kcl]B
�'Ty
'�A+�r@צA�:���
�'�䠢 ��rɋ6��I}�	�	�'��I��L?B�Ԁ��ŗI��<	�'�xHV�Y0� ���ڐr�'��5���A*�;0�=0枼r�'�b�3шA2�^)�A�*��8B�'�
��toH�h4 �w�'H��'¬�v�ƴLx$৏M�$:ؐ�'Vft��fɳI&�+"�(P�N�+
�']<𠃂[����ËI����'�P�ӧ){��a��l��F�v���'�.Tɐ \}˚⭉-߆���'� �[b�CZ�q�$��'1h�@�'ۢ-)�i����{x�y�b;D�<�A��hل)U̬��|�s*&D���#Ȕ�GѮ�d�N��h��L%D��Q���*,&�c�Č Ai&��D�!D��q�E�`^L��<e[1Ç�!D�����CVXH��8a������ D��K�\����H
U�����>D���Qiګl�2Z��D X��E0D��a�1�d9�_��
�3� D��Qj�<O^�آm�8�6-� �=D����m�5,��E ��.0�.���
!D��a��L�&vzub%S+h�"��D!D��r!��;c��iۥ���Z��@8t"3D�,��,_�xa�xR�V�=<�,�&H/D�X����;~`ؕhn�Rj�H,D�$@���4���@gm_�!(����-D�(�],N�"ɦ��:�B�bcn-D�`����?��@�rKI&���� D���\$L�1���Y <��2�E9D�T��N� `i�$�r�RZ��i�8D�$�'
[?FH��"`���f����:D�ܹ�؀l���R��W�yx�qg6�㈟R���B
Z<0�ڢ�;#[*��"O\�xЈ�1g8>D�Pd�0!zՉ`"OT�"C���V���Q#R�;r4�G"O$`�R���H���G���5�"O.q� �p�f����?y8 Q�"O6�(B+C�6��]��g��kr~�h�"O` �@R�d&piŽ�ÚYQ"O�1J�䍎"F�rlK�\��8�"O��V�̏B�p���	��=ʡ"O��ª�<{�%Yu���⚨��"O~�
���,�𬈂Ղ1܊!��"Of4�B�zr<Y$�{��y� "O4t!�g\E8����7P����"O�dH��	�Y	�<Ц�ϼ7�$��7"O��I��
y"�|�f�Y�P���"O���R���>HR H�`�<=��8Cs"O���C˾�(�P�������"O� ���_�!��Z�.�Y��"O���uj�c0��� �)p�XS"O8HCp�
V��W@�1~â<	"O��觢����������"O�H��o�.��űvM�*� 	*"O��9D�?�Ѩ�쐐3�H���"O�{�� �� ٲ�N�J,�)5"OH42R�P���8uȟ�FH�3�"O<�)�0E�8�ZR�פ'||�	�'����D�ԑjNF9*2�X	-��TH�'\r��"*J���b*�p�Y�'��i�t�X.fg�HJ"!O<w�.�{�'��ReB�W�BT �=Q<��'4�L���ql�x���x�N� 
�'���N�
GqtM8���qzr2�'Ϯ���,Y���4��h6��J�'��8p��i�v���&\0\4,��'��p��(|�: ���'$��'<,�����K,��%�(M�:͙�'�ށ�Vb��s�(�!T?�p�9�'��y�[�A�t8��=U���'m��`l��9Ǌ$B��D��-s�'��q�k"�P�a��B5����'�����ȓ��ء0a��7���2�'d���:h���#Bh��'e�A��'b>]����> [x�� �U�!�x1��'7��A��E:MȮ��A�1F���'["�ʴD݊?�9Pfb""��j�'a��@R/��(�"W'�XXq�'���I�)	�8
��@
G���"�'JP�s�$��	�i�@� �*c
�'@$��f�]�}8��Y���4�hY�	�'夕����"Ѐj3%Q�L��'�`�r��>k��S�c�1k���'52�(��ǿ����i�����'�n�7�O$::XK�ҨI�~h�'��-[������	4*!�'������M�ܐI���#Y�	��'6^Y �A�98��ű�R�Bˏ�y�O`�̍�����^���.�F�<�$�I2<%L "�鈏x	��Q�.��<�����4,�K�
E�k<��+gÕy�<I���'�B9h�Xp��5_���ȓE�,�rP��}m��Q���9�h)��^Xm�rGNX}��e��5���$D��#$���Ǐ+o=@��C��a%!���`�5�×���Kdq!�$I�'p�Lq1E	�t��u��/GV!�d8_a�ѭ�6�2,c�� x0!�RЕ���#H�ظ�mX�V!�ć�$�J���-��-�^�	M]	f�!��)��5�h��1�:|ٴ@804!���/2���r`
�;𪉃'��6M!��4Y�慰�'��H�qr(ǥ\!������z���7�X� i�0'!�d̞�^��G��:w�^��HY�5!�DԔpx�����+N�@C��Y=w�!��W&m�lYR��C:Bw )��FS�y�!�dE*�tQ���.��9#g虴u!���;��Q�V�U� ̑���:/�!򄈻%H�r���z˪�	��<F!��W7#)�e�`�D:dR��Eis!� b�a�	�uI��Kg�˭ �!�d��!_F�kv��+�؉
t儮�!�� n��g&,v�k5�Q1"O$�3���:"5��z҃O�T l�J�"O�C�տ[%@��dE]2F�P"O@\�R>%�8e:wA0T(1�"O��C���W\����ȕHpc"O�c � 	�g�Y1�P3�"O�V�}`a��G>� �)!򄄛1��8����y�ʄٷ�׋d!�(]�s5��w���j��S&S!�ֹ7���+"�͡��I��[)!���i/�л��ˍX}��r�=/o��䋭�2���4���s�􈤷%me��!�f��i
  'KKH6i�U�����U��@�v$�WA1�S�?�NM���ђ�.\f�E��[�#�����>R���I�(zw���r� B)1"�o��GR>ט'nq��
Aj��p���e
Q'75W�KqӲnϟX�O���M�Ц�%\?��p2d�������
y?�����>�4ɐ�\RA	S�gWдw��r�'8�7���E%�dkG��Ԫɔa��Ȋ&��4nta�$@��	�0�h��4ݰ<��J�to�	�����_��q�(�:�v��t� ;������,���On6�Ex�c�5�d����]�7�����BfAP(��r���Pm(N��誟^]r�(�^����i��$��Ä�|�d��!�>V��dC��T�?�glF!�?���i������OP�drӾ��1"؃<�$�Qi�(KƬys"O�k�͍,�~ �A�Y z&pj�X0�M��iL�'��d�O��g��%+�9:�̨ ��Y���ՅVLfΑ���ȟ�
�ZzFLq��M2T�V�##�j� � �#�gy��֪[�Szٵ�	2-(��ʒ웮VDf�1��$p �\x%��Jт�������
4Ɓ�nc|Ƞ��&+(&�$������O
7�Je�h��%Zv����"��iK�D`�4�?�)O�$�OޒO�Ӯ,��Ѹ�D���`����CզB䉚��"�AF8]�c�ar�ɟ�M+U�i������4�?9����iH�_�|��?x�>}���b~��	dJ��������<B��@��� B� N�~��>PD@�C�B���!�*/�r�(�� U��<9���R�����"��0�U�g�.�b7.��<���D7~`���#�n���n�"��#�nm��П`��4�?9���9��E�"�b�AǍF/:x�lc�I��Mk��@*��<E�N�{�|-��a[�z��H�2�O�o��M�40���7i�Pd<�Qf��>q��h�ޠ���if�W���?�%�����ŀ<2�,�'���N�BS�������E�(Gg��1���0��!�J(�S�?���AU��=�B,�kбe̛��R�"�&� 2!\�Tܚ7m]�Qɸp�a Z�:V�#�˹|�1�.�h�DγN�6��˝+C��oZ%M���Ʀ�`�4�?�Οv����oԳ3?���v���ԙ&lĕ���O���dF�i��n�/a�R�paݟMjQ� bݴ8?���|��O<��hY��	b)q�hzC敡r6�h�	Пĩ����^=��ȟd�I؟X:[w���i�d�ItLF=5N�#�N��b]�	a�/L�q��p[�V���(*�!��f�iF�`�!3s�|"��B4�S���o��Myp�U�o�: ���1�i��� �p�a��j���f��\�H�@�����c,_-����� .%r�P���?�"�?�?1U��3[L�gyR�OD��9��\�`�֮fn�1�J8Bp��G{J~j���la��	�!-A�'��6'6\⦍�I��M3�>�e����䧏56�
�] |  �    C  '  W  �  �!  *(  �)   Ĵ���	����Zv)�ll\�0R�P��
O�z�V ]�n�1���2�����ӊ�y��D_�~!�$���dJ��c@�1q^���)�!E�n�u �,4|�Sf�����ש�:�h䈋3�$��E�f�h���ҙAiص�c�F^6��5��s+�-xW _�6��a�$��R�2Qv�ُm1���	�RvFL@��A=AԄ8[�L�/�� KY�W�P��Nǭ(��h��3;���{��'�r�'�Rk�~�F+<p<�n�����a$�R�
��ɫ#ך("'��H��Dkd�	���!�(�~�)vB�(&'��h��
�<�b쎝iʧk"��C F�F�XX��d�����A"d��bMo���0�����LJߴT��<����~�]�-|ȑ�'!>%�Ip�HZ��y�A��A�*�@��:�:�CVS��M���ɤA�*���]y�m�ʆ�i�dE=�%XlH(/��d":D��1�ߥP@�+ՊX �$��bh'D���U�X����
�A�P��Q�P-#D��J�Gӟ[r�Ѡa��0@R��M D�pR�X�a��q��nS�|�*Ds�9D��Kdj��n�Z`�ʑ�ct�P;��4D��[6)Y =�
h� �k��{"%D�C�(�/-� D
D왂W�F�C� D�����<R�֌�A!�;o��8�%-D���A�T9�l��Ƅ1(-Ƅq�,D��P���v� ����bT�b�'D��C��� =\����1z��(!�#D�����;^y�eC����|3n���� D�DxS`�E?HI�v��w�hP��L3D�l���Q�H�rP��߹ DD[`G,D��
6��*���b�K_�Kv����4D���U��kcX!�Ƥ"����4%=D���nI�.�faڄ6�^ɹ®8D���fר`Qv���B�K!�Tٓ�$D�|��&��\�nՊ"�/\0��%�%D��{�儯	�v��u�Ǔ!o>���K"D�H2�dѲU����e邥%!�@�!D�t�W�Y=j� ���:h�%b�,-D��p��U����j��Z�H�JQ! !D����E�U��!��O1H�0����.D���ۼE�\���Ŵ<���$�,D�PaV!ԭ_��� �k2p�h�6)D��J��/Q'j�q�	]�Z��Cg6D�Xh�dZ�"-�9r��&t��X���4D�t��Kčl��p٥�[8���"4D�|�d��W^Z5�v͔�/�Δp��<D����kǱ	
�`��1cg��cn>D�����2@]�)i�a��^��`�?D��;�'�+c�.���hS�<�`��ԏ<D�|`w/�)%6�aQG��g"���G=D��Ò���L����v�Ś+ D���S-�+�Vp�}r��YW��yr�� 1��j���x�Lj�K[��yr�W<@$i���r��䪧��yRjV����wm��V��牅
�y�J ,2�
�KʏQR��`�&@��yRCz�X2k��S�(@���y��TNh����b=:�#�y��7.�n\H����J2��
�yb���� �T���`)7��8�y�M v��`��8o�Y���(�y�Wod�trGP3	&�`�Ĉ��y ��"�������=0��!�D �y�G�4����Qj�� �TK�9�yB"��U@�R2	��?�v���2�yBI�4��h�!5�<�K�J���y�L8_��2��N��{!���y҉�4	���r)�	^T�Ê�y/fk�Y*G%�WaP�h����y
� v���G69.��	/�N��"O�8;�/Ƙ
*���ġл� ѩ�"O�G�D��zhڶa^2`Xq�"O6j�Ӣ��U0��ү B��"O������ZE���J97W��'"O���$a��Zi�Q��mO��S"OL��ʇ$H������:Rd�� 6"O^a�W�׃eF�Ԣc狨b�|�&"O:�xr �1p*�"��C
OJ��2"O@�9I;Jά(!�>�L�"O,Y¢	^6h��5��K��4�:di"O���E�]�b4��)�Z���B"Ox���9;֊���`�難"O�)�V*����p��pQ\�i "O���F� �,&�Ii�$�"<j� "O�"V)P1r���%B��kxE"O��p��k�%���r�lM��"Oɚ�ˆ-JŐ��� u�R�!"O��`��(
LP�+�]�}��0CQ"OX$S Bgle��囷p�v��"OdX��H�r�U���27Z���"Oht
faR�[�̌>'�A"O:��r�(=n&�x�`QmF$Ч"O��;��W�/�^�9�J�:Q�h�"O:�Jæ S�J�
��H����3�"OJPcv�L�tSs�-�� �"O��w�Ӥ6Yθ'd�al�]c"O\�J'��0764���f)�d"OH r�m��|�a��jı4��l��"O�@�p�BȤt
��Qf$ �6"O.�BS�0�z�B�-dIB,�"O(Y�f;M�$�����5�Nt�"Ozt�R�ыe�B9P�^1-��4c�"O�i��h��c��^�`c$"On�Rpj��a�x���اo�iIq"O<�� `�-��0�u�U;m�I"�"O��Xp͚U.|��@��/�\p�"Oz�t��O��h�b]�	��"O�u8wi�.>)�����w��"O���#�= ��J�瓊
� Lk�*Oޭ�Te|V=��o�6��� 	�'�DͲ�B�o�*�֫���m��'��)H�7>XC�F�y����'��Tl�!r��I���;k�0�'Z��T*\��@30,�,��X�'�D�;V(��r#�rR�_R�c�'��y�ү�;�<�5�TPgށ �'μa����R��
�gW�9&��:
�'�0a�ȃY�D/��l���j��m5 �X	�'y�i�̎#+�m{��O!���\flI�jU�먁�5.E���aΆ$n!�'���E�,O�`�5b����l4c����'O��b�U�~� i8�I�$���*�g	9`�\�������$J\���C]�;?2���!��I��yBM�{�2��)��	�ɶ*~-
�)_�9*h��A�8�!�đ$a�����fG��l��RNU�S��4����ӭ��8'
8� D�H�������|��(g왂$�&X)""O�.��5��y����4Y���/�iR�Yg�ǟL�@�.1yq��'�,�3/B?:4V܀q`��5%��
�'M,�1��ėL �m�U�OMC~�ʓj+oL}� ��&���0�WJ��,S���}��9��Ϫ ��z��%O��y"�ؙ.�V�h�4�����!8V� d��Dlh&�y0�
1�!�������g.?���XE�D�1�剙���jR!����Pw5�E�T�ãK���t�Ўx�`� 6�ԧ�y
� Nq#a��I.�Yڑ�^"��{v�R��!��*��]�.�!�ʟ'��O91O��"t�F�3q ���*j�f�k��'k�� p�������,P��0��]!Xvʼ�4� Q(� qB� �azBG�=1`"  ��7��4��ɿ��Oā��"\@-X�D�'fn�S`G\��V�t��(6� '�^P�<C䉦r�x1���O��pA��,�ʓ�H����#�l������n����V�"����J�7R�eqJĶtp!�$ETK�q�A�R5������RC�L
7\�,T���ڸzl@0�Օ����1�z9�U�ekb�z3��}A!��[}��;�-���3vDB2f�RK��^�iY�i�#�$�ד[J�r��V��A�
�Q��ɰ�~�J'E�X��B�F�Rb�$3Ӣ� >DQ@��#9�Z�"O�9�u�Y�:�0a�A�x���� /�vEq�ん�H��]� ���ffĐpM�iux�+�"O��G'����
���Lk���㆑�>�-�4�N~��=�g}rG�	�UJ􋇹tl� �[��y)�kf�E[��8z{ �/�3�M#q�ܘ(k�p C�'�BŅU�3���1Ə�{<L���w����t��)]��C�!�e9#�5-��)qN˻k�!�$ςCS���]�8�*I����}VqO���R��k�#� C>���2�I y0�M�W��l�<q2W3qP ;��͖\y�g�p4�?����O��1�˸GET}��M4mЊu�"O��`�6��}1� n�4X�w"O� �B"��t!8�[�nF�4[t5pB"Oؽ
�)ǘ�*M[�MPx�\Yw"O.����ʋU�V4��G��ddX��"ObH�MFO��!S#gʁ}��0S"OPeIc�	� v0Y#�`�>=}Ȍ"OB��2���H��4m�c����P"O8�3�P�z�Dj��^�ZPs�"O�H뇡8��k���HҜ\��"O���DfM�-A�Q;d-�^�JA�"O$3w�H2;��;Sf��^���ۅ"O�V��; �d��ʗa7*;�"O�Ak���Q����� $"��0"O6X@B'G��M�P
ɼT!�]P"O~e�h�i��]��J?P���"Or�B����
ږUJD��:)|h�"O*��,�2t&a�q�ψpB��W"O��c��P2/u���J�XxК"O���k¤&$tT8 CZ�3P:��7"O�%xc/Y�0X�;���kG^�I�"O�,a+P�H��Wa��a�r �s"O��C� ���80�Z�i�4,y�"O�Rt@�Acr�QԉH�F\sg"O����� <n��Ba	52��-��"O�$��m���
K�v�`��0"O��z�BWᐩ��o�	�Z�"O�)�F�0'�bX�w.�f����C"Ov\P�˛�<s<q�爵b�d9Q�"O��b�l�$��d��9o7���"Ot�딣[=!+F*B.�9y*� �"Ob��B��%$��j�,TuZ��"O�����x��)Ж�M�5Oe)w"O���[#M%b�)2���"�DH��"OT�a�ȏ.rJX�&D��p�J�ò"OH�ib�]!H������X !"O���AVR�$*�հ�	�b"O����˄G��a#��{�r�T"OB1��>���7��0}R"O��!���gŎ|i�A^#X�J!W"O�D�aKR�8"�T���8Z�6���'L��҅нD�z<"��I5��Q��� �bdd��S�șQvb!i!�Q��"O^�2��QjAI��n��C��р"O@���Y�H�qt��K�f�v"O�D�!��խ�iײY�v"O�QZV*B�_�ГSC�3?���0"O�H�2h�R���ǣ��-�)�"OXX�m�)FJ$$r!�]����"O,0u �=��G�*"&��1"O<Q�ɗ<��Bƅ\_&��"O��:C�"j�����B�����"Oh`��F�"3�Lbb�$Ԏ�p"O�yТ	>;�
t1Tj�@��p�""O&�c��C��h��@���V��!�$�8X�h�G/y����b<�a��T�00��㕔tmر°L�p/d,@�'4D�P�4K�s%Ic+�:4�|�62D��l��$x���*��+fV0��lJh�<��-�:���
7f��xq1M {�<�v�X��X��>w��ز&�v�<���4�8)9�,/'���׍^I�<��
��0�$)N�t{&&n�<7b��6e["���i?�hq�N�m�<)1��,�&��9���E�D�<i *�#2\-�WfE��u1eCQF�<� ��E��L�aIS�:�ar��|�<aT�W�f'����O*Yl��+�B^�<	�� ���ٱH˥6
4L�W�@F�<�唄>��H	�%ΣJ�����NC�<���֊y��)�G�� r�!4�X~�<�f�q�a#\@-90	NT�<S�\Y,h� ����N2�h�2��Q�<�'�ֺgK�d��+0&4�LyS��g�<�G�/t�8X9��K�
�D�f�<�%bG�8��͏ k�� �
Z�<��kAvQ�'-�t R1�	VK�<�W
P���K�B��[�K�<�wgԀzGt�S�MZ8ܰ#fb_D�<� @�I���)޿s�����E�<Y���XT��Ш�q��"ƙ!�D$M���z�A�:��UJwaX�F�!�$N.��0�Pށ��K2�!�Dǡ Chu� %� ;!l*���z!�DOl�!Pd�߷�|0"�B��!�$òS|i"b��  �N(�k��5,4��z���2�\ ��e�V,���1D�Pi��L�d[�;��QR<00e�<D���7gƏͪЫ��ϗW&��W%D��)�ݥpm&\9g�L4 6@��#D��UI�qXx�S�.���*t��($D��ȗ��/yTX�I��:\"�	!D���Q������g@�#XN��db D���1]�E�z�aLA�� 选;D���@ ��	�ԁ�`�1 ��7D�,sv�ЛX��iqd��c�ޜC5k4D��1�
�7d�)���Q�Q[%S)=D�(����%Q��Hf��*i��f�5D�� �Ζ�3��A5N�r���pb6D�<*7C?@�!��LhX�� 'D��C�HE��"�JO��XQ+0D�H##��5�8G���%������,D�(pwN]�s���0�H �;t�+D�| !\:�"6�>p�ܽ�7G%D���6R#��8GC�wĊ�aR"9D� ��(��TX���+V�e[p�8D�� P<2FDIc���m
�X�ƈ �"O�@���;�NP��+�)h��"O$�pW�@�!"��wiS=d
H:r"O$���� _Ƃ ��#]E��6"O�4�pg��(��C���):�.�yb�^�t�E]6�%�f��y�L��9�D۠B�9=�TXрM�;�y�
�1[���`"��>1���@�yBn�y[��P狇�}l����ձ�y�
2Q��DHB��J�~�2���y�j+?b��P@	¥6D<Q*����y�)�<�����e��+��Ys�_��y��J�R!�Q	0��*=��Z��y�e�%g*Qb���+�4|�@�y��ڵ=-J��ӫ�B��>EȊ���'��1kr-ҹXW�UH�l�96��`�'�N���~�Xjs��3'�Ԁ�
�'�����B �B���G�V���a
�'u��&�
za �K�.7��e	�'�ڱ�g쁡�"�r���aB��
�'�%��h� p���n
�W��'l�,;��9��bu Z�Y�"hP�'_�y�!�UL��{DiɊ=�F�{�'�M;4�c,T��C�ʋ!��#�',��'P2P��G�޹Q^��'����C��n(�[�x%��2�'->x��K�!����ܝ8���'l������;��ܱ`$e\�H��'������<?�"��@e /1Ld@�'�8 fR�r�j�2@�P��|A�'��X��Ԕ��a�Ʉ�)�T*�' r-h�]x������S��`��'Y�4×	�U}訸�%�.?���	�'�MWNʎ<�f�(�`V>P%��'K�dC��ΜX3�B /�%�'(ҤPgl9Fe>9Ї"ְj��'�^eZħ�ah��ڗ6��3�'�J<)���%r��V�C�<ܢ
�'�4uk���l���/�	:��A
�'�y1vNR
;��	�98�Hi9�'^�i��n�X`�G�0V�|1�'�B��"�Y���xhp���@�a"�'����K�+L��DQ*g�0��'�C4��7 Bе��kZi3ji�'᬴�FB,b;^�h�+��`2�'n0���k�T�&��	/D�"�'�������Rn�����+�0�3
�'����� ^<534���@X+	��,��'R m�7���C����m�R�ڴK	�'��C�+�(���C"Dk����'X��k��� BZXqp4�C�T���'|F��
�m�h���<��	�'k�����!^��Ȉ�d��:B�I'=?Ҝi���(M�$(�%�?t 2B��T��4FV f��e��N�K��D{��9OT)
�m��IU�<�f���=� �9"O�P���D�=��ؠ�Lu�����"OT��`b��CJn0��ˈ<���"OT@y�V+}�C�e��I$�"Oa{AH؝^���Vʆ�I:R� �"O�q"����f���wH��4�p�bD"OHcS+�2G,U����0^w<e0"Of�[H�� �z(z3[12k �R7"O��I���R�8Ȓ�`-�Jx�A"O� *k�ѳd�n���v�f�*�"O���c�ETk�耆�ݘK2�e1�"O�Q2�I�#?ҙ���T)S'�Mc�"O��P��[�zP�=��KN�P<��"O����Àm�ր�fAJ7`S>�Y�"O虱�g��Suv0�%q�6ء"Oj���x�^��D��d���a�"O�(8� c9 �k��A*�'"O�0��KM�y�n9kT�+��k�"Oa��οg�� �p�A� <��"O�-x�j�9-	E�ue��)(�P"O���W}z0z"�TV�� k�"O���@g�(T�DHa��Q�2��aPw"O�9�gCX;)����QŪU�"O��r� �n�p��R��'�"�ۄ"O\�H%�c�&%��j��<��4�Q"O,ɣ��R�X,H1V��8�2��"OT��1�^���9&��$=�0��D"OL5SbΖ���`Ò�P�?�Z��""Ov8�������(�`��W�X��b"O,����M�и���ϱ{�>�{"O��q�*Y��|���תu�~]��"On���%D��\Ҧ rgPX�"O�I2m��K$0�B�Оrhrɉ1"O�yS��ށh�I�.�=[f%"O�=��'K-\��R�صA'�T� "O�h���/*��@P���J.�K�"O�S�RA7�`��+h��g"O"��"�P.w��eQ���3Z�8`"O�����'t�Yb2M9Z�ݱ1"Ox̩��!K��M(U
_!h�����"O��c�h�`��IB5	�t�F��"OPd�`)ʒO��Թ5H5�f���"OZ�%O;:ي�#�J% �4��""O��+�̜�l����heP�"OPT�&�?!��1�ή����"O�8��.��;F�� ����"O�M�!9�L����,�u"O���reF�HR� ��σa���%"O�l;�����
iE��yS֌�"Obͫ��؋/��,���Z�rPp���"Ol�XSA�a-�!��"a7��b�"O}�Vh�>y��w��"����"O�y�0 ݓh�FM�Ék����"O�`C�5@�J
��߁!��["O��S	�
+���Z������b"O�A�5�H�$��=�tC�6�Ƒs�"O�-KbBۧS�` ��k�<(�p"O���>O�T�"F�H��5��"O���fƅ!/\�E"���G�`�!�"OL�S6��&<���� S�]pv"O�8�vKھr܄��@
.�|ٰ"Ol�����$B���\�ܼ�	�"O���O�=��A�@R,%�pt"O��xAW춴��O��48H��"O��*���9~h́�M)&��Q @"O$yCg
C�1�Jy�LKt���"O�tj�e�%@6ܡ@��(o���g"Oz��$瓶_6!p��2bX|�"O�����J	o�a�C��<�H� "O�QKg�'BlD����`/��0"Oؽ�$��q�t��3���9���@�"OFd��#G$jJ����+q��§"O������I9W*\�ff8 "O� ڐ:*��|ɲ��`��C�"O�Q�+W)i���O��Q~%�"O�H
e��/{�ћ�-^/�h�*�"O�pQb�'J=x���(�	"O��A���"5��seN���D�6"O����*O$
ܹ9��΋\��(��"Op���@�9|5���B�UN�0f"O`�cr�O>Q�j�B5�Yt0T%H�"O�|˰&�R���2%���'�Y"OR�Z:J��pE�F�G��Х"O�T�aە������V�H����r"O�M��W'<�)g�<� �sp"O�eP�ʅ�E���Q7�J�Ibf"Oz��ˍ>�J�i�������y�"Of�q�W��hQIDK�"x
q�p"O.�;�A8e�lz���#fH*�"O��g� 
NSp,��CפUဳ"Oz1$�۽X)�u��C��lX���"O��ȓ�  �P   k
  .  �  E!  H(  �0  7  X=  �C  �I  wQ  X  W^  �d  �j  %q  iw  �}  E�   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl�
�;�>O�1"�'"d�D�B��3�91���b���IWov���W��;���nd�%R���?ڑ���?M�A��iκ�)���XP ����bu��;uɐ�_�V8�Fl)#�(�:w�[��u��S�����'�t(�!�J��d���Ae���i�EW%
��TfB�O�٪a�$i���Y��զ2�J����ß0����r���=ͬ0����ِ���۟p�I��}�4���O�@р���d�O8��jEQ������1�´0��O���O��d�O��SV��OH@C!�'�����4���%��u��)�$���5�O\�	_]�g�̿d�m�2�G	K���y��|b�ON�ٴ�����)�9|Y�4�����%
�������'-��'[��'p��'�������Q��tC���*UX�1��ڟ0�ݴ6���w��X�'-h7� .�@�nZk ���� �z��X�vrre(dcÏ2�F�h����r�9Џ�	¸
s4�����%N�l�{p,�{�ȩ���]H8�x�d�;��7M���c�4���3V�ؓ���%H��9'�DPj@�JO"R�(|җ�i�������� �I��ۇO�hss�E�.p�(�$p�hyo�>�M[���

f�"�)� N��M��
�����*D�&f��io|6����ёC�Ԛ}��jSn�5qE��k�oe�8���0v4�i �ʃ%}��!O�C �ac�C���6����)��4@��q�[�$(�DD�J6mU:V��Ð-��*2
	�ϴ~��H�⊇$"C����:72�děQ��3��G�	l"�`�� 9���>�Iԟ\���B��Xj�4��Iǒ�H��ڳ	  �p�F$�Q�d��͟�'9P��8Ⱦ\�#����Mc`�_������1�.Qx�����0<	$����`�E�&���� G�����4,��t�Gn�܆�	9&��$�O,�'^2T 穇" bX�X�mڡf891��?�������ON�IRx0�# O�,!��z=�"�j�p0�"�**��d���&<�xH��Ҧ�?R�T���'��T�V�>��7#�(+F��(ccD=�!�ªb9�BB)M#o�@�sa8�!�DO�5T:d�W�B�ȹ"�m�R*!�  �b��󃍬pl���˿D(!���z�H�JG�5(^De���צa�!�䄈*��o�^W��`k�:�R���O?����@-����>38��afOp�<1�nG>ck̔{�C��l��= o\C�<��kJ�N",���Y�A���� �~�<�1��9o�$$a��]�B���9Vōc�<ib�"`�2��*�
������v�<A�CҖU�P�*�\����9���kybEץ�p>�"D
;v�t�
ĥg�y�O�h�<9cB��\���3&�:RbR	95�e�<R�S77q;��E�i��I3�
Za�<���3Q��e.�Lq�e1�@E�<��ޕY�Vmj�j>���P�%Tfx��RCI�M����?3�Y(u�4aХ�
a>0��E��?��.�Dl���?���u���a�M��Ɗ�h��T�S��y��.*U�塣ǚ�|�axR+�dN�)*#	B�	�B���� 0Ku,��ąدQ4󲮈� <8��/�~�	�Cش�?�i#]��zC�=���� e؞���O�⟢|:G��3@�W�\��\��ǟ�Y�b�X�'�>���4	�z1*��10AR1 ���u��ч�i��'�`Q8C���9&�O���%V
�Bc�Ͱh씣P3�C�Iu[41��a�'|�|��h��C�	�Z�+��V#9<������C�@}��o� �%�Ǧ�?�0C�I�(�MZ�:�Z,���ǵ&�C��8-N�;&���T8QuǕ�^��oZH�U\��͟p��ҟ\�''X�.�?�:u�D�G3&LHw$	6�66�����P�ݑ=v6��O�:�8�i�7}��P�-��O:^�xf
��J��3�U�5�B|;d�G��b>�kwH�w����<uJ�ų&4���c+Ⱥdpj6-�y"-\��?�����?���4t��a���V��A�z�a
ϓx��O��B`d3D��U����'3r��4R�DI�4CJ��|�Oh��T���I͘n0 �:v�A7԰�A	Q�66Bl�������������u��'��8�|T�B�B�wP5yC�#�:a[CGƀ��x��Y����N?<OT�uA]�	��"s,��f���qP@M�U��]%��#e.'<OY��n�8rRt�����p��@��U��'WB�D(�'B&҄��̄�^��Q3�dȿ2�t���
3���R;�v])tnE2> Y'����4�?	,ON�W+�ަ}�O8f]�k�x/�hk噦nƌ������O��d�Oz�{�R�#���9����W�H�)� X �3���<�u�T�2��@�'�����K�Hب1UOK��y��j��D�c��6+j��1u#!�0<	'&
ǟ�[۴�?��hH�:�dRQڦ�N��B��U���?����?9����'��'�)�%�;�$�F`�<�p��O_��B`|y{��H�k�&��c�(�?q-O6�˶*��q��ß�O�.� ��'6Vٳw�ל�r�
ąT<����g�'R�_�v8��T>�'��Y�����Y�k��X��@�Ox���)§dT�5�a�36�lY��˳U+�4�'k�����ɧ����#x{�pԒÊ y�*@�"O܌1��Լo�����IÜ�����	�h�2E�v'�Lj��D	N=�`�s���D�O��d8���c��O����OF��x�yz�eTI,�8@c���� �'����@�A��0�nAc>A��T�&/� =�~�����vHЙ�d�Gv��P3CoZ�������	@�t�U�	W�p��\`�'�q��*��L��T M�R����in^�k��	�?����'t�2@dMC��BQpH|��'�>|@6��uWڽH�kA�<�+O*�Fz�OH]��v�A�W���)뇆|z�}@$��/v���p�ܟ��Iڟ��	"�u��'(�0�V�A����e+b��TF�"yfH��i�g�!�D@�SO*�0+�	1c6���o^�5i���O$�0p��3BbD������͘��ڪw���'�O� �K�+M�n��l�3)i��A�"O^1;PA��SD���9Md�Qe�|2�e�ʒO`�7k�K�T�'"h���˔\��a�f�K�}qh�3��'8�H�o���'	�i�e�R4�GlG�Y�=zuf�O�%��\�"���S�I�/&l^L8r�'���Ȗ���{L<H�䏋L��B���f��4A�:u0���)�0<���`��Q~�2�R@`�At��H�F�����?���:�Cg!D�(	�!�,���I��?9k�7��{V풵Π��BE�l�'�����`�>������l*B�$�4xmj1
ڮ�6������O����˕�]�0) r�M�:]d�kq!����_>q�Ϟ?v�L8Ѷb����`�KGW~���^o2��㡙u:���'���a%'W?J�}qQ�Oh%BH�_��Mr3�H��
8��O�����'�7Mܦ���l�Ol�p� �@)k����읳l[�`�K>Y��?������O��?7�1�(�-%���6	G���dD2�c�.m`��9=D�2�N<x4��3��eh8��4�?����?�qb�?L�����?���?1�;H;�)aׯ[2��P4��,�Ȣ�Ð�D�b�r���q������E�RO+���L)�D'�<m�Q�S�� 4�Hq��Z(vtT-Җꐖ3x�BE�<���z;(��a��8��:e ҹTOYDP*��Ϧ���4�?�cV��?я�,O��$ԛ$�JQ+�[�p	9�J�<>����O4ʓ�?���L�z��N��d�3�"�ҽ ���<�$�i7�=��|�,O6p�ֈ�B��)չ�N��g�����&�O>�D�O����׺����?��OG���Dc��J;2����S����K�gϗ`2�A��%�c�數���*������'�)�$LΦ~媰*��Ԓ��� �3`��T�4��:X䐭�C��{{��Պ�n�'�>욥F�/�6X��/�� �����L�?9��it�#=9��D�4Y#R�#�*�+v�,�3��,}�!�����e�e-
$hҞ�9��'-`7-�O�=Z�4+[?��ɤ����+��3_HE)�אvސ��	��h �ПL�I�|�5��1��F��@��}2�L��i�TY:�	�(���g��	$@!��h�8W�|�<�I��#e�l)��ȁ?H i�����ۣ�_���D�'��>0n��"M�&	E �<�`�$��43�I-���6膀m�R4�"��69Ŕ�Ot��$zy8��'YP`�Ц������O�I��/[-hw�Ѹ���ԥP��'��O�Uhg�ϼ�DU����iG%7�>Q[F�@�<�Wh�*qZ�)`��Y�-2l�D~�<aD��E}�@s���n�"$^�<�WK�&�]kת� &�\��b�V�<)cD��O*��� gN�MG���R��H�<1�[������n묬��ȎП�K1�S�O�|ش�]�O��Ex7n�^=\=�@"O0]2�)�(^$F��`��:�`:G"O@�S늉�����+I�h���"O�\z�*N�;ZĂ������[�"O����n�RM�g	��{�x�!q"O6����}�ƭ�u.^���1�[���@�)�O�8�n��VC�8PP��	��R"O� �0��3+/D§ϔ�s�:�"A"O��큼92�Q�nL@�M��"O�-ѳ�C�L���+� q�"O�)hL�:��ܙ�c�/�Nu��'����'¼i��T��p�Y�m-��
�'��tȭ?"�m�`�G�R��S�'NB�Q�A�$?n��Wm��kB5��'Q����@�W��h`��7�`�'榽�cŎ�)#ؘ�v��1� ��'80�)�I��ce����
L�!��@���±s�Q?(&�֕R�<��&V�2t*!�'D�б�@�# q|h��NT�;Q"����%D�,����c� yP��V�3�7D�0"���d@nx��$M-%�F�A�3D��6,���a�wFL�H�V��@B6D�Ĩ��đ-��qw��D������O��"�)�'2��;�Ȏ�l��ab�B�T���'s�<�� ��0�����>O*��'�\aXե�8k�ʁ�"��!�h��'��#��I�b��lX!-��|��'��ՃW�jB�[#AW)&.�I��'�0M�͞>EԮM��d=!���-O�@��'ea�
J@,)s��K&HT�pB�'�� zc�ǭ](�A(B@\�KJi��'7��2�L&bL1�a�pH�,��'[�$�@�\4M�\ٓ1���n��Q2�'Qg@EO�Ā A�B�7�0�H���%b(X�l?)���F�Ę�~	�ȓ���#獂�(B�(0�*�>W�p�ȓc�Eأ���;b0ś7�7��`�ȓ3x,<�B,	d�f"0�+_*х�]m��ْ�)�����mZ��ȓ9<@`3���W�b5s���E�
�E{��Ѱ﨟��Q��}���*ԬE�k�T��"O��p�f_�`������׏M�%�"O�3F���t������
�
Pw"O����h���M ��Y`t�)pV"O�#g�SA��:⦍�rc����"OV�sb�#eD%�RdP,;:�
��'������Ӊ F�T�L�`�� d)��thć�=�@E(�̖	<��-�)�J��ȓ)�Da
���b!Z$	rF�NW���.R�`�P����ɠ�C^3XU��M����tk�o@����N�tFɇ�EQ�����
�'�Z�����4�X$�'7`���%���*1�ױf�<8�����@�!�D�����d�>-��Q���&�!�$۫w���A��#�p)���+?�!�;�N�� &�c>�C���)�!�D�ZjZ$P�fW{ �q*Я�*��}"@� �~¦�M:ب*2��x��AP�Ŝ��y�&�'�pM��xӤ$���@�y�刵!�d�@�F��^��8�a�K��y�eJ�G�b���W<�i	a�ϓ�yR�@5�����Q��	�����y�ꞁ"��8�&A��奚��hOtEA��өS���q�U�|Ţ�c�cJ�C�;���b�@8������)�C�I6�jH�U��)3iT�� ۶q�dC�ɇS1&ap�
�euN�1��]�,C�	�	��0RC䟨 64��M'
C�	/}n��k��
Hb| t�J�0���)��"~B��]-r�xH��e��(���!��0�y�d�.���
�s]T�3a�A+�y
� ���chOUh�C���!I *e�"O2U+�!��'�P$���$m�(�"Oư�v%L%�z-�%�A4�}�Q"O��r���l/��SW�@_�uP�Y�@�D�"�O�<�Ab��I�$��J
�lT�	R�"Oș�
�Cv%��ߺ1��XU"O*�+�C\'�()%i�'%�;D"O����Z!jx�5.E���J`�:�y��eX��0枝2ޔ=B 
��>����g?AW+*n{� o�utpAY��x�<����J1섑|��%9��u�<i"bg�t�v]��s���y�<��	PG����cF�MH�}su�<ygD'�> uM�NV���S[l�<�!B�<�z�"�+v�k�Cd�'n�u+��Ɏ�-�	��Cبi�� �˜i!��	E��e�C����iк[!�ε3>��a�M_�M̌<*�GٻP!��~��0��ӃG��#VNM!��MN�1�G�/s�����f�8q>!�d#�>��uat,��B�Z:23��4�O?]�O҄30~��͖4���c �K�<��I�q4�8���7@٪�AK�<����lh�s�,J����d�I�<��U�D5�!��4*"���/CG�<�(*/|�KT�Xdm8Ј�F�<�d^�1Ө�b�.Ԅ;30��dh\FyRdJ�p>�%D�����ҍ��H�n�!��L�<q@"P�3ݎAzSɅ=!O d)�l�r�<�6�V�����S:P��M	�m	p�<a��̤���
�DT�f	K?I6�C�I/cBzI�k l��13�ج:~���DE���>�Zx:aE҄[;626�!R!� ��@��)d$���J��`�!�B>L�M��:��8�(�_G!��ٚR_������!L�(YQ���L�!�Dނ��I��w=�������!�d��?�YYD��0Q%��$��<p�ў0a0�'� �!#�B:E���1P��ȓR*��Pz�W� /|����o&�L���)t���;b���Z<��!rkҒn�k�	���Ѕ�e���YRG�N���׏��ߢ8��^����OLTV&����Ӆ'ǀ��ɶt:#<E�D��&X��,"7�Ã8��Ia`#N�\�!��'#"���$�'6=��9"�ܣd�!���pK��{��9���q����-�!�D1KTX d�~@���k!��6���{&�ϱg���o��r�!��ۏv� ̈b@R�P`���Ȇo��I�6^���C#o�*��1JF$M��a�'R?hQ!��V�(�ƀCˀ�a8������bP!��F�2�
"��;bm؄��n!�$ц���1 #���A�FVb!��O��T#���7�� �E\:^�}2����~¥O�C��wI�8n�
l:�J��y��HCȥ�'`ǯ_�d�������y�G֋<���QL��^l|�ȧ ���yZrvq)5bx��\�f�$E@A�ȓ3LI��f
G0���D�"t�P���\ޑ�0��/�D2�Mܴd�)F{R��>����II���Ha�"h*�F���"O�Y��-�EbXD�@�M2
��,�d"OP���.}��	�嚌m;��"O� <��sl�G%��Zq#�x�����"O�Qh�Nq��=�s'G�{h��"O��0�u��yPp���m^ Q��'Lp,����Ӭ�b(�p`ӥh.uyWLޖ	�M�ȓ=��pC&��4�r)��d��I�E���	U�V�<���6����d�R<&�������D�ȓ?0�i��ж-���4F�_���xN�!�Ԡ� U�ԡ��B�<x�葖'��P��S2�@�!����m���B76~����)��u�AD�3(@R����p�j̆ȓYI��W R@z�z��	*@�TT���R��O(N�y���;n�2�3wh1D�P2�
C�j����1qU"���b0�O�\cU�O�r+aՉ�FF�F^ddA3"�A�<��#ɵ8�P5�J�/d��D1��D�<	��L,!���aA�(_{�p�ERj�<�V����#'h��s��Ճ#��d�<4c��Q��Q�r��2u
(��.Jk�<� �3&ẕ��!�M+
,"�(�^�'��=���� �+h(3!64��\2GQ��!�dE#QV�@v��Gj�]&�9�!�
N���
���we���F�X'U�!�DM�_�5)N]�RWڈ�T%ޔ�!�C�Ft.!+T̉?'���B�ў+!򤉞~�����m������1e��F'�O?��(��:W&i�h�YK]U�<�Q�� �6)��ݘ.�1�z�<i��F k�� [wHٔoT�`�Ǆ�t�<��CV/F�fi��aM��U��`q�<y"���2�@�N'!km3�ph<a��۬\�Rx�1�H�B!��&�A��?)J�,�)O`�l��M��1�?q��#��<bv%5a��XL�S���
�2=������?9��X�F�k E �
�q���J�^;vO�;!Z�:���n���	t"�g&�Q��D�q�'Z�rdnΓY�긠���NC� ׂũI��QX����m13aܪb!��el�^�'� �Q�1��#"�I,�0�k$��[��)��@��Ix���G�Qd��b�k,y%�)�5#�O|ԕ'T���u��= W�^���"d  3�Oz��O2��ƒ	qw��Ӄ톷O��u"O��!���mpӋ�P�^E86"O�ib�_	m��J�ʁ�6��LX!"O�|�oŠK`��&��r��U��"O�H�u�Z��$�,1q<41'"O�,b%%�z:�@���4rjB4��K��O��}��W|,Ā�
Ř��)�1�_j�V �ȓڐ s��L��Hi�V�^=V��ȓ"Ȓ�#�
�Jp(�4��"a�ń�P[�iA��+-��̳EL	 hؼ]��'~��e��#�$PYY���}�<�G�`}0Af&�,<��yeɓ���!�<�OT�pfיA�r�JO9�P�P"O:�`C�Q�f��x��b%�|p4"O|@pv@�\��q��m/���3"O�t�AD�6fX�������"O ��pBÏFvB(rF���l��\���'벴2I�0����mB��V�K�%D��:B�S7/�|�c� �+H$�
 �/D���A$Z^C��2��N���� ,D���5�Ɏ��1J�j���;�l+D�0r����"�D������-D���B[�Y:�)g��X��p1�ɦ}��"<���-�%��B��q����D��@"O^(	R舓Ӝ=!��_ ,%��"OTf@��m�i��/q�	�b"O� J��AE�d`��N�vY^) �"OhmX��K5S>pP`��T]��U�U"Ot}��	�T*
�����-�6B���O��}��e_0Qz�f�5�x0C�[��Y�ȓ6�ʑHq��xS�a���Ԕ9
\C����D'62xA$�n�D��&j/D�L���"%��H���3W �*D�`;�
�:lj�I���@��u(4D'D���t��;)t��0��''ʎpi !�OAh��'&�D��H�3�Kgbי"iv	�	�'��h�A&��i$���������i�	�'�z�.% ����](!��afCN�<!rg�%�,<8��Ϣ!ET9Q	K�<����z��(�ڔ��t��h�F�'�@H����>�������-����%��
|]�"���?��O�?A��?��d���`1F��N1�)�R��0|�U�ƅ,NA�Y��U/nh||�d��1�pGyR��z.:��ѾT��36��
`^�B'�M�l0a�#�1M�ɣ ��/�F�Ey����?��ib���2�;1%؆'MZa�kKҐ��d �O@�Cm)8�ZU3��E�@�
b�'�˓1:��؂(�I@r�ǀ,��u�'mB�'��t�'��|���Ib�M�T;��yG���-9ʢ?	��S�>��ݫ�m���4q���&��⟈C��*����?1ϟ���@�d@Q��F�w�Lr����'� H�O���<�%���V�ìT�{vx��P��eT��0�O谤O\�Z%�>�����j��N��:p�� �>� ���Z��5�O�9���h��D"wZ\���ηvEZ�Tp^d%)��>�$�>y!X���w���_�P8����G�&�J����?��E|�$��v��?�P�L/j�y�4ń���0�����&}��1}�)Ҕ���0�M+������;ՆP�3�Y�q��sy������#�ȟ�$�D�
c|�����+���)7�i?����p�T>�	�u�^�"� D��<P��
Q���:�A���f(6���O.18���δ1� ��D˪'�.Y�� ��2��x?A����?�M~��t�3y��	�+"���RL�= `)�Iw�aRbZ� ��)v���&���;�y��Y(���
��Py<Qj��צ�M{���?�+O<���Of���ƺ�S��4P׈�$U24���iRP����&����O�˧�?�ڣf�h���w���1��?�؍%�L�	_��|�K�����(d7f���ϰM�$Ӈ!)D�����H�Z�����M��/��l�t�<i#������k�g�Y�i�\�<�*�=�����N=E�<��s�J`�<aP� ����q��G'��1��X�<�b����J�v�*��!�^`�<��W�D���w,ܯ&z�!��_�<)��)+B*��2�^F���0��q�<���G[� �M^�R��a��i�<i��+�d	�"D�<0��M�R!�e�',�"=�O�M7�@�^~.	�EF0v���'��� a�H�"�*}`AO�*t�x8��}r-�J��+��;&Ő@��������[ae��<.r@c�l���#�
����4@v�?Lؠaf,^:,�8,[�.ARS!�X�
ubΩ#�:ԁ��%$$X@�A7PO��Y᪚>�� s͘R�8$�5�M���	 ���n!��-ͯD+,|�c���T���	�M���9�U�!�U���	AS�Y��	��ݟ�A7O "Ķ�N>�O��	X��P�"R�E��5����O��r�!z�	݁�����>$�F�'�!�GÃDeTt8��Q�^�D�(�a�o�	#:�h���̦���4�?��aS�_�F��dV�\�jH�`@O��':B�'ՖriՋw`�d(��T�Y�]9�*�Q��Cr��"�D�P�O]>�.��e�K�(�9)���>q��W%�0� �6]�q;5f�V�<IҭW$	ε3*KX�!�,�y�<�U�K�q  ��Z�N&Q�cn�J�<�AAQ�;�p�׫�*��qB��AE�<1��J+7z�� �%4��ꠦ�U�<9�$����:Ê �W�� 95��U�<��LI,N���FּC���P`@_P�<� L��)V� p���" ��C"OV�`�J�9�a�6�>,txy�A"O�$�Gh�:/��`��G�FTX�v"O�-!tdD3�p$�4!��LF�{�"O��J��$���n���3"O>=�����D=��J�̌�I�tEkB"O���s)�qA{A�0 �*"Ov!�(�4}Li`P�ʒ_�d�["O�I9��6R?��i�-lI���b"O��4�?���3�JlB%��"O4���="$���!ՏU&i�@"O����F�5�|lb�`�h�Nd �"O���GH��� 3$��(�n��"O�l��7�#���n���"O^�"��ْ�Ҹ)�K��.�|���"O@�������Jِ+�jju"O�X�k8u�����C�8['��#!"ON�`RAV� $<!�^>4�8X�"O~<taƯq@) ᑒ%�E��"O�Y�b�K�_(� 2U�*i+�"O�D���^{Ү��R�D`2"O"Ai�G%t����
D>�!�P"O�͊tdO�xQ���S#� �"O�}@�V���r�f�7U�1"Oź�%c�"�1�c��	��T"OF�Z�DJ�j���:D�.`6i��"ODUb�սC�h�H�#��N:�A�0"O�,0���p�n5��ȹ
}��"O��%Eۣ��t��"͊mHE1"O�A�g־p<ȅ�Gk�b��g"OΩ	 d['/,�(�E�R���-��"OH ʲ�Ol���R��<���Pq"O\eC�
6Bς�3����2�򘈐"O�!aC�d$�!�@�>m�|"�"O�܊��Qh���m�T�l��"OT!��@3_P<PP�T�X:���E"OR�x�@�Z���m~&p�9D�����o��!��ֵ+���Xs&7D�Ȳ2�7k϶��'V�0����qb7D��y��ٳ?��KGaY�w+ �sJ7D� �E�*((m
��Y��AI@�6D��b��T�A�@�p1'�h;���, D����q����A���u���!D�0���A1�4��ӑ2����J>D����+ƥiR!�Q(�~M�%>D�H� "�?:C"!����d8�#n0D�(ȡ�(9��"p�&4�f��C,D���m�����1M��5>�0�F.D���`IE�2�Z<r���J[<(#�*D���ȟ�&ǂ���`{��B�=D��[`�%hd�0E+�*$�3��>D����c^<������Y3g�ִ*�.D�,`d��u��u����:eE\�*�!D�p�`M�V�|�*�œ��Y�En;D��A�)��dl0�L�
���r�5D�(Z��O�T���%�
�gǸ�.&D��y��X�fq[��ʸnĠ�:��%D�����O�
蒼��Ɓ"%�\s�&T��¦GW 88�� ��ޛf�HU "O@����X0b8LU�D��Q�ιH'"O��QS�B�e�*�K�D��o��%bP"O�`�g�:eܨ��;0[����"O�x��bO��c�/U��`""Ora+�^/d�NL��h�2fQL���"O� \XVJZ�J�~�;�B�")6�q�"O6X;�..0��\6�c"OD�@`�	�[�����a�1m�l��"Ox��c�(*Bdq�n����V"O<1a��>15��b�޳��1��"O�PS���X٨�̓�[� ��p�<��)�X��o[����]n�<1qH٪o�F ��l�u?
a�CF�n�<A9R��"��Ŋ$`�\�Pɇb�<�1��	�.����Ӑ.�F�1��]�<1���I=(�X2A�V �D� �Z�<��N�AVbe�eJL�8�`h�C��R�<)��/f���DI^p���gPV�<���X�l�" G�'+�P��Lz�<IEa8+ZI/%�haT�*xhB�,��0e��;cH�{�,B�	"�=�͚���12�C��+�R(e�.}�~%`�h�b�~C�	!�:eQω���x35�޽q�^C䉿!H�0xt�7��4����&.��C�ɣ7:��*օ�-o��#Q��VPC�I|B�3EB^B�S���VC�	�t@�p���E�� �.��hB�B�	)\AxȲK� @�̛ĥ�B��/���*���D� (�ž��B�ɔV�@P�fY�h�^` ��^8$JjB�I:yT$8A.\��o����/�d5��Q����� ހz�H<�ȓQR�J�j�G�l�D	�J�ȓJS���
� V����[�[Җ��ȓ�����PB�p+\�#�&��ȓ[SH)���V�N�ٻ��C�0�6D�ȓ �|ekբ�%g`b��E �:[o�y�ȓ6��ؠ.�4���"�
ceф�7�fX�'N1ւh��ˀ�*�N �ȓT��Xqw�<R���̗�?��L��h�Ȱ�t�5%�
X��	�xh-���I`e��(0�! �D�	��]�ȓhQ��A"G�<,��MY��Hu�ȓviڈ�wS�GΚ��G�D6(贅�eQ|��c��*"�4I�Y0u������	+9Z(��W�y�4�ȓ(�,@b���)�-��!�.̈́ȓd���Ф��'N|���-�|�T��ȓ�(����.ot�;2�7���ȓ	����"�F�ӢVM���m��x"���|�e��"!���|N�i@aD -�!��n���'Y��I�F�o�~�HRB�p���c�']�
@��_'f�sk�cj�"�'��x���m��L�r&��d<�\��'���QB�M��|(�J*�P�	�'��Tf�;p��`��� M��'��� )N�A�����mK��L��'��!����`-�4X�lʖi����'�0�k��� ��(�$�	�'����)�4x�d��lG�O0��'B����1<P��I}t����'�4z�̍`W%��C��G�`�2�'�4�H%�9��=�b�H@,v$Y�'�x�7�N	6yF��KF�?�. y�'L�8Eo� 8��}�F4�Ty��'�v�ђFO`�L��h�+/�QQ�'�D�BG�1�l�'�	*tFD��� ����
�O��AY����FN�)��"O��֥Q�)��\�,�S�p��"O$=pg�	��i�e�2ǂ�i7�#D��#Ŝ����i�$� ͊�� D���1kM�,E�Lhf��-?<*�x4(!D���ぁ�A������C�%�U�,D�07�C��`�ri�H�B-��+D��;��mb,Ds��}�)p�%D�$+"@��8��ڶ./���h��C�	=W`г�h�R�	���͝� C�	Q�X�S�MD�����6J�#%��B�I�Zb���-_��d#�#Wa{rB�:p�`��v�;��@X@K�-�XB�|�y��@�=Нr� '�B�	�LE��Y��'R�§M�jҰC��kǆ�1���%/7��I&)ܻz�lC�ɮv��{�C�|�`u1`��&�tC�I ڠ��(�bG8���X%$BC�I�r9�IؕO�-b�
 AX4_`C�I���hɁN�0�L���l��
��C�ɬ-;0@��fO�F��X���B.��B�I�h-�l����({��� ��7,٨B䉣'��cs(�Z�:D{��]!H���EN����τ�y41��3!�$�'Xp=�7*X�V�G, 9!�$�2g��b@�|u�6T+!��4KѼ�G���6t�	���K)�!��W#r���< U6����!�dG�	>�}�BԻJ:��A��$(!��ä �¥��̲{&bp��} !��@�B��܊u�Vo�.W�.��X�ȓY�č	PH�2�胑	+��-�ȓڔH�D�p�����ʬ6�N���I��d+���;�� +H��ȓ.R���B�LO�#��GWFb5�ȓ4���G�ޑ+��c�ٰTk|0�ȓn�`����<Q�t�kuF�[A���ȓ1F�hՇJ�Gz�S�m�:݄ȓ@�93��
_e�)�,�#g)t�ȓD�rI�G��Jl�}Ђ݈@B����4��q�-�<5���ɍ!t��ȓ)�PT�G�B�[�6�ȆBëeK�m�ȓ&/FUrc��CWXMH��Ok��ȓy[�� ��<Nh��#ΎP@=�ȓwX:����és�H�s�C\q ���Y젙PR�\�	A$���p��,�ȓ}y\���H\$-��`�=q⩄ȓ��1�nŶv.8�� PJ�͇ȓ�N�|	3���G_F%�ȓ#L�Ak�nо)�N��q��7rf���ȓg��i�7�/\�(��3�*�E��aԩ�� %b���Bۋz�\�ȓ4��ɣ�g�I^�yҀ��C�����X��0j^$ 8ڌ�B��D����PJ�L�9>���
�~�ȅ�n��� ��,}��b�Ԁ)S�}��`�9�F^n�a9���!���ȓ3�x`y���
�� �	�=Qz��ȓ�L�!�_�U�h��C/� ��ȓnwP8��	ۮ�ro^L0 )�ȓ3��x�U�˪I�=#��	�,?l$�ȓ�r9s`:fղ�:��"�h��/����F��*����eJ#]�� -� (�(� �<1&4�
ϓ|/��p�'B�T���A�:B.Ň�S�? ����	+�miR�)h](\x�"O\�bA�"�h@��:Z��"OH��&Ǐz�(�q�A�Dv���"Oz�x��:����)2[4��$"Ov�*�k͌�C2�KO��K7"OXHp�T�	l4IHP��z�� ��"Oe0����c�^mj�(W'���4"O0�s�ё g\��#�8d�<��"O"�j��ߍm:���B̊�`6e��"OՊĀ^�9
|�x5��0X�U�s"On�4��-p#��rC�nSVm@"O��1���53�q�D��x�`!"O�9ڐ�ܤv �@"�ۆd�Y
"O6���%W�T�#a꘷Kd(�R"OnM�F	
�.Ŷ|Q��qo�D"O���׋D�f�H������
8"O�=P`G�,j&��9D��|��"OZ���)Qe��i�N��bĴ�A"O ��R��H��Y GF�wR���"O
4+���<wb}��C�"$ M�"O�Ҵf�1���Ã(I�F�i�"OT��A\� 
�@�"�+�P��"O�pC����|����`�&�	q"Od`�kA�W�!7M"P�5�"OV�s6���:�S�C�U��0k�"Oh��҆��n]�ӤH*WI�#"OH��ՇJ xd��DM�J�h�y�<�+�T֕�v�B��1RcE�t�<�"ʋ+@Vm� ��r3�N�<	��RU��!hq'B��|�D��<��N�)~4c��U:W=��yeυ|�<���XӐY��G�1%���`�Ct�<	�fF��}`,Ԭa�j���ls�<����4�$��7׳r��1A��CM�<1�����<YcTs]V���MT�<��"���feL40�<�aƯE�<�ȓ�r���Pp��WC����D�<�#.�:H��+�!O/B�$�b�C�<��	�ISaQt��k4f��u^�<yT"a3�	c"��3���`�j�b�<)��Sz���fߟ/�lfLXb�<a�"��0>��`��ѐ����iE�<�G�H"G�F	��΁1��a�EM�[�<q��^�IV� ƍ	��jQ��lFB�<A������ҕ��720!C���y�<Q���6�r�S�&3��� ��}�<q2ᎋ�P����1u�{W�Lq�<qs
"7��:�j<�Y8dK�x�<1�̚9ZXC��;�F��w��m�<�&�y���AJ u�`@F��g�<Id >P�8���G���k[g�<9�g���H�'�6y���	#��x�<�%�J����S��0{���I�<yͶ,Z�=�K
�X0��B�<ɱF�X���[���|�b�+�KRD�<�1*�(i��K�d�:#ܮd��j�^�<1'�4�$�q���n��jfl�W�<�v�U��00%�����S�<�1MB�]oR�8v	��� ���Q�<��T�A�%"aC�x��Xu��P�<ie�Yڎ���E��� �w�<�!F�_8|�[�c�T��a�	J�<�!���h����f
:�h9����F�<9��W�6�`����=i���A�<� x��.�'3V��R�	?ef�y�"OT��eˑ����2�:D"�"ON��2�E�@j$����y���*O�uj�	�	a6F܃�ϲ$F� 3�'V�pj�!T�i��s�ا^FR�r�'���[�\�ԅ�R"��$����'��883�\�P�]`Rɛ���b�' j���i>Wޞ�{�a�'?ےm��'�2t�P�KbW�����P�ma"PY�'� =Ig�"����CH�`.��
�'�>4��)݂rd���
+3f�#
�'G,Q荄U���p�YB�A��'������Z!ې��5Dy���'��h�V�y	�\����i>I(�'�(U����M"h�8��K�&؋�'{^�!��*Gz0���Nq�ԆȓH�8����03>��@�ηo��t��J��B�.؆2;��I�0g�q��;0��RF#Җk�XfJ��쥄ȓ1��k3�^�9}����O��  �ȓ���RL���(!�C�BZ�)�ʓ2��3�+�©ȃCP"�B�I���P��� �:�N2ū�(�B�	�@�i�1�2�(]k1��c��B�I7��P��D��,Qデ�C'�B�,2Xٰ^>62H;t�:��B��R�L��0+S0I�hH���5.�~C�I5|�,��E4�u�� �$�ȓE���g�	Z�>e�`�N(d:Bx��`h�Y��,L4Z�w,��=23dMk�<"BY� �V��J�@��cIh�<�A��2�H�ݨ�&�6M�`�<9�h��C�xXg��hO�u��`�<!wjS6:E���T�I���0��~�<y�C6d� �D�0�Ji!'@�<A���{|N8�&J��4��Ȳg�^]�<��(�0g��Q����O�$���G�C؟�pD�A�a���� e(��W�P'^2^� �'yp%a�ŖC, �P�
 b��0��$�d̰��e@0�S�T�^�9D��'|���CNZw,B�Ik����r�[)B4����G([��7��ny�$M�����S��Ms�aTq��"6� {^��hvb�l�<��LF�B���s��=/���b�e}Ը[%�`zLX$W�xro�O�@UYӅR�)?8�)��4�0>��A\4�(�3 �nB|H#6�ُJ-�]S�I8�6Q�"̗��?Cb�*��X
�-ۛi�0ܲ�gWg�'V���0�� �V`��K�wS�Ox����ؗ#y<�Yc&մP���p�'dP��bV37�,�b��I��dH�}�f4q�)�"l�jј�.�h��ދT��d)��C${O�I���8!!�D�5t|,��d@˔�|���g�DXA�����M�D����Ar��ϨODD�� A�
DV�g�R��E�Q�'u��D"B��ꉊ4�Qΰ3�f��m=^� �-�	ƺ4���C��~�.���0&Aa�^�ɢi�6��'��i���X�L��h�$m���yq�~p)~�6Q��̖�u���
�'�P�<i�lǄ\�ܴ;���,��4q�L��fIvM�q�]�s>@��\3WO��F���O����Tp��\�aL�J�"O�!r�K�qC3R�c�D��Q�Y0"���0�t� T9�ED�]��8�S�X��MC=s���A�Nl���	w����ׁ�b'� �rʒ�!��R;[L����S',Ȫj�n��l��K�<���VI���@�5��+�P�A���1�~�HȊ�$̤�X��g�1H
heS���P�M�A"O�TR�ȇy*(Mے)P5Vt�U� bXE|9���mTaA�J��>��4PN:Q���_�PeT/$��
�k%D���ĳ6���A�hՁ\�R`�U�ߡ^J=��+倓
�j}���� � Z@�n��6�܅툱�V�'U��)SM���}Z��K,m��d�b2"-�8:5��G<��$U�Vp<���\�za��?��RTh��@��$?i0E�F?�)Q��ϥ88�����<D�ؐ�r��E�פʆ0[��z(����%��f�6��N<E�-�=K�ݹ�nT.z,�&�2�y��Kl�ͫ�ܘ-P��(�<��I�q�8�h�A�p<q�-�/���t���?�$�&]X�� �&�3.1|�C��4BG�T#s,C�YH��6	nh<��,�'.��xa!��"��z�I�'9<pkP哋/�\s#24;�h��!�1�fB��R8P��B��Y�#�7/�B�	�� �v��B)v���FS�s!�C䉆g
r=C�D	RQ
La��2�B�H<Ix��U�b6�X�D�Z4C�I�8������9;�DW.>/lC�	�?Dzm����h���٠�C�`�>B�I�Zm p���䴅��"�33�LC�	�EX��ՉG���9�ǋABFC�ɔ%��P�ǥ�Jw�-��B��8C�I'"1xp�DL�kP�ע>S��B䉣8�P��mB� d49%ě��B�	=md����%&aH����0�B�Ƀ`�xQ4��������J;W��B�I2�I�R��A2���
CB>B��,P/ڍ#��P�Qӊ�J��]/h�B�	�K���9p�̳;Tv�Q�7�
C�ɥ
�$�p�/�_�F�b��L��C�ɌU�<(rϋ:`'.L(5
��R�jB�	3]����d��'Mi(��4�  1�B�I�^���Q'e�<_6(Z�-?w�B䉝[TDIb5
\���,�u'LC�I*;�4;v��S�@Ԣ��(<C�C4�ؕ�_23�Uq���$e6�C�	�M�d�a�T���!��Bs�<Xw"O (bj�>3j�I�I�yd4��"O�ik`珵*{�Y�@�еEa��R"OVmZ㍓�x�Ux$�
Nޅp�"OȔP��-i� l���,D�	9�"O܍�p�	�W$�d2r)���`̳0"O��$,�*��95�S-��ر"O�Q���2�@p���Ȩc�� �"O~@A�,�/܄�b��;��%�w"O�  �%ю}ʐ���pX.ͩp"O���I���m�wlؠ1�rr�"O�{EƄ%6c��PN��-x�"O��J��֥4��us+A�M��Ya�"O~�Csl��w�"�:K����"O��2C,ȽW1�����tn2�"O � ��B�iK�o<A�  K�"O�dqo��3T�y+2V�9�����"OlF��O�����L��hY"O̱�sIV	 ���K�E5rA�T"O��1gn
�D�MXu�?,��<Z�"O(A	�n�+]%"�
Ӄ7�Lt�U"O�U�vmO#�(��R�\Q&Ь1�"OT��B�9s.�Bc�Y�Uz!3"OT��GF�G�T̑t�8d���a"On����$Ze�$�e�$`�1BE"OT����Y�����oJ|)��"Oδh��h6�j��T�����"Oh	X�
5`�>L��O�U�^"O��8�+ιB�Q3'�B	fY�"O�x�Hϳ&� ��9y���"O� ��*�-%p��5�@9r��A��"O]�we��
��p��޷���[%"Otdp��G�PzEr7��.|��!�NO���z�_4W���e�2<Oh� E
�u���P��`����"O��A�#�2��a�P��X<Z�"O��(C�/��$���fu"O��Q�H��lY�������p5"O���Ĩ�����a�;N����F"OP=#&'�{��Aҳ�Y�A70��"OR`���VzDh�,�R0���"O�Q�pƔ	o��@5��.n�Y�A"O�tAʞ�h�`}�di�+\Z�3a"O@4��$̚m&��dK�&p@��"O�(è�N&�l�S2 2H���"O@Qkr
�oe|�2��5~�I�"O���\�4��A'��L�8���"O̘�'��0F���%W!È!�"O> �gDY�A4�0�e �M�.ٻP"O�X�ì�pjL��'�0c�"O�-���΀Ӗ��U�Lt��"O�{�K\���]�#�^�f�K�"O�A'���0{"��R!T�w��l��"O����Gh}8� �1 v]�"O�q�T�N�+������[gq<�k�"O6t�3jU(d]�l��-�-\�Q)�"O2�b���ڄ��*x�"O��#��\zD�NO����"Oԝ�LK8�xS���.u���� "O��T	s�����Я2����p"O�,�c�P�{m4�F�T�W�6�t*O$@h%�U��l5c�����IC	�'�jl
f�ѻz�^�A��\�S��uC�'g�8�e1!1^�����5~o���'��y��+~-��2W��~�lq	�'�D���<Qj���LK�G�|��
�'�><; �G5�(�aQ�.S� �k
�'��|8p�
u�Ƶ�`��O���	�'�jY"��P�z?"4P�B�@�`I	�'c�L2�bC9d9,h{B�%;���q�']�YX��Q�AJ䵙��֙/�� �'*`�QQ��=+$��c�;,�IK�'���gE�{$�e� �&f�x)�'�^��'K[�T��L�J>T���'ư!4A�nYrGÆ9l AK�'�t<�� 8�J�����8�@u��'w���UD6:�X�S�G�C� ��'%΅`U��2H��`�.10c�d��'��U��q`t(#�
�.��e�'߾�K��)mC,Rt�S�7J�(��'�	�&*-l
dMM�  X��'dу4�"�ɐc!ݠ:�iS
�'hx�aʡT)�w�R�t4���	�'X ��bk�s�:)�����Hա�'à�ңoTpG��p�@!O}��'��F/Q�CF�-qO��Kk��'^� �ef�����C.+�U(�'�n��O Jez9�"M� H��'Z:�h�י���L�	B�
�'�Xe#�ӻ��y�&�0l���'�l{�)W I�|�[�*ֵ_�2I��']NV�ZUA�<��FI�D�;�'��ܩ�&ŋ,��	�B�D�m�H-
�'Ȍ���cP�7�����H�3�UY�'.�e*�b�'�ܙa�dǸ�|�A��� tq�F�]�y���7��c*���"O�'
�	s���B�l�>H���"O��؁C�DK�اɂ�c�TP"OLuH4ǎ\J<�aj� /�l�J�"O<��*�7r��8��$��<R!"O��s��B>�^Uc!(��qܺ04"O�-�W%)T��\!W�(��a��"O��R��� z�e��+�����"O��Eؤ��E͏-kР�u"Ozq`@��)����>�<	�"OXs�/�k��IoZ/J��()v"O|L��i,j2j���GM3k��
"Onm!�"��J� ��e�����A'"O��j����<$�dӤ唳hz�`Z "O@Ai�ߍ�>YHd�*��	"O�СWj�.&��QK��0)�
xb�"O�M��M�i(�pU�[>E�֤��"Op!��,	n��W�:S�@� 1"O��P�P�nLn�K"HP�+��t`$"OX�pșm]�y�RE�#c��iT"Oj�b�@ID���s���M�|�1�"O<$��jY�Ŋ��/S� ��V"Ox)QS���F��	���-^<L�{"O��A ��qf��i�ݫo%\�c�"O���'!p)*����|��Q2�"OpL;�@���AZ� #�J��F�!��M��-H������u*tÄ]�!���,����'5|��!B
�!��		M�����X�|�=y#��!��];!}J��Ҡʭ���"�K��oz!�ϑ/�ܵ#�ڇM�.�����	8�!�Dʲ�.y�A���Bٱ�ɻ$�!�[�^�i��8�|�*g���!�]TB�*QꎅY��q�"H��!�D�D�4z%��P�F4K4- 'e{!�\�cH��%��`��ʒm16h!�d«B��죦⒚�`��ɛ1?U!�C������m[.{�ִ�F��=
8!�2x�5K�f�2-�"�H�iH�I+!�d�	ޖ@h�lV��qsH_.!�r���`J�f��S0��!�DK� � M�4U��}cd����!�d44���s⪙;6���T�!�!��|�Zժ ͜�+�h�IP��S�!� B����"U�E\*��� E�!�$ʗ1�Z�� �fX�9 �K3�!�	k�朸S�B#�ԥ*�W�!�	���"�#HE�d"��U�!�_�a�x� 6h 20��;WƇ��PyB�7LG䬸%���6f���y2���|���A�,��y�����y��B(1���@Ţ�#-�J'��yҮ�mi�� ��Y� a��& ��yb/O�Hfy�����0+҅���y��JH��9�Gְu>z��%�D��y��==Cr��4<{|x��n�.�yA( D1�p��};׊�#�0<)��C�V�=a%���ڬ�g[:@�!�D˲wKD��(�0��52��Z8!��ѹZbT��� D��6e��H!�	�J��s�2����3�!�$M.0��e	7~��)s�_�!��/!;�E9f�֭ ��E���!�d��8�X4 g�,� 6��ms!�� ��Tȕ)%@8i`�F�  �"O0 	ç��n+n%A�)�`���G"O��H4旘_�-:"ȍ�0Hz8W"O�p�ԇƩw0���T�Й9\�eR&"OHI�B�ի5|z�;萢Y���"O:`i�oy`����+.,�5"O~t9V�G!*Zy�F甌c�`�$"O�p�U�8{;�e�bK�L��i�"O�]8eD�0-��)I���¥�"O���ɑ��"	�b&�y��i"O�t�J�!  p��PL�$�r"O@���葕F�$8�π89��cB"OΨj�[h�b��w�³D�D��"OD��5�����.��+7"O2T����JʢI�GǄ�<���G"O�K�D�V�4ұ�K
N�8�"Oh@30޽�t��8�fd1�"Ol�ҲiОi� e"4iV[�θ� "O<�� �4jV�+�ȕ��z��"O�uKd�q��8��fF"P�¤�d"O�1��g�T@آ�� f��%�"O(M�A�F�\z��4��;m�x�E"Oڠzb���^zΕ��j!�-��"Op�"��ֆ~���z����F��4"Or��G�V !J�d9�
���(��"O0Ih�ƒ<"z���PIߚf)�#"O�$0"�?JpK�V�+�Z��d"ODpA�'��AY!-݆�z���"OJ ���Z,p�S�숾�n9ZU"O<� EёR:fc'-ց~~x��"O��A�,�ZP����:g�p���"O"l�,]�@5lr�\#gxl��"O�Q	TA�Dv�	�jSm*�"Ofeb/H�p�X���G&9S�\��"O��kPf_n��pp���$I�B"OR4�u]�S ���cE�M��|@�"O��	V�D�?i��@�ۂk�Je�5"Oai�k�9,3&Ɉ���:`f��zE"O�0 ���t�
�;� `�"O�qs��F6���<�z�r�"O&��7'�5ܘ���_�T�*���"O�j��[�f�:��Ô�0DC�"ON�"�[[����`�=0�ZP�"O ����
�5v��cm��� (q"OH��!� io����n��^��	2T"Ó3�n���tT!���&�~�9r"O$��6��J�(���Y�~��EQ0"O�����Rg�Qb��'��)r"OF�c�JJ!����o��j��A��"Ol�8@��A�!\,��H:�"O�! �'�(B�(��7{h�T0�"Of���
O�m�|y���c�����"OJ�qd$ � �H���� �"O��䈄3-?Z��4B_'#0���6"OĴ����'6A.����6|쀲�"O��`���t�f1�����d� �r!"OJ����z��Q �.�:'�BE±"O��C'�߿gp`!�U/A:E�|��"O<���Dl�"��0�Ā �K�"OiR����/W�!*r��(PMp���"O�EX��G)B�*�0�&Ͽq8heC!"O Pː)M�P1ҙ�be�!$�%�A"Oj�`Ʉf���Bd�F�ډ0"O�i3W��,d�&i�"��&y��"O� t�[fE��X S�h6��A7"OZ��>&\��3�~�xQT"O�t��19F5!E'ܹM|.8`�"O���K�,Z����D��y���E�r��EM��>�z����
��y�hH��y�EL�Ƕ���#V��y�G|��ئ��{� �R�M���yBg@>kp��rɛ�ulLh𴫆�y�l�:?,,	3���s��8�'����yr包呂�S�ؽ~��� �)�y��%)�)ۇ(�_���Ye��1�yb(��z��r$�P�r<zq"��y"NU�~���S�Y�O=�p�$ٹ�y���H�U��c�/zJr�0��'�y�L8
X���.�'lP��8._;�yRA�m�lHR6��#f�" �e�U��y�j�C)��yC�g[,T�%%ݡ�y�)���nh�֭M�W)%�4F��yBg�y먉���3PY�01c ��y��^���h"�P�A2���1Y,�y�`5�d��!8�	�#N�y2n �=f<��@�b# ����yҬΎa�$ 1�6^qvlB�N�1�y���D���b5KZ��uG_��y� Z{��5Ι�/���HC�yB�[�}�P{�`�:h8��$�ֹ�y��
>a��A�ɖ����4ķ�y�JF��7�݀�t���)�yL�"L�����6���)G4�y��&BJ�m�g
�Im�=KBg� �yR��),q�`�\9zeP��3�y�J�.@�0��q(��<�5��	���yB�\"uln��
86@Q��a���y�/�v��d�ӑ3*f�����y�bF�y�<I7��}���b:�y���2Ge�qr&.4}�<<{���+�y�fõ��t��O�q�dad����y��<Yx�L*FeAc�q3�O	��yb+O�L���X�%B �T����_9�y�CW=���F'*xmε�	Z<�y�nL~���Xy�|�;�$���y@�h�&�0��P�nJHJ��W0�y��;Vnm���\}F�i	0���y���Q��F��/���梑?�yB��
,�f)s�j�%N6��`ē!�y2�X�ߜ��Rz/�0åJ�y�/NF	�����˲m��X�4k̓�y@V�:�0T�����` 8�ac�W��y¡�xf�l �GPb��b��'�yBi�<P��Tp�����l��yb�I�<��4yЂ�'=����yBb"$�.��4�C�S��sׇ�y"�ų.�2��&�J1A�^�����yR�Y�p̤b�N��9������y���G=��3�"�T�YЊ�y�Οxi�3�g�(|a�"����y�������sLX���Q�Qa��y���/2�P��ۥ?h�J���y�Z�0*�Q��m��$��5pℊ�y�F&�:1�J�2�4�kV��)�yR��2٘�F�&�J[�hY��yRMXj�8�fO��8��A0�yR➬o5�9���۞����y��3��1A�^r���9�	��y
� D��1/ʶj�Թ�6O�.dY��C�"O��G�8���yîȮ5bj8�"O�Y�gO��t�T��Cn�:D�v"O`���SC�*��T,@"|��"OKGT�v �N��V|�$qf��yB.�
@]�h��!�<B�`�2�:�yR�U�8� �K���8h��9P&�y�D�q�D��M�]=��贃�"�yr�u��+'���h`�`��y��������1nN܉-Z��y��κai�i��i[()^�{�O��yb']�4���5)x�Q����y"��#H���A���l ��Ɩ��y�C��)��|RX:{D�ʡN��y [D�u�Ru\��",�/�y2%_&	���c_r^0M��æ�yҋ^.���〈dР�Z1M$�y2���?�"�V啒Q��=���Z��y"cǸ-�Lѣ�
NH��q�T*�y��T��`�����;�J T	�y�JV�,K��J��K�Tpm���R�yҏ�7�A�RLT"[^���5#�'�y�Q�H#F\{$�)O��e�4��"�y��v�Dī��B�pd�p����y�P�sdH�jr�`\�����y���7���0�U�NQS$�y�dY�@�>츱ܵE��|!��/�y����LAЧ�6%l��Ɠ�yR�7|�0x�t��)�:h�����y2�t�� f`�&^1�V�]*�yR�	����̖�9�Y9F�ۘ�y2�K�m���2fCн
��݈bF���y�l^+o�a�S	�$���K�"�y"��=�}A.�>��a�׃�y��G�5��u{Q]�9����u���y�%'0�r �Q��|����U.��y��%���R�J�|�F����yR���<�!�Ň����O��y�`�;ko��D�(~~�4�W
B��yB83_h+Q)�a��]�'�9�Py�ˢ e4�bB�O�fʉc7�J�<	���P�Ȃ��*@���@bE�<!�	�yB�pz���J��T�h�<Ia�D���,��*/!��  L�\�<�p��hS<I��ޤv| q�s#�L�<A��� zFx�'C
�
�؉JA�@�<I��GX��-��q��1�>�����(q��ڐ,ҀYq�-w��@a�"OP)Ja�c�6��9#j�lʅ"O0I�l�&�s���7Q����"Or�K���^�`��w�%Cc�e["O��'�E�W6�I@��-?}�ubR"OT�wQ�o��	PЄ\�ku\`{�"O������l�ٻ�(h&�Kr"O������H��ƣ9
X�"O��g�!����ϗ�G����"Of��F�U�/��Yp�۳q�T�"O���კ�%?8�#��9��PRQ"OtP9���>c�!���?n�f��@"O�8�L]�&vرР��g'4$ �"O2�!�8�,r���)�H�"O���O�?SkJ�*�����!��"O赡��{��i��� ߦm�"OF�I���r����tL�w��8�"O� }�s�	�^8\�{G,P��rI�"O��s��۩3ʩ�Ə'O�b��"O�}�� S�Qq��A�¤@"O��F�N�8�p�����u6"O<���%�5�͛��	rC�h��"O�͓�Nn���b$�_;PY C"O�"M 
2Eh⼲hy�ESy�<C�Ľ:#����\�12��#�K�<I��\�r1�Ij��
0s�N9��Ä~�<�W���2�xْ��E�C��lh2�	~�<yP%ͼ,A�@��Zx���3d�I{�<y_X��#!fāA�CߍrsB@�ȓ)&�x���B�~h�P�&IIOr6نȓ]j��/��Kn�$�rn-#`��ȓw@ �h3阳�r!w��Ҹ�ȓ�l��ԫ@�_n�@�7&Dфȓ!6�00g�̭M����q�q���w�pM��Iʂy��Άm90|��wlH"7
��	��yZ#�"ybP��ȓ� P���7`�zdz�m�k�q�ȓ��a"Bm/wF�i���=5d��ȓ&"�A&�S߈����R��rŇȓ����]������%�`�ȓ}�������-�;���j��݇�A���t�W(nq����ȎQŚ��ȓ=��q@�V�N`����Y
�����u�h�j�Z�WR�*u�
}N�X��[�!���� h�l6��P����A���X1A*ġr������"O�]���ڥm`x�Q�+�"W�["O�9���
i��Y��&|3"O�db卋D�P��t��t8�uc"O��bF�L(+9�䒰狗
T�"O��%ϻ{
��RG�{ߦ��f"OP�s��X�m���*s ����"O0�RiY�.2e��nY��j�S"O�PS��>�hّ��&n2�5�p"OP�2�	Y�����x<���"O�-C�A� :�)B\_�b�r�˟N�<A�ܑ��� �H�6Z�h��,H�<��F];�B��"����q��S\�<��  ���` S"=����̚T�<����Z��cb��)ҖT5$PP�<��i��&�^����w4�I#���c�<��J��G,<J�֓}�0�#@D_�<9��$nv�1�o#���B5G�<�#!�.�@5j�U�����^�<�T�*`f%qB�
 .	���]X�<��ͨhh��㣣��,�S��X�<ٶ��"-��q���Q?��c�!KQ�<a�M\�J��@f՚6)��كC�e�<�v
���֐�� Փ�@=iD/^�<�P�qQ�x�5�*o2� �"�\�<��u�I�Q�Y(>V\��%�WW�<6�J�N4zh!�W�x٫��h�<y���8L M�wf�rX8�����m�<9PKڗg�j����9\Gt!a���j�<�D��_�$�J��ùy��L�T��g�<���#nTe�wF�y�ڱ1!o
b�<��D4Y�t�J%���&����m�[�<��G@p� � Ȩ�+Bi�Z�<9�KF���<�͇�M�����X�<��ݸp�,�@��O�K6�sba�U�<��	v��p���wv�T�B�U�<� ��RǭJ1I�13"%S�D�v�D"O�Y²΅�"�`��G���V���"OP�4d�+YȞx[�S@ڴ�@"O��"��U�@n��:�g��-Z��q"O��A.͒Z�b�X�ɠPR�|*g"OL�i��	�pcDM�H��¶"O�l��_��y{B�R-V=:���"OT%����d��`��@�Rȴ1�6"OD�j��>x�
mN�a��lZV"O�Y��?Nq@)����G�p�1"O��q�E	����m@�.�B(Z�J�ON�{`���M�O?�ɥ\�긻��מ6͈y�e�˶	 ]¥ã=:騀��k���#&�8h�6�>I���H��/��LL&�+��V�nJ1�g�i8����A�Rm��0f�n��b������4i��s��#����S ��3�I�u�i��y0��'�2�f�p��/���{�)�@�,��@��="���檟d����̅�==�xs-=C6uy�0T/V�<Q�i\&6�,��޺��B�?xP[�@F�
�]�c=+>�'���# �`2r�'b�'�םΟ4lZlbX�h�e� 豉��f���Xt��mpXX�`��/ �Õ�W��bUA�=241%��'��2�d߈Cs�O�,� Y��R�9��8����&�}�8C�ȩfL9��'̑9wn[�59�$J���#�%����O�QQ�c�Op8lKt��<��'����І�9��RW���	T��w!�dE�t�z���J=t��zD䊺@V���4Qd�v�|R�O��tW��BrK��p��e��`G�Iz�q��,�tCv��a�Fx�t�ɛT;�ģR#כ)@|c,�|AJ��L�:�X�R�C�
ƮE MY>����(�LQ/B��EB�!� q���ut�*X�.av4��44�QɒiN�^2��
4� ��_3�����?P -)d.M�i厞nĝY$P��M���������?9�ڟ.�aPH)C�@�@r���`3���q"O*(�
����[�f��	6P� ��O�lZ/�M/O�xBc��̦��	�8�O{*��〵#�x��B�	6�l���ݤk>�$�O&���0ݓ�E�&�����E�+[4���L�pa���Q,�)�c�DhU���]�'Hm����b� �� %���Ƒ?�He{��ش�"0p��H�l@K��*7[d����SQj�~�V�	2�M3w�&��i���K'Mߪm�h@��Is^�	$+�O@�"~���*{�T�3��4]�2��5�f_��$Ħ��զ]:�lӚB�:�(O1u� ��b�����Cۏ�MC���?�,���T,�O���x�\����P ք�F�t���s��E�Y֩ !� �jAh9!TL̯s�x�t�\�4
����?�����U(k�$��H]����:�G���#v��t��u
d[�j�$�i�7i����%���g\���5v�^2�@A���Ns �r$h��M{Sf�������M����f�s�ā9e�4:U�C���<ٱ��O���>ړ��'���D�ҴIa�����O�Q�ȑ��ĝצqz�4�?A�i{ҏ̐dg�0Rl�"f#��I.>�a��"e������s���mJ��IП�����!_w�´iC�M�� ͺ~0d0! �[֒�P�"=*z ��D�%��լ"A����4�}���D|�ml^�!ȕ�(���SGރ< H��4yU|�2���|;��S��JP�혹'M>\���҃$�dP=%�py��H(ஈq$o��B?���_O������M�b�~�'�BV��#���-Jp���W�L,��b���>ؐx�C�uC��z�NZ*�*���I�M��4 ��V�|\>I�>IѮV0 >  �   W   Ĵ���	��Z��wI�/ʜ�cd�<��k٥���qe�H�4��6_2<<�3�ʄmn���s:�j�����Q�e_�c�7-⦅3ٴJ~�*�	_y䟛nSt���|F��Gb��*pH�A�IP���=Y�D3n�d7M�0e�R�3C���*���)�דc���(�Q�d-�.6��ɓ	�����ƌ
=���&?�,PtA���wL̴_��e�6�^�A�����X}��
W��P7�x�ϓ���{�OY���q�v*]*�ʐY��\;0�I��y��& W�����t
�C���Q��Փ���$�f�jd��$Nt�;�ͷ���ec��7�F%a��<� ��0�x$�<�Q�d�Z�,p��"D�kt`��c��컑�I�}D�i�J�Q�Ra�e�\��m��O5�O��Q�O����$��������YK��>� �3�\��RUk�%Z��1���@�
�nӔH���O�T�ůC��~<��^q��ȉ�&�/*W�Oܬq������(o��Za��vl�b�":39�I"#�PK����'���B�
�XZ(�\�EI�O֨9��˚�?���'p	���=e��7o c�Be|"<YEH3�$0k\�0�n��
D�(�a��/��dƾ�O\� H<Q�OlA�[e�`��bC	�F������'�Dʓ$����=R���O��Ē��6�O�-uj�:�O'��� ��L��'�`|Fx�#�s��&��T�pÔ�M��z�	��@��I�Y��H��I!E>qq��s�<�3k�7#stB�I�e�l�  �5;vZ4��"O0��7��o_>��Ǝ]82���d"Op�Zg�U$�����Zf��:6"O���U�_�<yR1��$}���"O�@���]�0�B��jx��"O��4��9/����]3"O��r@"O��bFւSvh!A��L(yL�Ě "OX��"ၹP���DN�$��09�"Ol��4L7�qJ�ʚ�n��K�"On$  �
k��d�'H�P��u"O:���,,KZ�Jr׻"�|ّ�"O�m�FÒ "��������P"O��0C�؍���c�E/Q]P���"O�噇����(�M���
M�'"O(�U!��|�'�͜w5�3�"OZmyv��nmH����>{,$�x�"O,8��;]H�ۖ�ސPXш�"O��r�� ,~�Q���^����"O�T�BP   h
  )  �  @!  C(  �0  7  V=  �C  �I  ~Q  	X  _^  �d  �j  +q  pw  �}  J�   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl�
�;�>O�1"�'"d:t&�����.}�ȕ��4��DK���8pp�hICAP
;��i��fݕ(e"��?���?j��~��e#�HծW���d�9gCL� �+_�Z�SfF\Pbf�b��+�u�͓�(���'�b��F%��%����)Hk�xÕ��-4"r�+K�Op�J1OS�#�r!��������"L�����������{'!�9�a���9i������D����ɖ_�$��޴���O�݊����t���O���!��/T��}��#�
�#�"�'���'��C��&r���?)�'���D�{�H`��5��Dc�ꔃ,��2<O�m���3Ւy��Q1�"��U������~BeǷ~Z��O8Ȉơ�l�ft�r�s�p����?���?����?����?�+�`�65`� ���6[������+��$��u1޴=����>u�id��
%w�2I�B�O�������j.�J�O`��g�~�'.����iL�Odrx�%��=�]c�զ}��$ 	Ɨ$��� �̛�f�Ni�Źix$7- ��S�?m�0%?�$gFF'	5��)@�S 	H��Uƃ��M��fIy$|J�cH�e��x�Ǭ��n=|�Q�⃧=�6�s�<(oZ�i��� o�"-����5� �#S-ܴU����^��Mo~Ӯ�mچ;�����^3 9��Z���2v*R�5Jb�!�%I ?�3�+� �"�k$�AW�d ڴ7��*hӲ4�Û%H�����-X�$��4>ZF���n�z#�$K���>i�}�	�b��8%�K-]�ʸz��~-,��'C�O>��S�w�L��2�V�p�*�R�I�O����	��H7투�M�̟@4�q�\�^�����Yw���'F�I���	�|�%b�aH��!�߅1��L:�4+Xp��DM7,��Da�c@=3Q��9ÓZ�f#�5,p���I%�?Q"HI	�e� �A�Svz1����{���pm�O���XMy"H�
+��1�B�o{������?���?Q���d>O8�ȅ�&`� �a j�AX�92p�'(
7��>;��r׀��f�(��F
�b��l�Y�������OV���T�ѻy�����[�`��r�"O0��e+������;\�9��"O>I�e�<2��|��[6��k�"O��"�D�+�&�z&	H�����`"O�={G�Ӯr%P���i�s��Jt"O�4J"dV:0��s��A;T�e�5�'��X����(J!�D�=����9-���ȓ|��q��<RۆMC'�5��ȓ�X��wg�3@3ԥ�H�&;4$���{�*Qi�鑻9v,�:���!ժ]�ȓr;nqy�IP��>D��S�,�͆ȓ?1F�S�A���"�l)��O�<���Qb8�x� S�TǺu����RD^���$D� ��NH%n���@�,`�uk�C.D��#F�W��<��Th�'W���)D�DPQ%X����sJ$C��4D�0HDd�-���6�Ⱦr
�ye*2<O�H3������I�����21Y@k�����b��4���'���9�'[��'�\� s�F�FA�6i����j�J��t,��9J{3 U�?���D�<X1BUPC�7�v��a�.H%�i�6�Y���E{�o��-3t`3��'�X���?�'�iYR
���*SG��'��z���0q#�՟�?E�dL��'3r�`q�� m[�Az�b���'Z�	H�O��7m�?Av����F 8KЎ��2C�|�oZv�Id�)�'QU�����Z�L�KpD�uh�r ]�yL77:+�B�O�X��
5�y�M^W���ʃB	�t���1p���yX3�L�p��
<V��D�ˑ��y�W1Lv��F'�UC�1��V*�yb��7W@=a-V˞i��C1,>���|R��e_���' ��'T�+a|nԑp��n�����O�6����@��M���i�8pZv�@$U�S���'��`��cEO "m%-��«<8"�i��M"�`������O����ƛE?Y1,։lZ�Z3�6G�X�ʔ��M��R�4����Ohb>�d�O.��@�2Z|���EH��L�7� wB��DPG�o� Y���D���%�P"z���'�F6X�)&���?ɖ'�Z��V���J�^������vM����H������'���'	Үݙ�I��t�'S}�	�Pe��2�z��7�O%����?9F�P��J�.���Z�Y���"ANSU`ȥo=Sǃ Ww�捨eiT��ϓTt��E9|�Q�QK<MX��E��X��̟��?1��)��v�	�m�4۰e�&[k�!��H�'!��`+M&��p��c��'i7��O�~]rA��i��S�8��
s��D�Դ�e��.u��$�<9��?���<�*��"ա ���&�Ɔ�y
� ���S�?��$�્<�<@�E�'��y �#UlM�t�''��yB��a��+g��P�V��@�/�0<Y���ݴ�?���c��R�dL�s�y���?�@I����?����?����'Ø'�
4�d�"���ZS��./Wq���s<�M�N���!00,�u��[��?y(OXh(@!�ߦU��럠�O����F�'���{ծĶ&d��[�]�E��c�'�B�P�cB�T>�'Tp�r��t�كo�n<B���O�T���)§k�	h���6���ѳ��/'zB��'j�1��#Bɧ��qC"g qݔaӃ�ѾM�jQ��"O`|kǇP�x�-CC�$:p�r�ɠ�h��TQ�F�>^&�l���&^�B0��i����O��
�E�*~b�'���'��݉1�|�eA]�\������ҩh�(�HZADb�,߉#�"��4�S��%��'���UhK�7T�A�'��d0L��J��a�n����oL ��f�ĸƘO)�9�Ic?!��1B�ź���$4�4ARee]�M�dS��٦)�O���:&������*Z�#k��TG�\�a�S�<�Ed�2R����K�H�v�Vy 1��|j�����P��N��iM�R�@\!CO�-";��y��ڂw����O(���O\쮻�?�����!%WD���Oڇe��!�"�#x�iS�'��%�K�2kҍq�N�L�ĩ�C��xRcK�1�B���F��:'
���Ģ�Ҝb��tc����Sk�m��ɇ.�%�e�_��y�-(�����H>[x�������$��&�|R�
�YA�'�?ف��<K6����%RU�PU@�?1����XB���?1�Oer�R#L�-c3\�F�FD_B�la��T�q�ne��7G���e��0:��3e.�c���?�DA
DP��#�rII���]�L� ��Oz�,?�TH�fņ0��%�%�I�x�ܒO��)LO�=���F+FA��F#d�P�A��'���5��c�É"(͌T�2MV;;J�\��Z�ʶ����OʧU�4�1��K���c")C����C�3Q;�|h��? bQz�2���$�,P�[%�V��O��S�0������E��1jS�R
9T��'��u��',��� �Y���ݤw��{���3�TJުby���K��c���� �'"��3�t���wӈ�D §o���c�P�mJ~���j����&���Iʟ���{y��'*��,N]�p��oF�N��`!�9hT�?�u�i��6�.��2)�b,�!$Cs\��P7�f,o̟`�	̟̃�(�z����I���������yJd���Ȇ4q���<�4�BV�.�^�C��I�(���	H�S7~�'���m&҆�H��f�5���^s���k"��d�
��f ߲<��Q��Z>M�W�ן|�>�C.0T����eJE��j�85^�Ul���M���T"�������D�Oxxp#ύ4��#�W�Lr��O���<������I�-b�YSm�&B'��!�H,74�Z��v"fӀ�O��'���I���tQm�('E`U�G�1@�{�J��+�f���O~�D�O�p�;�?������ж��$��͗�r^��#�P�Lm���!�<уTgȀ7�Y�6	��+� �Gyr�O�Ks�B���,�iQ�S�|R	ہ ܫPK� qNߗ?`�A9��ب'aGyb�Q0@�vP9#���)�P�_�|������%:��O�q����^�h�:t�
��� �B"O����R
X�f��� �[�T���|�t���d�<a�K� |���ş@�Ǜ�&��IŦ��h5P�;������I�a������Χ�b b��Z�[�hZ`Ć�fVQ*ffT�|u�rd�x�R�P���:ʓ�Hѐ�b�/��̊��	�bbnm�R�M5�e&S$X��h�1�@�2��X� ԑN�Q� ���O`l�����4:ҖmIaP,<�!/σw�'Ca| Q�Nf���)��p2�_���?�4�'Zb�yfMĲ4�����n�аr����'�J9���i�%��@��<o4l�HQ��`�k-D�DH�kU\��b.�d���p��&D�X�qF�(#ؑ����0�0y�E&D��0!Si7��p�!wˈ`4�#D�<B�,�}��{ua�S$J8[�� D��I�ܽ7~��e��&���O0 ��)�sU���N?�y��|Qp!�'�r=S0暇C<d��&ʓ�o�z���'��HCV �hP ���e�`}I�'�p8&�%<*E�W�a��`��'��p�CFڷ:ڨ��g,6_P,M	�'���j�lD2F��0i��^�$R�U@,O��4�'rq���G�P�Ȧf�;�8ę��� ܹң��T���Sb8��9��"O2�;e��5�Q����_��Y�"Oޭ�&�*.���`̥>���c"OV�93��+#+�A('	N ���'���X�'�|*�6h�@1�6�N�"TL8�
�'o@�@t��S�L)a��������'=��%�j�@U��7%�X��'SX��A �={_�y�� N�*դ���'�8В��j���Z%+űMٮl!�'J��5�����U�D
L8��8- Q?]�D�;g���ဧם�b�j7D����N��B�X���9u���sPL8D��2p��:<+�X�0w��-�P$+D�`���(e(�dxǌS-i�P�f�(D�@ U ̋X�n Z@㎬��i֩*D�p�d���2N�Dz�-G/Zߔe����O&���)�'6����s��L�p�����1V��:�'�� ���9�41�%���.x��'L�św���<��9	aM�+���0
�'i�%����$<�J��`�κ$pU�	�'Q^Lj'����d��B�"�h���'e\ۆ)�!3��$RG	�	�Y�.O2q�d�'�)��ޭ~��k���4|��Y��'���+�D�;���P#�!oDd��
�'�`��5'��܀�B;q���'���xS#�%\�^�X�m��ֱ��'t���s�v�J���G��H��8:"����X�QË,\����P�"�*�ȓ�I� &?�ʀI��C3��m�ȓ\h����Z�
�!�EOl�Z��Pva!,[<&��X"L����%�ȓ[~e��`֧d�^�c�lkZ^���CL����Ⱥ.� ��1�͜-W��F{�$�쨟>̫ ��%d�[��"]r �g"OVmZ ��v ���T�.mP�H�"O�	#Ub�'�Z	[Q�S=v8�-	1"Ot� )�*�"X�#�
�G�!��"O�E�sϏ�*��i�BMY7!Q��"O �I�F���m@C	��B����'垙 ���08Ĺ��N�!!4I"a�U����ȓ_A,Y��R�d�t���6�"U;T"Ov�[�8�ҹ�(�*	-�=2S"O
	kpA�$I2�#s�I ��a"Oܹ8fnC������&'d���"OU;R!�?֨Ax�j�i�^�Q�\��X�"�O��k��?�,�������"OĐ� �[�P_N,ix:<�a"O���@ܑB�dɡ恇z�>��U"O�=�@["}��W�đ���a�"OޜI�h��p��+��u���c�'RI�'Ψ䙠�����q�@H
�'����U3Q.���c�:ix	�'�̤)3�̓~(Hܰ� �8`*�3	�'c�����`rT ֯�5y�����'鼕������*��p���>D��@�k_7Hyz�ѮY��˰�"�tٮE��NT�R����
N�$�y2�ҋ�yB��L�L�D�?9�T���O4�PyN�V�,�7$X�;L����C�s�<�G#9���A�]�3�0!7�i�<qB PB�z�T�Ʊwp`��AO�e�<�£�`Җ��N�(�� Q�F��т6�S�Ox����Y�ak�u�㠒$wK�y@R"O�=��ܦD���#Ƀ3%,\`��"O� p<����6Dct�C����U�8i��"O�T�5HL|�~����W�D��|�"O �8�N�u�B�R�G�+/�ZL��"O:��fƍ �\-)'@~��+�V�؈BK;�O\�y&��"2�� ��՗%�.,0g"O�$c�
+ZfX�ZqF�6��y�a"O
	�w��-o�� �M|g���p"O���v��:�����X@I�r "O����YpdB�9V���@�'�z)*�'9V���\��^���(�ܡ�'��5x��\� ���a�R,�j�J�'�2!��DH�_j���M�x޼
�'@�`�DT�s�}���ZX�6Hb	�'�t���'@!d敐�g̛Y�\q��'�8ؘ0�Z�6����ˎ$Y�b��dޘq�Q?�t�MCE��ÉH$V�\�K4	%D�@g,�;KWZ��B̴WV�a�#D���K��9Q�9@�H�7Jm���%'T��aEL>,t���B@�����"O�0j�I�d��T���h���"O>(@�
�I#i�F�C�%��Y���'.V}a���S4{��G�T|\j0��.�%+#)�ȓ9T��1 �h��D"T!�ȓhFZ� �1Ӏ���}�4D��+�R��#�ӧ�$,@��}i�цȓY���"��7�:�S���5H`&ņ�}���p�b��\��|C&k�3 ��Ė')�x��p9�9��ےDg��b�fر�x���T���h��\�bp^��G�	9�Z��ȓ�|DM�3s�fL��8���s�($c�oM^�@��фm�P��xo�� u�౲#I�!�����^i��	1B�����ćr�B����| �C�	�L��2 \'hC6��@�8��C�|	|u��Ɍ[B��b�%��C�	���䣵�ȅb�(���ªh�xC�	(|��[a�,�8�p�#���
B�IT�M�r���U�:@b"&A�H��=���|�O�$-P�
Һ-u:(�eж$�Z%��'�^$���Yz���mɞ����'� �!� ������W�~`�y9�'l�`胎;W�8IG�	(r��X�'�)����>k�xWU�k�T��'p����!a���"�5$9`�� ���Ex����_f�b+N�r|p����˅<khB�	�l���M*~<qy�T�D�C�I�f����&݄Q2vm�oч2� C�	. ��#�L�(��KL?�B�������ޝ@����!�f�
C�	�E�Y��Is�iB�R�p��ʓ&�2\��ɬ^�z��t��C���;%m��<RB��,
^0p�Qz�����1�JB� x�H0�5{��� E��M�$B�I�g?Ԕ0�̽x���O��Y6�C�	�iTU@N��F��['j)fS����̖����"-����%�9^��h#D�!�]�(~(���+-��Y@e�	=_�!�$�Wd&���
m�yӦeI�%�!�$N�C\^���� oXpX��ÀZ?!�W<<�DQ�I�&B�Z7�Q�!�d��t�nq(u�&Z��UpWh�5V&ўd#��"�'v��bE<6	Z̰��Y�"
Pń�)���%/Ja� ��C�I-O;�Ą�to��u�{f!����,��S�? @qHS��%J���b��F�Q�Fp0�"O��D��^��)����v}X���"OV��T�4[��T�P�C��*�1��'�нH���S�D�Xq�A�[f�t�����a� ���'�)��J�D���H���6��1��E���H��}sPٱF&j�0�ȓl�ĸ��.�� �B�̤��@��(�}z��ų�*�A�#!X����������GMȬ��`�"����'������j�RLL0dm��1,� KM�I��A����� �� 0;6&��d��nw���gP��T�'��H�ȓ(byצZ5Dƶ@"���� "D؆��<��섵0�������a�:����5>��	�}9��CvIׄ	��D��D�UN�B�	�"�d�ҧ��$���A&w�vB�I�d� p3,
�@�TJѢI7�!��W9k�ʸz0�Z�a�@���J!��{��
�BR�W�b�c�
]!�DCJ@�Ȅ�Z	R��h�587xў*�;�G4Ld�e�"S�lbsh��!���A��C",5�5�¤�5Bǐ@��Bm�$�cG	���IrI���$u��wHȲ"�=#�ةy��J�3�,��#�L��̶nTH%���?޺�ȓ8���?o`�30���A���	�O� #<E�4��4+'h�#L�1T��,t�!� �9��,b�v1�����!�,Z����ʜ34�!��\�xo!��'p�y�� !�r��A�WY!򤞲w��h�2#B�##�(ܡ��:/��H�H	�0t
�@�v��#}RH�<i&�^�IB6M��=����<T:%��=*u���<Df�¢�O8�9d��O�d�OZCf���t6�퉇-�
dS�e�d���s�J�~�P��'eT����`�Q�0sekؕI�����<+E�QH�L�W��i""A�4`���[��^�X1(Q��%ۼ|Q��C�g�O�o���&jVT�����!~t lKC
�D�'�a~�啦ciX��r�\;���ê�.��>�4U�țTK�93D�lQ�AQD���J��+�� /V&0�?��g?��IصsN.��DĆ >�^A)���j�<Y���5pRP�Տ�4� D�O�<1 �N��{R`��8:q�gSP�<�ǀ�wW(4å�ڃ1����X�<�G%�A����'&�@dHy�<�@*L�G�x�2)�_��l��I��u[<#<����O0Y �gշ$+F����o9"�c"Ok��*U���I�@I2J\���"O�5�#���"-V<�P3C߈���"O�����Q7Q�r�8r��2"O���.@6��ź��m���	u"O �7n@�\��h��$xٶ�p�'�I1
�0D��(�CO���p鈵jPp����t�c�U#TYBM:��ȗG�����N�:<)C@�*e��y�E�e�n��|`*<��慷_��`�ģ�vP*P��2�A�b�ME�y'N�?�<���I'j�'IaKg��I4t��g5e^A�'4�*�L�)�%xW�V�*��3
�'R@A�ft#&�;��F*�	q	�'���!"�"���q��4
�]!�'��-��׳���`���;��)�'��R���(�*�q����������Ί�O�;$�[�E�	P���55��ȓ]؄���E7���yd
��@��D��n���
�K�C'Ly��(�,�����S�? �t5Y�ZM2�C	 Q��xҴ"O�T����_#bm���I.�T=ʴ"O>-�gM�-\d�3�(�-���c�
-�O��}�0-4̘�<P\��.̐t��	�'<(x�$+�'�)�� �"]�F1�	�'@Lx���+L �"OQhҜ��'8���� ��c��rC� D
�'8����X!eݦ��H���T �'��QbG�W<)D�M��a��@]���	�8��I�y��u�f�ϼHS�ճ)��7i,C�	�O�du�#鐭��9�Cj>#�B�	�
 !�&��KhL3�*;U��B�ɀ��1�V�G�O�V�2�Mɱf��B䉧{�>��!��4v�\��OHp\�?�E+ڻ��	ٟ��'h�d�(Ï�@���`@n�=�(������	ʟ �I@Ɍ��Ks�@u�h����l��(|q�tk�<(�����?K� ���:�4H՚�m'�h<yרG�y��q�" �M�
 㰬�R��Q7�ظC���RkQ��3���O`�n���'R��C�j�l�燢BH�)5^�d��I
@���p�k��9���\�%�b��$�Wy� 
`l TgH7���I#Ǿ��$�O��O^���-?�a�1�,�k�'X<L�J��Q�'�*�}���O�P����B�:P�l��Ib�O�6�%�\b��'����N�0��w��|;�E`�!T?l��zy��lK�S��'�pr��)3��L�ո���W��q�ɫ��I�=�2�'d �j�r���	bcP�Ӂ/�~؈#,����I��~��s��9dn��Oq~�����9\5jcEM�.A���'�X�',2�J��Z���u���j}�0�q�Й���SQ�'H��PI�P��4�'&�lb��N��z��rc�Iǘ�@��5��O���Op8�1�>Y��i�4�(���0-������S:#,O�@���>)%�S�t�"Xxf \?�1��^
���:�'�l��H���<$SP~,6�i�W��O�L�H �Ǣp�8x�BS��Z�CAڟ��	�{��>�1 埖g�0QҊT @c8 sA��O�Q�'�
#�'���y��ً�~Be�*,�%��d��u f�z�Ɍ#�?�2�;�O����-�8���폙l�nU�"O`P�d�9>x�:�j��Iʜ���i���'����h�I_yRY>�XhZY�7�ܿxi����h��6M�O�˓�?��V?-�	Y���'aZ����-w���P ^[�Hy`A�*��O6��Sg��J�p����.��Q0'e�!��Oؘ�z'�� �xt�'���!�$��VǨdxd��iS(LK�DN� �!��-Q90]
v��'��c�cعq!��(�,Ta�D�jE���;X�!�D1!H�3ǃB/>�x�'G�m!�YPr���%�Q�Y��G�5jM!�$،f�����C�C7� ��E�X:!�dE�3 �(�S���T��1!򄝯F��q2I�6�,�	wDUA�P����?��TnP2 @�9�o6(ON4��<D�P�4)�	\�(s��x�(���<���
��8'A�&xA2@�C,�3B�i ���~="�D�X��P��)�Zd9��4va (%A��Ҡ9"+G�% ���TA�ln<�ӫ�ު��B�.B	̀i�[��RQ�N�9�EpT�J�l���˒.	�OE~�X��A��A�[%�ɜ�LY�g�!�6ypܴb;<q;aI F�V��5�T�+�X�)f�'�2)mׄU�P�;�T>�O}�5%�˵l�v�a�-E,,*@+J<�"WjX����b�<W�F�����?`	��\,���>C�Œ e;�z�ģ�i=�'����3ӛ6�p�d��<�SL�\��Ǣ��Q�CK�F���NX��04K� �h)��[]rZ� "0O|�Ey���	H�Q����Tߺ���m�"�nqj���O��Þ{W��
����}�"aK8B!�D �CF~�K6.^>E���WV-�!� �<�r��Q��{����eD!��T�`��=�7K�2�𣃍�J��5�r�e�E50�΁��hކT�v���L��@c툉;K���qBT4��h�ȓe�F=�6��(:���� !nm��S�? �Uc��@,h�~\�U��09��!�"O��J J&z���O�(�Z5�S"OR��k2�X����w�P��"Ov5��a�0�p�x�L,y,2)� "ONP���
vj�8�]0�i�S"OPC��l�:����Ě?��E"Opi�M�|�8���\e#F"Of�8�e9��!Plj�"O�|Y�!�4ji��)`�-"O����u�$08���+V찤[�"OX5j�dN�'/�a袧asf]��"O�$xp��R�Z@X�`�V�~�G"OZ=��+ pq�J?6�tre"O�E���	p>�P�m �M��av"O��)�U�h�0v"H�p�12"O���菣v6��#Vb� 褻T"O`I
� ]#O���z���,T����"O����\�J�b�.T�5*�"O��"�$ (]����uK�4p�bR!�$K6"ǀ�
��Ve��MGŒ$R�!��&ƠE��HþN'�i!�.Ob�!��"ߨQC����@4 2o5!�$�	b�p�*T��G��
4��@`!��ʱ؁`��;F]2��@��!�$�V��aj��˭E�u����!�DE7|��r��Xl�)���!��y�0j,U�>O�ai #Ϸ'!�$I�My�<h�Ò`A��K��!�D��S����o)M#Hp±�6-�!�� pĚ<K�JV�)P��˙!�$�/7vn�r�
�U��H�b���F�!�d��Bp�dZ���;�P�;�-UN!�dU�p̘��Ǘp�<�O�l1!�ہ�T��t��xv���*̨B !�� {�La4C�;Xo��ժ(8�!�D� ���cR�,E�(U�C)�
G!� �(e���U�ma�Ѓ�2!�ѷ
�ީDB�rΕ�ֆ��!�d\$���bƍHk*\sGƎx�!�$�\�L���9P.,0��d�%/!�d/�f����P(�C�$�%}!�3@ٲi:Ҍ��8��+�A�3�!�D�x"�!�IͦA/`�2�� !!�N?o{�]�p/	Yv��րB0F�!��?C�J4��[6g��rB�ТS!�dV=^�����鏪#yj�)�O�1�PylF�]�T�;�,�a7�a����y"��2P��(�"a��Z�L������y"T2�ܕ�����j}R���y���3��Jp�@{)���"�y�(K�eGn�� 埨y;�u�����y,@�d�R�An�j-"b��=�yr,�*)<z�b��Eb���ɡ���y���8O
��ҧG�
]C��E��1�y"%04��)���N��0��&�y�L	5S�8��OR=Nčhtş�y����W=2����Y9@��
5%ڷ�y�+]�25�c��@�rUS����y��Վ@� e���"
����/�y�D�?H��b����	A�k��y�i�N��!�2LLi,��`�틞�yB`�)��<S���<Z�5�b*��yrM��m ��4�>S |[ₔ!�y�*ϙC� QQ��Z)Q.Z���ā��y
� hX�r�L��N"%�O.y�mCW"O%;�� a�Ae�7v���"O��)F�JYRf�RD������"O2�/F�5���CX�N	����'^�b��dVnUP� ҷU4��	�'�����٫.��l�E�XK,�i		�'�������^+Z�x��� C����'��6/�0H��GC�4vI��8�'��5���R�m�N8���aid��'����չ^~5�,��Rߌ!�'HV�XBR���9QVy��'�^��V�T�s��3e�E0]�(u��'r4y	!�x�r(�*e�v�
�'s��A�o��G�Z�{W-_�'2���	�'J��F�Y�d�@}��ѱt8�4�	�'S�r�Bq3`ͪ�gAh���@�'+��
q)�_pe�N�$a����' R�ygc��J��%��,J �}��'l��SEI!�@��0�X�:��\{�'l�y� I(:�)�G��9�ڬ��'������=0�p`���,@��'�Y��e^+#! p�S�T5�����'�F�$�.����U�E�)��u��'���(�͓3i��)@Dߋ �FI2�'䬂Pk�KA���[�����'�����D��7&BU����'�Xm7��Nxz��G��*~2T��'F����Iܤ
���7�EzJ���'UP�b�F҈R���(t��z�d���'�d��Ǎ�>v��0bD�>wY���
�'���C�s$$��2ɉ�y�Έ�'ֈ�SbԶ!���zb��DZ<��'��0��Љ9G�x,<JT���'upc�%\�Y�^"Sm�Q �
�'��y+ߦI�Hu�r�øs
 ��'���xc��K}��ّ�Öj��Q�
�'˰����!�np`4/X5~U��'��Ź`L��/2�5��7Vhĳ�'Ϭe�f��}�6 �����|x��'���xB�\�a�Q�ËX�"ف�'͖4�� K�D �B�፲~�R�'݂�P�f"C>�+F�J'�<J�'�9����1C�.0���ӽA^H��'�lH&%�Q��K1�W/���'��I�(
i���g�Vv6��'��5ʃQ�!G!֪NK��S�'8e�%ND�L�S�AɰD�@��
�'N`��ȭ]�����g��q��'&�ىQ*Z,S �ჁQ�7NrQ��'�`�	�6 �1�C�I�>H�D��'�6�I0(jn$�� �� �����'��!�u�Z$@��b�%	�	�$
�'�r�'H��8He5LB�y��'�άҗ��^D�kT��K
�ن�ls���R�Y)^;����m�/�i�ȓl��u�%��}1�x�Fn�%%�(����iAe�Y�L ��LΫ>��ȓt��c�C�/n(��)F�0ϊ��ȓU���L�\.�e !#�B׎8�ȓk��u˓��w�����ؘG�A��D���[���;��(dS`���ȓs֤�w�	0#�d�EO�f� �ȓ>��9CKȽst�$cW���9��]���t'N%M? �K��҈(�n���S�? ����(�1W�>�y�O��
!�iZ�"O����#�*V�^t���x��#�"O����A��@t[�,ʝA�Z��"OxIr�F'~*��:ˀ jA0"O<�� 	ͩcv�3A��"�<�Rr"O�E�fJ[�o�jAT���fή�S�"O4a������9$Ҋz� հ&"O��qΚC��X��Jt�
y�"O`a��_)3��!+"P"O�\���O?V!��DϜ3*���"O�p��	˨��3-��`�.��"O��jdo�4�e;׬���� C"O�I�M#b���Q�5�ॹs"O�����	H�� ��*$o���G"O�5
wa�

<y�\�����"O��:���8!D��Z%�h1��"O�@�W]Mb\9z���A����"O��{䥎����kdH����"O	�A"�2J�VXK0G��|i2�"�"OFI����ÄD�����e�"O���%�΢P��Y�E����a"O&ŸEO-?etUB��Z$8&�e�"O�����$l��|�B��	L�6"O݊�园{h�su �a���*4"O�D���LK�*Щ��	���I{�"O8	I2�
_(A�cD��x�Y�7"Or�R��"qL��Bc�9If<��"O~��b�>��l3���8A+�xjS"O�ᢖ-H9i�^�ñ��2p ,�34"O��jAU�9��� ���q�"OvkY%r=  ���S�>Q C"O� zr����iC�>gO�x�w"O���L@�u��Hyf��8�@h�"Ob=ɤm�)\�8����P#n�(�P�"O$�:P�]"5x��A�ꗤE�21G"O>-���r� Ҋ��\9"O�C���gZ<�� �<4k�"O�L����.X�gԌ4p!��"O@���Q�9A�k2�Sv"O���ȎG�jIz�Ee}�XQ�"OJ��2C�@\���Ƥ({��"O{��$,�f�M״N�0p5"Oplc�'Cw�tY���Jp���Q"O����L�=�F�+д@��̓F"OL(i�.��Z�Ec�Dӽ��]��"O@��fVkz����ď�E�0� D"OIX�a�[ߺ)���/�@�"O!@�T�0V�(4��q���w"O�"��f�j9����Yt��"O.��2Řg^ư����&4��"O����f��M:$˷��$[8,�Q"Oj����E���8�VA��m����p"Of]��6顐��7���)7"Oи8r�ݟYDT�h���O�X!��"O>��S�d�(իsm׉
[�D�%"O�Y��j�?�&���+pY>m��"O���C�,Od���R%��2"O�H�֏ͲgI:Ÿ�ؗ]�Jx��"O���0�=n�v�Z1႖(�Y�"O��s ��7<z���/A+��x"O�M` ���q_�4��/�3"9:��"O�H�K�/h���H��M�u&4��$"O"�HP.��x4�"�C|�pZ�"ڛ$�b��O�	"���%e'<O�0P��6p��I� �ҽ	a�U�%"O� ~��B��q��H�*D�7Z($��"O��J@"*Ta��h�k���2$"O���@�2��I��Y��5�b"O���C��x��ZHI#r��	�"O���2JH�y��a�L���KG"O����#ٱNؘC��=`�x��"O��k>j��H{���]jt|x�"O���HΪP��Y3���7b���"O�����, �n�ʁ�F�oB�Ĉ"O�r�+��^�n��
ݶ="f�� "O�h����(�
Ae�C�Y̌�#"O��;t�#�^�9SM��Q�ze�P"O� ����k�Lr��S�s7@t��"O8uY`�ʽ i��!@���i(,�ʣ"O�p���E�1ب�����!��{d"O�a
��N�4����
��`����"O��R�E%?�X
T�@&�(Z$"O���iT)1���fi� ] |,��"O�d�6k�Ґ��h�#���"O��x�D�m`���I�]`I��"O�ThQE�!6�i����.`��i�"O�����*&�sR@W�8].��u"Om+��ݞm�<	��Ǚ0Tx>���"O%`u��!q�{p�QV�Ri�r"O(x�0*���i���O�2�0�"O�ɇa75�@!�c��̐��"O�lx�.�"a� �lg�5�"O��%4il��R#I&_�5C#"O�0�7�[���`��7G>�L�%"O���� *�+]	XR];g"O��1p�0Bu�U�i��k�"O�y+bEK��ip�NN�m��"O��P���_���6Cɉ*в�"O���q�� �8�ա�h���"O��Cށ �\P��O,~��2�"O�}YFo����0�0�HQ�"O~1��4h ������,���i�<i�+V�da"t��B*� ��Vd�<Q��� ��Y����t���H�<Ag�T=o���K�+�&�C��G�<!���,?�ʢ�ީ|�$)�J�_�<aĊ�1���r�)F+:��b�P[�<a�f͢h*�Y�
U�^�����S�<	b�I6u~ �+§%�F���d�S�<fG�*H4(����<>ҝ��G�m�<I�j̐ow8���L�)��XE�^�<���;:ީ3�(��
�J����S�<1D�N7N��V,�2"b ��]s�<1B+]8Pp�/�ub��i��w�<�bC��AK��!���j�E���Sz�<�r�SN��8��ɝ�htd��A�y�<��	*Ks�Y���� 
���\K�<�QM�\/.���&n� �_J�<�r�D�}XbM�3��WX�ԑ��AP�<�6d�(\+dp	������ N�`�<��)�.w��0A����Q�M��< ��bŲ��W0m��I�cw�<��d�8���Cg�&@
]��̇p�<��$�;�L�� !� x�F�U�<���7f�6����� 9����f�YS�<iE	��"`�ӳ,����
�H�<�phG�W�VB� �1N��s�@�B�<o�=[ݸO=Ԙ�b���Y�<#�FE|����M�<2Utu@��Y�<� B���"J-r��fGQ/7�qR"O� !�J<��� ����[�j8""O �%��+���e�W"x��`�T"O�����	z�Tۦ��U�����"O4��dH�/c�4��"Ӹ1�BH�5"O��C�'Ů\��cb�\]Ψ�t"O���q���i/F�K��Ϻ~aN�X�"O6��u+�5Qz�8�a��HAR��"OD%pa�0t����b��ZD�I�"O�pb��;OV��"H�"֬�"O<APu��&dQ�}^��A"OT:ŎIv�I4�Q8iَ���"O�@X��ޔ�^����A��=��"O(ٚ�.J��^E��G�6|V�!V"O�����:?S.����^D��D1�"O$mS�jK �y�H2yR�("O�Da�E�s�N!��� G���T"O���7&�tAjg�6M�j"�"OV�;&f��,�z�C��VP �"O��#S����'F a�ա6"O�=3g��W���ƒ�FJʍc�"O�5�3�"+����0�R9�*�Pb"O@��'��8.B����*L�I�"O ���(�&
Б�.�U��]`�"O&i!��l�r5�k8m=FѻU"O^P��֕`�Phw*�"ԂAC"O<�Ygl�'J"� �P�=7�))�"O��G-�Z_���D�W7G!,�y'"OVI5�ܷS�t!��H#h����"O�A(��\?�
����(�tZ"O�X�f�!vk.�##�� Mx���"OD�Th�YQ ���(�9?~�}��"O&@��ȇW�M�b�� �j� b"O`;艵-u dђ�Cf��@�"O�x���.x��`�LG���E�""O�p�G�J�!�%@ᖚĆ٩6"O&� ��)-_!��@��-�҅�B�'ѨM "I��>�3҃�)'�� #�盳�jC�	�:�= ��'�p$��N�H#>�UKדG�x=����.N�Y�#%䕥/�8���+�y"bA6=�Y���X�y�tl��Mˢ�p+ґQÀ���s�$٨%G�n����9&��ku"Op���D��<��F1x���p�R� �3��\������c8��	"b	3LEFE��V=(�x	w�#�O�@C��[�+���̖+5@��׬�z
�y I$^l�P�	4�O��a�$<�	��g�q�Y�p��+�n��ǄY\�6	D	�@��<��M�R��������7&C�	�Y�n9�\�E�tdS&��7�$ ��䆓Q��tY�GW%r�|A�N2�g?�V�щJL<�!�섔)ڨ���U�<1�k�aF��sCN�Gi����%NC>6pb�Iw���{�N��	���3�"0�ea�kAd�Dd� \�l��,b���[�-�`�ɖL�C,*��]�b5�剈IT=3���B��l���7h�����A�_�ty�4('�	^$ȵ�ƣN\������/DI~����p(0�0 ��L�'��E�Q	7"O\4�  ɼe���#d�<{hnqQ�U�L���iUn}�6ͱ��1�>��3���D�F�(��IH�	�SJ4m�ȓO�ҙ��F.g��룭�{�&��P&��oh`�p����~Z�`�aRݺK��6=�R���R��"%� -�3Xa{R�J�D����d,�l`dg�R����_؀I�A��V�j�'8�p���*]��e�&�F�J�}��Y�Q4R���ENh��u
�)c��'<T�y fZ >i��?_��8��4D�����K�W	nj�Aނ$�P���>=߸%{��ƀv��,J&Şq뀣}��Y�T�R��Ⱦk�Q�׌�&`�Y�ȓg���� �jP�x��}xC �~hG�
��ɓ��Q�� ,�'������dB"J�ܕ���'�X2�G�4)��,	�-%�|R����LH����r����CM"le00h�)o��C�>�{��%�bI@&C&�$?��g�'yJ���ҁ$��("�$1D��c7�Ϝj���S��3m���5Ű�T��HT�R��h�L<E��/Gh�'%���F8Se�J�y�JK�$I��8�O
�}�l��gNV���4\{��Raǌ��p<E�@�q#գB��
��f��q��1��"�b��E�B?z�H�3�c��{G�XOh<�#��;VD&��p
��7���y�'�ް 6�Ӳsɘ�ȕlu����#�C�I�����S�_��9ծ�=_��C�I'6Ԓ��d�F�D����u#�C䉽wJ�]�G޸��&n�*t<B�	�J驢�C�yN�eh�c�B�ɠm�i2�ϗ�Y�*�3��$C�I*ZV�� "۪�.�`�N�a{`B�.V����Y�A aK���2�RB�I�=�@��܆/k��a�LV(RB��v�a�dǋSwjЪ�	��B�I�E~��ZkDa���q��R� (�B䉧���[0���3�̸�D�^$P�|C�I"B1�m8��0��-��.��~C|C�	6��(%��tP�F��7m�B�Ɋ�fĂ�/�:������q�`B�ɕ��S/�_�P��良(|C䉼<�d��#�5$���aċ�>�hC�	� �J��É�=(���	�.�{��C�
1��B�$L�\�@�ևOA�B���J�zQ��j�\��f�.��B���N�{��.	Ud�RB��ZC�)_D9S H�?Y2�
�-ϼQr�C�ɒ��,Cg!�#'5�w�Y
-!�B�'x�x�cŊk���!�R!+�NB�ɂ?�D�X�`Kz�`Ժ��_aC�I�e\�2*�3ZW4�q����0��C�	8ɼ����(:L�y�ē�0��C�I$dTe��a�C~q��V9idB�I5[���c�7��(�}A�C�I(0�@u���%)������O�6��C�I�)ʶ�)��ݙA�]�w���7`�C䉚f�tY�B%�'lے��č�70�B�24_����,��/�TS��A5W�B�I�=gr��� �!j�<��Όz�B䉖E�h��ȁ/�JPD��rC�I���y{��A�KW�ׁ	�>C�4S��@k����Q�T���K{
C䉝mX��C��>!\�c���h�C�	zS�L�d�K$�(y5o��
D8C�I�[�����+N*��X� ��+�C�I(x`�L[!��
L�y�iJ���C�I�#���٦J� �lU!'"�-M�fB��O�L�G�%2V���'�'b�DB��%@r�(r� ��M2Q��
-�B�I�tܤ����6H�3	
�.M@B�I6 BH��M��YڑS��֏'TC�ɁO�lm�֭Sfj�I�%��e��B��
w��D�`�:|1��B�WR�B��9x��`$�\��& ��"JdC�ɍ9�إ3�*Cp ��D#G[�(C��v�nYy�EIZ�� ��o�,B�	12�@�ƪ�yv����(�bP�C�I�l����9���ڔҼG��C�I?=i�p��j/�L+D��*'��C�)� ��1�ݫ6g�%� ��̖��"O���VMB�A�H�{F�_=Z�*��"O>a��Ā[�3��áS��Z�X<��w��!C9�;�M3<Oz(�q��0�(�biF�<p�"O8ĺ��G�V�P���,�,DȢ"O�͒��D5h�بKRe�xi�R"O�L�R��[�P2��S	�y��
�ju�6�*G;�xB���y2��Iᖕ:�"9�#��yre�<;D����z��]�!-@9�y�N�u����b��m�!␱�yrG�*7ӎ8P�E��a�(8�S2�y!�2��bV%+ �H��,�yBg
�`���Y�(T*�>��/���y���Q��A�I�#*f�ff��yMC;t���0��D���YH���y�-E�
ՠ�]�u�l�%��yB,(ܮpꄎ��r�N]
���y�%�w�DeR��s*�����y��!u	�Ճ�kjPYF�@�y���'���r�ݬ}�~!	��y�l@�=���9@��v��}b����yb���\5�u���:���8Rb��y"���X<�# Ժ5Ꞁ���yR���#,�xp
Ԃ�Y{p=�y���.^*0�*T"R8�v'V��y��ز�d���Á�'���*墄��y�ŁEڌ��C��0�}(�+���y�	X�~lr�m	��9�qՆЖ�y��^~Tv4��+@@o�,iŬ4�y"��Z�Ř���$���t�.�y⩇� �����g+���D&�	�y"GҬ=��E��X;K��Y1��)�yB�8t���ڃz�H�� ձ�y�.��7:N��f��X~�j�OI��y�e�(rD�}[@bG((Ԏ5hBl��yң�p�c&O�
Twj�uCL��yB#.5Q�Q�޴S��D%^9�y��K�e�P�eA��".8dᔦ���y2�XA�����	@P�ħ���y��Z�}�������r
� �yrk4s_F���(��n�t��G��y�g�4��1U���*��t,V��y®]�D;�C� 0�Y���۝�yҤ_�m���@F!s��Hs�Y��y�N+6j|qT�����*c�À�yBe�v=���0��a$��)b���y�VP���ؑ��3]�t Ґ�W
�yeK(;L�Y��KN�,<���ޕ�yB��N���EJ�ur`)`OT��ybi@��x�����hF\��WGA(�yB��/����Ma7fE��yBiSd��9��	�>FD�f
��y�j�Јk�Ă�/l.�I�c�(�y�瀇 nl��FF�.��x�0��>�yr���{ݚ�ӆ
�rADa!�ʂ��y��C�f��4��lS�!���
GCP��y���&'��T�a��9���&AA/�y����Z@	��D@O���$%Y��y� t|T1A�錴4��pc`F��y�������B�,1�xZf̀��y�O	�M�(˃FV!&�`�����y�k&;VFlX�� +$x(�C��y�(G�lp��I�$7���reZ��y
� �HDㅵD)@��gEKya����"O,)�JP�t�*Y���HM6 �J�"Oҵ �ŀ�yI����&�j<t��"O�y�P$#z��8cHΊ�e~�<i�kܗ6	Hhz�˗�~�\� խ�u�<�eo� I�(�Tٹ~D.���n�<�F��$]�Es�\�A�Q�v�<�!�*w` ��ɲT�n(aѣu�<��F0?y�x���)&X  ��i�<	uh�G�Ԥ*���.<J��rm�f�<qP�ӸS�* f��->���0��{�<�.�?o�����;o���P�a�<�̏%up�<qS�Z1��a!�^_�<�S��J�(+%#N�Ȝ1��!^�<y�Dʤ��U��?e%(T��N�E�<YP��9&��s��##�[F�<BeH�[<N̛� �&ـ��1��m�<�r��~ �(��+�!`M0Lh��_u�<y5HI�hz<�f��N�tE�3EMp�<Ѣ��$|M�eB0k
4�$�COAB�<QR^?j��pJ@�Er��i[sO{�<i��Si:��c�B
?��|���u�<	7b�8|�p�FR-fC����gIm�<!c�I�U�Fȸ�*�+�t�8ALO�<��	4^|E�m�3�Ȕ�E�<� Ȇ�l^�[�Gt_^�`�-�k�<IG�"<^ܸ�C�^��Y�N�N�<B̵5nL�[T���ZAf�k�� G�<�w���#�b��A`�6�����'�@�<�c]-^D$0�N�BX�A� /�d�<��̂l72�ie@C�(¦(-Yq�B�	��Hs��ٴw�P��/�B�	b(40G�ƞA)d(K �:8)�C�I�W�
��C:�A���u�%D��	0�!Q:, ��l !�A�-D�
rG���,�����,�&��1#0D��	���v��SR�87O�84d/D��0v.��9r� p��.���c-D� �&9b�E�&D��]b $,D������%{!D ���[�8I�%�$D���w�>X1j��!#S@Q�m$D��"p`^���(;l��4�g$D�D{0\	�y�'�6-2�"&I#D�4���W&f��3�dy[���ed D�@k���*`�}Zv&Գ2����`!D��c�i�Q�'�"vLƐr�K>D��A��1�Fa�ЉaĦh$�:D�L���L"
lW�i�����7D�����D`9�k��
Uk�`J�7D���P�jt���j���ڇ*D�������;�лR�	 {$j�� �#D����Q�m8����Y=��b�%D�sRM>sT��q��$S��X�ӭ!D�xpb.��	��x1b7,�D)AP>D�X0f��#���"�E<)8���a"D��K#�Z�U.Z�hF�7.��̀��,D�0�a�)P&d���B� �ĵj��*D��PG�EB�`ٰ��$U��-�V�=D��Ӕ-A�x��"�����p�??����ӠD�09BV��"kȱ���"C,$C䉮:����p(E
b��P��(:x��C�	�*��r��Sά�a��T�
�fB�7v�����x@�(��	�TB�I�5�,1^�t��D�J��U�2B�)� �X�j�[���%�%]��Q"O�"�H�<E����ߠ3�*E9�"O��z���}W�`:G�3_�V���"O���.؏F]8}�1c��	�`y�"OZ�X�HW=b(��5��i��"O�)��
�x�p ���06�tS�"O:���+��0j ��+h*b�c "OƔ��昒PqDac�.?)V�0�"O�+ ��	bir(p$�
/|��س"O>�9v�L;&f|��2���h3�"O"��� �ce��顭�H1�� 7"O� gf�(�\	���> �b"O>aA��Ez�X��(eM� "O��2�B$))�H����;N�ʵ�"O��B2-ӴM�F��MY,�}3�"O���I�S�䘀CƏ ��H#"O�M�TgL�_�BqrWO5w�v-q�"O�M�5F�)b<	aHK�N�.��"O��� >9�lh3��w����"OZ�a!O$-�hH'�1#�� �r"Or�c6��0�l%xU��h���"O�Uhe��+$2�!dh��Êq��"O�����2I"p���L&gH�yE"O��2��@:D�|=[`W�Z>6�k�"O8�+�*W �����%,N�i�"OB̊��j��J4
_:pl� ��"Oh�� �N/Z�~�2�ȼp;����"O$-� ���^�rň]."�� ""O��Ps͓�w]�i�`�S�"�(Xs"O���"nQ���D�(_�2��c"O|2E�D3zd���4"ɸUkG"O,��b&�6[�%[��WAP* ��"OX1���E���Մ�4�P�G"O���a-$�n���՟xe��"O�M���..��m���R�E�`���"O,(�BE�p@ ���ךP5l��"O|e� A������ ǜ4&*�{t"O�13�E� @������"OL��7��70. �ɡ�0S�A"O"��֒x(؀���H���6"O�h��ضnvL)Bf�2�g"O�H��bL2j�a#���$b��"O����S!*���㖗9p$�!2"OB9K6�I�4_4m���͗O
�i3�"OlmcQ��!ZB���Q�9�8X��"O(����NV�5�O�tb,`0"O���JV#s6��P=�t�F"O��c�����Iq�,LM3P��s"O�1�j�=��aa�KLG�R�"O��S��*?"|i��j6~Q3%"Oڀ�q�=U�L��E����"O�pР� >��4�)�f��"O�@z���=%�8��G�)c`�9r"OР�׬�$|��q�(E�����"OƜ�a�,C�2Ykd��$J�"OC�ê{Ԟ$��5 Ξ(��"O���_>N@������ +�pq"ONi3	�#Q��� e�%�,��"O�A��r(J�gD0��e��"O�����ڢ!�����G�f�N��%"O8�jw�:&,�C�;9��4;a"OJ�@�
�>NE��2B;t" p"O�E��bȇP~�= \(+�([f"O�����S[-��;��" �1e"O� @�adjC Fr�]�h�(Ȳ�g"O��bj�t�V����ȔRa����"O ]*ч�9
���	q�&e2��s"O��ے(����˴�)har�s"O@M����Z�z��t_�{2��e"O����F�2x�p����0f��.�yBEZ([��$;6�Af������y�fӄM�aX#Ŏ2��b�>�y£��ZE��0-�,�Qc�=�y�ͽ �Y W#���EmB�yRIW"��IKpHY=f��Hce���y⥓<z�����)�v��ŀ�H��y���O�>��5bD*_�`���b̚�y�EY#2�b�+�V��a�F�yB��:h1� �%��Z:< ��+�y���*aj�OGb��b�.���y�	��9.� Foٸk���#O���yr�D3+�D�#�:k/��&�0�y��L�nM�mQ�c�7Zd� �B��y2��+-�^L��D9
[�!p�]��yrG�B}�f!�����7 �y�� Y>�Y��v��R�a���y$y6Ċ�'N?;qZ������yb�]sx g`&��)i���y��X�FfH���ab�83�B,�y�CB&1�܀n��A���A"���y⍟�$$�t���� J6h��9�y򫐍l��K�NUoI�M��[�y��55V�p҇_g�L��B�6�y���_�x\��_�>E�A��y�b�VI.�b'�9$}�T�@MR��y�'�qL] ��)�4T i��y��pEn�Z����Z����N/�y�ԇ>�����I��J�;��!�y�Y�BN����%��=�����yrh˄P����U�.O�<hV���y˅J1��*��-Lbzxc �F �y�.}�L媄�?B�6�z���y�-� /Ո�*U�):\���aOO��y�F���MBԅ�,cl�a���y���"�x�D�μyff��0K*�y��O��"ū�C�);���6�yrbжaR�c@͞#�����X*�y""ۚhFmz4�Q�<`��^��y�tA��
ab�PQ��@Ӷ�y�o�!��4c�Ȗ@��)рM+�y��
{!68��),1�VA`NJ��y���<���K�M�.@(!����yr�S�=�EC�N�5;x�q��ߊ�y�$O�\�tp 2��33�x��2/�,�yb�_�;.�����f��C�̙�yb�^y����#�9ք�
daR��y.J$n������R���D,�y���<"�`N��ypT���Ґ�y¨�7������vF~@�"��y���)��{aC��strEARlť�y�܉3'41"���{�t�*�!�,�y�Ɛ�-�$���EՉ~��q�·�y@I2���k@��8=Z��U=�y��&&�(0P")�'Q����7� �y�7ƪQ�#��8��*w��yb΀56g@��f,��<��/���y"�
�C�q��%�&�j%L���y�% �5�BD��@�!�����G�y
� `�hT�E	��t�٧@l�0�0"Ox�L�s�2�˶F�
R���"O�Q��ƺ-X�8(c�I��.�j"O���
'NYvl�gd�� �~��P"OXer�E��lZ�1T3S�t]��"O�1
�OP5zT\(�"X�Lj��(b"O�h�\
*�0�i�Y�k�<,�7"OxT��j
�(�10�c�Y��	�"O�US� ���N4�"��& yW"O��HFVsnJ�Z���U��hӇ"O�2�iSRӴ�:����*�"O���"9��X6�>шL��"O�]�'��Dz5P���1lȾ)�@"O�,�Tʖ  �Q���R��l�"O�ԡ�J�y�q�&��bD޸hC"O�aV)�Q�d�byC�d�d"Orи�HcJ�م�<K��4"O�	 �ܕs{ވn��M��$@vL3D��R�A�(q��2����Q]XY��3D�Ȩ�NՅ,���:���@�`�)�6D�X󢈖'4�����!Ǥx:Ra��"D��$*��Ǥ���D?(
�� ��3D���A��~)�2� ��\��4D���eNǂ�Xƪ�,B�|)�0�4D�� !��QP,��Q�_��Fm+2b2D�$�L��Q���1�ʒT�����2D�X��:6�N�kP)���v1D�X��L�&K�L	��<1b©
�H-D�|;���z(2����)F�r���i.D�l�$�H&��(�B!��m{:e 1�0D���^/T��)Y�	�g�f�Kf@/D�`i1�Bn5໔d��^7T�K&+D�@����$�(��EiT�viHըQ�)D�d��%S�@��*�@�7~���.+D���@�/j��,�a��6c��Y2�,)D���%dS�II��%��''��ba�9D�؃2g�
S>��K��N�\4��L;D����3�"��N�=Pj�+��5D�� �
K���2b�H�o�4���/D��C!s���!�[�RD.m�'o-D�p�#� R}�y	҅T�E�2M�G7D���2'�\�nA�����Uk$%�5D�p�BB�|�Hi�R#V�%w�!@g�1D��9Ӥ^�;�J�p��R����;�	#D� �Մ(�\�������j�	Ũ3D��
 b PŎ=�g� g�hɊ��1D�`���Ș$�s⟚���
b�*��䈟��JЁU��HbS�؟*7
��1"On��s�A�[�X��M�
 O>(�"Ofy� ���%����l�48�\�b"O(�����0� ��?=V��"O��Q&K�4h�ci�#��r"Oxa��
j��0����/��Q"O i�$���Mz�t�`т"ODՀl}L�i0DCS$�Љ�"O�lJ�-��kw������jjp�C�"O^Bug<�}J���H~�A�'�г`��b����(�J�!�'\�;f'$&��H b�U�~Ux
�'��pd���q�ds�� Y���
�'�f�9���V\���V\(����'�|���Z�W�d�9��=��t:�'-~�{�M�7����`��9��	�'C�٧k �8�hHSnA"������ >%���kЈ� ��&QF��C"Oy"WᗥH�(�I���ODl�"OP�(�m����'S3��ZW"Op�� N�+^5�m�zy&%�"O��T��LB����b�xa��"O�8��$����`�ukM  �±ɦ"O�����J�(J�S����G���Kg"O�����Z����)W/L��F"O�ceNK�F��Uy�Ĝ4�xA�"O.�S��H01�H�;p��0�����"O��r!���\�ǏV>b�V=�3"O�њ�G?z"@��ߞP;b\�w"O0Q#��7K���q�P,�\�R"Oz9���$jVLI�%@ N��pq�"O�����X3�]9f��3����"O
d+"�A)��t+���M�p��"O�'c�3Gȳ ��39�n�J "O�����'_��WaH(F� ;�"O�܈�䅫�Ĝ�Ŝ%1�*�:�"O���i�R��%�,x�@�`�"O*X�7�5!q����R�4��<""OPIkF�`�����J�*arT�"O�)�cK [5�A*��8P`R��"O$	���B`�~H�3I�.j�51a"O��sꎉ2��=�egƕ" ��5"O���cl�%1sԘ#D�k�9�#D���aר-ִS�A8_���m!D�Ԉf��Q�R�9���.T��B�3D���b���v����΢"Tn��3�$D��+�H����3O�qu@u��6D�XZ�$� A�}9�b=i�Դ"5j3D�$��퓊�j��DM�]�Ę��@1D����$F�S9�H�o�\Ia�#D�D)bi�>�t�Q�Xkڸ��#D�\Cu��9��L
D��u�d�� 4D��Pr�.Kl��'�m�h�"g�?D�8����,��`��C1�"Q�� >D�����ʥ�xѳ ��`�60���9D���H
8�Z-[F'��mV4k
6D��xv!Ή@u�R ��K(2�kօ7D���R��@��T�$,�h#����3D���cHF�Y"��ğ�*�|�`��$D�(�(�S'ک�*қl�z9@��.D��6DD�t���F�.�${7D����۟]��L�#;e<L���5D�h97*���|3����6*��VH�d�<0TQ�f�آǒ�MMҨZ�H�{�<��χ� �8�1��6������P�<Q�!�%m��� MI Fu�- 6ɀa�<�b�)^��:v�\>j 2(�1)�H�<���ٹ6V��1�i6u�A�@)LY�<��)�#�v�����!j�]��%AO�<��� @�ԓ�͔<��{A+Kp�<�Sb� �"-�K�~��l�<��H:y:�Y+�3_�l���l�<ѳ��b ZQ �������Юq�<�׆��:bR Q4�͠lR��n�<���� }@���H#^ �U�Ѕs�<�ѭ�~M�1C��d:D�<5��n���*eͤ0�~ 3�K�B�<�� ��h+�IS�Ō IH]�.�}�<�G5 �,Т�ɂu,aS1a��<A\5 �E�R>q����/r�<ad>5rIP#�ϐ�G��qʣ"O� f8RL�� ��/B�v����"O�}��l]�Q�Xa����s�AV"O��r�#j��)��cM* �
�9�"O2u�0Ȅ;��B�BH	i5"O���cE�/*� Z���ne�"OD��T�ϗ)�6��� \�/��X��"O8a��Q�qT�t��H}|T�c�"O�E�n�z�*�DO/=G�B�"O\]�D�N�#r�����9\�1a"Ob�s�хt��iPƃ�/��۳"O�г�(��UF�X�Ϟ]�MJ�j�Ot�Ce퓉�M˫O?�	!�	HVʬjB�UF�6���EԘR���k�'D>f��R���bB�>����d�w�S��d�� �U.(Mʣ�i�dd��Џ�t��J�IYv��3�D� �@]��*��s�A+��N�ȑW�'~�]�ig�����'d�u�2��-��)�`��N��5Pՠ��HT;c�����쟘�퉖�J�C$���V��s�\_f�<ᕹi7�1��ɺvk^�c�rAH!TY�ģ^a�2�'m@Z���L2�'���'+DםΟ,o�+͚H[9��i�u� %�V�$� �v<��Zi>�Q���}��	�o�Hi�v�|ri
�a4^�k%' P��S�G�|3E#K4QpDba%٘�s��h1���<#�Q��k��$��.��@�F�J���!�(\��?��o��?��i ,����� �
9.��
+tNX����8e2z<��F�0��%gSL̼�N�9���a��u�|�o�S���?���sy2�U�B� �p2J�r��u�BS��v��H�'��y�'��=����^]�!��Аs��`��F�]~<���@�T�E~� �hR`�P/3 PĚ��Mc$$j`�<�>�#�k��y��tn~�ڤFS�NOz�ڤ�'��p)���]���m��_oa�����>6��O�� ����DB@Ϗ�!���e�H]��E~�<	uY�x�Xt0d� �3�|}���w?���i�66͵<�4튠7���'�"R?]�� Ť'.� �!y���� �%U6�M
��?��� aX�s&e�=k� ��=Y�Fx��}�%�2�<��K;(�d9��դwQ�H�F�"c`���l�"��������O6p8�^�j�CD��ϒ&���&\Z�cFiP�@�����
K}�j��?Iиi<����67M�8%"4�� [%ZMa`l�\w���	J�S��?A$Ȯw� ���<�"��΋W8�,��4�?ڴ7C&L��G�Ag ��}j8���~����i-R�'z�� 78��	ן�lZ�� �C�R]��ߌ�X4p�+���̌�#�U4�(MpC��,�ФC�l����'�zYc�����.�""(Q�s�0�P�Q�4ZmZC̾1U���gY^i���!17�P�Aʭ��Ƽ �U�V�4J�1εI�p�r��i�h�z��?	ոi�b�~:L|n�[���s���2s Dt2�C���I�G{"���K��×�Bjyz�d�@�Q� ��4��f�'7M�O� �g�|ݡ�W�H7U��L!�ݼ\  �T���?��КIR�� �?���?�	T�N�O�6�N���NC~��U�V ������%61>��� �m���b�L�?���C�|c��OJ��a�U]5PpӀ�F�ZZ�R��[զecHo*큒k �T�v�t\������fmZhS�' *ܨ�ϗ��`�:׍^�9�*�I��OT���O8nZ�-���<q������z�$$`�
��1�����%ò����iA`u!�	T-a�4RT�EYf��m�Ӧ99ݴ�䓹�	)�	�nOҖ  �   X   Ĵ���	��Z��wIJ(ʜ�cd�<��k٥���qe�H�4��6_2<<�3�ʄmn�.(��f̅3V��(�87�ݦ�+�4>��$<��uyB ��<�Ty���Ѥ������G�9S0��4|�0�=���%�1D7�Q\�:I�Ň��<�c�p��	��v]XT�ʂ��I>�.P�łN�:(���&a��֢s�LYʵ���^!�c�J��-��(Pl}2.�#<$Tz1>����%�ε:@cA�	�j�F�.Ar$� �w��I�yr�C�0A@喧�$�Z�"�PsW�I�}��7|
H���"8<Sþ�P�`eaea�
�˓9� ��nQ�}��Tkp��������9���y�d#<Q!)W*��)E0a���AO �d@YP�I3(���h�Z��Y7j<C���Ci8,|�)h�E&}r{�'.��=1UI�jR�IJ�!v�V�"2��ʦ݊�ቮ[N�dхĉ� �����I4]q��P��8
$b�TS�I�j��I�5�A� ��܅0�cL�*��� |�#<�`0�	�O�TaAFS���bK�#���t�Ɉ`�X��'�bh	w�N�[�:}X�G��>(ybHJW�'��&�t1�f՗,�<�1�� <dXm�������	(S'�'�����h��OB l,����b���xy��Z@?!�l]?��	��� \w��H�A�
h��'i w�)����;�O���H��b#��KF���Q�6�tD͢>�� �4�"<���5D�ThF�H�_2���A�<)@�� 2  ����C���q�.D�l�#�8d�l���R�{�LC�i,D�� N�{L�;@�°�Y�XAs"OT�j��R,������.�I٢"O�l�A�D-
5��2�NΒ"6��Y�"O��+�ƙ|�@=�t͋�
��?�yb�����x�,48� ̛����y�D�v��s���g�J�;��4�yB�Ƚ#8�a� L�`�ĕ���L!�$�"G"~D�ԩ��S4���«_�!��m�e;��S5��4�ӭܮd#!�deB�гP�ߋ	����U��6&�!��]��,=:�f��[�~]��mT�t!�dC=2݋�N�'�e"rbׇ|�!�����s�*07�d��Xu�!��_6:\��3Ҫ�7".�t	CDܐ5^!�DZaj�BVU#�4h�U�X�4m!�D�(>}.|[Ӡ��id�#�N?    �  *  �  �  ?"  �(  �*   Ĵ���	����Zv)Cll\�0R�P��
O�z��1Qv�i%��/��Qlр�yb��Z���Jc��?��J��ߪs������I�<7|�������ݚ�-͛J��j2@Q66�X
�ڠo��	�����N�9 J:��� �:OC��j3iZ�5���c��&h�St��� �����O.:���3�0S{����ځ8����$��A{�A�/� _�D�H�&�&3�@U�u�<�Iߟ��IڟT����$XM�@
i1��		sf-c��gy�AM�$����'
R�bt��^H���S$FlY�I7|��tŎ"d�$I"�擽���	�p���Հ���1!��K��Ξ��@	�\�M���'!��ٓ�'yB7me�,O������b�&�vY&�#1�ˆ@P��r�3D������H�֡Y�!�spAP�fl��!Dz2�H��V���bF� {��ɅcL	�b��)MdU��!�П���؟��	�u��'i"0�阁�'Hre�����'��l�.&{_r���$�O�����OD`���xl �,��dw�Kax�x;w(�O�����D��Re@\q�j\��QR�<�c�,�[r�5��%kg�x�<a7I�,&�6����"9F��f��J}B�{Ӳ�O��c ��'L	0(�a@աNvH�a5�i�j�Z���-q���F/v�:�r
�'܀@�s�іt���P����'�� ����2'�
0K H$����
�'3�tۇcM�=ņ�Jc-�!D9$�
�'��c��ƚEۘ���� p��'X<�g�+vc|�"�NNt�����'5n#�GMb�zh�c;-v���'�$�[�Ki�� `���a댼��'��Qu�	�6��	K�⁑;���'��y���0��£LD��)�	�'H���v.ɿl�XH�ɕ��P��	�'�L����I�c3���ՉA�1R�]B	�'��A11�%���A�#�h�'��$�ǚI��kL�X�Td��'��PA�	�p�a��Tj.�3�'WX`	eM3sV��� �9OQ��	�'����A�$C��$	c \�@\���'kn�
�ޠ0�ȉ��㝞���y�Ϗ�d`�W��[k.�����y�b�;!��`�&��i)��s 	*�y©H���ƯP��eQ�fZ��yrm�qNĜ1u���9�]0X��y�m��^�rP+���6"<�b���y��M�3n��7/Bz1t]��J��y2���xy�w�5l�^����O��y"m�%pQ2=둡�r�գ�f��yr�<	D�[�J�9e���5g\��y�O�� ��!���@
�	x�L��y��X�����N^�
�����;�y�Ȝ�U�5�g!��s�&$!�˔�y�R>H���c��{J��)��yR�!gh�a�d��yCO��y��N�K�
�q�gKЀ����yҏ�B"�4Ip��F Jȗ$�y��C48`����� >?�-h!ŀ�y���l�Vm�voT,4dx�C&���y��ME
5@�bO<@pܙQ�
�8�y�� Ű�����M�|�r��=�yB.ʑ\�P�j%nߩ��Y�_�y��V9� (Q��Wy週�VM��y���5B�lj����t	�q%!��y�kӎBQ�"a�!Znv�;�b���y��A�^� ��`���)�%"c̙�y�/"צ!��[����O#�y���4"<�U2�#��PϺx��e�=�y�$�(̥1�&�8V
��D��y¨�,(m)�H� R��T�Z��yr�1�v�xp��$O���G���y
� �(��d�$�%1���2Z�&��"O�e��O�?$�1�X�&0��"O�L! �/+���c���9,>��ٵ"Oܹc�#_0�\`���?!$l��"O(%�ԋY]L�p8�㗍+�2�1�"O�h��wKD�{#��4�c"O$u�R�$�@��R<�ƕi�"O�d��͞2���I��tv���"OF���E�t(<I5��\a"4[�"Oh�YR�]!t�5f��^��Њ�"O�S�նuF�B����Vh�"O�)Cn�:L��9R���
��h�"O�d٢��.�����_��
�"O�h�5�}�&�M�c
����ݍ_+!��!F�&};�����hh�G�!�!��_�p��7�(���[O�!����l��X�v��(��$լx�!�䃀]�� �9?Sx��U%�-{�!�.,m�����G�iך�J��0�!�D�D�ް���
>�(�EĐH�!�DA+�2l��Ϛ�*����SY!��:dzE�DFEl^X�5�	&0!�d\��^�'�A�i�0�)B!�$�<yhD=;�՞n^f@��&��e!��[�
#b�wBX ;�E��D~!��оn� [R΃2F�Ɲ�p��{o!�$�!��a��9D�ire��Ux!�$׼u�T��f޷;��91��2q!�dįEn�hD�H�|��9�2f�*:�!��B~�͓�Aί�0EP��!��]�\�W�̲2}x(UJ�b�!�Ĉ w7ލ���Q��TY!!�$J0�= D��{,����Xq!��� Ak�jg��[F*�"�$�n!�$�:}��cm�*`�L��b�6Q!�$ľ#|����,��<���-�!�R�F'z�¢�@"-�TA��!�61�!��L<���c��	�*N�G��7!�dt*�i��ʂ�~��� �_)!���K�2�[5��@l��&��QF!���b�2	��c�?�T]@���F�!��3����79�:�Δ$�!�d�(*.�S��i�(��+I�F�!���TXh�#5�L�du�i�W�[�/�!�ږ	�f5ȑ̕?k��ȗ)�7'�!�$�2 X��̗ׄv/�����
!���(��:!�<4+��7��gq!�ϫ.��,@�C�<y|�Q�#H�/N!��ʝ7G�)a^pd��� $BK!�ėl��nBP4)dD�P�b�;t"O�tٖl̛zВyq$+�� o����"O�����v�P�	HS����Q"O<�V��u���鍉q��qʃ"O�Z�k�~5�w�#s�x�xs"O�9��Ss�]Ru�R�/ؤ�[#"ϱS��OD�}�o����	���2�:v"O3&N��TV��.q�E�."|u�v��Tֆ�0�%��a}�ݼ)�1r�Θ�E����4����<q�ƈ�'���0���yrPF��#Q��Cn�P���y�����ӏ��.�
�5).�R�'��1!R$R��\��D��˘(>#>�1��V�J���r5b���y�Q�dņ8�K�%F���u��&��HRd�.0���@�G�h��L>�w$�+g�茢�ɔ"�HSgO(<9���dC��
qS:�)rl�U < K2���PG0t�թ��=� �<2����d!��\�<�!��'� ��t-�w�v��	�E�I��N�]���0AN.��!\W��B䉕^l�r2�5I��p@�+�!
:z�*\�dG��t��փ݂Φ�|��C]��y�+C�'w��� �F�<��!2D�rG�D$V�4����.h�,&K
7JEb�Ah��i'?E�<ِ� �Dt١��
�4����u��Xٔ�!r���fWIVL���*2��%OH�z�v$�`�ԝ�p���	�-j�� Vc� +��J�`ˢ�?!f
H�}���!�"Ѣm^YZ�k�:bZ ��fX������a�1(tn���'=�d�g��_����% M�1�Tr(O~�懇�t�6�ZV�Q�w����'§.q��ر�w#&L��E_N�D��.�5j2�O6v�a���>q��y�&�K�f��ch6?��g�g�y�G�N�à"ɯ��<��XxnԄ�I-gN�Ѷ��1Gb�g"E��Ycv�-��q �� 1�R��`�U���C�-*4�J�;Nv^�{�8O�i�T�Y��p��"�3WE�芥��	C�N���O�0`��䀧�[\<!�D� 2&�F*>$� %#rA�?1�I�~rQ��	 WiR��(�X����D��I �d��"OP��v��)pQ��	Z�Z��ۅ	E;,�X���
e�#�g?�ǄH	Ȟ�)��O?v)h\�Q��{�<с�� L��@���4A�X)��Φ=D�Y�[(�ԑ"�+lO�8#M��u�L���E C���u�'r\��h��1:�	�v�S�{�XB0#��`��C�V_�P��	_�xH�3-�*Rvb�L	����]�X|��I�>k�T�Gd�L�B'��4 �!�$Y�~V�	(Y0/J���A�����c��P�I�F.Q>˓�RMbՆ�;$_8:��ٹPW:��ȓ�r 
��2N�zI��K�����	�p@N,����S��Zӂ[ 0�H��F֢k�B�	9���PAÒ-8x�T��k,RC��( aP����
l��Pp�$�7>*C�	�C���τ�I.�1��F��7��C䉸b�&�s�o�:w��!맣Нox
B�I�9f�1�5H�l`�`�a�ЋS-B�I�ao�|�S�T�G'�xyfi̲|L�B�ɐ����5�Z�����"MTB�	���i�G�"�2��gB�8kRB�	 -�N��W�öQ2.Ma��,Z
!��Z�t��d2s� <���Ӧ��3!!�S�l��0SF�3lQR#AK�9	+!�$}���a�v���hSlٹ!�d&S��M	�Ծ�$ 0#��#*g!�W�`��)� ۶1he�f��-W!�$p�t`�L|��,+�F�!�$�'�!����70舠��N\�`�!�R�:KD��� &0x.x����!�dV�>�:�ˣ��yk��`>!��Ք(�Z=�P%�L6�<1PCF*!��
��� D�.BX��@�D4!��P�ٓ"��6u����5+!�$��[`�l�`�so4DJ]�D!�26t�t�� ��,rZA��鍜=/!�d�9|r�ȖF�#ZP�$J�m!���� {��ҽwq���B�	e}!�Y��0��@e�!S2Y���M{!��A�p�P�
5/\X� e$1r!�$[�~B��	����T��2b� f�!�d�!r�0:�Ħ)�b��-M(!�D��k�x�r���1��ɤ�i'!�DY�0: PQ�� R�|����}!�d�W��j�%�1P����,�y!��U�E����`��;�bY!�d��$���	�iø<��/0�!��u�*<B)�����уR�!�� �i�l��&	��S�L���AE"O�8q!�8LTLڄ�Bu�c�"O�]M_�73��ِg_j`Q�"Oj��G�ly��q6Ɓ�7B� �g"O�ԋ�ɞ@`1�3D�)X�` �"O�h �$�P}�86+�8�F³"O2�� �+RT0z��E�>��"OZ�q�lV0eϊ���қ&u��"O��h��	 �r�bA��.��c"O"�S'�.C�J=�&	�f�4� "O��C�\#g���3��,F�%*�"O��xP��<=�*%Yx����"O��Z��)9����o�O�,�"O*�X�KE�=�|���9�F�t*O28�K4_^��D]<w8��K�'�젊ա�#Y�P��@�ךhfܰ@�'��!��U'+~-J�+K�TȔh[�'\&���#F��`k�D]�S^�@Q	�'�H���-t��Qo��Ay ���'9J��V�]HbX)�T�������M���@��B���5���׼<e���A�ten��2�)� ɫfo���yb�\7`n5���67
�bGl@
�yr��#�J�Qo� �4 �e+���y�j q�j�(Q,} !����yrk��r�2��p��=/�M�+�(�yBn�< �A��{0lS���y�cɪw��,S6O^l0�x` �y"�Ǡ4i0,�vN�6\�ب�F"�+�y"��{?^���DO,R�D���`[��y2��+Mg4R	O1Y2r ��y"�+�]{V����Y���Ȏ�yR�C?X��ע�>�<�QB͍�y"�\��%��C,`��1�s�Z��yb��*f��5r�(Q�^{�X+C#��y�W+C�����BR+]N���s$� �y��!f%��a��Z�~�H�+�yBC�D�t,�G�֤U�"�2#P �y��:Iq>���)��G���k�/��y�,ژwx]���_�o�E�TL̂�y2�+>��q�l�}mB��� �y�J�� (
Y�WGW�Q����9�y2�ƹj/�j�Ò^8��D\�y!	�wEZB��uO��CG���yR���I�xY�"'oǨy��l[��y�RR����K3jB��2��)�y��R�r �BK�v�
d+�j^�yC��� @�o@�22��*'T��`�'S���!� G�|$�d�(]bY��'�>��g�0�DhJ�Ĕ|<1"�'�J���l�#�21Q�	{T- �'Q0%�S�A�Tz�8@��˂�\���'#N=����	�fչ�關8�h�'�Z���@}t	zgL��r;�@�
�'c�m�`�\'qP���;>�H��'&8)���G>Fqΰ�R+Ą3�����'�<,�f�$츒�A;|�⤲�'�*C��E�6Wl�{� ,zCp���'��0���D��u*��n؀(�'\*�8rˇ��j��c�Y]z<a
�'I^���U".Kp�b��	g��-�'K�Z�C�k.@)�A/.��
�'�r<���B�t��	+��O,5ܑ��'��9[c���b�a��L�0)�i!�'�L����FM!�).Z��:��� ��	��XVqY��Z�h���3�"O*|h�C�$e� ���z,�f"OT�;,E�mߤ4��-��%)��R�"ON�襅[�xe���t�I7>��"O��1��}FD�9���x�"P"O��	�;\����T eR���"O*�8��]�&M�{" ��|��52�"OF�haN�n�0Z�.�2��h�$"O:�+w�[�@`���&���Q@"O(q���ɾ}�$�Y��X���"O�8q������^1P��yb"O���kW�I�Hp����|Z*Y��"Olp"$mL5VLH��jҔ�F,��"O�i4�C��m���_!R�0t�C"Od�;嚃Jd���glS�?r����"O���Rc����D��9�!��"OD���,���!���4S��]��"O��j�$�[���!�"�*t�<"O�5k�f�#9� �Q���v[@"O����c��P9�������"O��ksi�<��J!�)�\ X�"O��X���~6>�@��
z^�Dr�"O����Y�"<+�oG>3��pq"O �ThB�7C�aQս-h���U"O,d���
�28��2GS���"Ot$��Q�܀�BG�B7���W"O��HЉ*9�0�:��=(5v"On|� �)EUR��A@Ȁ3���%"OH�3B�ˉS�
L�D�u?�c"OJ��)ح`Ă�`�mU2p��I�"O��Yg�X�Ȃ|����=w�j��4"O(�VE9��l���1�9"O�9��ȍ\^mk1��6Df��"O��;��
o����E/j)�XBa"O�!�e��+e��x���ՍO��(�A"O����T�iED�(��T$B6
e�"Oʤ0N%ubR�x�!�= 1" �R"O�V��-9H�J�`Y�a0֌H"O����Gf"��� Y
8 "O�����l���D�j*P"O0P���4MKl5�7��6�� "O`I�e� =&�j�� �K]�#u"O�( ���6�Ȃ�ŎC��"O�4BVM0n��h�1�P�6m[�"Of��F��x�$��u��(��!��"O`(�(�1IS4��c�A���	�"O�|C���{ڶu�+�(���a"O�������BH� ���=d����&D���K�C|��C	��`����f&D�Ȩ"��40q�j#�>������#D��µ���UUH �1�I;JrRB䉅;�4P�c�1ZzPI�*�8�HB�	�n�l�"o� i���1Gi�~�@B�	�N�2�Ae�O�)Jt���(5HB��,>�$��N�t }X��S0E.B�	8�`��%@"c"��9���[�8B��wo�,����-�x���T�(B䉲f�X��l�*6�-�1gzq�C�*� ۣ�0�)`g���C䉞$��T�W'�j���&Uw�C����{�n®C{���W�ޭ�>�{��x��aH�2�l���d��a��3D����d]�y�6	r/D�������4D��1U�2i��"�"Woz�q�2D�� ���S�V��
"+�?˴���"O@�*�@��ุ�
�4A��\K"O�0��^Y8p����l>U�R"O�d���3��ibec� 48��R "O�mr7Cu�*Ca¤g8D#�"O��B��T0}>�{�G1.-��+"O�S���}#n=j#.&_
R1�"O򕂴o��B�s&�1���f"O��R�����	����6����"OX�w��$kG`�
��@�E�X@�1"O��jE����*� u4�1&"O�rG���g)�9��D�'syZMH���I#�l��"B��J��B�N���C�	���u!p!B�_��)��L�[�B�	
��l��9e�Qb�L�,w�B��i8
0���+I&���V�H#B���6ě@�A�P��3�#��coPB�	� 6��@7�E��z���L�d�C�I7.�6$�vft
�����2#C䉼+�i���&_��|J�Fև9��C��!oj�t��3`�UXg�3#��B�	�	�nō(�0�p�n>��B�I�tǞ5��'۠�.�iG�w0C�/[����3&3D�����;�B�I_�tP���l�0�;�dD�|��B��{+����E]�����sD����B�I�k�h	5�N���mj��=ԔB���8 &�
k�͡��W8%vB�I>#R!@vC�B(�dp�(�:%.C�2f4Aq'͒nL����Ä�(��B�I)p�b�@"k>b�P�n�t!�ط+q��F
�t#�i����)m!�3Q"m��ϊ:v`5 ����	�!��X=�}'�A�t���R0 �!��K�f�a���J{��C+��!�D �_�9��2��y�G�
-K!��#Q�EZ LK#G�0限A\�_-!�]I�(�(dE���PSt��7;!�$�*���t�,VN �_�`!�9njH	�EJϗJD�xهOůO!��΋}G�����9,@XrU(˦V]!���3pMtȨ���~%�%� �̑UV!��N�N�ك뚇B	�,r�Ε�5�!��7-^��pg^Sc� K����!򄄣��aɴNR�SQ�-(��9�!���g�`!!�%V����4�!�T�\��i��惵"2hQ�OQ�!�(IN��&A�"$���A-O/`~!�d��6ukU�G�
��'�6pq!��J2:��Kf�s��=x׬W�0�!��9Kb 1g���fLvlP&��hC!�D�r&xk�kO�FCZXzPl�^1!�^�,ai�i661J��ӼD!��`dh���5��m�
N�	!���}0��]$.r��R/�!����6,(f���I2�P�C�9Y!�d�=�.���%d�p��l��
W!��!`�^�z��ƄR�C�� /I!�K�r�tY�È#T���HΩI)!�Ćt���9�Kǎ~�Ӥ&��?�!�D�/��I��,9�������I�!�$���&ȓ%����(�HE�$�!�L���|p���(o�|}*�h4'!�D���\�mȍq�2��3e�1&1xB�)� ���Nh�$��&  ?L|�t"O"5��D�K�p�9��S?\x�f"O�i��eǄ
���P�:"O^����K}���bg�x⢥�"O�A��d����StZ=�ч�b�<Q�m�o6�U)!XO�y��ŕ[�<�` ��|��Ca��=����Ą�M�<q�-D&&8:v`9�vHs��@S�<I7��M )�o#,�3
R�<1���������C�<�MJM�<a�(��m��9'�[:� %�`�S�<�0#�"$�h0�KϫvP��K�h�<	�C�	�(�"�⎐rc"ٛ�"L�<A�M7�*){�gK�TW|X�1��c�<�����G��ԹG'D?+�X�ʇZ�<1�(K~	��xm�9R�.�qmTQ�<��i�13�h3$-'����͊H�<��#�1N�`�@#E�Lw)�1
�^�<���+{�j�葬
�G�!�D)�Z�<�p-�:� ��ݟ!d�[�*@�<R�������.�$m��*�y�<)�D��� ;F���`��p�<��L�������Ȋ(@��P�u�<��!0s� h#Ŏ��;|	3���Z�<��# *  �   V   Ĵ���	��Z�wI
)ʜ�cd�<��k٥���qe�H�4��6_2<<y��ʄo���+�􀷅�5��l��#D�#7�6٦���4Fs�*�I\y��7f_��k�D����ة�L�G�ԁ�%�vJ�9�=9��9g��7��,#�U�ϐQ�8"�'�Ir�dT�smÄ3m�"A��y����
0���p�2�NS"bzpw� E��0�B�w}�%�6f�^}����
��zל���G�a >�(%\���b�c^4)E&\I ��_?��?OT� KU�� �82�S	:��	�4{D",�@�p��+��I2���S����9_�PL�'� ���*���'�"pR�Ƀ�,H!����6���'��GxR��m�'cj0����y�6���"{t0Bed6�>�r#<9��>�c-�%X"��V$�(�f+*�-�O�J�{�)OJ�͜W�L�*WCW6�MS'#>�C�#<c�B�p��x��Ĵ41
4XU'��L�>���;�E���.<��{���m�us�f�,?x�'���Dx�VI��x:K%��@�雕�ا;Q��s��/��#<ia �O�8�h�5LF�$�ӎؾ;�j�*��d�>�O$� H<�O�-���Cb'��3Y&D�ѭ�x?��� �RxHOFL��b¸	�&c��1���w�R4�I4���f�DGn<N�'�~"Cg��w�t��3MX�Z�Te��W|�|�$�6ቹ!�$��B�g�TV6�k%B�
&����'�(XEx"��z�'NV<p�K*-�<a��%%ڍ�'�vݳ@ ���W��o�<�Go�� J��Խ!��P:��Q�<�'d�rI��B�j#��U���UM�<�B�#��PK݉iή�X&��K�<���\P���ɤ���B��؂��H�<�R
4-h�8�'b��QiKN�<Y�NG��Ǫ��fJ���bEFG�<��L&�.t�Ql�Q��pP��E�<��#ܮZ&���g';7V����<��'E�k{�d�0/��I�4XZ��}�<��d �E�� �L�Rj� �a�<�B�E�`MVM9�lF�N��F��a�<�� ePP%@f�ϞV���xR`�W�<�4*Z��Ɣ���\�5���"��l�<�"��2]���'	��2ސ�+�H�C�<y�6Q�\��q�z6�����W�<yF�ʎq�jDʓ�> ��W�<��	�&-�2�{��t@n9Q��j�<�HC;Ģ�1��I�J�(1QQ�<9v��e�pRDC�9�b�
īP�<AuퟱH�R@�5���K�z���Q�<���7�&�#�͘4ǎ5���F�<)V�QJ�A*u>Ƽ$��]�<	c�F- ��
�g� ��u:S�W�<��II�)hL"��ε�Y���I�<� ��#��WR~����/(s�5W"O�{��Գ-`ô�V�E���"O���'��i��e�V&(d"O��%!��=}N̻�d� /FX��a"O>l���@9RY��15$�uB  w�ßXx�fP�v����'K��T?�{�%R�$L��BF3.�IS�ֿ��� ��?i�<��5�dN ���r�`ί~ʽ��+{>9p��
k���5���D� ͓�O/ғ]�E&��%0�`{�G�h��ᤥO�\(֩�6�� 
HF��>[��"��0ʓU�	>�M#���d�icą0�/%ް��CV37��7F�O`���'ATm0�+K0Tf�	��-
��ɨ�����f�R7��{,�!��iX�;G�]!:���(�l���4�?�����i�0�����Ox7���3Pd(����c�69AeH��e%Z�������Jj\����V�H�k|��A�t�O�kF�9?�I��0� �ɱFK	T�F�ʃl�5{E�\���Mf�TD�\c�4�C��F�D�8� �>���ߴuJR���՟X+O�4�s�Vu�sa�9\�pl��[���P��O��d0ړ��'�NhX-Y����$�=�	9���^轢2�4��O&�n'��Dto�"��#�g��g����	ğ��ԁ��;�fE�	ҟ��	��c_w�R�iTЋ&�ݔ<$�ZN��,�4�$&X��ӄ1��M��şLT��� �O>�����1��4I�b872.Ta���%jJ����ɖ-�rb�f(�SY'Db�Pz���*w,���R�p8c�h�>y�L�ܟ��	���?������r�8�/e��A�r �7Gt|��'�"�'�ʟ�O&� Tf^����!�;s����l±�McR�i�ɧ���O��	#E8��`TF�	vb�X#(
\	��
 lѽ<�ĵ�	ğ$�IꟜ�A\ȟt�	ڟ�J*�0aQ��` L�R�iS
�,z����b�H�z����o� i�d�Ij(��
�Bذc�n@�Rs�8�Q�קV�6<"D`3��   	*	A��k$H�xeb��{$��O�53Ц��S]���So�9|�&�����im`%�x��˟`�?�O{�h8e��R�Nx�G���pE��'4�"=E��_p&��k6��y4��&��9�~b~���lZIy��2(,�7��OL��~R�M?mv�rR�:LK6��RM U�)Ц�'���'�B��瓊L���I�'wN�8����|
�BٴYt�h�r�.2��b�UX�'� �(���1*7��8v�V������@�$�l������p���Q!|l��(N3c�4����On���j��)�TFݾ�8%���� ��<h�D�2�?9I>��S��?�"L΄���ҢP�8����,K�`�'��6-�o�)w�ڝh��ªP�T�dd�K> �*@�iA�DC���>���?A��x~�U����?)�4{�|���� _�������w�y�G�ϰX�V��V	+ڸ���/A���'�����ט0h[hxe�S�s@��1mP�tAt6�C�?ǔ��S�ND\�;����S�ll���s���磖�l�%p� �wS]KAcc�~���'646��ߦ���~��M�Æ	�O�H񪙽��у�m?����?���$�Ob��4�IRm�F���+�?]�L1�u�Vb�Q���޴؛V7OB7��O��%�g݁1$��lmdMPqL�/f �Y6D����=��$   �   J   Ĵ���	��Z�ZvIJ(ʜ�cd�<������qe�H�4��_?8<�q�i��6m�M�X\�W�]�Cqj`�Jʦ�Btm)�M���i��F쓄�ؒ+��I��+X�
)�G��چ/��3 �"�{b@f�'4mZ6��h��b]BzP�{����1���#�-��#�@�� ���(6�ٱJ�\�E����A�eLIY�ĸR�BXC���l��&�ğ�� )O�i�8_��	P@��V��я��s�H��,�M�'c?��L�Rɺq$���튚R��ɋjt(����Lve(SMJ-VX�Ih�@i"* �ɿL�D�E� �	B%��[�J�ℛv󤇠�O����kG<��ga�8 �$Ւ;�EFx��\�'���'�~]�0��H�`�QDR8Q���cI�<S�ɚ'�qOz�� M�'��,�GE��"�\;D�i�5Ex2%�K�'B�xx�o]�,K�HbLD�-].�D����'::�Fx�N�X~2@�����! �'���q���� �O�BL�7e�� 9S��#G8���Ό;ĀDxBlGg�'̈�ɇ�T�ҰP�;.�m@W�	�@b����IR��'&2�cJJ�r�̓��[�6 ��'�*iDx���Z��9�~$�! 2-��E.1��p0�̀��?�լ�>A����e��s�T�O���;^n�5B ��1Y�}s�4��@A�{
�}�'@��O��)�!�:b��G�>�.IµT�l���I�m��8�f�A6����5�؅Č9;fe2D��h�   �$ J](P�y�~�i�,/D��R#ř"}l����B$~it�"�.D��XvhN*,.��Á��f�F�r�!0D��"���;���s�Ɋ � I���3D�`r�� =���cv)H6V����d0D���q�O�H`��DoS� ���/D��ZU.�1@�|� �Ȣ]y�\sq.(D�h[�F��Yҵj�h�S%�'D��y�e�C��\�g�T=�=�v�!D�D���ߜW9b�j�#�8 �Yڔ	?D�ԣS͔T�J	��ϑ�r����c=D�p(���'TVl�����20�t-pө?D�\vF�FxMa��E!R�45K*?D�lcc���lqR�PB'���[�D;D��a��M�_��H��_*I��|#&�:D��z`O�}f�"̟6���ˢo7D��ʅ��YF|�����	`��5D�1��Ȕx(�ڟ�΄q�i4D��(Q�\�j�    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �   Y   Ĵ���	��Z#tI
)ʜ�cd�<��k٥���qe�H�4��6_?><�'��4f�V�R{�4��#��:��Zׅ�J�7M�ܦAZشIm�$=��[y�!+3��	�� ����摹&~a�灑� 2q�=	�((��6mۻ|\Պ����&��8zկK"��ɦ>���í��$g�	�Es��{��o}�<��H@�,��X��g��"���q@-3�d�#.8�|Rc��r/8H�tEL2td��Ҝ`C�����eӠ�y�����?���(S���	n>��8s�&�#�K�.�kLE����`�!$&6܋��[&F��D���%�1�+���ʎy�e3��|`B��#Q��� ���y҅x�'���Fx2,�!�`�J�d�!;c�_4M��#<q��,.��
���sՍ�*s��5���8#C�%�O0����$���'�b�8'��%&�֡�$�[_�)�4d�"<q�#��n`@�j�%�2���/9|:�E��{�q��"<$. ?ɓ%N3	�X�h�(�Y�8�k�D6?�..i�$�@+`k .dlNXAB[*8?�Ai��ċI�`{��Il�b)8c�9���,F�I&��'ݘ'��HFx�-Wb��	���� �E��qS��Ԅst8�	(f�Lu�x��Q�<�16Nv��y�ƌ�k��X�Y��� ��Oȥз+r�3'lę���E?�d��F����4^u@lI��X�Sބ�a'�	���X���>	�㐏%��p����#F:�
b�G}��a�'M^�Fxb
�!.d�|����.L�Q$�ڛ�y��A d  �'w^h�aC�qĜ��퇾<����'\�t��t�Rh"0'�"e�����'���ɲmҬ]7R����Ö��y��'LpD9���G`^� ��!����'���!�!+����O�}2���'������@�Vx�	Ѡ��sh@���'�	)ad�	��]C!�ޤr%Ƥ�'�����1[����CM��byT�0
�'���@O�l4b��ܞ%H���'q�i(Q ��ݞ��b��.� ��'�:e�%G):����ХF"�F���'��(�RL�"JB����Q���'(62�"��0�JiC���4`,
�B�)��,Y(`XfmQ�g�]� �B���<���ߟr^�[��Ѽ ��ˢ���!�Ĕ,,� �i
&]��j�� M�!�D%��P�MB��5���K�=!�,\    �    �  �  )"  m(  �*   Ĵ���	����Zv)Ú'll\�0R�P����=9pn\�Ёba�#������{�<I�d� �t�Z5$��vT�aN�!@ i®�,]Q�����E���I�A���0�2rTƌ�&���L�/xP�A�^�M� maf�E�m�];g�0'h{G��PZ��xv�Ӳ]m^X�S�a���N�y�D�{�e�>;P`���H�F���;;��ac5����$����72>���)ӹ-#����O����O�e�O1a�Ta��x)���g�%i/J��T��<��F;�"9��(�<1�)ޗ1	4iY����@���DƎ� ���ғEt���0 S���?i����l}B%�iU�`('.�(���x��[=�M[����p����.�|�',2�O��j��֝'9ʙRF]]��e"O$��nں_�p���M��Զ8�D�iL>"=Q��:�?a+O�q�JV�W�`,�5�@���#Μ�q�L|��,�O����O��������?��OYy����
4ɷΔ;o
$�06�P.�Tq5�'i,�P�'	�@ƪͷqº��f^�$ X��	�'X����fB쀀o�~a@�/j<0P	�'����`P�����cb[d���"	�'�PĂB��qr��C�[
_�\Q�O�0o�{�I<H`$4`#ϫ�>����%��6�(]�΅Q�.ų.pA(�N\�;�!�F�a?�d�t�Ŷ32��j2#�8�!�dQ�P��5&��O*Bx�'���!��P%V�-r�*E�����1�!���$-�<��)[ lzP&<p�!�d�Z���bH��O�%�UJP}�!򄍲a�ĘJ��Y-D� i�&�F�A�!�$o�9Іeh�4sƆ�2.!���KFB����7o��Az��ѬV�!���(Z��E	�Κ��;L�!�d�Q9�Y��Q2� V	F0�!�^��c�.$1��¡�$_5!�_7r���R ��9HH��wa��!�䓢.P���f�7}ĸ�1 O��!򤟕o{zH���3b��u�k�!�� +$���BP:�ԩA�g�7"OL����TV�ИSD# V��A�"OB�16K\:[E襉P�^�a����f"O���6O�W�x�A5��&�z(@�"Orqh���?�lP�B�m����"OJ|Q�Aקh�h4A�k#z<��6"O 
����$�!�*�
0kx�"O<<N�K+P`�)@(fd�$P�"O��1V����&���I�J��t�"O��3`ţq�`��3�L�g� ��"OX�2�,E���1��]$6�5(�"OΨ�6�W�x��D�@���Iv�@�"O��*�ON�fX��L�\�r��V"O���t�>�BX�%��X?��B"OnqbG�3 ���΅~-L�`v"O�����?�H�+Nʋ!t@X�"O�h#)Ux1�/adܡ"O�a��ኌE�@I"T@�08V�*"OJh┈	� ��I� -n{��K�"O�i�Ȋ.Y���'��Hq�9��"Ol� �T�>�kS�B�<i&œd"O�3a��w���`&� �D�-�P"O2(�VϜ	��!)���y��ږ"Op K�d*���cN�h|�b"O��Gi�E ���G�&wr�y"O�(x��Ї-��A�m7:Y��	T"O��4oW:Ikp��&mݥfhv��"O��2��$y�P�Gb��!e�0�g"O���b��n�ި��a��b�P�p"O�m�G�DaL�,�T T�Q�Y��"O� ��F��2q0�a\.gLh4J�"O�STB�'e�z�ɤ�^��4JQ"O��Ұh��3�x��R�L���(&"O� ��qC�k*�N�b񺡊�"O⥓��,6p[ P�몠q�"OЕ���n��bv��,�,)t"O6��#�ϫl�4	I�@�#4&4J�"Op5M��]���A��Q$����"O��#�S-?Q`S��!@���"O�L����)l��Z��p�| s�"O&�i��ϊMܑJ"	+:�@�d"OnؙJ�h|R8ѓ��ȍ�"O�*a��q�F��al��)���"O�l4Ɲ8920�qQlا1���1"O���NZ�����6��}��"O��dlL�r�n�x'��XN@ڥ"O�Xz�턚ؾi{�e� ��u"Od�!�%�Y�r��2x,��e"O
�ݝw�>5�@՜*_��ӓ"Ot�[QꌁJÔ(�v��[U�x�"O��{�L�~�ш�!'F@��"O�*�C[/P��a��e�VAh "O��9��G���Rk�5���Q`"Ox|�! B�Ed2AH$�}�\غ�"O�̘uBÉ7�H �3�X<8��qp"O���"&��i�L�f�Q���8�"O��ӂ�O���}*'�N�\�]��"O�X�`�Cq� ��%�4�D�F"Ox�Sq�>R�`i���\-�4ye"O� !��C�P�TU�E@3N�ࡁ7"O8�a�P)�0mN�lJ�Ѧ"O�����=&{��tɅ�3Th�� "O.Ѐ�I�$4n���G���P�"O6�@��;YS^E�˓G���:3"O�D����cJ�hr�<Fq�u"O:�3l[j��H�f)N~���J�"Os�6�9�"۳�L���ի�!��C!=8��#���l�ZxJ�^�\�!��7N}k�PY���`RV�!�$P4v<��O(�h�3���%N�!���'�E�����ĄA��M�sD!�D�,N^̀¤Y�1�.��r�-
@!�d�$}d��"ݣ`L���N�-�!�A�JH�zvm�i�N A��De4!���.:��S�&iތIrs�W�i#!�Ï2�e
3�^�|��a�R)�!��3O�S�a�$���Ɇ��=;�!�$J+$�X��d̆f�Ya��$m�!���b��}Cw��.X�=��$W�!�$�Z,�PAP�ۨdX����'ƅ!�!���,�@� #S8~� ���QzY!�ē�ex$�����O��7�/F!�ě���%��F��ꨈ䪁��!�D��(�@`ؓ�ϫd�\y��*�0�!�� Hb�8���O'E@�-����8�!򤋩;��xuAX�7�J��wl<O�!���q,X�ת�8E���ee�#�!�d�'P�D� V�	��*֗�S��ń�d�`8�JS�#u♘u�k�ޱ�ȓ+���P����|,�F$T�I-ez
=���E�$�F� (�|���<I
���_���*!�>9�IǉX;�,�G. &j(��2eP[�<!Ѣ�5�ʜ�o��F�@Y���^�@X���>R�z\G��%�:A0�璈F��X�B�yK_�# �u[�A��
�.SD,Ir1�8JI���D�d���?�'�b��5h�,yںm	G!ժ5��
�'1R�Ё�
o  I ��R(A,~�au@�.]h���$�*����� ȁ�Wkӯtq�b�L1�����'?A��!�)x�0�Z��2���FR�Ql$��f�Բ5��K2��2�y�2F��܉�Iь L�q%�G����Y���+�BܯXF�<S Ʊ�(�@����#y$���.X��	�"O�R��Y�rQh	�&疇E xe�g����+�� )rnxZ �G�:�1�1O|H�R�רW�<(���G�+�n����'{|I�VV�"��혰ژ� Z$G B�`$)�cͮI렌[t���az�I��|�:y:�!�� �Na�Ƣ]���O�t���L�`NQ9��
�6]�`�c,�M}���r�F�6�ؠrE�ځg�JB�ɬ8;��f����T ��k�˓i2z�V�@�#�@��3#ޮpg ����)E�!�!��F�d���G��!�ӱ^�~���Aԣ:���O4Z8���<�D<U���Z}@ᤝ�T�S�R,��Jݶ%(���H\����C��R�@��(y�@�9��׫@ެ�5)ŎH������|�P�'��A$l�^����)Hu.M��!{��B�̠�ʩq%`�
W�!�B靚>�"d�!�o��d�"�G�<!��.?�1G��.�u"�aUl~bV�t �iER�XM���>ʧ Y@��F
A����F��
�؆�W��\I���#)�Iצ�<|��p�ܵt�X=p��>����O������	S7��@F8�����"O�MI�5-� �Q�~U��)��ii ����8`�p �
�9�4�ԯ9Ft@��:YGjŇ�ɨN��C#�X��y2G>)�� �c�FS�z�b&���y�I�9x`�)� K��^���bq@	���'(XRF��Ef�"~�T��#
x� B��-h� #.�d�<�`
D <)(9�&�(eZ�����L&@�|���~���$�-in�R�B,
��U�󭏓E�!�d��|�	AF��h�-B�|��Ǘ�`�a~2�^�w�R��1�D�@Sr1���*�y"�\]�� ���0L�
T� e��y�OE
+D���&DO!P"�����y��B&)�VXav�@'Xu�� H�y2�άN��y�ՠ'�VY��͏7�y� ��H�����xI���y"�I�q$X�P	��<_f�!2���yB�+T&�(gA��7Ų��e�� �y'��q�	�-Õe��Ȕ��yr�2E3��P 睹(���aǥ�'�y2�ռ���W��q� I��ǟ�y�mS$����lM"6X6�:�+�8�y2�Ƀ+|�L2��-���k刎�y�ʈ_���ң,(y�na$�ɴ�yO�0[ 
c��e �y�`Ҡ�y���-C��#q!�/y�0`�I��yFZTEz�1D�E���Yf�B�y2�̱a���+��S#!=�ʀ:�y(�6A$�p��W� �.ɻT�&�y��̄Q��,Y��V�d@p���y���r��x�d�@�K4	��G�<�y�A�=P��j��Trh|�V��(�y2�\:3h���feїf�!F�G?�y��$`���v�`�И����y�K&N�d�
	a�@��bѨ�y���@S>a�5�S�X:�yR�ĘP���P�#S�h��	��yR�U�V9�����H�����N�yR���H9�d�XW��M���]
�y�K�1W��&�%N��jq�Y�y��Ä j�Iy�Ћ@+bQ����'�y+�3y樢c�/�`@ ����y�Ȉ%,�I���w�5�/	~pB�I+<�4��ՀG�y�� �ψ5<pB�	���E� ��?WI�a���EB�ɦ4pv����:0�j��Pe��N��C�)� X�0���'�f�(�����$�e"OЕq�/��<̈́T����5T���3S"O�5��۸�)�eᗕT��-��"O���!Ȑ:E�� O�7�uC$"OFЁbI
 �>D�F B�*x9y"O�к�E9)w�Ժǭ %T��Bp"O�Aխ�	\��U$�:�2�i�"OޱJ�o�+�L!�����ՙ�"Oh���O�����Dハp=�� �"Ozap/|��!�B�@3Y���"Oh��M"� |�d�S`"��s1"O��	gZ26�0Qk2LT:1*lr�"O 8i�	�Gm�QAPC��5���ۗ"O� �"KƧ=�(�[�'�p���"OTU�ҏ�d�PP�s�Å?��y�3"Oh9'��x�v4s�
�-��@x6"O�⇨��H
��XҦ�2�Ɖ�u"O����l� )Τ�c�sS���U"O����۴�R�Q�J:!I���W"O)a�jWUS �@J֋B$�)2�	w�Z�� mXr��$ �G��6�ǀ5�ؚ�O��etDMs�nģ@!��N��Zb�Å/i��i%L-H	!�̅]l񕂉�Wb!bL
�!�Dϳk�|�H��حy��!jY}!��>�����S'Mu^�q�)�9_!��A�{tp]#ӁQu�4x�j�!�Ė�1�\�F�^�~7�5��J�!��Я`۰@��0�xh���f�!�dQ�o��q*Ò+޸Qss��!$�!�d�9>�H�a�{Ί�B�!ʶ4�!��«@C�{��ќ����+0!�D��N�� � Z�@�B��s!�D��`q���wM�%�䎅�[�!��i�Iy��6n����-L�!��.�<�w�DՀ������Py���"}ΒD����fQ�u!��]��y�NB� THq ����;0�Z��y"�
U�+��٠ ֲ�xV(]�y��?��h���a�̉�����yRM�:)t�B*�,�dR��O��y��� � �h^�!`�[��yү�!���Rf�	d��������yb�;C���!&c8RH�@��y�`�iM�AP��mn��ke���y2o�~�̔� @I�bm�P�e���yBeOt��Y�LٸB���-Ԁ�yrϛ)O���k �0	�B��t�\�y2)\٢\�D��*B�rW�Y�yR�$o8��ІO�{*DZ�L��yB �	n�H�C2 [I���7���y��V</v��$h]�����M���y�O�U$n=�c[�R�hSV��y��&��uQq�4L�du���?�y�A��I/���G)�I��䳲�S)�yr��#�T
2�C
l ǠH��y�/Z�t�z|�v�߀:��uZ���y2��o	thl�3FƠ�#��G|!���a�"e(��I	)W@`�Gڠxq!�Dn>��(0�M[��I�̲o!��/q/v����&�b��!�ܓR@!�Dݤf�����Z�SD&D �ax"퉚4�(eХ��6�pm�bP~�jC�	VD%���U�$U��)2�C�	�
�pA�ҮU�Y4�qj7�KJ�0C�)� �@�RXw��J�lء0g��`�"O�a�nS�)�>��kX(b��t"OfѠ��K�Om���R77�$}�$"On;��%W�@Y�d�[y$<�f"O�0��/�2�1ƦP�Pn	�"O�$*���0t�[�e�}pM�g"O�h�eo�4uxD�%�I
p+w"O���)Ā~�h�0u$�8	�RS"O�,���jt��	a��]��"O��Qd��`���&j� �S"O�����M�~>T�[�B��zU�H�"OL�*�.��c"[�qR�E��'J4��[�x*�`ܙA�l(b�IW/�y2͖+[�t鑦b��lr�ډ�yR��'x*0	�o�5Ka����P��y�F�>
��!
7ni����)�y"ŉ�'��-�u��k;��Z`۽�y�"ˮ2�0�	-�j�2�ϓ�yҀ�0P��1�)�%�n(�!bF �yB�� h"���g�	4�`]���\ �yR�D,�� *A�)+^j��yB(ݤ=�DjS�o}UP���yb!�_6Ҹj2�ЭV�FQ���,�y�k�8Yh��#H&�����'�y�-ֵ!�`|�0|�r�A�8�y�jX�o�0��PȷGT����݂�yѢ>>X=�� ;�����	��yB�C!X\=�w!^�.��Pq!D��yr��t�<�S�"�|(�@��y���]"$�hhL�	�kL��yb��놌�c��5YShaX�݃�y�J�A��c���M9xt�ĩ��yB�վ d�s�/��GY��Ʌώ��yr�<�f��0J�n�n�zE��'�y�i����u�\0w��ЄdB��y�@W���D�w�� o�
�����y2�7^$Jت�
R�g�θ�-��yb�G�8Yxʍ,m:��2���y���<'R��O�7-VH�T
��y"��=�`�DL�p��1�y�)�I�	��[2��Sţ7�y�JL K�p=�C/�?(|D�����y� ]�p/�|ۡ��62�l5KB��y�	�WԌ=��#�~Ad���ŉ��y��.8�
���4g�"��ܝ�y�e[  a�@œf��@�%dJ1�y��ǀ?���Iϊ����3ujʂ�y�2)�p`N�:]^�"�FV��y�!c	T�b���B]�U��+ �yҡ.k����U!���h��"A��yRυ'��9i!�^�� i���y��[�E�|*�K��k�̽BB�#�y�Ç�m'U���4;�ɛvFԱ�yB#�8)���
�<a#\9`���yR�UR�lH��D�ѕ���8B�I0Ba	�pe��#*qA�璸]��C�I�.�(���˻	������I5 B䉴oTP)s%X�|��q��@U'
��C�	�>�jt�W��?/�,`�'�onB�	 5I����9#"d�c�NbB�	�.̄ �I�j� YT�Q�P$�IR��л�'��Cz��
����*خ�{g=D����c[)o�,����RLA
b�(D��F��XKh���/�ٹ�I&D�� ��f��=�L�T �9&����"OH��3HH�"�4�a��iʍ�1"OAb7� 7a"<9�F�&qN�UPr"O
٪���'�L�
�Y�D ��"Oz�KC��$A��)��(�'�&4"O�d"�D)e�F�sC�W"L�^bQ"O�00�NN ��"���&X>x�B6"OdT�Q'�<(���BU��}A�}R�"OzmI"�^��,� $M#b{P"OKۖO*��wD �"�̉3n]��y���}��F�6"Xx���K��y���
�`�7���Hp�z� ߇�y�!�;n���R�-;��XS��y��KZ\�s!\�$P���-�yr#��<a��۵���	#�?�y��H7r��-K�J� �B0�o
�y(P �����$��ٙBA�)�y@���u��\ b�񨞠�yB�ƨz5P�H�D�7,%��
�,�y2J_��h��U�'2�I2��C��y�j_�wvJ�Pq�N�1��Сc @6�y�N=�RH˦�>����� ���y����q���S�V�3���;V���y�R�?��X�D�1��D�d����yҨ_�d����W,O��A狽�y�
J���9 �d�	��x1 ڔ�yrj ��^#$
��mE�@��y�DY<�
7��8\\B�{T��y"&��;w�(��hG�Xjä���y�	T50溱9�,�7R�*����y���%����1P*b�IĒ�y�
�Ա�_6m�P2'�&�y�e�1pəRIH���@y����y"�ݬ:&MS�b�87�D�CI���y"J��q �4
I�M�R�-�y���_^�H�/Z�'"q�g��'�y�o�"f�´HU�Ң.�537�P�yr�;���H�G$	�Å��y2 ҋB�8�����&f�����ybX?y�v��呄�8����y�O6eL�!�"�~BP:�Kέ�y��z������ds�͈�y���Bt,��a��`���@��R��y�k̢Kh��C��3X��#�+��yBlE�_q�X�+�
K\I")� �y��N�[�^@��G�1DFMB�o�2�y2HD'`��<{�dҷ,�B��2�T�y2W�]u6�с$�#�]�0� �y�WD>HɣG�ϴ����yNE;Nv��C�
�
�RC�V��yBF�� �LzdF�W��B��yB-��[� ����|�D9jҋ�y�O+p3�42C^� q*q�R!�yr��j���a�2X��p �4�y"O+��@b!�0��(�����y���<Ѥq �F_9i�&$��e���y"k j��l)f�Fc��MC�K�-�y��&P򩺴gH%[��YA�j�y2EǚInQzᩝgB^t�6Ɣ�y�gJ�F��ьv�f`��]��yre��F�H�"ŤM'$�NYҵ�@��y�B�8I�<����Fi�5�G#�y�i׹I8,%#qC���d:%	�y��F9K� -j%$�fd�!ʺ�y
� �x�k��E^&{p@�=F(�X'"O>�#�h�JC����)
zh�|��"O�,+o[�D��Ѹ�.Q;ZSZ�[p"O�|�O�1A�� �홨L?���%"O^�!�-�y]� Aި%���+1"O8�8t���su�Հ"�Q�j�pV"O�(�p�݋�sd�X@�$%8�"O$	;E�()4̤	��@8��P�"O��*�1��Q����Tn�X*G"O"�[��ԛz��y`N!J�%��"OFt[B֊~ܸ�A!�#���"On���]4s�ASB	W�\�18c"O�iV'�
^�ܸ���O�t��"Or�ɴn����51D.��AFu��"Of	9Ń]�2l�X�Ы�!W@$��"O��z�nU�YKl��o�kT�:G"O0�u�ƛd�Va�4��?d���"Oҙ��G¤_U���nPQ��s�"O,�9�B\;~i���.ŎW5���"O&�IW��:����L�0F.��:f"O0�"�(�'|�E���P�0�g"O�!�3*Y T+*�  ��7n��Tb�"O͡p�9%�\9�>(P�3�\|�<���J�"���kW�ԅ)�te��ds�<�uc[# *  �   M   Ĵ���	��Z cwIJ(ʜ�cd�<��k٥���qe�H�4��6_?><y�ʄd�V�k�,h"�l�A���օ�0267���հش=�D8�IBy2 ��E�@F�4mBԁ@�ϻU�,u���:$c �=�G�"�o�6�"eZ�p��7O�|�	3��
;2���<&f�J$a؏U�Ɂk*���Ȏ;q�I U Bd����:~�(��(�,{� .��O|p$)
�=��'�D��*ʟ?#�PȓNUoO���$DlPN�o�Z��ΓC���͡<q�O�e�P˩('ąm��6$>ax��L���p,O��*��J�)7�jC�䙲��Y�y!_3"���Ƈ,5PVN��yb"�w�'�L8Fx"c�J����f�q����w����#<�)T���%sp�����T2����&�W��O�)ێ��J���'�L��I�=f࢙R3#���:ͩ�461�"<���9�@�&9;��Ȕft��CV<�����O�H�� "<A!?A�͝] ��pON6$��s2�Ly�B�'����?9���JU�tȃ\��~t����2ܒ"<��a$�L4���H1*
�i��G�9kp��l\= �1O��	����1�ē:,�"vɉd
�yY� �%G, ��4NJ#<ف&6�[?Q�L��v<�k��o�z��%���\��P�l��O*Րg)"��'H*ם�f��`eύ$�R��Ʈp8��=	W�(�S��'�$�ޟ�B�kB���<���O �Ȋ�� �O����
��~�z0j�	Z�iR"O0�p�  �x�"OfY��IE1{�%���L.P]Z7"O�Y�D�1 ���)e��H��"On@S���9Y���s�ıS��T�#"O�$Ѐ#�Հs�a�Y[�ъ6"O�d��J�:�I1�E�$fИ w"O�)�9R�� pХ�\�հ�"OHu{�̓Dm�1h�d
<q�z�{�"OLx��Eƾ( ��uW���qȒ"O�8�"��V�9�2k� 3�ڑ�D"O��xs�Պ ��0Ѣ��/�u!w"O�D������� E�5F6x�'"O�1��/V�F8��Q3E	 "���S"O�li6�z0n� �_�N�P}�"O�QP��s��k����	�4�y#"O���c��0=v"�'�+���X�"O��ۦi6��yXtf��l�h�(�"O0�AE�(X2�9�c�D�.����"O
�X��Z�h�xQ�)*�����"O�}rd`S�tC19F�5uk���	�'<6�c���#�XI�@]	E�| [�'��Ĩ�� >1��bc�+,lII��}�65���1)���
���x�D�1�x���K�Q��(��|iL���E�'%��a����$p!�}��{�Z�@�J�8GR`����#����ȓ^ځ@��<����R	�Z��ȓ2�J�x�d�[m 0�M��M���v�����L@�+�b�{�Hs�⑄�N]�99��K|���g�ѱc�*���AfLZ���4�*Y���Js�@�ȓV�b|9���>3��c��+�D�ȓ8{�I�D���:
��` ����nC�O]�H��jR*�>G�B8��[ݬ��JB�8!���Jӌ��L����ٕ~�lHI�g��gl�%�ȓ	�^���)"�>P��I�TI�T��*�4{���1���iE-SL�&��ȓnf��jWdǠ<��v���ڝ��y���v@�H�̩��f�yҲ���^�5��.�!����з=����Dr��bR�Y������0��ȓL~zP�g� ����Q�܅3�>e�ȓ&"���oH�w�L�R�SC6Y�ȓS-$�K�ʈ�x�P<�3 \ �"���f�`T(�� tX����"�h=����k��EAd)E�m#"퍟D8���!̪d��<Ԯ�btGA�Mآ�ȓ!���Pe&���f/¬	�"h�ȓz��iҡI[���Y�͒#e�Դ���R��ī=;VX��oWH�@l�ȓ.�|i�2o��R���a�&97�хȓq��з	7_�u9;Et���'���wnƕ����V1B@�ȓc�8Eǘ�<N�� �$ձ\�~8��L)�I��)�f4�ɐ��*|l��ȓf<�mԤH
da�p�j�t�&)��� S�LEB��'�8�L �-�
4���� %J��X�'�\��¦�v�:ɬ�'q�Hs�.�4���[e"��H�(���� ,�� y*zX �"O� \m2�-�5��\�Aˍp��Ȼ �U��,�a3*H���)��<��*�?`�����W �6��l�E�<!�͊6 �t�� ��.��)�����<yC�M�Dy�­=\O�����9�
�`vm�y��	��'�����O;3�ra�E YjN��'�K�f�^0��y�"@�lQXt���T���`�!�4�O8��f℃\Ӭ����)�3d��c
�w��Hq! ҠZ!��77L��r�8k3�I� �*X <@�C՚*�`��N�"~Γ^
T�
�W/7:��yqJ�i�Q��9������Ϙ ThY�p t��I�y|��i�'B��$��F����
�J��ez���a|��
#Ḑ�e�ӣD�d��k�d�5	�F2p�a��'׮���AQ�W��-��������䟁?��u������(�8PI�Z7 �h g�]�>m(q9"O2h*B�\�^��m0F��7o�@Г& �Ĺ�uH^���)��<�Q O/OK���8*����\p�<�B�Sx}� ��]l��t����l?�3`E�-��h�e���G�EU��� Wb����	��"1��'��r��>FP"��'��P�<��'�l���%�	N��Cw�I*���'��mV�B8'����JJ?���S	�'�d�"J�"h���8V癈Bh��'�~(�����<�P�됞w+bɲ���^;�>9(��W����S��0d�]�oK�!�$��P_x�T]�d��!�n2p�]��A'O���hQF�S�R('��O����6Kv��(.�~��7"OD�8�P��%��x H���@@��9�s��Y[JT�'�T/{��I�^�Ԉ��;M�� "pD�8l�
��d��E��9�m (���Q�F��"O��`c��)c�Ԥ�sB�`���'�ea��JSB���AMGG�ȓ�}��2 ���K�e��( D���79�O��b3�_��$�k��D�2Vz͙	�'�L�
�͂0Jz�p��@�(^��ao�+�<(�$癀�A�����7
�,�I.�\�șw��К���P+Rh�Ј5q�X	�']�L��;�7��i�����!ʗK3N�p§<D'�u��-L�T�d��'~2�k$�ݗ��	=l���Sႆ$"�KfD��4�4��d��9s2���}��!�L�$S� �i��%����T�\�1Кt ��H��B�J�K�I��q
�'�M��`\��� .� |���B�y2N��~�����7h�4��h�-��wȏ)7�e��[�I�a�$O��CBڇ#�Y��'/���P!�z�b���J*�0R��Έ�T�'O~�ҙ�AB�#-�����|�l���j�(� z�w����5F�h}� �G�ۡ�i	�'����Ռɍc��X"w�Y~��e����Q�0��H&t��e��j�_x��H�,�a��pz�
�y��M��O$��%HBaJ��׌Ϝp�D�	�v�<1��]�\;rAS�B���%C�+'H1I£�.C���b�ه^4�͂"�$>��bĬ�+S֔u��	�;�6|b�˔1n"ɚ�����RjȘل+וO
�eKpi��L�r���J�nu������� �ѱH�y[c���N��AcJ�sH��'�� c�؏wZ"�&#���s��06Z�� w�D�@mօA"�9��(+EtP:�Ɲ% �䑛wo�U�A�'X-(���V0$�~�K��5j�}���C; ��q�РxP`1R�M�^�$�c�A�@�1��E�"6����O�r�(Ѿ,��'��)��Y*6�����[�:��э��d��2s�O�iC�hj�DV+pB |{
V�t��4��2;�:æ��6v�b˓>���`,;,O��[��LUߊ=9!�E,����V�t���W��+�nK�#��1��ն`LL�>i��'�M^�0���i��(D���Ñ\��	1��t�M;�-�H7�������s'N5 �l����c7�>���I�F*B+�? ��K�*P<�3$]�|���H!� "ZM ��UJ�<T����w�^	W 4�����X���۰<�D(�2zz���g��n#s!�J8����j��x�2h�L�A)8���@-?���`5B��7�е� �"O�5�6
Ͻr��m �B��$� �Ap��S�I��h n��Py�#}�k `t ��������
B�<	D �8i��xK�i��;��ġíѡE���v+w��b�����H���G3�Y$F;Yy!��H���j ��n'���f�F�W��	���,���Vb)|Oi�DꄖVy�\��3a[�j�'n�2�ٕ �V)��i����NS�R�~dpG�(�6��	��� "�zv!���Ԉ"�O�rU41����)�Tҷ�Ա�h"}���0@|��70x�y�@Q�<A�jTXP@�`��3$g�`ƬZ7�RE��EU�dC�I�k4Q>˓��8;��8�����[�&����ȓS0R|����l�F�rQ�R� K^�l��u�rm[�T+n����O�]C�:�d��qmH�y�{r�֝۞T��g��������TO �ք�`l��+D���
W>Z�^-qg7p&��@�+�I$V�Y��蔯~��>E�	��}��KH8RP@d"�L)D�����P�����K�_&n Q4-�;}_�"����	N��~Bi�)H�M�1�[�nɚ�dņ�y�k��(JDO�Y�X�"P%ƍ�ybI�#F�=���'eĂ��-
�� Ϗq��x�?L�9��q�$��P7Qф0�W-�7=� 9��-D��p3̝���,��/[� ̼s'�&D�$����r��8�X?�)��"D��:�,�
1�����?zٔ@
C�>D��Hǝ3^μa�`�fN�ɛd�>D��h4(W�s�� �Q�Jt����+D����$f|��f!M:L�6'D�l� �$kVӃ��.��ܙ���� I��eta|Riؕx30q	AK D<�u.�0>)�`�.A�xa��L\�{��4S)����ۢR�\Ʉȓ=�B��� zg^9�4���`�|������	�g�O6�#i�|�ӌ�i�:���k���y ���G$!B]B�nSL��3+-i��5��Q�FĮ8Ѷ���=�Ъ�ZL��~�� �u�+@�؊��U�U��K$U�.�H�㉒V�R�3s,�Uܶ�sPJ�<�h̀6m3~`p�A�V�W��X�!�'��`#��`���I�$�N1�
�+���@�+���W$��W ��V.��+0^�' \i��8|�B=K�N۔Q~�H��^= �7��!��]G0-��&R�}��ɂP�ڠ(ƴt�DҁXa6��G��-@����X@:%��O�"�+���M7g�q�r�U(:� �  �J�5�az�j�A�X̓^j��h�DηE/���d�Q�0�~iI�״SC�|;��N
�`�ח�?)uϵF+����!����'���t�է,��"�h�Z���L>)��CX������@RU�2'ت�2ԐթK���	�'��<��Q���l� j��G6�?��l��$4q�FI�G��y2�9��xV��j�Yv�J�T&%Ё�ì�1U�L�1�H��b�'2b���<���iÌ  �tR�R�z�rP��	\�2K��j6$C�ɽT�.� �GD�wdA:\XK��ζi~<����dB������r��d�V!��? Pp��z?1Ǉ��=�9X$�O�(�x2�݆Y�=�`"$,O^�0��S��<kܴ
i��T\- 	� �0��K����^}��ѳx	,e��Oqy��W
A����Lr�I�0a*W������5�8Od=ڥK��`e8�4E���˷��G�b��� M 'X�]�I�(��H��1��dQ��K�:�Gr���
�FY����آ;� |�b�A�\Y��E�Ơ���K�O����N�R3d$���S�|�Hَ\N@ �vb����?�Px���o�2�90��4��"�+1hn��iқ���.�,��f�n�>�) �n�D��|�n�7\�
��Q�R0[�4XE%FjX� �c�$c�
�y�Z���
Z*:���.�-��)��Dl�^Q{�4q�ص�M�"~nڮ/,� {Ce	,���@�
x�O��!���z���	Wed #�UNJ��#KY'��I�l��lj��\X��y���K��ģ���en�(X�ě6k-���=a�u�'UN�u���?K�`c�Θ	9�<���9D\�%��'�MԋόO�����,L��C����h�~����]�tY�� E�%n��!�CA"�!��ŗd�`T!wj�( �sR�A$D�!����`�pP�
�����NS!�#�ڝ��I�O�
�����%!� w�y�$�.Oٔ"t�)P!�dӃZZBa*QkRC����c X�m	!���+z1�(I&r��d�q�@�K!�$�φ�H$h�03�� ��34�!���~�0��6.ǁj��\��n�>}�!��
Y�XXcCY�f���@�^�!��O5��e��H��S�Ʌ�e�!��Q�Pd�O� t�,�!�� �P�c�P4"i�Տ�mX	�"O�%8�mR�#���0D�٣[�T�4"O����BOS$�q@!4��"Ot���B�*�3R��K�Q��"O<�����H?��� ��Z"O���K�#b��S`�C�p�L*"O,}ᔯ�N"&���Y0X�hٵ"O6���(��:�c7cP�P�XP�"O` r�F�M��2�m��~��4"O�i�ӌY4̖�a6>�%lO��y��ا[�����Je��f�A��y҉&0���0�(�NW�����'�yBL�=�f��̩~e���b$*�yr'S�I�v�C ��8`�ĝ��y҇G-"B�D�E� v��yF����y��{��er��}b���(:�y�Cԛ3ʘ����t�i;�H�y�䞁,<���˜�\�*�:!�R"�yB	�t���Q�"��U�>i�`���y�%�u	<k�њ������D��y2�/'N�,rC Ս�&��Rh ��y��I6O��2���3}�e:3���y���7ܮ%���
5��(٢ �:�yҀ�j^��CP� ����=�y��`��aϾ�����&5D�p���70��d�68��-3@l5D�hj�藇:�%�Y�^��c7E<D�p�bF��\v���f�U3��L=D�L{b,ښ,h�
�'F}�)ju�=D�8f�66t�k� �[�4�91F;D���2��y�ұ� �U>4��#6D�Ъv]�K��Spd_�jt�27D�D�2�Ջ@(�1�?�ѐV�3D�x�1)�h�EJ�C�	��a�#:D�����6W��+"ݍi����%<D��3�IǢK1�\8�iO/� ��(9D���ᄝ�nM�A� �>�ꠘB�4D�ԋ�^W�����	Z����S�2D�3�N
h�N��`�K?v����2E3D�8��4�>���"ǖ{r-
�#1D��(��&Tg��9��ѿ7��(��.D����dE�xAK��6�zܠa*D��!!��DX�X3���8�T�r��5D�8sB�'A�$T�C�^�^sD3D�����ɣP��l�q��.���Z��1D�أ�hK�WX.3��D=D�� 	T�"D���a�v���y��^?Q��QBn5D��	�Kфej����Oe����$D���M�\�x`�R�(�j)�c#D�h����nn���e�!^��1Po2D�Tf�alHU{��+*.=��3D��I��3s(�ّ�E;7P	��.D���𤘋+	Rܱ�dB�y4F����.D�$1��Þ*��ذ��/�:��d�1D��{w@�C���� 1T�e!�5D��qnO�e��&� �Xc�'D���N�9Ʊ�P�S�<^�`���0D��١�.�R���]�~zu�WC*D�8����&OC�i�O۪|i@�o+D��x6��	"Q<�i���6�HA��c&D��&$%=T��Y����0��Q�3D���A�G�7k���*
2����!2D�`�І�F��XЂi_+���ڤ�'D��h��߅>����%�ڷ-{�)׏(D�� �I�F�"�S�]�xK�0��'��)@ �$*CI�&g�H�@��������rd"D�h[5鍽{�ޔ1f��<Fl�\���"�K� |sei=�H�(���n1(��q���$�ʅ��"O��� 6��Irp��H����oذ}g|Y����)��<�qN�xd-��/� w;��T�Mx�<��%A0��k5\6����U�<q���)���a�%3\O����#ˬE����F<�)�C�'�,���X/�L����fA�A�*W ~e 		�	� �y����:ij�l�6l4� ��OM�@����&�(��Ă$	B
d�^�13��0A��S�"OY��� ��!�f��()��Z�Qf��`�H_#��)��<� ��1��E�$�~5"(��G�<iW�^�x�<��w���e�����`��<�g,CzXr�`&J=\Op�z���i�C�?	X��q��' �U�r���!�� �C��"�����m0Bԓq-��y"BʒY�H
�k��b}�q����Oꤢ�� /����$Xk�@iU�4#2p�R �Y�!�X	�����L$T���ψ1(����Ѐ��*ږ��L�"~�|�����U P�j,$�@�ye�]�ȓ_Q��X3�ʀH��L˲(H2f�h�ITP7��Ű=�`���&����!ȝd���
ҥFX���5��	B�E&,���L1hQ��,�$�y��؟z3�]����3�����ą�y��,ݔ���'Q9#,��C��y"fɨQb�:ƂAA���p�dѥ�y�Nʊ��6�M6.P�@�K� �yԀ)��MΫ_�`�Wƌ�y�EM��J�ΑLHμ���A���'Iʴ���R�S�'9
�*�̜<?6�H�HD~�Є�"�R�ʔjR.��cA����FQ�o�m�ɱ�LE��Oq)�%ά0���Ɖp�IjdO�t�&B�ry�s�,�6d�!�#�Jg,���_���>�0@'6Z����i�NR��rA��wX����RM����R�h�Ԣ�=E 49�a�0u�i%�-D���ǤK
��[�	ξW!�PL*�S~!� "�Aؕ�M��B4�c?����t|�9Q�B�#x0X(��+D��dM>Q����F���~�᥎I���+۾Bjn諁H�[�vb?%�Odhk�a�0c��x�5
'd�HO^tЖ�&]�򙛣LA0m�SÁ�n�tQ���߸8�P q��<0l��I�� �ʀ�ߒW�(|`j�"F!��D�>&�lm�� ��D�J$1c��$/�=��"�Pn���Ԑ� |��\s<�󌅠>�f�34��k�(T	�%8�\ ��-����Y�L��:U�ܴ��D���%8t�	���%	��n_�T�t��-�S�r��B��!�D߄V��;�lK�(ؽȥ��/��!y�� �θ��`�	YTX���o��% � e^@U9�NE/,�^p��O�������y�<H�E�-�H��I[wZ�)��]�r�hR�̣i&t��Ռ�iq2��$�'3r��C��^����v��	aO�eb�'�;1)���2/����:�i��Ǻ:R��.8L��M���h��ǉ``�(��ďi߈i��.�|�h�o^��ZQ��N�-e�bL�a`֩
�ꥨ�'St: ����UA���d����V������^eo��za�W{Sv@�O=��]Y�F��|���w�N�x@Ư~a&މ|"�=���h�@�@$F�d�b}	�'�Y�]�և��QKz�+��gv��eˑE�I�fr���%�1��S�~����e
/���[q��*=�џ(��"�/��aҖ/�2|�������@cœj�>�����$�h5���|��]$�l1��I3+������<r:0�E囚g�\˓C��`L�j`��#u��j�|#}�K�P��u`�"^-vl41y�<q�H^4{H�r�)R=Fp�	��E���yy�G�)6�"�sTg_�)Xȭ'?�ԛb��)zc$���lڨ�`c�)7�Ћ")�kh�IW�#3��U��ʝ��=��!Vv� $S�e��P97#Q�F���	Y@��ݰ�O.OA���fw�3cF��y2�g>�3ǓQ�F���A	��y/�q�^u$_*1Ķ�X7-Y8��'�n��6l|�G��됇@��8�Ԧ�4,�Y)6��5�y���-b���y�m�.[�`�V+H�+B�B6l�����:PQ>�S�? 4i���2u�Y���S(~��M��"OHI넀�) <)��,P8.�>4�4L|�R	� ��ă�|��qArخ��r�z�"ܷ.q�C��c�X]�� ւA4���	��y�ꝌG�P���/?k@�ywa���'"����N�P�t$��Ӿɪ񙗨�f`�8P �I�C�I-+�.���O+Q�paF�5N��͊m�X����*O:�K��Y�TA5b¨]�s�Eܹ[� ��!/D�Ќ׀TZ]A���1�lӘ�2��@(,$��J!�'���5S!`Z@ڥ�9$���
ߓ\_T�S��^-(�
6�M�cOZl+f�4t	���� X�Be!�d�t[�����P�S��[ i�O�m; aL(�R����0�`�F�uY�2��2o!�ċ�ٰ��jVH��C뙉'�̋��J�b��OL�}��9�xd��M�હ���,�� ��$B�䓼r��K�F�MB��ϓ|B6����>��=�B�CJ��yI���N%fmb���C8����Ʌ�F�d]��Z���n�=Є�G��,2�!��=w�A��@��!Su�ǅj�!����ad�@�G�T��b���!�Ę�}`^��ŝ�D�{G�~�!��L�cU8a��O㪬�T@D��!�""�I2bo�7٪L�m��\�!�F!L|ꅩJT�i�aPSU#|�!�DN�!].@V������Y�K�>X����VP�0��\��@Ӗ]3�0�$stم�0o�*����̟��gJl��%냯K�l���Ǐ,D�P��/����$q�M���4��O q)`�ϒ�~�eϡR����G��A�O�B�QG�j�)�)��n<Q��"OHi�dI�0�$0�%gG�e0��7�O�@i@sJ�Yw~�Q�'Q��Pb��h��Sq�{�+
�TXђ�,ON�����`�*z��05	�`�E�5,�M
pj�aB�$	 �&�?I�Y��N�)v�/lO~ęU�(d�#��	/s��a[��r@��\�����ȍ=���0�����)�Ŏ^3j���[wb����s�,"�
4v(h�'۸��@k��`pC��P6z\6AX��
�.���F�U]}��eaנ��+C�|J��y[8Yp�w?ęz�^!6F)ф�v�p�(ӓ��`R�*f���A�U1~�~m�b�Q;��QwkI(�q��ו)n��î�p�����'{�nu�Bf�
>���<a�c��98������i���Aov�h���/Q��P���N;O�!�֌@
�Q3���*Bl]���J27زP�s�^+-`M���x��8K���$?��]�
�8�hy5�?ZA�b%��pf�8�S��M��ȂX�<Q N�Gx��r�����
R��h�g/>k��,<�y��E��CL^�1�
O�%��HD�RV� J��J:�L� o�m�T�J��ȠO��{A��#���ʖ�ĬQT���z?�o��A(~K��M��8:�F8��l��F.,O��IԨ��v6��48�]�ʲ�����[��0�$k�K�S!�K�I��= Q�Mcy2�E�+�8�� �a�~����V03�@���oFwVO���e	�<����4k��=�e,��R�:�q��t��}q��n��
���S5Z�j�@��S�\��e���I$�'^:h*��A� \t��#�Kuh�� �B'`i��@�z=�ԉ4�W��h�0�ӼYa�ѻjP�6��m��_��ć1�A�fAV5���u�B-v�ب�E�$b4Pc|��b@g�z[I+���V4��'���S�*�t�@SN��*]3u.�9@Z���:-I�Jܶ��V=9l �$�Kc���!!M1Λf�G�	��� Hg�ӧ������o#�#d�����R�@������z����0|J��ǺC�l����}�̭+���^}r���7����4.Qx����S�}��9"�)��;�M0��P�{�qO$�p��@	���S���\J�@�{� %��i�`�B�	't�`	T���qKʘbC����">)��N-�ȣ|T�<(��S&/��?hpP�,RP�<����7 ���)��w������E�<�e1)�2�+�$S�R�١�%�}�<�a��F��KvC�K2�a2��}�<��JC����j��MG�%��a�b�<���Y�FE6��dɚP�P�
Z�<��k�$��$C�ޛ0��@e�P�<��8y��@�<��UX�+Q�<� �10W�'%jl����ш,Z�`�"O�"�S2�|�2�S�6� �i�"Oޠ���n0��a�T/��Aiu"O�����ОMU�-�BgM �X	�C"O���nV�>�y�#HA�,��"OpP��İ*:�X��S�1�65!!"O�#AF�1vq��"�����"O��J�DL�ð��ʆ��I��"O�\Ba���B`Bn �?�luӴ*Od�Kg�[��=���27�8�	�'��]�df�/;Y �*F�%�"��	�'�EG�D�i����/,l��@�'Ǟ)Q�(���L��ō"e�f�#
�'mx /�fz.��@�>^�0�p�'�
�p/4
��p�G\!y>�8	�'��i��W�� ��g���49ڽ��'0f�	.$r)L��e>Y����'�(���fϨ��i�Dȣ;���'��ar@Z�,� ���5ː`��'�t�����]�T(�A�.[w�Mp	�'��,	��R-Zwba1�W_����'�j%0�ƈ�3R@� O�W����'à����/�8�d�E)�)��'u�x��"ε��*P
M�:"��'m$�Z�Yuj�R��F�2�6���'����cH�,���fX2%$ٺ�'�6T37Jͦi4"Թ��(:f�'�~-���$(�F��$C U�&���':a[�$��n���\ �����'�~i�e�֓M���1허)����'��k��>E|�a�`���_�4��'@ �*�͂c��tBӥ֟C]��a�'����`��7���z��;�8I�'�L�鷈:w�ā��$֪S���
�'4���V�^<�%� �I3��˲#)i:��Ë�1-����|Oȝҁ@�Up,M����<u?�]��e'
�y�헰+�����������L���fɊ�ohy��,�D5��ȓ<�p0C7HY�{@�T�Hr@�ȓP��%��^� ���F�e����M�����G3V%�-�"NQ��b|�ȓ*T�ƭP���ӧ�	����<�ÇGI���O���J�)V�@Er�Dd��
&��'�`7��؍�'���B^w� �3?�')�d�$�4J�f<���V\���kFA��E�,OrE���O=L��W%]�,(�hT�g�B1B��T�|T�	U���(1��	�fǓ0��	�M�d�8 ���@}rh�6i@!�֡@���	Ll�OE�Ub�H��%v�u��h^B�HSd�V���Rr�7��%���O�?�yPƋ4%�А�œN�	�1Ad�L[�@I�A\8�'���	ׂl}@��"l�,xԜY�)�ZQr)��'�,Ô���Mx^Ԃ
ç)�R��G��jѨw,S�R�x��Ż�~B�=c�P����+����O� J��p��cyp%%�����8=|E�X^M%�����۞r��d9�����d��K�UD��!7(�<a�kFy��IZ�a�J����w
L����تΦ����,��	�'�8<'?-8I~�6#�20eb� �q�$�6"
�h2И�0#�V�m�;a"��}n:�+	�{Q��B���=�4��/O�V������������|xX���S�{��@�b�*wU�  BF� @�h���OV��'@�2S�W�?����j�|_�<еJ�xg(%�@K}"��.U[��3S	I%���Z �\ �+ZGjX 5l�	C�D�$�����x�f�E�~�>q(7���>sPF]JY�@��`��S�p�^3�ݠ��Tb�ѩ��\:�!�$-]��J�O 7.5ry@p��
%�!��/1�X��AӑL��(c�'�;e�!� 
g"�9��L�S�Z���O�i�!�d�>.(*yJR(�8φ(K#��2!�� ��S0��?iT���J��p��E��"O�)pE�ڸ��q
���7����"O��!���o�T�ZB���8k"O>�`%o��%���($���mrX��"O�I��ŨN�@"q��M���ɐ"O�h��K��P���	��=A���"O�;��Έ@r�� ���0/2F"O�%�`����	�b�:"W�c�!�ٳBl⸒7/��>i�	�v�ͧN�!�_�S��`��-4hf��nE	2�!��4d!�Հ�m���P�L�!�FY�<=�;U6����"�!���I#���'��I�pxQ�B�[�!�P�R��A{U@V�H�P�����&&�!�dUz�>�o"Z�&H� ��!�DX%=��b��&Z܈c�.Sk�!��-_$*w[�byI��"!�=~�,���@e>NEZ$��'p!�^�@�Z�0��L����-z!��2�`�"�F�SH�!#g�<r!��3WO��j���a>��B#&�:gp!��w`�t%R=r{7JB-S!�*W�|{���-�T���F!�%)�����_�m{�@�fA�$)!���{���;rT$d ����>Yj!򤌆@�T�3b����E���]K!��[�R��!S o�w���(r��y�!��-?���J>|���T%�?F�!�d�.���g#R�tx�U	��aK!�D��_a(��ԁ̏P�ĹQ)B�#F!�כ[� �k��(��	1����m�!�D����4#P ��0Z� T�A"[�!�W�y��q����O�@�	㉈�!�L:o�.Q�q��6�D9� ND �!��0-PZ���ʅ
����Т�!�ĕ�GjLfB�Ut��qɅ�!�$=xޑ�a�: �r��6)���!�d�&@E��
Ԣ�F*h��P탄b�!�D�>|�t��$�Ux��<�!�d�F������'���ǂ���!�$)3��c��-Y4Re)G�N�/�!�]%o����ʰ*w6h`�R�y�!�$�?����ӛjZl}��`	J�!��͒Lŋ�̃{���@" ��8.!��LJV�P�b*��e��rr�̇%!�DÁZBJݲ�	�r���3��|�!�o���`$Z�t�0#� �!��4E@0�#���4#�aD�!�
'��4��([c`��+VN�a!򄛙R�&�3&�8nC�11�lS6rP!��VG;Pp��M�P*Z}��J1%�!��Ǟx	�B�3��*�jѵF�!�D[>Y��ģ���0FըQ��O�!�dNcs�HA`��� ���*�!�d %-���1&a  �0�RW��*U�!�Z�4�& ��LSX���g�<q�!�d:9<�5q��4v��y��Z?\�!�č��b{�M��	�R��фW%�!���}P� �`߇�4M(���G!򄀃=F$`%FP�d�8����ZIV!�A��� Ʈw�y �\%SS!�$������-�-a��7L����R�5�r�!mڹ�lI��y��֬P��D�!��}ɦ�9&ڗ�y
� �D�g�ʁgF` ���!j.�#�"O����Z�<M��$�UW��Y�"O�a����"'K� �C�<o6pI��"Of8{�C�>�j&�<`%pE�7"Oj��b�Ēx{�HE�]�5�Ekc"O�)���\&0�@8����2�`"Oz���ߋ�2��v��	� �r"O:����
)��|Z�#	Q�ؘU"O��q��#ҭ��E%Җh�2"O,���/�`����#�+)$ʬ�C"O���D� �TK���d`p�"O�)sW)��Z��#\K�l�"Oʴ�P�&�>�I��k�`���"OΉ+��ԇX���X�^]�~@BW"O��D�ϯU�����KW3v�� ¡"O����n7����٢#��	b&"Or`z _�
�xE�s��r��a"O���&-L���A��_1R%09"Ob<�'gq�0&j�1��I��"O5�$�B�E]�e*ѹK�}��"O&�xD
N�0i5d�xS��i�"Op�P"i_�1��0��P�'<L�5"OJ��t�V�H�� �%[��§"O�|ђi�"rHhׇ��pҐX�"Oа��C�$���ǔ$��u�0"O<���gÈP����2&�-�x�W"O����
�HO�Ar��W
)��iB"O*���ܧ|X��{��Ü)�X��"O��R%́�#��cg-��#�V�iD"O��qv��B�Ѻ�픛"�d�S"O
d�d&�6��X�M�d.�qW"O5rc�7>l5!���Ѵ(�"OH Z� ˕)��`+2%��[�t�"O��`��8��ph�a�z�Q
d"O������(���OR����"O*��uAH8^�~9��d	�\�R�"ON�"(�;��	t)�._�,5�"Oެ���3�j��'y�.�C3"O|��n�r~���`��;m`Z�@�"OB�+pD�>ڌh9�k^�r�z�""OD�[�N�7'��y��a�t�"O��*���k���U�/b	I6"OȰ!�f�,J�COQ_���V"ONI�S�ޟSs ����g��%"O8���K�{�������|�� �"O0TZ��H�sm����K����"O�%���()���F� 9�(d	P"Or(���f��]��Z�7�P�q"ON`��c�d�YC�k���*V"O]���H$"#j$��l�E�z"O8���ӎ{���I!0�d�a1"O�l�kȗcGb����kYr�qC"O֥�U"���Ait�X?�ũ�"O��{��ѯ2�@,	��̵P�0�"O�;���a�U�� ԛ=A� A@"O$XV�v�� 7�1|���	�"O�`�ǟvg�t�U �V��e1�"O������4C�,��(Ȱ	5�u��"O���#�X�{�����@�&y�D��"Oy#畑 ���'�D� \{ "O.Q�C�Q3
�� �wE�]1֕��"O�9 D_�"����]5x����"On\�g���p�L��N
��"O�FI
�phQ���
Ҥ��4"O� l!pa��	�d ����/��9�"O>�"�[:J�0�"��s��A�"Ox 4
�:|��1uDFb"O8�1�˞I���&��d�)�"O�n�*��Dh3I�����OժD�!��Ƞ@:ݙ�l�j���0��!��Je4���J55�Bu��D�!�ć�?Qr,�g��*�	`d�!�D��V�@кA��"*�j��D�!�dD���1,�!�F��UÁ�_�!�{G��6AN�/^Xj�!�H�!����@�Bd"\�f)`���4�!��V�j��M��-��`p�E/�!�$�L�Pq��C���=;�D�F�!�d��Y� ���
-'��I���P'Oޡ�d�$5�
�p��:}J�`Z�A��y��� i��S��O�]k��i Lӊ�y�Cݽ|#�K�,C�H�ɛ��V0�y(C�nhct䔤R�tH!d��)�y��]1�̀a�ڟ���
����y�%����9�ԥu����D �yb��r�ŋ�'o(D�5��-�y"'S���p�sJ|H���d7�yB�NFP��e�)<m��(�	�yRlZ�r�B6E���!�ϵ��4��'���@eD�1=�A+&Ɛ+lX���'�4��̗�xO޸be'�	r���'�^�J�V�9�rk�/�+�:Uq�'���QmѢG] �td�3
z��'�*B�@"�@�3JC%����'w���fȀP2<�B�+U��(�r�'t�����W�������Y��)q
�'^u;fE�9}�0�K"A�����'��	�n�?w����B��<C,�J�'����a�Т�F�5����'3���@�1��`"6��,&e4p��'��ԁ�Ɍh U��X3�Xx1�'ǾMA&���S�X!*����h
�'֌����+U8Ȑ�tO(u \0
�'�����.Km�D0�	^<t�X�	�'Bh%7��w�pT��9 �D��'p"����X&���#]&Q�;	�':�`E��q�<P6��C�
�
�'Ѹu`Qfխ	e�l��4�\�	�'a�})΄1l��A���W���\�	�'ox9��j�T|ma�\�_���'�x,���	
 W���b�� Pm��'J���e杹��,bả�f��i�'$�����6^����C&'���R�'{�E�biB�{�0��#���P�
�'�B\��c�%#� ujG�H4���@
�'�Ι*�@Z+L%�D!��-#�JiB	�'�xe����b�~l��-ƍ!�P��'"����L�e�h��2l�
eI�':Z��aش"*���e��j	�'l�idA�O���A�0$�i��'��4�P�	��+�F�#@*�@�'�D���Kj�^�"��Dh5��a�'JhH����L�Re[W⑴p����'Lb�"�	qF�]����#��Gy�<aw�'\��UrU'\-p���AFPt�<� ]�L��@��E���m�<�4��0�6i��[0ޘ��#�	f�<�2�����dE��)Nq��hM�<�+w�   �   �  ,  �  �  ,*  u1  	8  "?  eE  �K  �Q  /X  r^  �d  k  _q  �w  ~  W�  ��  ې  �  c�  ��  �  '�  ��  /�  ��  [�  �  J�  ��  A�  ��  ��  ��   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C�>����鞿6�!d��x�^��I��~�!��
�l����v���:�9a��:uZ!�L�,Ƞ�#g��UԀ�e��t�!��v.qc�ʁA�P{U�C-h�!�DD�x>B��cG;c�lK�,��"�ayR�	� Q2���F��u�t��� �/��C�I�Ld֘8����D��T�U�#�fO��=�~bh(e������M?��m���Tg�<� �������T�����R�g��dR"O���ѣi�A	�͖<|l��"O�ȁ�N��SO��µ'�#{u�L�"Oҕ�sGY�>u�0@�'B>]ԕ�b�'I�O 5j����)ɲV�л�"O"}��J]�P#JLa�׊R�Q�֓|��S���O��Ḡ/��l"�88�n�:!�D�	�'X���P��u�҅� D�l7�<��'{���6f-虡4��	.�<�R�'L�Q8�C d� ��욯zA��'a�l�3�F!C����4},0|ϓ�O�4 6g�'���z�h�!�P�R�"O�$Kue��Vrl��MΈӲX�S"O�!X$�ZD��z%��B����C"O:0���b�V�a@���VĪH��I8�\��׆pT����Y)i3	=D�$�&���;�#!a��9��H7D�|��BP���x� 脖~g�T�#5D�H��
�Kh��Fo�Z�s#�'D��)F�^��$H�/ǐ'��(#D�8�\�.V>���bYO�9�4m%D��3"�Pq�f�2P.p���(B��$K
~%x�b1Fb�la�CN�.��C䉮T��[#A�$I����(��AC�C��H�XtN)qH�!!��A��C�IHh,����s�6C K�R�jB�	����#塕��Z����}�B�ɥ~�� 2
?<�[�"��nZ�B�I)&�ĝ[uj	�%��a��;�hC�	�f�-� ���=��d�E۸a� B��;}�܉�e�1(��1��ġ=JB�I�!�\3�oԾ�p��C2h�C�	FxXz�g��dp�Հ	c�C䉇>�6���a9yVa�W�vdlC�	�!2,ҧ�?U�*�����5�0C� XwZp''�q�1c̀�ThfB�I(wM��+����k�I�@�ӽ	LB䉆���F^�=*Q�@GB�	�4�ܵ�!�� (Yv	`s��7�B�	?s�r��d����hj��I(8�C�	�g��d,�(M>�h�h��q��C�	�TTx�5��<�� ��&��C䉿[.� �� �a�P��/ԌV�tC�	3F�!wFY�b �'NV��C�	>=F�m�FǵxZ8U�ց�	tLC�ɦ:�p�n[�u�ҴY�!ӣd�BC�+;���U&�<b��T�@�����C�	<+A����Ǜ �R�I�.ݻs�C䉂Ԫc��T/T.nL���ܴS�B�	->�N�9�N��T]@xËZ�a��B�I�E�Ĭ1� ̮j��� A��'�B�I8[�2�r ͫ���TP�]`tB�$�0C$�!O�偷ƛpuNB��]EdP�o�4'��m
D�ُ9.2B�4$�t(*d�8X�}cRd�+DB䉷L�T���k�2n�i�CE�[SB�ISQji��6��{@��/'�C�	�sϴ�;u
�?�X�:b
��~/�C�I�F!*t��N�:�0�h�-	NzB��<�C��3}"%���CW@B��&`H�ܸ�Ζ)��p��+� .fC�	'�n�x�$t���2�I8�^C䉟2�F�@�╧Nt��q�ŪXtB�I15D�"� 0h},�H���yA�B�)� ��aF�H=�`z�aN�'b��v*O��xc���2�~�0����}��'���� 0����
Wl��*
�'��ԁH>pxcG�o�����'\za�2mF�3��H��ˀ%o�����?)��?����?���?���?Q�=�q���-xpB�ѧ�B�j��9��?i���?���?9��?a���?i�vD�U����;�Pĥ��?P����?A���?���?���?���?q��S�x�+��� &�h	���#OVlI���?���?���?���?���?��j�$X�գ���l�o�d����?a���?���?����?A���?��(b���[tu��+�B�h�J�2��?���?����?���?����?a�I$>�K�m�����Bl����?��?	��?���?i��?��,�lyGm�1��x����n��,���?��?���?���?����?��g�x˷EǂP�C���'�
�C��?����?I���?���?���?�7ⴹW)>��
A�������?	��?����?i��?����?��s��A�N &)*�n_�a ��0��?��?1���?I���?����?a����*��)[�|��� ��r�J��?Y��?���?���?y���?Q�z�(��P��
^CB�ve��A�Z)[��?	���?1��?)��?�c�iC��'�:�i�ƩQ+x��r-dԙt��<A�����0�4)�f����s�P�p��&�:�S�C{~��nӘ��s����9��S�Z�A�u�_�ƚ-��՟�R�(����'Z�	P�?�����uc2&MD+0�ѯs�du�����Of��h�d�Uk�19�A�v�R�q�2�a�����#1!#��L�'Ad��w1���G�[	7��%�ECN��xM9�'$�?O��S�')����4�yR���B�@T@��)T����pM��y�9O�����ў�ş�%�dȌ��#QV5���%`�L�'�'67��-�1O�0�vg��k��Lץ
�ؑ��/�����d�O���u���'|��Gw��Ȃu B�}{�O4�DK�1
>	���I.�?��H�O\�p�n߲iM�:Q�F�Bc�m ��<Y(O���s���$ޑ6��$ѳMyE��uOv�`�ٴX�t-�'f�7-+�i>�ꖉ Q2�8��Q�'�a���o� ��ß@�	�ED�n�q~�=�,��&c�<hJ��~KL,�&ş)���#�|V����p��џ�	џ�Rp�N
W,
��IV�LH*3��oy�u�mIB��Ot���O̓��d^��%D�8Gr��i���Hb�Ʃ<����M��'L�>���O�;5($s �� �h��MM�Kx�S� �>��@jhy`�ьO�ؖ'c(`�C� ��,��D�	H��'/��'�����S��ݴ`� 	�@F��	�/􁻂�D3`.d	�Z�����g}r�i� 	l��tK#�^�p� �G7Y~���D�Uo��m�^~�닥�ܠ��w�'ojk�3=� !e��!'2<)�+�T���O����O���O��$9��b�.Iy�$:?F ���>/�(���՟���9�M�$)Y���dNߦ�'����M��d�di6�ώBb�(CUFN:�ēM���Fu��	]YD�6�7?!g����(� 
����s���?�Jx�$��E�F�$������4���$�OX�$R)�e�5ᛧaU�l�FnUd�$�O�˓Z>��.M�\��'erZ>�05#�+$�����LDA�=�l)?�_���4 ��v
&�?]SGKE!F�:�tB��@¸��4u T0h�I3���|��`�ONd9L>9����IF��Q.2�Ψg�ކ�?a���?����?�|"*O�$o��Zm�U��h�r����L_!h��I�������I��Mc��B�<�4w���E픧��=9� S{$��sǿi��7mC0H+�7�??Ae힧����3��[�j�x���,Ү��qe\
�y�P�L��ܟ���˟(����ܕOΰ5���m��eg��$��XXmq�(x��-�O��d�O����dD٦睈B]�a���q#~-�
ӈh%ډ�	��
O<�|z��0�Ms�'�ص 7���NcHLp���A#��؟'��)�4Ǆş�$�|rW��S��k���FTn��"��6%�Rw�\�������	hy2�{�T�*�OF���O��.���P�C��Ii�r�Э8�����D�O�7��]�'e�:D�P�1R���i�d�	ǟ$#����2U#B|~��O2P��	�x���0'��(e�(ј	h4&ז�"�' �'E�����"�!�3����^�qo6`x3�C���4.G~�S.OBl�l�Ӽ#����Is�y	V�A<e�L��E�]�<���?��i0�a�ia�$�O���WJ���!*�v'z���n�4���2#�F�RUp�O���|����?����?����>4��D�5����LN2,.� )O�o��+�m��ȟ���X�Sȟ��G/�-?�н�d��Y�b�*�(C����I妹��4Sg�����O���H�3U8�UY�� Q�YggI*Ly EY��d�*\�n����*h��Of�(2��2�K�4�X�d��蚘���?	���?���|�+OzUm�
INL�ɺ/?� IRa�8:x(�cC+��H��	6�M#�2$�>��?׵i�\��R�*1ՎQ�G�N��Q3#7��:O`�d>Bf�Z��Vb�	�?��=� vmS��A%1TCV:l5t0s�4O���O6�D�O$���OZ�?ᘡ�.n�Ȉ�ɇ8�Z�#"��Ny��'_F6��+5�)�Or nW�	&P(vă����j�*@M<	���?�'hҰaش��d(<	��E�ϢiR�|
��G{J�#�C*�?�&�,�d�<ͧ�?a��?�U�O�"ߘ8{V�5i���Y�	�?!����������ٟ��I�� �Oh�I���.�J�*��6�&��Oܘ�'R�i��O�S'Y��YA`�<1B,�!!���t�Dy�eo�()ں�s�:?ͧZP��DH���bd��q!�M��1��ɮ�	���?i��?y�Ş��d�ͦ5q���$u��j���v_����+^5A�X��'��7�>�	���pӄ�b��;L��6ʍ[=���EOH��P�4*;r�4��$��X;~���'��5��]�5ɂC�5{��W"���Iuy��'�R�'���'��[>uP�Ɠ�e���QBOϫ�j���gۀ�M�Q�?a���?�H~j�v}��w�"𠱩�
,��(�EC�g�ԵSv�b�v�l��<ɪO1�0�1�}��ɡv�j����W�Jq�偄�qUd�	�js~q��'6H�&�����')n���J�X�����V.TEK��'��'m�Q��"�4h`Bs��?���'�N BT�O9z�*q��@V���i�B&�>Au�i��7�WC�ɤi��9:R�II!b��2
F���*�#ϟ�t�D�|�c��O�D��0��#�d@(5�pBvI�(]�
�c��?1��?���h���$Λ<�f��S�[�8s�Ao҉H���Ϧ�P�B��D��:�Mk��w�t�d��3[˸p�WlI��`�'F�6m�צ5�4}��`�ܴ��Y L�6 ��z�v-c���m��!�@�~���cB7�Ľ<ͧ�?a���?9��?���1]lM)eeA�S3���r�U���dW��M"q�ןX�	ڟ�&?�I2de<��4�E_@�y���إ
��IY.O~�Dr�>]$���[�Ş_4�ځ��o�(M�wӄ#��!���\����B��f�	cy�
�nH����K$t��Y@��f���'zR�'��OL�ɪ�?AE����@g�ż'�� Y��'g�@H  ϟ�a�4��'����?���fk�QθZ�K[vhrYyA-V�2�h��iH��e�X����O�q�d�N�& S�b�ײ�0�����Z>��O&�d�O����OP�d1��R�L0B��7�^	���->t2��'$�ix������?�j�4��7����N�.6�6�`F���\0�x��'��O �Ҥ�i��I	T�{��&L&�`��ǌo�� �p�ؿvn2"Lf�	y�Ob�'�Ɍ�J�4�A()8[P�ԗ���')�ɮ�M{����?A��?9-���(��Ģ|.��S�D�	���8ѐ���/Ot�$g�\$&�ʧ�"�c�X�n-�HA��:G�2�#��D�$�N���"}~�OT��I#z(�'���3V��VT�[r�ϊsjV��V�'sR�'�����O��	��M�1%KmȾ� #Z/��
�!��zF���.OT�l�`��/�Iݟ�w��	[��ٛ!ǆ�}�\E
\🸠�43�pڴ����H��Ÿ����+Z>�$��2�r�U�1�D�	my2�'���'���'��X>�WDF3Ӕ$��,%s@]A����MK����?���?�K~�F!��w�h9c�[	T�V��W!�_wZ����'�2)%��)��+��6k�� ���M�p�!�'аC��б�$r�����#|B�H]�\y�O��Dؼ�p���f��سQ�Y�4��'���'3剸�M���I��?���?�sd��l<dK�C��L�2`C�����'��ꓬ?I��H��'V�Hq*��Z�,ʳ��)+:(	(�O4�ٖ��(J P:`�IN��?`��OF)x$$�3���Ԥ�<�l�`&��O����O*�D�O6�}:��4&Te*��4k�t��0FS!{GR�(��K��f�ɸB�'�J6m3�i޵����u;����$þ���i�j��������;ش�R1޴����(oȤ�'|�8��6?��H���9$i��*v�7���<ͧ�?���?���?���=|&�u�aE�L��%9uFY����Ӧ�1
	�,�	���'?牝T�d-��!V1b(�3���>�P�S�O:�mZ1�M��x��t���k�$	׆��l?�0Y%ˀ��T�aH����Q0�����!"ؒO��.Ɋpk�@��#J�����|���H���?����?��|�/O�oq@v|�I�E
j�!�J�� �VA��ɺ�M3���>����?���i'H����?U�zh!π�(�S2aWd������lA�S!������ld�Beǡ�썣+��H�B4Ot���Op���O�d�O��?���E�`�8����U�3
d��b�Gϟl�I�d�ٴfy ��'�?��i[�'&黳��-������
�i2O�W웦�q��\|6�+?q�ȆD�ШB���3#7�#�윀r���H�O�9;J>�-O��O��d�OĽ `�����)��� ��E�g��OJ�ĩ<�'�i���<��柠�Oz��(�	�H�Ĥ� d�zX��O���'k|6MS��i�S��du�|B�I�Z��"�F6Q��	V'uSB�RS_!��4�P����ָ'?2�h��M�8�h�A�.x��	�'�^Dt�/ƺڂ� ?tI�	�S�~�-Дh"q�A��Q=�P
�e��5<��@�쟃�С��B�ncn���@NR�iX@���HvgĐd<��6错;� Q3�O�R�\� ��e��oP�yh�͹pT<"�̟E�V�Q�'��0��̛���4/���H�B ��A!"��*��Ap�,�8���f��[���,o��kf"O��g�F8�(0_XeX��S���pT&I�c��'v��f�7��ݫd�L�y �E8F�F��q�Ȳ ��k�� ��D�F�[�|��`�`�����N"r��4���Ŭ<a>�F��e�A�!��F|-�FDN&aI?:<z8H!E�bXlaH���-H(5*��.$���%"�K$�� �c�O\uP��� >�6q"D�K�9C6�9Å�O��d�O�,�@:Jy�nW���y[�IG��������X��#E�k���Jg��)�(O�<s��*�� �	�Y�"+$�r���T<E ���9P��a�'Ot�'r�D����?�O~����t�z�c^���´c�:��$K�����?E��'��	�-��`8��`��,�>`����'�'�����
Roâ:�&����O���D��P䊦o�m�R Y`+'4!��թ	<��!�1Bz<�ꡨǽ4!�C&��A��;W Q�pHߋz�!�$�2��|�Df��| ��J�AH�Z�!�d9�Z=K���bg��%��br!�$g��e��m�� L�9�4BƃXh!�$Y�f�T-�5���B�XZt�@�y�!��i���`1�Q�T��
C���,y!�T�{V��%/���P]PP��H!�D�7Ul�@���h����Lև!!�䕘6��B��Q�چс�AJ�r�!��4 Vl�$J(P�x;6�)=�!�ě�a�H�8P�%�9��$�x?!�d�/&�b�F���l��S7@�!��+ێ�(�NA�+"*Q�� �2r�!�d�Q��"U#H�a:(PoZ:9!�$D6~=�UJE�N% Q��՟;!�6NS*���	� �'�n�!�$T�r�p�ra@A���u�<&!�DQ�.o
��'�Z#'���׉�2�!��� �@��A
B9��-Q��|�!�$D<��y	d"F�b�^1"�m՘x�!򤃪q54����YXX��l��r!�ĝ�[�6��GBY��{�K b!�DZ%�X��_�8�x@�%��uK!���*N����(����cӶ28!�"z��Lyˎ��jd��O�_L!��?-h�D� [5G���V!�䃠��(z�SN
}S�f)R!�ď�{��S�'߳7J���Q�T M!�&>�$����
n*�U��O[d!��s�<�)��?t�l�ir��RL!�){z���n�;u�>��Z~�!�$M�17[Q��E��yұ�л�!��g�A��{��I�V�z 衇ȓL��air�O�E���Ƃ�4`�괆ȓJ=�!�*w�x)�JB�d��"O��bR!JZ��݁B%��g}t�KT"Ov����&��)���)���z�"Oh�wM�0�p!��u���(r"OL!	R@>R��a��f١��R�"OvL�7K�e0�����ߘXՊ�s�"O��%� =hV��U�nӪ�2�"O�}x���ј�cW�W�N�V��$"OR�ă��3`ٰ��W�N]�a"O�Ps��ϻT
�#
6`��m�V"O:ԃ0-� &���cJ���[�"Obm��a������#��BGJ�k4!�D��N;��h���)eF��b�>!�d�#"^ �B�B�B �͠���EG!�l���k��W�H̢I�'d�>?!�D��Ji`��Q\�,�QB�?.�!��C7'�8.)v`m�7IM6 ������ i!C$µu�p�n�30���"O��A�a[�F,,l�-C&�nyx"OB�0d��2HL�x3���eې�"O&M f�G0
8���.I�bl�q"O�xcGE�X$A��+�|�"O�ѣ�FG����Q�N-SC�q�"O�B"��@=�H!W#�+vEp"O~���X61���g_�"l��T"O�8I2�й_Z ���'˥����"O��Zu�h�挠��� LN-J"O:��чѧD�9�4i�#7�t��g"O>��C	}_26'Y�<%R�94"O��B��������ܪR��A�"OL���"�=p',ac�Ϗw.c�"O��!��8M�H��/#����"OR,ٗ�qIr��:E~0U��"O�+��"���bg�'5{�LJ�"O����n�S��qq�JE�MD��T"O��
'� 
�Xx)C%'�UI�"O�p���*3`�9Վ��.�Pl��"OD8���܇pI�`9�&��T��*�"O��Y�,���N��e/�g"O�yg"�/v�$�H�#]�*,d��"O|��p�Z�1!i�R��A>�y�"O(	榓�]3&�+rb82�"O��sVk� j�M��K^�K�j��u"O��!��r'��:3Ii����"O���Ǘz�A��s�^(�"O����o"*469 G�HXŪ��C"Oĭj�DI+!����'+�=�S"O���0��zڂ�Y��Y`�y"O�!���>^��)UD�_\]P�"Ob]��HV�+�\y�RC�]�։)"O
�fE$ }B�Ŧe���"�"O���5�V�?�,����Xئ�	 "O��2��������#��9��"O$)ht+�0Vs!���'=���A"OVy@oϦb$ ����A���"O�E�N�`� BfݿK�zE �"OP�A�'8Z�����	�$;PLB�"Oބ2��ԌPW�p8������"O��� �]�%�X�* (V!�@��D"OLb׹�V�ز@��*_�P��t�<A%���}{�ms����"i�4�]G�<9�/�2q���K_=b)x �fQo�<1�4a����ڒ!|�4��Q�<�LT�P,h�!bU�P�:�[��q�<	�	.XP�S��ňb�y�"��q�<a��ݒr�&)X��
�d��f�[l�<�I�7 :fa�k�8���ʑA�<���6N��Q�g��V}�`�+�{}�Rx��	���)a��FF�_�����%8�O������<�N�LѤ0�&mj+1�o�<qS�D�;	�-�DI�D@h(0�KZC�'�rHi�0�k�uc2�1*=
��� �2���O�����G��d$}�ek�.����N�i��O?�ɝDB%�� I(�:X�R�2"�JC�r�($K����
�2#/�0J�$��I�D;�@��$��#��lx��b�ߣRt�Ň�&v<�p���A	��$�\4 ���O���b�(@)*�!�92A�Ѹ'�J�D>�Hr�'IH��'��Ip�/Y!*��E��Oƃ��<ȶC �@=��D\��yr˔;1l`5��D�zH���jS�W7L��&�ņR/>�ZmE#)�M-F��é��9�����S�? ���Q��
/3j80�(�7 rg�i�JX�mV-ǰ>���(�$ً��:O���x�@K؞�Q�aǵR/p ��$��z����Dd~)b����w/v���S����c
�(�b��iH8EDx�	׃H&�����T�9�lyU �4;Sn�b��E�T!�䄑(�� ���L�H��+�l�N��b�/ �' �>���8�pv��~��(�c��*Z�zB�ɜ+~J���Ϩ]�]�Q��(BP6�_�`zZ��R�lCP`\2H�8���I@��%q�$?lO"1K ��d���~h}�1��0��q����7�^��ȓ�$�s��JzX)� -2B���?�AN�Z��H��I֜4�ԑ7'Z�M��L!�Cě�!�d�%/ND�,�$�l��C������թH��b�"~nZ��ҴB6��a�
	+�n�vC�	��`��=%^� ��j�L�@��+��'��xb��U6W�B�`��IM��u1�D\�d0OD���64����*5���r"O�-��/�;l�����!4�)��	�dm���):>@\�a�܄0��IBᏑOb!���u�<�&��?A���z��׬]�����p�=E��4�p�C�\H�I:��N:;�&��s/�x�ph	�K�E�G@]�#�U�'��[D!��=�0�ӗ:=zr�- ;���c�JX������u��6m�p�\��E.k~X��K��^�!��,&I<tXf뚾H��@�d�Iq��H�Ee�D��>���!��Rq�TKc��D�e�*D�<�U�76���ӵ�!.l�`a��tӪ���
LK�S��MKCE�4cBᲖ�l��)Q�Cg�<��Ы-�E #�^�^	�`�g�WN}r$(a6���d��U2QТM�8X@=z���)~4a}��3<��I.���e�Q� ����G;6B�<3ꜰ0&EG	:�i{�Oq�"=�!L�)�?�"�D�.@1C[�t֒��<D��I��J�5�<��Z�G�8T�C�d�4\����w�S��Ms�F	����B�_.Q�Xm���[�<I���-Sr��{ �. ��f�Uy2��p>yA�\�V<��KթH'9bA`D�PN�<iDh�c���#��L0lJ�UN�<A�nX�����*	(�}���J�<yG���'Lx�D�E|�lp@�_E�<�5bz����!b��{�����[�<����m�V)*hj(�S��S�<�Qn��6����'ԦN��Kf��L�<y�Ē�7��r�*�96�飰��l�<�`�ƨ!��I�愜��A�Ġi�<Ap���/�:���J\��xp��l�<�ҦȂ[F����	-[<�ي1̇e�<��f�l͚l8c���j¦?�B�	�nw���#�Y4U�2aCj�i��B�I3&�I$,
�-P���_�`&�C��8c2R��E��x���T!�C��0,-��ȿ4i�ZV�Y0`zC�Aih�@�G��BU���=@C�ɑ*`(�j>>Lr��?��B�I� p���+9�d�x�N�a�B�I��h�;��E<� ��&L��Y�6C�ɷ������( �I�C�	*n͸���e�	^&3C䉁?�b�r�o<!���� 7)לC�	�Yޚy�FK3e�l�h��`��B�I�i8��W�5=���;��B�I�U��Y�v�?A���HԤ��L�\B��`���JgIka4�Ǒ_!X"/$D��� �ϠVbR�gL@%Yܼ���/D��  ��nR5W$V�b��b.Љ��"O���a17U4 �0́�S%�	��"OPi��jY�W�<�d,�?~ZI�Q"O�`�-Ϟ �R��g+�5�@��"Ob4z�,I�U��4
�)Z�3@"OXM�1��X%Z��6� K�l�s�"O��ƒ3>�
���a��I�:��'"Ov$ ��2j���f(s���R�"O��Y�,ʙ�
,1�%�YkX�F"O ��'/̀���CϩR~i�#"O�Yڄ�ޘ\&�\Ygτ' ��sP"O&ܰ�
5Y]\��c"0�&@J*O�S������sV�1�`S�'��񩠄�3�1U���K��XJ�'A��0�*W<@� ���ِ@ 4�
�'ۆ�RO�1`����OH;᎘r
�'BYʴ���V������I,8�ƝS�'�^գr�[�k��Ea��ڢ&@��'�ڙ�D�2<���ϳ~2�!��'����F֟N�,�AY���K�'�R�!B��YD�k�i8~�V�C�'5�y���΂2��ᓢ�Vs1z���'[zDZ*��z49��4l��@P�'چ��g�#+VX�q�[�d����'m
�A�#�~Y�P��,1��`�'W���OA�J|h"��<�x��'͒�R�f 6'Yb��`Ç ���'%��IEOQ������V&��'Ȣ��g �4b8�	�	��}Q<���'8�����'�� J� ��@��X�'#�]s���|��Q�eEm�X=k�'�h̹!a�ڎ�C$�� TT�':���ʃ��,z�i�)i&���'�8��w	�>lܴ�C���̴��'�P\�e-JBg&�h�]:!����
�'�z%�S-S�H����s�ܸ
�'�2�Fn��'�&9�v� .�ab�'-�)S�N�Q�;A��-l�έ��'-´Ҷ�N.@�q`#�ؘ\��\3�'�q+���S�9+��T"?3\���'+n��iNb����8��(C�')�xpi_H�\�h�JP�/a ec�'
,� gV3A{&����(�$�Q�'5���˖8�vDQe�-ml��Y�'�8���"L�``Q�
�����'��2&�Y�2��{B�]�;p��'o���@�6!iQ����*���y	�'���b�# ,M�I0�����I	�'4Zy�AOP*L!z�C��N+9æ��'<�:6�TE u�&��
i�	�':�(g�B! ���R)�]!Ԣ	�'�"I����첢k�,�F���'ў��f�46A�[�&���j
�'A�8*gC�Vݦu
�ψ4#�<z
�',)��	(%)�(���t�9�	�'��XC��O�>	zU�O�X�`S�'$��23H�x��q�����v�����'�xY �#�+�"itO�$�@	��'V�]3�EE���������'���{��& �������"�A:�'�v�9r�
c`�0K����;�' p�AAǌM$��06G�=Z�'����`�pE��b�ŋ�'���	�'$e˓�S�i��%*�iZ���}���� I�F��&v�"�R�P#
�[�"Oj��nC��X�Q-D,u6Mp�"O��V�&���;����"O��R�l�b� ���#h����P"OԚTm�)=�@��bQ������"OP\��&�	]������L�$�D"OV="u��BRx��qC� �����"O ���aֵ���K!�Y�?��Ԛ�"O�@� �ʍRQ��yCAʎ�ĸ�"O�5Xp��_���Q͕�K��ՙ2"O�8��&ڋ��	P���cܤ`��"OJ���gUHD��p��Ы}��X��"O\���])X��-��c�F*a$"O����7
NLm* �_�/�(p1�"O:�!�'vH���l�(V,�4"O,���ۈ	5�pr�˅Mv,��B"O6�K�ʚ20[�l�-ɚG^�l:"O
@1�LD
J��h�U�R�ոd"O�9B��O��KӬ�&8Jص"O�=���L6D�B�"�N5����"Oܘ�@ ��P�N�"F�S"O�l�0N�"��9����I�1��"O$�s�@9jEBT�@�r!^���"OD�r%(T!Cv`u��hs����"O���H�r���P&�V1'�fi�&"O�a�Q��!zZLD��ǈ�A߾��"O|$��K8=�d���۔a���"O�	�#F�h׋�iqL��G"O���piX�R2�I�kÂ>il�0�"O$)Iq���!�/�CGt�JV"O�%#ծM�mBdXc��Qb����"OFk��N�WP� I`�/O�̊�"O��;p'�r�0(ʣ�
 ?@�p�"O��@L�"Q2�[�14��p"O�;3L��(�����:@�y�!"O(x�b��!%��l��0�y�r"O@�5圐i�<���L�;:VFA�P"O"��Sn��`((m	;<h, �"O���af�g�Эj��J�Y"l�"�"O�hT�\10Ą�ɂ��+#"O�l��0W$I�E��P2�"O��t��@�R�3���(��J"O���jLo-������74�,C�"OF(�UGaJX�!Ƣ�C�]r"O��YR�F6�
�i��B(�fd��"OB���cT4(��e9��9æ�w"O�Y.�1%��b"%D�N�Ľv"O���Ǝe�����CM'��H;P"O�i@��Ff��$BɳC�����"ON��ો�V��a2���T�Bh@�"Ot؄��W�yC������"OB�[�d�0 ;�92 �D�g�%��"O�2ri�I��i���oؔ�""O�i
�_��+��@� �|�jW"O
�{&�P1����V��
�0��"O�M	6#�*�N`0��2;�,�!"OtQ�Z/�6����
�Ŗ� �"O&�`1"��.i�gh6�fe) "ON��e�F'U�.�7�¨B��P�6"O������X͊5
C*Řw�40xP"Om9��+�Ui0�_�R�8��s"Of9SV(���-�!� |�"O��*d���P����qm�r��s"O�����4Pz,�r�oΌ��"O� �H���[�^��R�ΎF�!3W"O��Ѧ�;&�
�ٳ�(�����"O�́���P�����b�$�i4"OZd  ���&�9�����F"O��Z5t� ��۵62���"O~���'�uN�� Ê2M0�)�t�'��D��(��h�$ �O�r�=�ȓ;�$	aTd�V�4�PR�6��	��y�Z!�ܬ#R��R��?4"�}�ȓA�ָ-9 a���]�H����aJ4D��u%;\E:��CA]��-c�*O A�T���X�n���n�{���D"O��#6A�JNԥ�$`	�Iѐ��r"O��@���1��(q"�;V'��ا"Oj�:" �>e"͐�A�u
� ��"O�l�r#ʴ<�L1b�<_�	�"Oh	�I:6<f-i㠎�;��u�"O�-�T�Oo�i�f�Y����S"O|ܢ�ˌ5�~��u�ژf�e""O
pA���T�p ���6"O�����K�AA���dR�0g"O�����.���#�N]��r0�W"OFU���&�~�K�B�~Э��"O`T� �B�q �C�CK�"O�T+3)��|�U"M8[��-Y�"ON����.EcDq�
B��d��"O�0儋�R�TÁe�p�ޭS�"O� ;���f�$� ���c���X�"O$H�C��A��U�BM��/N�T�"OJ91$ܤ	��X�ۿD8�x�"O4P9'k�G�������MJN�`"O�IiFg�;D��d�`G�}��"O��@��Ne�%"ǡU
M�*D�Q"O����B����a�����w"O��" = L�Kp/E20��"OVԓ�I�|P�=�)_�Q��"O����Ίd�� TB
:fni�"Oֵ����@�^̸g�@��h"O���CBT�M� �����"O�!�MX-P�fPr�^]�k�"O���D-2rc�V��T��"O��k\/���
�k �5Kd"O��a$��>ܡ���%T��"O�q��b�b�nm�w�[B�4��"ODmQ
������� Q
�I�"Oڬ��@V.`���
T�9�I�@"O��9��\[&@��R�T�D"O^�y�]�+@��A�;Y�0�B"O($�#շqæt���܇��y��"O2aԩ9� 8��BÑ �~���"O���a��Da:�h�n~���D"OxB2��!@������"nl,y�"O� ��n'A|&�BP��P_\�rS"O��>y�bG_>S"��"O*@q"I�l3���#��?I�#"O���R���`��	�m�F��"O��	��̑�nА�핳M5*$�"O����ڦR@m��˕Y n��"O8��`I/M����*��jT@$"O�1�E��d	�
4�J,W�H�+3"Op�P�ˬ�ܘh&��&>�(��"OP�Zq	�Sb;�抣e6&�U"On��g�K�j�BE�P��7��J"O&��螂(�J@/���p���"O� �s���v�F��4�i�<�cD"O�I�$�!0��Q�#G݄}�&�#"OQP#֑��y;�^��:�h"O��[���d}Ԕ��>,$��5"OB):_2L�!��_!:>�0i�]��yr�4͈U����(�l�w�Z?�y��@ld��0拷�쩓VjP�y`����Ҽo��정��$3��	�ȓ"B���R�%"�H���L���ȓ,{r`�3����t`X��_8��ȓ��@cA� �X�w��;�l��ȓdx]p%�C�uH 8�I�b�х� ߆0;AGQ�t�:t҂*R�B����5Z'AV�&d����K7Ji�ȓ˰!�IW��l�Qj7�^Ɇ�b�D�l�!((�֤\
��ȓc��U@�G�t����T�$���m�(!��$C �L��%��(�9�ȓ.�T������`)������ȓ��S�gU9��H�&��[�x�ȓ6̨�cង���Q7-�k}4���POZW�6)F ���F)xp"O���D)BtH��aID�� �q�"O����k�Z	��u)�#j稬82"OR�y�F%S����t� ���"O��p�=c1���ǈ�^����"O޼��-*�� ҡ���\���"OZ���ָU�^�� �ȟ(��͊�"O䰊$j@.K� �ׅ�$�|��"OD�Dm��U��d�#�0�w"O\�`'L��{H�Y�գ�?�Q�"On�Q��؂Y$<�h���;:mA�"Oq�3����}��- �"O~�	@����Lb G�*e~l��3"O���rd�D �{@�P�� P"O*A��OȥoX:�"Q3���C�"O�J�r�X�2�O�����"O$$c��_9>T@��:��4��"O�=��qk������ 8/L�Z"OF��Q�.~�6�!WԌ9(ܼ:a"O&%!����|M"lJD�ۦ$P�T"OjĩE$.A���ظL��|�@"OT|��9MR�b"c��E=L�+�"O�H�񮓯6��H��E;̹B"O�@1�ޚ(��9@,�S'N5��"O���e�9F�ܤS�JX"^�ٻa*O�Y1T	�Kba
���}��y)	�'w�Tѣ�D?8]ڭ�S��<�ޑ��'f"�Ig/њtb-1$E�np\m�
�'&��s ��#w(�f�S�_���	�'d���cԋA��j60T7	C	�'.�C֕B٢������FrB		�'����.�2�r�dK.>���Q�'����6Nͮw�x���S%v��2�'b �����)A��a�NIG�)��'ly�%�ͅs줼S�n�	b�8�'����*)����+�$K	z@��'���H�+�.��8 TI��B6!q�'��@�+<7\��-%A(,E{�'���q�œ?BG����8����'���#��ݵ{�H=+p�X�B���x�'���@�u)���@΃DJ�q�'�j�!C�yG�a[�셞B�ȩ��'���@�ɢL�QcQ\B���S��� �E�$D�yj`�Bc��(xx��{T"OX��a��=3>�)��R!No(��"O@�x��2������MW�@��"O��[�Cѡ}@Uk�$n>T�"O�l@�O��P�����vak "OH��V�c,�c��h��y�"O�CP��c��4�;#���`�"OD���R9"nB��w떈Y|:8�&"O�b�������Z` x�e"O�a2���Y�T�CҨ�!ET��3"O����\����-h1��b�"O�d��	�.�dd�m�
�*p"O�`����tۤ-&�C
�����"O�}���8<pAx ��F�D�6"O440��]3C� GD��3�|�5"O�����DIP��`��d"O��YW��l�a�T�.�xYې"O�����T	�e�3��&\Tlp¥"O4��ꃪn��@�B�F����"O�-�r�W�4������K	1^��z�"O|(�fm��V�6AW�0%4�%"O�R3������!ǰxӈE�c"O������
�z�ՠ�&�F�#"Oj�bs� U�x��o�~��x��"O,�"���>@�$����� ~~e+"O�9�^:(�b�Va3zY��#�"Ob 3eτ�	� a�t�<K$(qQ"O���p K7Z��H�5C��2DT"O��� �E�_R���X6{���X4"OP�+�j]3X*
�`��3��4��"Oh�i]�M���WFP�q�d��"O��B*�)�\�H�l�hH�"O��fhϮ*>,p� <am�5p�"OʱӅ�V'i��J�O�_V�T �"O����2Z|�K � �[�@ �""O2�SƬ�I��`��O�O����7"OfL�UB�%Q�:@1�b@�+����s"O�	*�MVj�q��׋j�޴�@"O�=�e� b��1���_����"O�=��,�%�
�C͂�_��1c"Ot�@`�H���Dk�
�Y""O!12��{����I�y�8��"Or�b�F'uK��qۓh s4��ȓk�����7x���9dN�r
&$�ȓ@)��pm�;���%�г.;~��ȓjhm9�HU�D��Ap�/T��8��ȓr<���ä��F��Y�`e�zهȓ/0��sa�Ia�Qn;ꅇ�&4��(7&M@�	qe�M2*$ҽ��|��}�G��&�z)���O�*��ȓ����9-�)�RŖ=E�r�ȓi�J����o�й�A� �g$��ȓ<$��b��3?`ģ���2#EDՄȓN�B�[��+"��}SU�׬��ȓCe�[G�:]]6�9�_�c\|����BcO�>etT9j���!UVh��#3UA�#�63^<4�H��ȓj��<��@7/8��i��Zk�����a����1LB�m�#$��-f�`������2���`k�9����Ĥ��z"���.а*u���AB������W�L�z�MĆ\ڂ))�-P<Gt��ȓ�����Ȝ�7D�u���� ��@rL3�O	�)�,����Z�D����S�? �4�El^%��1�5�K�
���e"Ojt�7A�3W�<��!�;z�Ѳ"OJ��'B\��i11*�2K��"&"O6�k(^��lC�iY�wH��y��E�D���K�V�"�1D�·�y2N_�B�L(�í[G�,ȓ�'�yR�0�p���DU.	|d&A���yR���P�z�z&�S"}�r�b堆�y".�v��Hۧ�ֺa�]sD@G]�<�al2�ꈚ���.)�]ҥ�}�<�h̰/A��/��p׊��W��a�<���U��h�G�	�t���5��t�<�j�=~J\,�A�Ğ�j4�Wlp�<�d瞽"��#R�v`���p�<�Uf�.>0�B�6^܉�NS�<)`L���z`�Γ[(L�+�Q�<a��	��lɷ%�n0���`NO�<y3�M�i��h塌����eEO�<!�Ay��8���?M�;a!s�<!S!eȆ3���2u�EH�<q#�'LCT�PSU�|�l9��N@�<�VO��ZTȄc�~8Șb��u�<�E�j�����z��0t��t�<᳉S�W��D���]�B=���m�<PB�']Vii�eƉ)�d��c�<Q%1Z����^�t�����A	E�<�w� )�x�	���`*�H�d��e�<�&S2��8ɐkK��4hRi^�<��@��N�t�Cϖ�f4(A�$S�<yeK�Jn6e�o��a�N5��*�t�<�sg�=c�`�'��c�=a�o�<�%�3y�*-�Dτ�6����#��l�<��-C�>Q�JX�n��]�3 �s�<�ӌ�#�P� ��I�tlj�kHU�<a�Ӽp�ذ+��@�1�萫Ӂ�M�<A���O���DD^�v���e�o�<��i%~.�`�ǋ�4{bPk���g�<�v�G8ze:�b���h_^�(�_I�<I���8Z!�ѤX�`+n8xdF�<�P�Q��2����M/��1��-VI�<�nƌ&����큈G� @�Z}�<�7���`9��ˡfQ0+ʰS%B�{�<�1o�D�U�s���P9�9{�k�v�<A�I��8hZh�$��X̮���)WX�<1RK��l���Z2�K�̈���Q�<�⋕{����U��c�:9���U�<y҄�=th�!j�fW��F�`4D�O�<�W�P$b$ք^����aV�^I�<�7�G�*�<0a)�)pnY�BO�D�<��I�6j8t��3J�2�����@�<�3�Bj�zͲ����*M��Dh�~�<)6�" �V��"-ON�!�À|�<YSN�>�V��	ؐ`5>�q�kSz�<��(X�Kyl��ve�"�F�+��vx���'LD+1B���a2U��i��d%O���u�~R�"�ܞ����"O ���A[>��X`�DK�{�La��"O�A7C��}�D���D	U�� ��"Ol��� o|����B�R�|T@�"OВ���3ZJ�h���7x�x��"O&��m��c&Nb�� �"O� 8��� (j�|Ç䒽pC�d(�"O�P)�l\��J��7ߠf���8S"O�,���!���a��3 �LI�"O� ��*w`з,�Ā:�D}�
���"O����Nɼl�������E��S0"O��b OԿ4���a��܆&��9��"O��p� �w[�`��fҼS��=��"O����I��$	h%�랖D~���%"O|�X� ΰZ�� �C
jN؂7"O�9�
S=k����d*�Ch�|P�"On�y���3B�P�Hu��}(��"O~���)œx�.q[�	E�m�"OY8��	,J��PfߋX�e��"O�u��H�(��a�ܳ��("O(�!�&�6�3$�0i�؀��"O����$\���t���;�"O8�ã�+|�L�*���g�2�
�"O@a�vHc|�dC3��|�h�S "O���6![�g삡�$�&���"O���'D_� �WD0A!��z�"OD8�1�Q�!,�TB�$<�L��"O,��^�K��L8�&O�B�09"O~i0D�"�ZX�ͬ%��$�w"Oj�R�k_�
]y��X�U��0�"O��R��9x�t���mI!I���U"ONA[%iEo��t����F�0e�t"O��4��uD��	8*�Ќ+�"O8xp�G�^��uږ�\#�*�J�"O�<kQ�ǒ&����A.^����"O��@4�Z41F��p@R P ]� "O�0J�$��f*T�ϓ.Cab�S"Oz�P��� wΪ��mΝ����"O����ʰ;2�ē��I�߼�1�"O
0��D�5��������c0`��"O���g�dNԴ	0��F'D|�"O��C'��su"�B�Ȑ>E�}���D(LO�YQ#@�	R`���OL�~��pI2"O����\3$I�yXh�f"O>�86��L��xKfΔ�_Z ��"O��p��||<���9iC~�S�"O4��I��"$��l�>O*��� "O21�P(8�rt�LҰ5z�A"O��A"�Y�T��@ ��-qX@Qw"O����홻%�Α)�(�̄$#"O�	� � �BZ�g��d%
�"O�Y�
�8b`XR�o����!��"Oꉺ���BC:IN���uH��|�!�$���`u����={B�h:���!��ğ��q�.T".�=��'_vz�y��'�1O��p�� /�U�5�?pQ���"O,�**��l# �85�I�(J�k'"O�d�D�m7p�����O=D�)g"ODLi��ЗA��UJ�8_�ԡ �"O􈈆!�@�V�����y��"O�LS��J]b���f�lp��I�"O�Jq	�.i�r�`��n=�I矰�	çrwR�Z�!�i[���G"Ht�ȓ]T���\�"�T%#�E]�^h��*�~%��H1DD�q�Ӌ���ȓ?���TJ(
�.�Ag��+�ʐ�ȓI&���C+|���x�$ɉ�p��ȓC@`R��}�"�
 �̯J`��ȓIW��7�LY-��{SL�@�0��NNl�j��2G��	q!I �t��Wԍ���?ٴ4`�%��!��ȓt��k�cUv���OU0�z���}oj�"�拍��S��Lc/Ć�S�? l��5�\?�!J`HYgܽ�"O>% �b|���  IN��"O.���п7҄�SL[8 />�q&"Ox%A�#κ'e�]��N.X&�m�"O0GD�.�t}hւ,X�+�"O< �s�W)�جw��k`b��'"Ou2�o[�\�D)�gU
\U�� "O�Hx�ϋ!V�N�B2G^�{��v"O� R�c��{��P��&U4��"OƝ٠"U,I@ �PB1n+���s"O�����	/6�;�B	_"|��"O��U��,�	إ��9�T�0"O`�S �Bs8���DJA(�"O�e���B�m��|��@�y�n��w"O:�����
.����!J�ē5"O�TA���$�|�*BׄAН�"O��ub�R0�};�@C'�b��"Ov`"�,C�h���@���Je��T"O�<If���%0$X,W�`�)�"O�y{�/�Nr��A<y��t��"OTH���=�l�ʦ8���z`"O�����%�Z� >9ҒU�g"O>�Z�Ǝ�W��@���:�B�2B"O�q�5�[
~�l�o��a�i�"O�P�ii�J��-�t��I��"O2�b��]t��X���M�W"O�6�P�k���z� � h�~���"O�d(	??aDٳ�P>Y�>a��"O��X���(�lh��،s����"O&�vI`; ���"ĥy>�m�"O\����[��<��!ޮN/0��%"Ot�4�/}t�z�� W�HI�4"Ota�s@͔=R�	Ǭ˨#�$�j�"O:�q�횋P�E�ԋO�S5V���"O�t�����Q8�%`*O b���"O��kM��0���2S��0la�|��"O�9J	޷T�
���ac�i��"O
��e��G�ةq���2va\T�"O�Lx�N%t�D0#�֚"�(�"O�,�C�0����b�,I���"O<�āU�A'0�:Adçy�`��p"O2�aɂ�^��[f۷NYf�i�"OȰ��$O�<ĔAS���-��u�g"O�,�B�)�2R#�.��hiw"O�������)�7�U5-��Å\�T�IK�S�O��\@� dB��qgX@+.%`�'���`��оRi�8Х,�=�2uK�'6�=b Nؒh�E��O@��;�'C��bBN�T����\i�'����,�Z����#M��6ܢ�'5����A�.7ɰycE h�|8�'�RAGӏނ	�2�ŚtQ��Z/O@��)�)ʧ�B���ΧYT�\���]1�\��`�L�¢
*(�)��#!�\����Ar&K>C�f0Ɂ��8a��ȓ2�(9w�D3mvI�]�UxL��ȓ7��X�e�.����3O�J�d��ȓ 醨��))}�� b�#4�ȓ|d
2�ġ:L\d�t#�$t��a�����1Vz�@ �I�g;�|�� ���j����Z�.�#���)���0��I�5C�T�S���i�l���.�X@�򇉅n�N��e��%je"T��\����:�� ��"byj%��S�? �y0��]�N���Y��3jq����"O��p��p��pJTA)k@����"Oa�	[�L����t�� \949`'"O%�C21Ը�Ue�8s���"O昀� �i�`h���!H
�"O��i6!)ekL�F�Ն)��
�"O$}�512��C�X�x�"O0	g�<~n���`������'o^��Rl	�<�݈��Z�ER$�'Ђ�Z2�� %��T���U';Ҭ|�
�'�t�ä���P@^�9�
��g�2�:�'�6�P��W������oM�S���'5j\: '�6[\��q@�$��Q
�'8��*EC�#��ps�,��t�U0
�'d�esv#�R*
�1/��a����	�'� 0�	�<Q��a�0h:	{
�'Gb��U����|%i�	ۦg�e�	�'X��+X�jy)��C�k���G��`�<�q&��|�d��̄/ar��w�`�<��0��@��,EK�q��I�Y�<&B��6EtM:3��#u�X}�֭�O�<ɗ��8V��BL��}*ZQ �g�<I4˕�>�`� V�V9�eA�^�<�e-td�(�7��^R~$��+b�<!�9�J���R/k����/�u�<q�gȣg��Z��7��{�TG�<!$M� )J��7�LZ8�q�Jh�<Y��m���郞��u��m�< dY
.���՛v��"���`�<���T�k��xVd�C=h�z���[�<Q5�
6-~B�&����dB5�DP�<	�L���p���_@��r'&
u�<Y"O��'�p��ǖ@�䙥��i�<q���VQ��C!7�v�Y�UJ�<��U�j��J���b�(؋#@I�<���P]�ڔ*��ܲEQh\e�Nx��'?,�(A0�P����L�t��	�'�:(!�*1�^]���L�3 ^H*�'d��j�%�	-�d��p �~���'� ����\�ntc��_6�L�
�'�@�!�d��	�4�i'�F8.�F���'t��%�A!~�J�f*�= >��	�'{���,Y�?�P��2m����t�	���'q�}��-U�{�Z� �jQ��:	�'e<	����%>��������'���R�ѺH�r٣R���߂���'$�+���"K���pO�#un`��'��쁣��
K�2Q����!V����'p�y��B�3d�-��%�* "�xi�'�%Y'h�(@���kR����бr����F&L���qf˚M@l�b	�I�!�d�>w/.�㔦J�tD6�"�d�L�!�@e�Y���8�1��
�g�!�d�Q �%������g�&_[!�$[�9t���_8i�V	��b� 1!�qt�4:TW�U}^�
�AG,# !�<, Q%@�@l�����F�]k!�A!��	�a��wX�m$ �`!�d�SH��3�o�)BFpcc�݌Q!�d0g�QX��@�E�Y��o�?H�!�$�#"�2�ISbB�u�,8�h�%T�!�W�A/�=��مg�j��:&�!�i�jYZ�D�� ����B5�!��Օwa6��2�C�V�z䇔�5�!�� �᳗b��5ߒ0!��	�HQb�"O�-�C��;J^Y��	�6uԴ��|��'`az2݋v,�(j`L#S)p��"`��yr�Q�:���H���`�1�F���ybg�L��Q`��]��0�@�yB�."q�[��A-���k�i��y�ᗃz�%D��y��Q�:�y�ʂ8621��J�=qo�)������OT"~b2���K���"e�,v7LP8RC�K���0=�di�:Pڈ	�"פO�HX�g�G�<q���^4�� ��"���P�B�<�!I�P�8���5x����z�<����r�`�u�H�H�@Tq�<�M˕R1�9C�냒QK��v�R�<q�,:(l�h� �3��0p��IJ��?�	�'6��ɰ��B 56\�^�VA�u�ȓ��h)�EX�k���k��H:l����Q��ab&g�HR<�9@@�l{PU��z�P��J�W�8��c�<@�z���J%`������(����|���ȓA2ĉQ�>&�pR��2�:9��a̓2�B��n��^`�Y�Bl��s���G"�S

��4�֛�Nu��!0ԨC��4A��bG<k?}S��Ò;��C�Ʉ����hU�`�1�6�O��JB��<U���Zf#��)JDK E��
�FB�I�zx�} ��(5v�hn	�c�0B�ɸP�$i���@4A@�j3�\W�ȣ?q��)Zݶ5`��� xr��v&�"�ў\��	�h��@��"��e��Y��H�C�I �ιc�E�K&�� �K7 TLC�I/�␙EH 7L��U�E,N91 C�I8g�ʀ�+n8�%JᏜ�C��2A����w+��G<��iwꎲL$C�I <>�� ��ɿ]R��gE�����d*�)wHh #(��#�8}�"���4B��H !&�����4#�@'��F{���G��U�
e�DBG�������yr��L%��j�W�y�t`���ybAA�.���9C,6�x���OX7�y"�@0\$4������&FB�Q��y�&@j������JG�$B��S��yRf]�l��j��F�@# 9䎏��y�)F-(E�Wh�9d�RC˝0�y2��m`�i��s��1�@ŜpI!����Х2��P�V�����I1!�Ğ0L���A��޼>��qR��#00!��&:b�Kdș�l�8,r�&ײ*!���]U�u���� 
u2L���; q!򤟦j�F)�4k	�+c��g#I�:�!��P�pi�a!�*U^�ab�*�!�DǑP��(qb��o:������~x!�$ԭA�R�z���@1��ի�rh!�D
�\�D�!��*�Ä�
]!�d��aͨ9�����F�I�Ĥ�(p!�d�=�vթ��d' ���eD!�D��=���#���rg�}�g�!�$�'s�ࠃ-H8v�%���!�
*&�4��k��a�@�;!�$#p��0hС,w\���b�5�!�$؈��D[R)��|S��^!�D�^FҥJ�Ê*"T��.� .�!�$X�t�L���iǷR"dU��ݖ{!��DRm �h��jb�\R�� t�!�� F��eG�]��+r�P�BߺQ1�|r�)��;9C|eb����}Ė1B�N�=Pq�B䉡;L~�Kw�Ʌ$����&U�b�rC䉍>�4ɑ�b�h�A�D�h8>C�.6ta@�8W(��2.TD�JB䉳OW0a��O۩b�I��b��H}�C䉬,�%���_ݞ��Ev�C�	�
�n��%#%W��sD����B�	�>�~ɓT���,����H*B�	;��4��1QɢȰaKD�2�bC�	�@|d8b���M�dI� ��B�I���Ű��@�i�((�%!��_HC��> ��`c`�v�(|��e�?@�dC�Ɉ>2|�A���-W�8S��G,Z C�	�1W�0$퍫]]D�d�<;hC�I�_��8UK'Z9\!�w쑝Q��B䉒,M:����O�Y-D�d�B��� ɝ���E(�p�!�"O ܓ2��,Nɮ�	�f���Ca"O������6�L�#��o�ʵ�T"O�:� L�s���9Ab��v�"O`���e(Ǣ ���Y�#%���"O*�����p<x Y���!��`"O��CM�R�.mbBBW~826"O�Up�(��
1 ų�(zYj�٧"O��!��q������qQ��'"O�#��J(lb�j�)?=x@"Oj��GhO����J�wN�Y�"O�d ���+��ݪ���vM��h3"O�%hf���5�6D��M_�>���Kf"O�YKV�-4�Z|a@ύ(%���`#"O�Z�Æ5�pq �����L��y�N�&n��hs�Y�5@00���!�yR%o�U����.��h�Ȕ��yb F���P�X/Q�*�RC���yR�O�ѣߵ7m���n	�?��ȓj�l�۶�?z��}k&ÒGP��ȓ�|��$��5V�I��N�P-�܅ȓ7�*��(�i��튑˓3+¸��ȓsن8��׆G����E΃-�<5�ȓ�|�)�#�R�"!д�]�f�4��ȓ4��3�-�B�}1�ȜHVDH���t���A],�$=c�ѠS�Ņȓ#��Y���I�NRTc����fQN-�ȓ^�b�	�lQ%<�"��p��E�d�ȓE ��
��XP'V�q2� 9x5�����l_&=a�t�ӱn�0ͅȓn{����C��$C�
!���ȓ�T{�瑒2�l��.60\�ȓjt|�gP5
�����pS�p�ȓ)��P����]3�@nRY�ȓ��@���;J�0;#��/hB��ȓ4ƜeK����/�4��Ƣڭf}!�d�20:�k�F�[����E��/!�B�kq"5*����(�@yZ�KM�!򄈱�$�JP�ݯhu�al�	!�d�9mԖ;oO��eHG*	16�!���.-�m�L�$& ��)_�*�!���=,qn�����{|��G�ڟi!�$ܫ,u8�:b�Ѿ���P"�,-!�ǌ�
I�7��<|�4��Вtm!�,:�*qm٧/�|��ʞc!�ɇ;�ҕ+"� B�8Hҩ�<a!��(V�BŨS��X��C��!�� �Ũ�kɚ+b���6�Ӡ8M<MYW"O@-�Eh��GKv9�rG�2נ���"O��i�A�~H�po�����U"O�	���U�� [�+��<��#"OJ���B�x���j�
v�,a3"O�@�D@؎h��p��RchP�@�"O��w�Eb�xDk�K��;^raH�"O9�S��TՖus�HB�~'�u;s"O��kpH�(<8�ၰ�]�I!�I�&"O8-�嬅d_&I"�e��8���Q"O�,[%	� �!�V���H�x�"ON�c�	�vt�aI�0F�p�4"Or�#v�ӸVa�h��4-��P"O��ÀFO7j�qJa��C"`��6"O�\��I�5�~�� H#C�d �"OD5)�(C#a�J�Z�'��{IV1a"O(Y�Ƣ�5b"�e(� `���"OZ�SKX�Z�L�a��Wۖ"O��Վ��!.�"v��=~��Y#"O���G���X*w�3n7\��T"O��B���72h�]��)��J��k"O��ӲSt�&	��(
�cb"O �Y����L�"I�3�^�S�d�QQ"OBM�Ph���)r�ֳ%-|�P$"O���Q��r0Ec��� �|@"O��p�o�!F��Q��["d��"O��sda��%5~�`U,iV��z�"O:	�Ɗ�8�dI�#f����("O
�	���PW
�2a�2��$"OH�J��
3����hI7O����"O�m��LtP�Q�Ι�Ol,�&"O*@� *��@��y��5�"O&�#���u��Y��?�:��"OސZ�I�8=�ԐR1S�c��I�"OJ-r�䇓HV��S�(����[�"OL9�J	�<���sG�$�0x�"OV�@�d��4p�#���hն��D"OPq֬B�G
��T��I-�	Y�"OF�"� �5r�b���fܬӷ"OĴ+$F�f�*B�T�M��z�"OzyX�遛b��+u�����"O�T{�O� ����G1Wt0�"OzH(`�'xl)��_�n>��#"Od��!�3�0�� g��u*��[S"OhI"� #D�p91���h�1ZW"On���V�r�d��hȝ(�vT�"O�]�4��X�,���fٝ~�Dܘ�"O��y��ٿ#.t|ʧˊ;*T:�:"OL�C��,�LT�mְgO��"O��4d���M��,Ǻ2O\Y��"O����W ,D��
C�s���+�"O� ��,DE\d���JT����"O���dE� p ��V��3r5��'U����H�\"8�W焊G.�"�'��;զ� qu.��Z�j�6a��']�E�#�I�h�<qc�� ?\M��'�v�wr��[�a�-B��e��'�V�)�咇�L�iT8<*�Ը�'$f�A򨃤y׬EA��1-��L��'H*�k�j�2Cl8�ʐl��+����'����P N!�00�*Y�[	�'!��8��
/`��2�� :M���'匕�. ����-"R.��"O¨r�'8b@�y��Ǒ
o)�e"O�  �8���a��m�fm��&Er���"O����e�z���8>jZR"O�P��k��t��cf׉G�x��"O$ �g,E5/N���E� ax�"O�Ay"�B�gߞ�sd��RE�@A"O����J��<�h�JtC0JC�Hk "O�T�`E�S�4�b��S>H3a"O�}�� T�D��騐����M���"D��C�`2K������`���3D��ƏZ��H���G�����*3D��4AŏJ�"P�H��K
�Qx4�2D�����/�
Q������B��/D�|����P��e�Z-@g��h �/D��e.ڵh��LcF�� G�4i�f�-D�(y�OZ8<�zq�U#�$��1D���� 12�\�k�`Q(���e,D�$���8z���a�S
����(D���l�|3fK��l[�Hj��!D�����R^¶���%> �����#D���qkA�ل�C�(M1�$����7D�@�#�8q��,
7��:M�����/9D� �5���]���pǆah��9�j7D������%"�̹7�Q]xHqAIb�<�C��4KO����	ژh��嘥�IX�<�dK��d,��tǜQT�MТ�K�<��"Q�l��8fbN�{ɂ��cŖI�<Ag��������ܾ!O�aA1dC�<��fJ9����*��I� !@�A�<���3�xx���]��]� ��t�<��KM�=n	(��X4�셁D��m�<���A?p���8�������`�FA�<��)N�V�nY( ��;H�`Q	�A|�<��סFDv��@!�Y�||q�)t�<���#$WH�PԎZ7w"�9�t��m�<�1d��[z��33��3 ��1��Z_�<i"�Ȗx�bݢ�hX�'>� ��^�<	4N�n.���[�0�3��Z�<y�[58�p0��_�:��SG�Z�<釉*k��ɓH��8\AYcG�X�<1�@~,ze{�Q�Dw �j5�X�<���ԪNS�0� ��&,��i*p�RQ�<���9Ąl��`	";2���b�<���-�*ɂ��8�(��Da�<���V:v�N"���\���`�r�<Q��U�=@!�R/�G1T<��cIo�<�SfX1_�t��$�!��aE-Hl�<yA��2"�h]�Sh���ܙз�A�<A($E�JT�6���9>�Ҩ�t�<9�!�0Ĭ���}%�蔌Ae�<p$�(taPo�WR�YHԯ�c�<q�j��?]d�!@��8�#��Ut�<QuCM/xn�:����B׸ZrBنȓ4A�¯T�$E��Gɝ���ц�=�����m����F�%*��݇�i��A��HE����b�j}��S�������HT�֖�<�ȓ�X}ÄK�.��V�ۑ ����ȓa�B���i	�z��ro��\&���ȓ��\@�ΐK��岷�P����ȓ@�~-��%P��Ja�R%�"���J+ � �\�6��cI 3x ń�L����L�#�&� ֹb�&�ȓm���Q(�7y��<�Ңa!2kKG�<!���ް���ܸa�rQ
��<� L�3��\�N�6�0���
@�*���"O�\	��T!'wv=�6�S�-甬��"O���T<B���$I;ֲ��"O�qQ����.�4 �Ï�K�=C"O��S a]�`}�QJ������"O�}�qg��H��t�#m^5k�F�Q"Oh�86C+%B��*BϳYE<0��"O`hHa�F+M��G��� >rX"O��y�,rI�.�'6,�B�"OPu��G&��{�C����"O�8R��< ���C /��&�T�`""O��JtL�QJ���sC�i�B��"O���F!DV��1)�!A3i��
�"O\�`5䔉S��d�b��A�t�Z"O`D�s�  �<�#Qg*��"O�}���C�OϞ���AF
\T�aP�"O�:iƲi��˳.[�L��\Z�"O,����
U_�di D,�άZ0"O41{7��=h��\�v��+M�����"O����'ބX*:l�R@7nLMB�"O���P�#"�pCD.O�@�az�"Ok�*�T ���,�(`� �"O�0S�쀑*���l�)!��3F"O@}:�����(�j�"�X��"OZ�{n
'?�D��3�:���z"On��T�X�M��<�2�H*�ZA� "O\T(&��OA��îP�sr��8""O��	P�Ln"J\���> ~�L�!"O��j�WfT4 �/�Cw���"O��	h�d�d��\q@��"Ov�{�l��б��o´e"O���)X�G,d��&�ΟCC�i	�"O� :RO�@_,q�Ǌ)d#*�Ї"Ojh��Ę��M�G�;��ӕ"O��r��l6��@O,�� �"O
LP��e�<D@��O�I:6�"O45Ѕ,g�	�1@\! ��� "O�@yU&
=�H�6	C%-�ŉ�"O�P�M�8 (�k��L�G����yB 	�{��k&n�>i�ⳇ���yL:Q�V�X�M)`�@����8�y��\+%�\���]A�q9Gj΍�y�/���>4`#.�V�����n�'�y�aĘx�����B�K^b}���y�MG<l��ٺ����7 ���ì�yB.S�"`~m�2�A�'^h(B��y�c�Jp �V�ܣ@�)�w`Q�y�˓X�|�`*i囶D\�y2+����`kC�HfB(�	?�y�cͷSF���$B�\�������y"hZs��86G�4Qh�$(6��y���2%1ܵYV��Q��p���y�D�PY��1q�F:r0���ǋ ��yr��pv�`�G�ΘcH�j���y�n�+����_�	�V�CF�Ȱ�y��4y\!��/�t 􀸶�ِ�y��V!+,���M(�j�UHO��yR�2�ޙ����M��0(O��yr�ɥn0�2 �ģ%6 �CJ�y�I��P�yO��V�@�P��y�ؖ6�je����V�V�IQ��?�yr�S%{�x���Fz̈��C��8�y"F'F<�d��	ۛx��+�Ɛ��yBoW��ָj ��s��Њ��[��y
� �9A���lm(�"R�75�V"O���b�
\�e!���/2���"O P�2��3������y0 ��D"O�J��U>/N���2,T��c"OB0"|P�8�I�$�����"O.�#%L9y쑢�a�x�� p�"O"u�"	�W��qb�5f���""O �Y)P</�\���}`U�B"OT�p$Ӯ$T���Hp]�I�7"OB�2U(�/3	t�1g(��L�j"OĄp�GN%���7�˟i�(�"O�dQ�\�D�P$8���&DX�0"ON`���ȈR�l%���q��� "Oੁ���%'���jg-��z~�s"O�{Ť�.+bR���KN	�\�
�"O���`�ܠ���{Ɗ��z�|�;g"O��C��;a���ĩT��8�"O��ZNV�IE�u�%�{{4�@"O����!��K���7@Y�0��"Ot��gM���9cK�J����"Or�#��V$��8;q�V�}��0�"O��&�Ӫ}5��@C����"O�qɢ+��f��t��*x�Q�"O:ɚ��W*o&�!8!�Nr^� "O&��1���&�����4�>��"Ot�A���BA"�3�6A�P�"O�嫓A�[�������s�T�a!"O�$v`P�Fm�`.������"ONi��j˧y�Vŉ0(�Q��p�"OҔ�1?hd��'H�&v�>��"Oր�F��Z�z�S�蝰0���C�"O�)���eu��*��|�bT"O^��1�[>Z�X���*P���Ec`"O�`���JL�� 8n��L a"O�<�F���F���j�3�(�!"O���AG^�Wc�ˡIǊ6�h	�2"O&AP��
.mP�9 k^�t�5��"O�%�����[;~490����z-�g"O��cqA�p$�8'`�=,����P"O��`�T�=~~�#�nWC�DP�"Ox"�Ƴ&�RkI� ��U�7"O|H��	�	:�t�8SJ<~|yb�"O�p��4,Y(,@�	���is�"O^��6�I-�b��k�}��	� "ObyQ-S2�$M�$
S,���0"OD����u�Р 	� Y����"O�@Q�NݮQ�ҡ��D�B��<�"O$��ڸ|}�Y	Ą�	c�p
�"Ovc�Z�l~�	w�E�Z��"O��fa׺n\��P� 
4O�a��"Ob!K�����\4�y$y��"O>��W�(6P-0�ȊA#x�f"O��z5O��[�����Q�D+S"O��b��w�y1�/� �@���"OH� э~��Y�Go�?^@���"O�!Aō�O↼��]�r��"O"{��&�`���];(7�՘�"O�A�@��s�j� �_A�yj�"O���򥗦#��Q�DH�[2�]+�"OΨ`A��!%��1BÒ�*x��5"O�!���#J�	�C�
����"OV)FL�0��8CU���V^�:�"O8�Yp-߰� ���r��P�"O�-�T�:���m��b����5"O� �HqQ(�9k0�qZ��	:�i�"O0���MW�t>�JCM�c��MXV"O�T�b��(7>�k1�,	�h���"Oҵ��ӅFO�(
�㕋\�} "OjD�r���h7��եL�"�@u�a"O"i�'(�6ڪ��n[3qў���"OV}sv��;Nn�ڱ��:�0�{ "O�,�iب%\�x �g�?,���"OD��iG�$`kw��W�PH�E"O�9�B�^�&!A�A�n�Ka"O�� �@C�$���o�RO��"O�i����0Ce����hs�h�+2"O2��(R�~�Aᐭ�7ۜ`h�"O�A�� �Q��{b���(��"OT:�ё'���b�k�;y�0��"OP	D�Gˎ�h7J��pLu��"Oz��fI�B�L����Q �}��"O�I���c�� �bIV�:�Y�"O>\[Q��`�~1�*G�V��tڤ"O���҉DN��3�*K`aZ	��"O4ub��ǡH&�E�C�ܿ(�
y�"O.��5/ ,:��S�³T�|�zU"O�ɲ �T�]��K3Q��"O,� ���BG�:UdM��㛝M�!��Q�e�)��2<r����!����,bqgI�V"�9�UA@�)�!�@�z�����."�<�QV�\�fF!�"sr0	WE�e��A���&,!򤜎T�,$k��#LlZM�$D�h!�DTi�ɻҨ-u0t@�c	�o!�d���F%�G�!~�(p-�u�!�:��I㋚�$��ݘ
�!��A6x4,�td��tm����2U�!�DK(\1���1�����	J�!�ė*U 	��ᕗ^Ķ8���e�!�D�&�2- '�C�0f%��i��=�!�$��UL!Pc�{�|��)���PyR(�2hX�Ls���oVZt[b��y�K�-Ҥ8���� ^����� ��yҌ�/KW��Ӂ�#Y1Q�R���yBۭ�jԙ1#���^yyb����y�o�(x�F�TjW0��bsB�y	�=P���&��7b�R�U>�y�BϏ3�>Գ��.�@�����3�y��G�^�����J�z1�ᐅ�y�N0
0ir�Q�t�0�
�����y¥A-G_�e�Ǔ�@jU"����yR���Mn]�蕊����m�y�	�n�nDj��T�xϪt�&����y�D,K n0��_��iㅅ���C�ɳ;6+o]J"����=М��'����,��;Q(pk0���a<�-��'~�y���[= ( R�l�V9�
�'V�=J�a���5c�
QǬ8��'��i���0�����J�n{�'�:��@4I�5�ț1�3
�'�̜ia ʔa�j�3%A>�L83	�'�� �/3����`K?Nꈫ�'�j�b�ǚ�a"� ���=X���
�'X��j�>��P)�$��|h����'� �çh(}�|���ʿ��9�'��X�Gc�"<� �@Ջ,%@��6�\,0��
v{R�{WFMx�t���A�S.Ze������
9Tԅ�S�? ��� P03�V�Y�ʥ~ȢD"O�]Y�>Cf�="ֆ�,��9q"O�U�d�'4Z����W��aI�"O~�fiH�A�����?4V$�aG"O|qiT��~l�Y�D��)@v�&"O�(�F�2*��lY���
GL
��*O�Е��h�\�2!�����
�' t�Ϙ�Bb�R�G���{�'�F5���TG+���Wn�D��EH�'@h�ȝ2�}�PKM�oԎu��'�㍐�j���V���a�L@�'t��S���0�^/X�ੇ�=�z܉A��_�� 9�)̓\8���ȓe�ĳ��ݑl�<J7�&k}� ��H��} Ǭ�?+�.4HS��1$���JO�(ɥE�a���a! �B�)��{�kƎ��@��F(��v� �ȓ:7I�D)?Ρ�lV�3���N���9�+� +�6\ G�
ݜ���7}���O	�AA,�Ud!��@$��H��|�ׯ�*���`�ް�B�É�h-@�={��ȓz�� ��2N��ȓ4�K�7,�i�ȓ'>�X��&�.��P�7�(I�ȓ/�,�:6ףg���#w,ӈD��H��#;�8�V�ɲA�sá�WFE�ȓ$���FB��>~l�ȓ%�RE�wk��t����@&ي4 F�ȓ#\ �#/T�� ��ʚ�=�޸��M��Sv�- #���Eك&�0��ȓ2�b����]�Hf@�k�ޣ:'t-��TT��2���@�"mN�ϪلȓdN��'e�6)D��B`��n�<�ȓV�Py2�@%њ��Z�&X�ȓV���H䀅'��⡦Bv�&��ȓ@&��e�
�E��D�ԅ�i�b̈́ȓ���[��U�vפy+D��a��M��wܱ����	x�����	�lhD-�ȓ6��zRh�i&P�
)���ȓ����ȉ�>�d�'AZ�!��l�ȓq������7�PAx�aF �q�ȓo���qM�4i`�mȥU�VT�ȓs�FH�ŬC�[��҃�|�p��PU�U����%�ԉ�K�(�ȓ{EN��Bo�%����b�ԅ<�@�ȓ?��p��/�aB
09!� �:����z^e���pNl�(G�P�V��ȓq�0 #Տע4�����]�@���$����
�$�3�mQ�6�����7,.�P gC�:� � �f	�Wo���:Z�x;�� "
�@1@��ދJ��I��t��a%�{�8 `�/e���ȓK��1����>�\ccL�S����,�Ry����9j\�����[X�L��x����#��<1ؔ�#B�ftZy��g6��glD�&�����iiL��ȓL��-��I$;�2��ӧ�1H�8<�ȓ8��,�&m]9Y��{7鋖Tr�<�ȓ�|#��=R~�!��̝'��)��&x��&kϛ�n	i���7��ņ�jb(W�q��_`���ȓD�\�����	KO��	�J��XXY�ȓ|A�X�&
(	r�
DK�+TH��g���c��d���"�)NC�)� H�Cdin���ʇ@ƚa"���"OxM�E&Z���ŠL y�]�"O�|�7��.z�`�`�C���"O�4� \�s��Rn���"O�M���źdp*����>/YĒ"O(L@�o%r*TYc��.K��j"O���w)w� �	��ݕvWʬS�"O��	��6z�Ljn,(3Rp��"O��4�_0}yJ�X�M�]�"Op��ԨV�7�6 ��
���K�"Oxx���ʤ��"C�<d��d�v"O�XS� /;r��t�RHan�b�"O��0�zD@����8b�����"Oha�7ʀr��Q��c�5�Ї"O��3p)�	>��V��	v6�2A"O�y豍ƓEk"���HT�kKr<k"O
��玨~Z2&� K,�%�"O:\ZB��	={$��"&�D� "O̫�Gk1P���n�"1l��'"Ov� Í�}2���  y�^��"O
E�I\�p�|�R�"�2p��"O�0�@D���u�P�z|B�"Od�����#���`�\�
���1"O������%ML���-�f�D�0"O�����\�f`C�e
�Ph}3v"O��a�!�5[�$5�%���d�K"O���E�B�\8:�8�ҮO�!��� �zQT�V�mN�ř��%$�!��6i�5`%ɔ*Lڑ�"��M!�dC-!6h`�2�*���nĊP�!�$Y�5�x���VϜ|㴇��^$!���(<"���`�8
�E��G�T!�H*o�j� Ì^�;��<��Ǖ�b!�7O�h��bV��zi�A�p"!�D��]�p!�H����$�s!�d�#=��;EF��U�8�p��K8	!��?%J�ɷ&��tg���虄n�!򤁯7-��!c�X���>�!�D�hC��#���4 �y/Z�(�!�$�	��k���s�t�I�!򄍧.0�Ei�A�cj�� ��^�!�$�2]��C�MV2HR��s�σ1�!�� �aN"��$GW?�퓐CE��!�dI�H��!��ܣqB�I�#�g�!򤅧\��тӮ0W��%¡��+8�!�dMH&�2'�
�Z2U� L�n~!��֋	xt�b�C�ww��(p�$2w!�dC����PWIi�X� �H�,w!�$I�"�z�x�	 R�X-�al!���Ȥl��#����'[H!�䝬=��q�m72�P�0�O��x-!�$��j3���B�� B��j�<��N��k�ŉ�f�:��.���ȓu�������r1��+~�*�ȓ%[.C��(�D�"� *-�`���th8�J�˘�f:�*��@?9C���A��=+�F�9ڎ���7T�B5��@�R�����Vd$�+pV����dUf0���9�0L����N�ܥ��-�d�t�ӇWv��ۤ@X��2-�� �@@�gI�L�J�I*�LV��ȓ ~J��R7U^�9䞼����a�L1�`�-���r�ݠe�\��
��j �øG���j�"^��Ȇ�S�? �=���� w��\��:��(�"Ol� ��;gj��#Oэ�&�P�"O�"UA���r�C��|���"OPD���� 6)2���U�4�A2�"OD��@/]"<�"��6�ˏ1 �ʴ"OH�yA�L�$��f#��B2 !�"Ol96(}�2���#M�� 
�"OZqɠeF�9��[�,ܪ#�jK�"O��d����h7&^9!U�
�"O��"���ifB������K`�rS"O2�$K^'1����}B^��"O���G&@=����±)b !�"Oz�
r��x<��q��f	l`��"O�bk@�^�na����,*��9�#"O��ؑ��d)�B����t��f"Of��5�Y��`���#*yXa���?D�h�@A�$*�h�3i�.-� K*D�\���5�p'ҝ)�6��'�&D��R��EN=���c�ì�(��!D� �Ѕ�g���BGhB5����!�>D��:gA�OLT�DdV�U���
P�;D� ��	�&gP�C�O<B�\M���9D��Z�/�ѸT;� �<�~�h@�8D�:��ߣP�^�q"��*v�p��G<D� ��IC�s��$("����<���$D��+�AE� t��(ǥh��z�f8D��s���S���s�:Fx�p�#<D����L�S5AH�o��&����9D�<2'$�D��D�����b%D��i2�H^%���G� �ɤ���7D�H3R����V ��L� px]�0�4D�ء�ر�6m�#I�>f9�w�0D�P��G k 0�	F������;D�����y]�ah�1V���$.D���Ȃ�Nd:|��aA>�d[!� D���C�� k�@q�dA�ckhQ$T��r@�Ymmh�9�-Q��8�a�"O�]��m�C�*�@&�E<�0���"O�<�o�&L�B�KS%˹8c,��'�(]"�b�-V��a#�P'iL �����!����-�4>htER�H !�!�D�3/�DC��|G0A26#�1�!��V�^&Д[�͟mMLu �i�){!�G�����z$vx�&�H�!�1 ɡbә�4��!�DK0~9N��A�ث6-��A����!�D��
,+wl�,SPa����9�!���k�"urF�	�L	�d��6*!��XlN�SQ!c�h(i��W!��6庵�d!F�p�^�z��Y,d�!�dS
��[rW<���H�H�+�!�䚥N�z�'$?G|$�A�Q�!�D�?C��C�,Ɲ!�����a��!�d�-#:����-(ʮd��C�:+�!��$An�ȃ [1{�����Q/Za!��W�/B00n m����!nİv�!����=D*�"��7(�����!���z��9yu���������5�!�$FzN�M2q�I.W4%y�ϑ�
L!�ė-'�.)����AD!��	�'�����ԬM"�p�"a��R �3�'�����"v��e�"k�U5����'pԁG:=���AG�ZM$�ϓ<��ag�V��D&y���$	�e'��Q
�qs!�d�?0�����=s�ء�j_�1��'x�\���?	`��� ¤��.�b��tp�f�{�2�Yr"Oڸ�j�((4�
��t��SPbͺ)�B�,�(�9�`$�3��ۗ{2QU�?MH��A��T�E�!���y��2�PR�x�yeÉ�A|Z�:˚� �5�XX��(")�4�HX��G!F��ط�(�l�ttᥓ�A]�)��jb7Ÿ;��@�0�2. }x�!p�<9Dh4`h`����`�sy�ᙇwPh�#'���i\
���(���sM�x��9�!��8yg�`X�kA801�EC��(u� ���
���3#޵Wq
�:�Y>�<�Q���ű@��+��Lkc�UHX����F�0F�ɓ	�6�]%
֣�x�Z�I[���0[@y9E�Vc8�:F��� �n{��!��Q�$�q`P�3|4��Q`D*it�=�Q ����ƅ�m�}��K�+�aҴ�y�X��z5:Ƨ�
���!3���I�"`{T�	1	Q=Lxu r�l��ygA�h�(y��צ�~Ma�.�yb�Fo���*�e�}����BX+�|���kX*AP��W��2$��Z��o���Fy�D_P��\k K�pǾM9ҀS���=GL�'.�7$��U�:A����v2Z��Р�bt���]ݮMr ��a8�	�g��ed���tn�uK�����;�I�Rq�U{�F�����3	�j��0;5G�?�°"�m�:I��ƑP�qҮ<D�4J ��p���I�MK!>�ٳAi\����bg�C֪(��iѾ��-j ������@ߙHY䵰"�=4$Q�4�w�<!�.Ҫ�q�#j׉(���g�֮$�6����P>�h�����-{�r�"�Nҫ|��<YքR-xh y&��z�Z�*���i��L�QC�������M�P|+��c@��'�Q�]�p���4U�"\s���:�p>��	7�8�RM��-:2�ã�b�ũaϐ�H��6	U�o�"X�a��I�qQV0I���6y�W���!�$�1\���C�e�,�p�E�H��<�%�^�SU|��2�M�qU�U��0��O�*��;�Z�����8����ɞ:
8D�ȓ|���Y��Cf�\�RaB:q�,1�7)I��* �)�.0�K��ӡ|���aP�"ʓj� qK��ͥYIH�yb��9b+�!���j�|��.��c���JTMA0m~�����<C�(h��
f� �vN�-ւ!��"\X���6nA:�I����	�=�h��K�<�r�F�v�m3� N���謟FAY�R$���@g�6#���D"Opzt�})�!�0+O8�a��v�|  �'��)��D�0@�P�J'§�V��MXa�c�#d�n�(p���6L^C��-�h=�#$��$�nM��4��l�R��=E�s�5-�֘`n�ٺ���N�.:V����#'	P��ӟ��{� ��wj2�9�M�,9��D.� !=�A��@��.A��c��,A�	
�� l ���(��Aѩǒ8Kh	Ex2�-#�hɑ"����Xgh�����ah��oOЄ�B"OH��&j�>���Q��V�{OF�T��)m�2��͍���S��?tR�5�Y[G�\�VM���Kv�<�R��98�N� �EXr��f�p�<9�*ÈJ��X��A��\1AM�q�<3�ސ[�����QQ�t�E�n�<��k=\��)�i�?�`��RC�o�<IM]���yqh���e�A%�d�<��+7~��W&�*8���Dz�<y�	;m��*%a��e�E��`�v�<i����j��+V�!xvB�P��]l�<��Y$n�: a2M�"X��U�� �D�<1ǌ�'ǘ��T	�=��9�	_A�<A�L��:�F�R��W��ܼ�F�B�<S�ױt!��0r ��4�L��M�{�<�Ģ��d�!�Αei>�C7/JL�<�CG�*F1��޽r�4"� O�<q���6eFua����%˕@�l�<��\5?���WI���T[���T�<9�+��d�0�`ې'��H����<9@�ǈg�(�b�ě�88E  ��m�<ѵ$��t�)�:F��DX#��j�<	3���Nu���7�B0MZ ��De�<	�f��$���� �,.�n��i�D�<� �LsE��L����_$~E�T�"O�(Bp�ߡ}��;uF�"x>��HT"O�,)����r�`[�f;7��@��"OS�%�7임 �ޯ*����"O�ڲ�!H�<٧ٕ(�� !�"O.�f�A`�
A��#�R��Pq"Ol�b��9:�c����SV��"OB���N�3�hX�!\�.F����"O�Yє�P�_r�Y:�[�i� �"O�EZeH�3~� U²�4@G��92"O�@��·W���B��A����"Op�ۢ͑(`�,U��ѓ\���"O4|�r��$?,�1׫�3d����"Od�I2j��c�RA�F�D���U�G"OT$��
k皔 @�PZ�0Y��"OLU��ɉ1�$�YBW.(`ڒ"O2�[G�܁`�H�(�s���e"Onњ���b�CF�ߠ��D�U"O�U�����ؚE�<1����"O�$3�ț����yb�5�mk@"O�P�ԯ�'���!�G��d4�@� "O2,���8�}k�� �"��"O�Rab�,C"���1�
��F"OX��Ī$:>D��d�=gPI��"O|l�w���Lu�����ˉqH��;�"O���M�:5�Z�{� Y8O�ܰR"O������>Yu����τ�s4d��"O��yc�A�[(1*M��f?��T"OԠ��9K����퐮z� "O�<��"]3\�j�P5LK.�IY�"ORLr�Z��Y��k�#1^`���"Oh���"3hȹ�)!p>zź "O,Mkp��.%�V��F9Ctp��"OJ�R� �v�����G�ok��3"Oƅ�.7DQ���Z=�0xg"O ����?10�V�J�L"�["O�t ���[�$���&חV���"O�TYюW2*h6YJL[��"O~���Ht����#*�=	�:��F��'w٪�ڍ�	�Kd�)c	;D��1�HٲJ!�d�=j�����˵ l*p��ԁ24@ѻ��I?��gl�|�'�$!Ă�V�`˅EA]3���'@tB�eV�X_��4�I:W���b2j�E\n5��刡LA����	�`���!�9yYDT�%�խZ���d�*r񺜀D� *Y��ۖ L�.�![��P�4���0�l��*���!��ېI$
���F��f�'�$�G��	<"ђG��3t4�F��)Pu��h�+��nO<�Ò��1�yBh�X�vq�F*��t��1�&�U�x��8�厗�n�t�CG���i6P����L>��n�Mc��i�%�v5D"�(<i��n�|P��B�p�9g���Sa���&��pҘ�`T·�q%���G1�������!,�!��Φ/�axR�ߦ<� �(�mX�z~$])��a� �`�T��h���� �̵!�Orh6Ι	\͜-JT眄wU¬�Ɲ�<C�N8澨9��H��!���s���xAAaKG�]0��IH�~x`݆ȓu�HCu@Ŋ-�b�&�Qq�A:7K�7R@�ಯ֟[k��(�G�f�'��.Gf���EW$B\F5y���KV��.Dn���*݌?�n1�`�S�6���X�����C� =(5QC	��<���(D�`��ƥC�u`tp�Bs�$�F�6*��kC#��w*��ʳ'��w�u�%�]�
�ڡ��-��\�Ɠi�0�#f�\��%���R4cS���'���cDMZ�m;D!�m^]dΜ ���L�`��� ������	4�!�$�T���x��`�
t��(q�dG�Q��!��0LƠXLC1�ĒO�`��iP�l(��u�$=�0
O4]�$"��v��9�J'�%��^�8
�c�N���0=� �PB0��=`��ls ��6��@���'���
�A9��T�sF-����4�Aa!�;{V\[�H�I�<��g��&�h�Rp�7
-$��M�ɃoR\v%[�}����$^m�Ojd�d攈c���6L:f�����'�(9�Ĩ	��`��Mv�6*ҒEJ�b������ � ���ē� ��슰(�@�"^sBh�Ɠ�*y��	��.u���ՐEi�y���R�yԒ0
щ��
�Z��䒠pL��/�I%z3v�zr�z�#�	�Y����<�g+R�X��<AR� ~HiR!��Z�<� 
:>��T ���,��g@J��@�c!�v��d�!(�B\8��^�y��.�>�I�)Cy�~5`��ѻ_y���ȓw�@��"{���×0*k\ ��_��c�"�$h�"��%l��<�ȓR5B�+�)n�+-"n�`�Q�"O��rA�I&��óLs˜u:&"O�ѡ��՗r�`Q豮[�w����"O����D�?C�Z�;6�]<��m�T"O(��q�Uk8�R%�
2����"O�)�'f��lF��&*B�*�,1�d"O2p� �(�X��P���w�1�P"O��%�47�`1C�,B
M
2,��"O�tt�2T����A��q�	
v"O �Y&k�<������&h�Q"O�)3a�)Q6`	aC/�zeb=��"O4%����302�{�,�#zEΉ�q"OdS�l�s$r)c녂G���kG"O�p�����*zpu�j�8st��[ "O�}Y7Q��R��d�Ot֥�W"O�̓���o0~e�`�!P�D���"Or�C�ʁ)M��l�� ��p�Cp"O�q1�
�z᎜c�H� dy�xr"O��8hB�о����/fb��"O�a��SC�F�pǫۏXfN<��"Oΰ��a�;%���bQD���� ��"O����C�h�:T+vĞ�[�z%�V"O��r�N�0��X�	Q�a��8�F"O,��r`�#k����ȗ~���f"O�u�VC�;pF���7a^}��"O 9���t�Q��V	)g�ċ�"O2|�2%�Z�8k�)��at����"O�EPT�D�MZ�И�'6P�{�"O*�s#�V�O�u��ѯd����"O�,Z�M�:\�,p�Z8iT^Lq "Oԉ�c�����r�.��N_Z4��"OvuZq� wƴ�'��%ʐF"O��!ਛ/n6\X��ſP �q�"O�]�Q �4	N�� �M�[���4"O|�
GEU�lf�8�ϳy |T"O���I�W���J�&ů\QFy
A"Oh���zҥ�g�[=*�b�"OP)CD�B�iu�\�a/y*�$��"O�cg���>���J�oT
P��"O���P�Φ0��уM�7
�4��"O JN҉�6�Q��D��.�"O^�8�V�Z( @8t��ag���g"Of�7`�*�`�)���W���4*O6����ܱv���
�V�s��1�'e���C�	���cϝ	�f�S�'E��1A`ʐy;Z��1fye����'�Lِ�cwJ��PPѱ$���z�'�81j��p��m G�A;���'��cƊ	#JR�0:'@";�$�H�'|~�DI*%R2��fG?�h4I	��� R�Jt*R�|.DT0&�,)c!y7"O�)�k��v=5��C�?ri�t��'<=��׿��	%I�.IC1�O	6xձ��� C�I=7 ��R_"�8M42[�O@�ib��jg�t��Ef*�0�g��p�y�o��g?�B䉺�Tͩ�)�?H<|9� iU�(}��Cq.U\~�a�+W�T�}&��W(��'���"�1g�h`��+����Ø+}N�H4�>H�Z��a&y�h����GE���K��Eʂ]$t�վ��b�&�w�@Ah"�Ō��]�J�q
g��V���o�J�E���W�<Av��8sD�!�w��*��d�Jgy����dL���"�>,�����	�;|:%q�Ƃ+H4�`�C�f�!�����[d���o=�с��D�I�t=apAڸD��p����{�Z��]>�<aa-��u��Y��)V�8;�Xh�KsX�H��D�5d(�y���G@�F!�g̍.k��s#,-X�`xxU�|��`��	� F���+�e���p�.֊YJ�<١%T�&J�ۥ�c���(T�����O��	�@�&�����6VX���'���w��9\���-�8ĩ(��x�ց[���1%vd�q�I��E��w�rd[G�hW����Z[(�B�'��lĄP��* ��/��u�h�BI��A �#I��R˟4���o�'�Fi��#Z@���j\�t_TX��n��Y
W%D�n�PE�+�!l����@a��q��i��d��%j��^�I���P����&�]�Ipu�fb�f���D�l3�v�c���8^�:܂��51�l�SSY�@�C�^�(�V�%\}�PC�I$	��`��b�K�耺t�F !<U�`om�"A�F&S{^a¢���.Y���4�sޅb0�U�Z�b����u�j�#'=D��hB�+�G�4���$LV�a[^�8ⴍ�t#�/�J�z�cF&G���0��J8 �Kt�X%�@����5���d�9,Wfܢ���6 H6��t���c��y��̒�{�Թ�L7nH��Cv��5Y�$!��I"c�(��F�Q��q�%W�DB㞰����'�-���j?L�j�L�)���0�O*��R�Y�8Ć��k�?T��yC�'�8�"4��mA�XId�<P�zlƩҪDL ��$�B��kE���a�0��~��x���T��sƞ��vg��F�D�b �,D���-̸v�]����(0��A%i�t���;'�i��\Ӳ��Q�����9r�Q���'�~<�
f�XC��b�7\O�	A�%r�����D�thVH� g�iؤ�8��^)d�,�AFĦy��-�K8���q�_�jQr!���U�Sjmke�#�	(����`�f��}�����dȨ�k�t�]�E����ȋ���@a�
�yҬǙZ��BF��Fw.`['*5p�t���.��`͸5P'��v�:M;���k���-�!��
$qiJ��nD�M�!��G�E-D��3�%Ji�A#A+E�3�v�S���<�@L����5�Z����D|�EA�JZ�#%AC�Q���rPEX���=	U͟/S�����AKx�Y�͔.J�x�t���WZ���	�N��	a@v@;��Qfѣ�I�+id�#<i�;.ƈ��F�Sy�O��Q��{�>4��f�!FX�];�'��!q҄٩dH"���Y'7�F��qO]&O��Z�Rz�)�矼
��%�����_�q��\��$D��+��<,��9GK�h�
ݛQ�"D�P!���s�v��@�eF�89�� D����&Ǽ_v@��n"tMR)� ?D�\#�FݏB,�u�p�q$}�cd?D���E��:�\-�fC�S���ڷI1D�xB�ٰJ�=�[��40��L�!�$�PMz�Q�Lϔg�MjA����!�dJ�Oc�)(e�ǝ	�����x�!�dӪ}G
8�D�=*Y>ݐ���*De!򄏛[ǆ�p����x@���&�#?a!�$2�	����7DT��(�84U!򄜫YP�@! 6�������:G!�ĝ3��Q�m��<����-�I!�$<vpƱ�5J�7)R}�흽P�!�YGB�뵁9?�@�\%�!�H�Bx�A��� f���oB��!�^X�u
�@�N�>՛�?V�!�� H�8#�Ϩ.�������H��"O<�YS���@6`�2��<���"OHU�A��_`��,*	�}S!"O��#L*RL����!��n���[u"O�YA.��U���ˁ,전�"Ovyc��ppSS�I49��"O�x�/�t:�h��%/�Y��"O�AbU��eD��
Ts��,e"O�)�V��/)�(b�j�3��J'"O�aCP�2�2H1		��!S"O��0�ǻ�P(r�h3�a�R"O�3 (D�/,
9�ѧ�M��@JB"Ore���L�D0 -8�������"O0DR�����|�*�G��w����"O�����$��xYW&A�T����"O&)�e��x���%�����"O���ូ�Q�O��g�d�q"O�<�P.�DX��J!a����"O4��B��}*8y-ȈD�����"O��FYp���B�M�)
@}Y�"O�i3��$+,PP�6&�p�\}��"O�u�b�ށBl��)��J�
��!�"Oz(c�_�}P�Z�gU�_StJ�"OĘ8@��T$��D��@���*W"O>�s�cI�1R��PD�rQ�X�"O��P*8&�,��Gʞ		@�qA4"O����ZTX��2G*���"O�T8ң��/�QF���]�D"O�,)��		~Z�$SV�F��rA��"Oĉ�J��^��c��X�A�p�&"OR��R�!Z���Ыk� �I�"O��"�ŽT�^�:dM�/r�6(ʒ"O�	bu�R��J�.N_UR�h5"O���Vc#����l��s312"O\m#�L�6m|<(ؔs#f r��>D���,�w�	j�&Gu� ��"�:D�X �/���Ƭ8��?
y��ɶ�?D�8� ��#~[1�2>K���(D�䛃�[�^(��y�R�F�����) D�9d*��/,���BM/~HD��s�;D� �a�Z�H��5���)L�f�2�9D�xa`��b��[@\5B|<i��:D��ۖ�nz�8	d�� i.H؋b?D��I�eĜi� [��W!FdLB�N/D��b�ؽL�V��'l�lE*D����.F��Za!�d��F�z��&D�hI� I�6�J�k�*L�
�����$D�x�����T���3rf̂,D��3EߏN����K�B���� D�$�A��2-��zW���8��<D�xs1 鶴�5&ݝD�
����6D�4ĂT�-�-�]��0��8B�	�z��L�k:@�J e۶)FB�I���p�W�eB� x�W�$:B�s��$q&���8�p@��9SB�	�H�vE�C �Q`�����Q&C�I�� I�bذ�d�b`f��C�	1ne�zs�é�����`�=�B�I�q�D�1l�96eHAk��A�O܀C䉩��L3S͜L�N5�C��m�~C��f��LD��~���&�6QMjC�zZT
�3M%���o��bgvC䉟s��3�-^3k�U�@�	/~W�C�/?L�H�c:&�X�с�8�<C�)� ���T´C�uC�m̊��l�C"Op��3�;v�;Cl�{��љ�"O��Bu�ҏ_o� �,�p���S�"O�]��MތH/tS�!n�x"O�����,
�Y;7l�a/�ę1"O��hW��(F��Cu���[!"O\���C.v�I�'*<���"O��#�P����"�$6.�2�"OI'$D�z�x�x5!D�h����"O8k�@<DZ�$����<k�"Oz�J��;|C��r��{G�!"O~)	��F9k��|���SJՋ�"O<)��G���6a����aZJ	Y�"O��B2�;1�A�a��"���
�"O��{`@�)�\��/iwԜ��"OVؚ�+�b# %P� ���2"O :D�4K�tض���9kBi��"O��jo�������4m\2�ڇ"O,ܰ`Ʌ��89�����9ؔ�"O!���?^�ҁr�(�Z��<3"O`@�C��6}�l��B"5���@"OF���2 ���K"�A�!���j�"O��ѱ*�+g(8��oB��� �P"O�}��͈���bcy�"O�0ʷ�3�:�b,	#(_\�HA"O@-y!O	a�)4="D�[�"O4X���}�RHt��'�]ʢ"O������Lɘ��ۋ�I��"O��Y�A�|�*�8D�� #��Mb�"O�\:U��+��m��'�(�� 4"O�]����`�ҥt�ɉ�X��4"O^�Kd`�,��m!0e�F�V���"O��"񥆉|��,P��FPt�xA"O��' �:�Zm��E%29���"O��A!IQ�����4]-r90"O��V��'�\����w0�{"OVɋb�-���c*�j�$*�"Oh9�Ř>*�����
�z�����"O�ZÐS����rE~�\��"OL�y��Q
��ue ]�`�D"O��4͵EO��aD
 0��k�"O&�$R1=t.��֗S5��� "O$Y�a��6xA���1<�
�"O�E9���$(�9�nO$_>.<h�"O��8g���M����a*ļGJ���"O�E���Lrb�8��U;D� Y��"O�x6�ҜX��a㗢��� �2O2���ٵy&$��1���$�1 ��ɫ*ϒ����,@�X�$�V�f0B�I�.�BMjs�_&?�����('3ZB�o�n�x��=*}�����L�h�C�	��� o\��Z-)��Ȗ����(?q��U�~}�5��M��`�<1ԌˊX��-q��UQ�H�1U�
w�<�a�¢��@` "�k���S&)�l�<�*j.g�=�.Ԫ��_e�<ɶ疼KpxH2'UM�ܐ��J\�<�rُNHcƝ=S$pZ�bRX�<�g,֢?%v���G WE�	��nJj�<���7h�� ��DP��	d��b�<rDث��E�2�r�,^j���E{�G(�����"	�2��x����u��<q�����'v���yU�C�2LP<����&WQ��9�V�4I��ا(��$A�أx�}z��Z��76O�9�'
1��?y�>0nԐK: ���E��E�f^��D	�����?� ���Ԉ;?.�Ivcէm���Z���H�'
v��i�'`��p�A�&��Ua�.��Oڹ��i>��\�`y��S�/ت�����!pz��%�P{7��o�S�.PX�g�ݺ>��S���'�%�'���a���ӟcԘ����! �x|S`�ٿZ�>����(O?1�WDϺd�	�	��ł�"ac�<��?3mZ��kMe�2]
4*^�<Ys�  ���'eV
K��,jEq�<�%[�M̆���d��#u�� ��v�<Q�O q���A(��(�6��G�u�<��d��*��=�t�zA�^p�<U�K�N�0��q�5JӁ�v�<���%(�p�ڇ�w�p�³#�r�<A�čA�Mh/	s$��+��s�<�0�\�P�2��@�߂��!BIW�<�� Й-�0�c��,+5�CQ�<�AI b��e�,j�x��&h�<�r�S��Hf
�*�T�#ĬNb�<�p�O��t���n�"t�ƽ����C�<!4�TPj�!]:�����=T��J�M׊GP�[��(1`��,D�$��h�4���CF�0_?��;�+D����n�?U��P�a��t)�	��(D�v�i�ê���j,�+^Rܘ��'c�0�����8�ʹ匊+j��x��'�\	/Cd'���Tˉ8_(rt��'[D��@�1~t��3����2��'��Ĳ7�ù^�003��%Py�i��'z`a�� ����oV�xXҁ"O�Q��R��m2���e{�"O~���
Ւg|��f�OV�8m��"O��{�jP%H���S�|x�0`b"O��"��t[r:�o#O�\"OT��c�޼G�D����G��};"O<� "Q�Ԁb�G�K��9��"OF,KՇU>�\tq��2\{�"O�Dį��@�y�i�6)�NܢT"O�3�Z�i�D�V��D�aW"Oz��S�L� �q�����p<�"O*Ⱥg�?}�x�Zu%VT�\y�"Ox�Z �I3"\���� ,:̪w"O�$U*.�:�c�@�#m���@Ot�<���4\ܦ�S��R �e �iF�<�0�<QLxPc��X���t�C�<i���q4�rD�O�S$BY��|�<���W|�qhEF�	(�\��NJp�<��-�8vA\�����f3�4��YV�<IuaN��{&b�*�n!s��\h�<���:H
fLЙ�4���Ίm�<��@'NO�E�D
H<�!�:�	���S?�b��v�C�!�d�;�Ԑ˄HG�a�Tat(��=�!�d�)U:,hF���p����>�!���f�p}�$+̀{�d�<D�!��;�p��C�� n��i�cܓn!�1y�J�" ��J�����4x!���+�ΐˑiBS����T�'
!�B�=^�yжK��+�>i	��I�X!���(}���#T�2]*6�1a͌!�σ.2 ��ߒy���cj<'!���x5f�s�)^�+׊ZD�C�{�!�$�|O
͡P#�M�E���	>�!���
�3qO��e���1%�ՐF�!�� �,��l�0���!"�M�!�� �4�se˥H�N�s�)��aQ*��"O�ɘg�ωS��E�O�{1Δ�@"O<4BfIE!g��0���DЀ#�"ObT8��Mӄ�x��>�@��"O~��@��Jy����(��+�"O�ܱP�GC�0��0[ɪ1�"O.��"i�&E��ð�>�.�k�"O@з��&/6��j��LĲ�"OX�C�jB
8��i�>��9;@"O�ҥ�%HcV�۰g��i�DQ "O��`Q��6Yd��(��[�B�Q�"O�lySǅ\��j����\���p7"O&��`�M:����83��ɉr"O¬�0�)[�X��W �F"F1��"O̙��A�"_ܲ��ɪ��/E�yrN)
Ll�����	�~�� ��yG�L<b��d�BVI�`������y�
ڀe�$Qum+c�<ēE%Ԍ�y�X"�YG�C-^Ȇ�B%O*�y«��l���b%l�;f���8 +@�ybM�2<�LAbq�-
^�,��
�y�i�d���r�9|�´3G`�?�yr�7|���8�h�KB�K:�4�ȓ_nq�1�ѷ	N$萦�+O���ȓh0�"�����['Z�9[�̈́�~s��b��!�r,a$EB�2�:Ʉ�,,x2V
����i����%�0نȓ �%8�mX*���V�R�5����!!g	7~u�����ޒ
��-��{��T�&̂��ʔ�We�)-�l���$�.y�p�֨Czm�f)�r�L��t�RI !��+;�4�F��ni�݆�7V�m�"��Q�F��e�%���|g�� 瞹+�A�SI��j �i�ȓ?�*	A%r�lx�Ğ�_v�����s�K�����E���i�`���-��1 !��R��72)h͇ȓP�Ј��ŕpf�u�i�	hE���(yy�B��WQ�|�'���8�ȓj�"�Y��XZ�P�(�*n깄�~�*����	�y���TBD<XSd�ȓ*q^��m��h!<0�&��k���ȓ���1���{��)��ί>M(X�ȓf��" Z�h�b�[�wX���G����׋E�7���$Ҽ~�怇ȓx\t�h`-��7P$�s6"\"h��@�.��b��	=�|�U&�5��}�ȓ7b� �I��T}��	WKP�r�J�����QCːx8�6�3A��9��b�� ϞY�at���捅ȓyŎX�s�R�q�X�x��A�5����^�bd�d�@ ��bBi��<�F���elv��S,�gꌨ*��� �Ą�a7�$
���T�,l�րB�4���qr|˂̀[w��!����y�ȓ	>ژ:�I�es���.�(Y���ȓ_nD���M�8�%�P�ը�2�����cGGD�J�, �Rl�ka*M�ȓNX�z��߁	_$��jӔR�\���0���g�TE�4��c%��sC��ȓ_=4�RDwfe��KW+E���ȓVs�T[��?/����R/T��0��G�r�J�
aĐe��@�7rp��;��Y!	�01�A���S4de��S�? ���O�>+�TMc��	3LY"O~��#cP�Qy�tP�h�
N4Y2�"OJY���N� ��8�i@�dhm�"O�e#�AYN	��&ޮh슑�#"O0�a�k4m�~�c(ҳ
s�}��"O,2��D1,a3L�:;�Q� "O�u�L�� D��e�"Qƭ��"Oޭ[��/�>�D��RW
̊A"OX| f��&q�8r�M|<\�P�"Ol%�r�-%�uʢ�!4-"�z"O��pʍ1m��M�D�A � C"Oބ�IJ�,a��Cm޲|z��"O>�+�(Ē_d���'LJFRF49g"O�8�FJ�{A���*�<1�=�u*O<e�#���KO�M���f���
�'=�Q��#�o���D�r�ؕK�'*|H���M�5vјU!�>�&P��'��%� �!z$t�����G��k�'��G��%�����a��P_�eq�'�����	Ю6u�� ���I�H�0�'���Bl�=���1� ҕx^��z�'njQ�#�!=�TE�F(H�;�xd�	�'�0�ڲ R�,\�+#��?3���A�'��[�l�;ޔt钣%1�XZ�'}d=q�OT(+l.������(Bd���'H60���̅
�;�!V7%:&���'�jh�C���&<0Hpd��(��k�'&F�;�Ζ�5������$���#�'8
0��j�c�m��5p����'�,	#���d
d}8��ye�a��'�ӄA �"G>���mϚ{��IB�' �����C��V8��d	@�G[@�<�&�t����7P��A��x�<�b������(�i��8��ae/F~�<a�fG�`Ɇʧ��
7�N��ZA�<ԅ:S�6}��A�npj���g�s�<A�o1p�u�0
8�l$au�Pl�<��N1Rm켁`!�%V�p��	B�<Yq�D�06U�a)N�q�v�#*ST�<�E
�
A�]hP�L+"pP���P�<��ŋW���	��I�x���+�g�q�<7b�'Z���he H��b��Øm�<9ԅ��K�\T�F�ucd�`��!�yI.~�8�I�G_
���
��y"�,7Cz���^?B� tH�hܒ�y��7C�\����F�"ȑ�V��y�%SA.���J2Bi� � �D��y��b�)��CR�:����ǆ2�y��D+v�^���AL;�ptYrb��y���	�@ب��S�d��ac�B�y"	��j�Bd�T�^�`J�J񫑈�yRf�.j�1F�G�j2 ��֪�y"Ɏ�=�e���K%��M�u���y�fD=���S�H*O˒���I��y��$����hKS��� �0�y���[����$Ets�ّ����yR/�=��Ҥ�O.W2�4�_��yRf�D�n}��K�op �	��y�j�)5�n��FJa8��K�AR��y�Ȁ/I<�0eŔ�{�`��P�y����f1� ��M�k�hI��ˋ�y�oA'!>������dq��T�
��yR��zGJ�B��n��1����yb�?%�R �7.������y
� ���ЂE�'�X�+�.;��2"O0z'�T�[��U�K���6�"�"O�dxV��	�^A��*ɡe��I�"O�A�VgV�m��u��	�$DB$� "O�=��E�#���
--�\ �T"O���biQ4j��-�t� V�z�1�"Oaa�bU*�RP;6�� ��٦"O��X��ǆe=@
�k�=� P��"O�I��6l� A�0�
, �JQ�"O
a�� �Z����g�'g� AI�"OĀ�f:M�T-3�
�[�\�"O�����Ǫ?��^�D���4"O��x�
   ��     �    �  �+  *8  BD  SP  �[  )g  xr  t|  <�  �   �  D�  ��  �  /�  q�  ��  �  ��  �  ]�  ��  7�  ��  ��  "�  i�  @   * �! �0 �7 LF U ^ Pd �j �p q  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^r�Bэ]lr"����Υc���!� �u�e|���ȓ_�}�㧟���\a�R�i��p��>�
H�?Дk ��t�Tلȓ*��5�&5y�d q%G�=QG>ĄȓGq�E@ÀVV�p`!��[�H�h���s�`HqH�Y�T}���ńi��=	�G$D��@1ib���eG�6�,�r�o�0��I�&��p�W� =O�AH�� ,P����D֪���8"s���G
�oºap� *}�C�IYW@	Pd]b��10#_� ��C�)� R"0)R�o"\�"e���v�X��"O��� ��)" u�g��w01��D|���On"�q�Z"f����m�,v�M��'�n9Z�HVYڢШw��)�8���'EИ�Ei�
G��Q�L��Z���'}�ݹ��f�i�6�F(]枅�ݴ�PxBjTWNX�Q꒘L�L�yV���=9���P}r�'[:��ƌ&)�D��h�X�� �'#I&�;#*��iYd�&ъ��Mh�OaV�������W���hc�!
�'�0��L�Hz1G��o2&R,Od�=E���N�T|v�8��?q����bI,�y� �+v�.m֦dVA���8�O��󄏊�j���]�,�̭���M*ޡ�/sj�=z�A��2oB}s��>��}�ƓJ�L�@&O!5ʀ�3�μx���G"=OС�~�q��5+�L\k�,� 0�~�q�'�z�<�U�2PI��|�\��s�v?���)�'^���k#��_3���d�ђD'�����%�Y4hD]��E�g�@���>�4 3Ч��!��0�f�y�!6D�<B�	A+�XE� AUj��R��)D�Pе�	)���q�Ɇ�`L�IC�'D�����R��$�� �h���bB�$D���-���|�⃌�b�t��&D��[���� ��Y�5	��3ru��`$D�7�=%o\�B���I9 x�@�7D��
�.�ag�� 2��7n6�r �4D��$Q�>�0�*�y<0l��0D��I�G�yPz�1�� }�q��-D���m�����c��L2�9I%,D�3�
_�B���#d�{�/�y��#��Ȱ?I����� ���.��ه�	{��t�M>QUKI�p�=����d|� �)�b��?�Ǔ�L:�D_"9&ScdɈ0�$h�ȓi����f� +m�n���k�2d��VϊI�.�yt
��-�;0oj��=�ۓD)p��S�XW����%ٳyyJ��ȓ#JJ�{m��:N�Xj��sb<ȅ�.�0@֦ӏr\��e�K&���w@�#g�^�;�1���V�?E�O���D
�n\@JP��Rð���&ء��hO�lT�f(�)���j��.5��j�"Op�s�Oƞ5`r,A�
�M���6�$#��?�,�J�2�)R�c�p���Yf<`�ēC�v��Q��T��t`w��2QϚ��v"O���� C�F��N��$����"OH<i��LC�(�sƁ%X�䝑�"Op4(!�EU@V�Aĕ�R� e�',Q�88�,�v�����oy�AVi%D��C�L�/H��t�`�F�H��y�N#�IM؞\�P
x�^<��žs;|�Te!D��Z쎏Y���y��^ :H��9�<D���� kf,򠠛�&�N�`�:D��J��0Ќbա�6��6�7D�h�s+��i<<aY6@Шԑ�e5D����}���1�L���0��0D��Q�hݞ(��DKg�D�*�n�p�E*D���T�R`@$���u Z���E(��o���(i���Y�5�H���D�C䉎L�10��$3���g�..����<�II����u�Ŵ
�.Q�� ��#^2C�əNBz��)��'��| �
?s��B��E8rJ�Iȑ\� }�N���B�)� ��SRk�6.��� �T�V;���6"OT��2��'@q�a <���"O��I0"Y&; ����!̈́KY�(A"OZ��҉ۼ9�u�@��~�h1a"O8|��42F�93�HO��86"OT�:�$�9P��v'Y9+�|1�"OB�Av���Q<��)�%�3B��ɖ"ObEc&�� BP%�f�͂c���Ys"O�aq�nƂO�j<��N�:��a�"O����K��h�ԭƁ/.\@�S"Ol�t錵x�Y!�Ưq���c"O~9��da ��c��9��O(.!��	1r�t�'���LY�2�I&!��B���D�+�m#2�ǽ_�!��)U"DL�7jݳAqrQ0'
!C�!����_���Y���yo�4���?6W!��ˢdjxEP��L�
��6.Q�|7!�J+#�|�X�I?"Ah0y���P!�Dp�L1��aߥJN|0Y�C��z-!��(
]��� �A:��"��D�!�DùF=��f��{�9�g�ڷH�!�H&+ڌ�aW��*J��� ���@�tG{���'��c��.L�H"2�J�:I�@0�'ת��Q��5H����1��5`,��'��BǬ5R~��E��*G�N�μ�p<��4�MSs�i�� qGX �wm	�w�V�  G��n<FC��'>�TлH�
,�Z�(�) D�b��n� �{��D'Y�ar� ��3t,��5�Ђ�yB�Ds�c��J�:�9�s���y"��@q�C�V�{8�	�����y���M�\��B�; YJL�"��y���3��=0��p���R�c��y�K!0t�Ur@���@آud
9�y�	��� 
�@3f�0�k��y��@2W��'C��9 �Q��g:�y��ˣ5X��{b���	�������y��M  ����P|�*4�����yb'�&D���ʌs)BM�W���yF��aH�	C�@	!�p�f���y�(�+x��6��a��q��H���yc�	'�� S�B���A� �>�y��?0|I�5�ʗn6�2����yoј�Q�e�i��l��͞��y�c��QҦ0rt�	�f�������y�I�2D��G T�YHD���!I��y2��>G��8�O'M��ث�9�y���JZ�	ِ���H��D������y��P0%`Ν u�]�F�v�AVǐ��y�ҕb�(J�	��`����y�m�1�����j�UJ(��
��y��0�*iPFE,�V�g�Q��y���_��V�L�w���Ə���y'U�H��"��	6m2±�W��y�!ײO��u�'	�:c*>�I&����y��	V�f%B��΋U�������y�mE"\�cQ�H%S�IL��y2K��&H�@K�A��Pe0���y��[*�� �VP��w(C��y�ʖ�Sh�����$i(uX'O��y2[�@f��F	��>X�1W����y�B]<l~�T@e�D�@�|�M��y����4HsM
12��	0`�:�y�gÂX̠Ke��6+�<Q� O��y����LRF`���RY�q�f���y
� ��� �"i���"�ҡ���Ѣ"O�9��#I9��� �J	td��"OT�ׂ�w 4f��TƽYf"Oz-���ˢ8��Hpю�E���!"O���ƨ��?��
���6/�#f�'��'qB�'�2�'Wb�'M�'��������"@�H�S���%�'���'Fr�'�"�'�2�'#"�'�%���B�'�ܻeHY�E��I��'b�'b�'�r�'@2�'�r�'�4�`�Q� ����d�Qj*�'\��'^2�'p��'�2�'j�'R�{�|f�2e��y[�1� �'��'���'o2�'
b�'Q"�'��y��k¢	���]utR� ��'�R�'pb�'�2�'
2�'���'r6M���a`4�a��3`6�H3�'/��'���'��'�"�'?2�'"��p�S�R��|VjD�yM��Je�'_2�'���'L��'��'rR�'E��2 ����t,�&�C�un�i���'jB�'���'r�'���'V��'�<2�M���N�X���P� �d�'���'���'��'z��'���'�أ���Q�j��G�S�:Ed�1��'r�'o�'YB�'�"�'OB�'4Msŋ�7$( �ők�]���u�4�?��?���?	���?	���?iE%VH��H b(U$��Hҗ ���?y���?	���?���?���R����'�c%Hd�T�T�Q�Ԝ^��˓�?Y-O1�����M�
�_X�1�A�#�ܱȧ�"b�l�'�R7?�i>�ݟ�h�i���|�B�+|��+Ю�۟X���ynZr~�5�|��Sl����?]@�8EH�]x�� Pm�,H�1O��D�<	���ݞP� �s� (n���,�#P�L1m��b���j��yWۉ���w�ؘ[l���K�^5b�'B�>�|�c���M��'�9t�T�2 ���)��t�'��$P���B��i>e��!H����aQi����D�L�	Jy��|"}�*A�����@����CW�]��c�aׄ!.㟜�Oz�D�O���W}B�%g���� +����CL�����O�}
����#31��y�#3�����23�� �+B�n���@��>,������O?�		��l��W�7��Å���6�N�	4�M�Ԋ�A~��kӢ��#�r0��/�	Ha��zLP*�H�	����h"n�Ħ��'��)��?��QB��^�↤V����
�.$�'��i>1��p�������>��0�*l3�����Z���'��7̈́Dj�-�S��O��$�������O�DF�F���1��3u�|	0��J�`�t���d��xmZ��'���'@L]�+�t�hs��:f���`���h3��%G
�3�HI�4|p�Yw���'K襔'G�9�	�,x�Tk�eZ�tꐁ2V�'��'	"�'�\�!��R��I2h6i�bi��;d�ը���O�X���ß&��ByRr�.ln���M�!K�z�X�h�y �X��T�u( s�4�y��'��E�#a��?���O(�	��k�ƈ2�R�*�톈��E�E�<)���?���?1���?qK~j4)W(W���� �j��y�ʥk&pb���?)�%M�f͌�N��S����uy"��k�P�S�=(���0�ā4��7�V}B�a�.�l��?�1&�֦uΓ�?�X5D�̼�'���Ha�5*�+=�����O>RH>-O�i�O��d�O� a�H��w��ٳ��q	P�p��ѯ	sbT�p'�<ױiLZ�j4�O���'����w���V��65k��Z�֦e��'2��X��Ҧ-8�4��O��d�&�|�ITd˲USv��7m�!��{"�­\ٶT3�O�)���?YfF*��H]H|k�E\x�ؠʳ�B~A
���O����O��<9w�i>��� �QV>̛A�ܡ6}��z�*�;��	9�M�����>qS�iypi�g�?hdE_���c�aӂ�D\� Ί7y���	�5L�h���O�
�
����)�r�͚ G�dy����D�O����O����Ot�d�|T$��)X�**��Zv�Ss�Mdr�6̎Q�B�'fB���'�26=�86l�i�Щ�L���1;s�/�M�w�i��>�'���ci(���4�y�O(3� �A"Ö�8w�8��*�1�y�R�$d!���l��' �i>���;Aծ|��/H�a���UhΒ"�F��	�l���@�'�6mY+ZnH�$�O������3Eʚbp�u� &�*�0k�Om���M#�'��	�$��1�M~ƽA�LR�t��I֟0�$K41X����4?!��lv��Ω�?�/�Pݎ��T�A51���[�(�?����?����?��i�O���'�
���ը"�M/Q�Z�SJ�O*�m��-渕'"�7��O��O��z���s�ޠc,�qDl�;a>�d]�Y0ܴ�?q���M��'T�a��b��!�7MJz�3��r�͙Z�����|RR��S�����ݟ��	Ɵ�����8!�Z�b�BE�C���CŘ`y�n�O�!6�'�2�'��Sx���||n��DO�+��9RE2j��	��M[��iZ�7�Vs��?	�ӡF@K��Я]��`���H�`L�5a\�T!���T�Уk���u���O���O����6��c����-i�Ѐ1Q���Zy��'�b�ҧl��Q2�'(�?���]�T�h��>��-��E�$↽"�7���	�<$���۴q�Lk��w���I�p�m��} �Ӷ�,b�Ha��g�	�d�'"�a��M���íi�e �@[�J����Z�{�? ��;`��Lߘ�)3A�+Z�(B�i�O\�D�O�$�O��d�O����OZչf� |����7	�&~���c��%>N��49O���OF�n�2�$�����Iɟ�Iޟ���`T$8fv`R�,8l�r���-�?y���@�۴*-�V�O��-�e�i���c���p"���(a�k`30kg��_\a� �'�F�$�d�')b�'�2�'�a+6!͉]V(uC��T�4z0e���'9"Q��x�4;����?���򉊮-�eY�[ g����DK�|s�I���D����4}Z���t�O[@�B��e����dܖMa��ҢԀ!{����a�Z��?i��Rƺ���'`�	��8��Q��<+�W�Y� �	ܟ��I�`�gjwƄ�	�L�	�?i3Yw�L�;��ɘ'�(����X���*3
�D?A����'���,J'�2�lӪHR�,�]Z,�c�%fxJ9�d����ڴV�*�ܴ���3_s�'��J�Z(J>gU��S���;Ԥ��`yR�'���'�R�'�2_>Uk4O�[΀Ii��S�Prh�'�M{�Q0�?���?��'��9O�1lzށ8�F�.hz贸 ��#Vx`��� �M�P�i+��>�'���� �8x�4�y򬞰u�ݣGI�>]������y�َz����	6��'��i>1��4p�6y���\ju!��p��,�Iן|��ǟ<�'�7�J��8�D�O��E�J�0�W�-�$٧C���B�xk�O�=n��M��x�-I�{�D��W�ՇxG�A���F�yr�'|Xݘ7��h��Y���S�/�f���8��͝:@Vv���O��UhV��L��T�����ԟ���Ӽ�a.݆L��wdιx�`բR&�.�?�F�i<�07�'W2�|Ӧ�O��4�Q{�
:������G4�c��OX6-\ঽIڴa,
۴�y�'Y��꓃��?�f	ߺ'�z�Y$�FmhH�s�׹�b�'c��'tB�'��'%r�'�2����!�	N"n*j�&�+��'%p��J���y�'���q�ܩ�#1O����1�9 L˨�4�U��4.���,�O��nZ �MS4�'@���O*�i�v�C�fb*��`*A=VW�\ �fҞu�&��s j�X�O6�9qo�?�?��!�$�<�U�3]<�YA�I�/0�����jń�?	���?��kT��������Y0�G��\z����x(� �A�$~���P`N埰��A�i>9�'��7���arݴs?rԩ�h�*[k*%�n=�P?5wb7-v���ɼgפ8���O=���"��f4�ME(MTx@��;~3��g2OV�d�O����O6�D�O�����"�*. ��ഋ�P6v��Sc¦'f��?���i��I1�'���'q�Z��Y��9\�$L�3 F]9Z�1��L�M3�[���ݴ�V�Oq��3�i���O�1b!͌6+V�8/��$)D�ap�Rv���"��,�0�d�<	�Ӻ��Ov��'��˲>�p{�!� ���SG/�=���'4�/�Ms��F����O��������K+P��Ò*��?4��rF4O��Or�$���	�4\���=��8�(���Ӊ60���Ob�"�����$j��'?ͧ$@�����
�R�P�-��DE���-'�`�3���?����?)��|R!���|-O��oZ�w��CE��7MmBc��?�z$���t�	�8�IQy��'��I��Mâ�A�#6��KE�g@��C`�.l_���f�"�* �m�� 72�ԡ����OL��XwnP�J�V�I�l��4@��'���x��ٟ����|�	i��aKߤY8�����#��D#S6�\����O���⟼�H�?�����O��]�� r�D?�(z���Fm�M��iG��|��'��ώ�M��'��l1T���N��@��z�2�'�*p��,^ş�k��|�\��'C��!c�	�9�Dt��>2<��ቁ�M�/4�?����?)�(A%e��B��S)J���ir�]��'�2�U����y�.�'����o�8 (z�Qw�N�f�ѳll�T��u����M<=�\�'?���Jğ,sU�'����&l�I�t����(B�|�4�'���'/�'��>��5T�2,��AV�]�N��Tg�V�Fh�	3�M���	�?����|��y�ė5:����iD�Zh��梏�y�mn�|�l�M[c#X��M3�'"F�l�@�S�5hvhq���"��mi@�fxjYxW�|RY����ܟD�I���	ܟ8�caߟ_�pi�`�  ,r�adF�Rymd��;���O��D�O.�����74��(Z�%�"��)�gO$g�jE�'Y�7�Ѧ���ħ�Z��P;L�*����VVz�9��4`�HxI��.n�"/O�a�Å�'�?y`�5�$�<��D �Y�@I�To��7}<�(���(�?���?���?ͧ��$�Ҧ��^OS2��8���B$,!��Q�H \���r�&�O$��@v}�z��mZ$�M�p�uMhT�!D�JlTM�&�@�g����4�yB�'�DYY�T�?��W�$�S�߹T��>`���B�
ſW�Υ���q���I�����Ꟙ�	�����j�4s#`�rwkYw�.�r�@�8�?��?9�i���'���'��'~^�g�0��H��C]�D�vq:�uӎ��'�7��1�J��Ln��<���;����䌑!jϮL���a�$,p�i�*X�8�$�4�?.Od��|
���?���
�*	�� W�.`X���1���9�xa+Oj�n�Z����ڟ��I|��F\)�\�C�A�/�HPi��8�y��'��П�l�	�MsА�4�Oz��Pp%m׳N�����Z):@q��`��r�vE��O����:�?y%=���2�v��F��=a�h�'fMQ.�d�O��d�O�4���D�O�`�vJ�<!Czݺ��_�t80#����'���'�'��R�|[�4� @�tys�+f���Ў�T�i��6�J�O�*7�u��
� �&3�l�C�OC����� B�����Lh!���)=H�%iǰi����'���'f��'sB�'��t��h��O�n=�Y2����a�޴O`��Y��?����:���?����?�;\h���1��#9���'�Y�o���׶i{�6-	Φ��O�	��i��K��6�e��ȅ�Di����\���9J{�dA�A<kb��c�IBy�O ҢϠh���C�bЩjՄT��'R�`n�'n�'8剶�M3�E��?���?A��s�i�U�	�f����+��'$>����%|�.'���U�B(s�@(����)ZEL���l����k#�A̓�[R��'s�d��2O��.U؟,���:9��`��J"dH�ƩRПx�	۟0�	Ɵ��ɂFAU�g-U�]��21F�0ƀ?{2���,W1R|���ɟ�Hڴ$P |�p�B�ͧ�����S>{��|Z�m��q��0
���	��؛��n�*�nZ�}	Dm��<�ڴ*FA1��1<����Ԁ��hU��&mU����hq��1EM�'��	ӟ��	�L�I埴�I�|���0�̛��I�ԅ��q�<��'%6MX-h�d�O��,�9O��엠~�P�S�� y:�cU�Uc}�dd�
�nZ��Şn�z��!N������B>iJ��8@�ܐS*O���i��?�CN!�D�<��	X8ظ��	�]�����B�2�?	���?��ӲشIc~H�*O��n�yǖE�5Uz��s�kU����s�������MK>��}��	��MCd�i�R7͜A���S$Ŝ5R�QR�=O쌐#n�>�៘�g�I�%��DI�iy��O��%5zD\��bJ�	��4S�C� R��'`��'sZ�v�'��ϟHs��Z�t�2x�d⟠sF���mΛ�@̗'���iӎDC2�8�$�Or�Op��䇉�SX�K�����Z}��'��6���=�Әgq�tn��<1�40���S+�&NӔ���K5����W)e�XU��\��'��I��|�	����w�(�r�KԹ@�d}��C㐁����8�'Fb7�һV�����O,���|b���W�ap�Φ#��A�a�o~"ǧ>A��i�6�UC�i>I�?S樭���׮)'LH� ��A��3E�ڞ$$0���b�wy��OY������M&���Tn�>	Sէ8ɢH��L�ٟ,��۟���؟�ӎv�<	�	Ay�uӦl��������D�]���+�hOS�d�$�O���>�d�O�ʓE���3� �"Aa�1]J1�V��;[�6-��iʀ ���M̓�?q4(����QUJ�7��d�"	UzYZ�,#s�i�3�,�<����?i���?y��?�)�nP�`L�x�V�;A�pHP�T��Ȧ!y@*Y�d���$?�6�M�;W`|�P͊�U�At����IqA�i��7-�U�i>=��?��7�s�P12��Q�i�����
�C�nH�d��p�p���rȰ�Orʓ�?��^�6a��*B�j�D
5%�y��4���?����?A.O~an�3X �	�8�ɧY)���c�ס=
�}��{	lQӃ��~}B/oӎ�m�&�ē]<��3����f����4/�z���?q�k*c��ūn������y���^ft���	(f
�P�I�8D���>6w����O ��O.��4�S��5�	�7u"ݡ�1#'6@���>{�� ����?YaG�ğ��	���$��s�}��e;�2 J4�B؂7���=��ܦi�40���gސpE��>O ���-C�:�Z�'!#��x�)��f�vH����K����a�=���<ͧ�?I���?���?� *�6)����ш�6T���������������ן�$?�,���$6W~uzI D�
��O0ilZ��M3�'}�O��$�'y��R�oE;_* �2�>^�� x!	?�V��OR�!�.D�?i��+�D�<ɖkA�.v(���+D(>��k��Ǘ�?���?A��?�'��DL̦y�����(Q�FɵIXșYGH�Gڠ!�v#j���4��'�&�
����{Ә���x�h �$�Z}2��C�v�T��,mӞ�Iȟ)�\0��K ?y�':dk,^�<�|�#�o�H{z`X-;#����O<���O��D�O��3�*h[L�	ӎ�N����)3>����ߟ���;�M�7!�2������'�TH`A-/�r��

a��L��<ɪOT,lZ��M��ID��޴�y��'h��i��!���X��9b�x�c�N�Q�.��Ʉ%m�'��i>��	ן��	;�v�*��!Ԥ����[�D�K������'7��k���d�O���N��Ǿ(:�9����[�l�i�䔥;���ON˓�������i�6��	�8Lx X!)�.FM~P[�&��\���s��M�8���<�S?���O�I�;�)@���&�����A�%B�8��şd�	��,�)�SGy2
h���{��c���iA�A�m�����L_�{�˓o���d@y}�#s� �fR�g��
��2���+���I�o�`o�<�O�tX2`��Ft�'�n���o�#O>��!c�:6b��'���̟D�I�p��˟P�	C�ԍ������1�D(��pA��(V�f6-S�2���Op������<A���y�ɗ��!S)��Tys�eU�U�6-��EH<�'����_И4��4�y���>���$�
Y���`)�3�y�-Q��v�'!,X'��'���'*��� �+[����Ŷ}(��'+�'�P���ݴh�X`���?��6^�%p6��K%���&R�h�N�0���>qb�i@6�z�P�'�TL�p�J0A6$UX�F���t%�'Y�FR6UI�.k�B��'e��G��$rQ�'��!�DҬ=����5ɘ�8�����'�'�2�'��>���|>��S�
B	 p�W�f�F,����M��K ��d����?�;먨����52H ����X�p���e��!�M���i�jŹi���O\l�Te���R�� |йW��	7���OE�n�`��3�/�d�Od���OT�D�O��D�Ob���L��i����A ����[g,�D�O�P��a�>���O��d�����1�v�d�ɣN��<`�I�/�½��ԗc�l�B�x�ٴg2���x�@�)�|*�'�@� �����R$���(�ب2�-����dT����Ofʓr@	9RÍzR��qEaѠ@w������?����?��|�(Oj�lW�����fg��ӗ��x�5򕊛�z���
�M��bO�>i��i��7͟�؀e7�\���ʜvi�eb���=(�n��<��Tx+���0�j-O@�i����AX�G�� ք�>fXyf3O����O��$�O
�$�O:�?5P�$�p�@���JT�:� �g�CyB�''>7-�ͧ�?�w�i/�'p`�c�SF�J �R��&By�}R4g6�Ʀ�8�4�b$CL��M��'�V('�x��A�,�Re�BƏ;d�]Qt·�x�Ҟ|B^����П ���|�T�)	��lP�ʹ}�r�8����I@yjӨ���O �d�Ovʧy����'`**��Pɖ�~�&�'��N��6ic�8��Y��?:F"��ḗ+_+�����ϱc��5Į�{�*���W��O�UhM>����oolyh��ȇ>5�ġ2��"�?����?���?�|�)Ol�l�-=��3F_��감`닰
h-����zykӔ㟀��O��l�1a�h��5� C��D@��M�0�0޴�?Q�Fڙ�M˟'R��c�u���DS�U���U`[�m�3B����O����O����OF���O����O$�D��@��Qa�ֆm��M���1bDǍ9f;�?���?ɑ�i ~U˟'\��'?"i����H�P��lt�Ua'ϊ�E�i�6-���
������?��S?X�(o�<�L	�]��Zf
Z�r6�����<�/D+v���$ù�����<���Fp�b|;p悋A��u�"�P��Jߴ;�x�8,O���(�>�[4�?{$╳t�G��t⟀;�O��o5�M�g�'&�I)� �چL{��P��	Ӣ�	��p����
�>�bЌSzyB�Ot ���4N�rc^~5=3��݌zDewG<e�'R�'e2�sށ�'+�[:Qk�+�(Y���d@P۟�	�4R�$�0���?i��i}�'F�w:Ј"d�C�]�왑��*fN�0�'06�Iצ�2�4K��kܴ��d�9{�v���'^�.�z��QV�̈jT�$m�[�D;�D�<���?y���?A��?��^��h��IW�Kj�؆(����dM�]9�Z�;�2A�������uJ��'��"�a��mC�-4��d�Z���Z�PߴYa�f�u�X�'>��S�?�BQhD�<Xj�r2
��:��<��gÐvE��c/?1 �A7���䓵�Ce��yP  2v^��8q��� ����OJ���O��4�ʓv
���t��R�pH`��U%��$�B��\��n�^⟰�)O��v�n�$$ԋ
vQj���h�
zԋa�٦%�'~|`�1�C�?�"D��$�w�����	 (�
� 6DS�|pe��'���'��'�R�'�r��(�����'Gby���������V�l�d|�r�'��' 7-��~R�'��|��[	\DT�Gf%�T@�-��/�Bh�֏�:ab�e��ql�*�M3 jA��M;�'�2�ḫ�{G��-�FH���/t*h�c���`�b�|B^��ߟ�����Y�i\�HOrZ8]�0I"���៼�'��6M��e�H�D�O�����t���2g��r1aC�Tv2���Jt���O���?)ܴ|��&�.�I���q�m].��#�G�:!�:fo�;�z�cD��=M\���?]H��'���$���6
�>6`5 ��	,R��5������ӟ���������}yK}�ڡ3�,��VF���&�@1b�F�+ʦ�$�O\�$+�4�`˓J�����.Q� ��p�W�n��F&E��6�V����0��ئe�'�x���V�?���
��lA=dW:�(%��*]0X��U1O��?q��?A��?������T;/YZ�+�d/L:\X���Ǵ�ioZ7�D�'1�)\��ݓ�^����(\r�w��<[�4?ߛ�B'�4�������G�z���|ڤ8��  �LL)5j�<h��!Q�z�(��'�v�$���'*R�'�t��^k��7e�"N�(x�1�'x��'B_���ڴ.�"�+���?��m��Ī��'���qÈ��c�F��N>)������M{ �ig���>��o�!*Z:D�&A�Z��Rf'w~BM��8�~!��Ι~�O�t�I�3�LÕՎ=�ǤCzc<�x�A\�u�2�'R�'M��s��� )O�B̉`�Ɗxr�<��,��Kݴ���x���?QV�i��'�we�%{���0=�!-( �A؜' T7����4!��U��4�y�'����
��?]{(S�f��Pu�I&A����.��{��'B�I�L�	����8�	�{�DsҤ!8�X#�D�y ė'Ύ6��Ӣ���O�����<q��;^|�A�X�a�J�Bb�?)W�	"�MT�iN�*�'5�rmJ��2�`S �7�nE���Y�N���'g��vb�|;��|"R�X��� �q�b ��p��`�3�Cԟ��ğ�����SRyb�z�lȱ�`>iPg��za���k;\�T�� �O�l�x%�x��O|�n�.�M��i�"�
0MXp� �ȇ�$)=���L��;���2O����?K��M��'�˓����b"M���#1\�ͻ�H��.�ϓ�?����?����?����O$�тnA9m��������c����v�'���'&6-ӳ,����O�nZ@�ɛ��hK�o��z}��
��ijt��I<�S�i��7��n�e�e���៘�!J-� �����˙h�4M�C@�2�P�J��?��:��<���?Q���?��:t`(���,ԂC`��'�)�?�����DUɦ�z�f�����㟠�O%>Q�1*^{����,�FH#�O�<�'�B6�T禁�O<�'���?�!X��2m����`	ӡA@����G�N���,O�)��?r`;��_�">�8��ڿ%��c��ʜ7I^���O
�D�O6��I�<�e�i�8$1W�˟"b��hp(���;Ҁ�sv2�'R6�;�������Ǧ�� ��1bN�!>\�B�=�Mp�i�����i��d�O�02,	��r�a�<�a ѧnx��ے��7�� ����<�.O�����5qжIq��e�����5��oڪh%օ�'�"�	���%e"`8���:��ۗA^�>���q�4|C����O���|�������+�MÝ'��H�EO*O|�l�6`���'T���QfA����|rV����ҟ<�V�ߦ}�b=Ӡ�!E*��0t�C�H�I�rU���Sm�Yy��yӺ����������O�<I(�Oߴ"r�ֳo����O ʓ�?��O�$p�p9o���Ă�2M�i:��F	S��&(EX���O���04P���T�����ex���ş�{�I'8�pV�8�f�X��S��	ğl�I۟'?��I����I,ib�)�CNW�@mT8�	C&3�0��I�M����*�?�,O �O�9�B�-*�>Q#�"�y�(�� �	��y�EsӈqmZ��M� �B<�M�'���k� ��8h,���H˫I�z�cP�H<P��2��|_�b>c�x�.�!~��QB�H˝_j�s��*?���i��xh�'��'��Zrb��/m4N�1&f��p���!S%^s}r�oӦ�mڛ���|R�'���ږkG���[ M�uqᑦ
�6a�r$�����n�d���s���Olʓ�v����>`���#�XԄ�	��M��� ��?�E!�Q�P��e�(�^�����<��i0�O\=�'�7m�����4kN��D�����PB/pn��AE���M��'^�ˍ�1�0��1	I���?I�Xcs:(C����n	�s�\�Z%ؙ'Ob�'��'5��'��6!!�HFr�8�pt@ e���5��Of�$�O
�nڦ�D�SΟD�4������L�O�n9x`dZ�%܈�P�'���#�M��iA�ԂZ"�6<O��$��S����U�K� ,Z����Z]�R����?�0�+�$�<���?���?�b�߄5�6|�Q!؆S�p��AV��?Q��������ˑHBʟ����̔O�z�����4����
J���O�=�'��i꼓O���OoB���&�NLI��%U�H3��H�"�н"V�T�n�	�?�Sg�'R�q%�a-�
S5D��l�u��b���}����O��4�����O��f����
�N$�v�ۚ.��}��/N{��h�@�'ub�'�ɧ�^����4}�б'�˨Z�!��A,IB��k��i��6�Hn�7�o���	�)+Bq�g�Ob�r���'�w�fQ��҂R@��ϓ���O��O����OB��|����tp�������˃4��v�ٛL��'~��O.�s������3��W�W,�H�u�=x��L����-s��e�`Q%��S�?���0ZLT�o��<��G��}�`D��#[XB��&��<�WÔ+?���G����?���a�	��両�ݠ섬X�GB�6�h!ء�>d� �6�W&:��)��Ο �'�u��О�y��' �b	_���h��]�qy:��1�C ,r�'�2C\%d�����'��7m�����Xw��=����B�1C,�@�eA�k�e���	�Q�b�q��5�'t�tc��;!0�۴��d��@jB�M�b+z%."A�Ji�N	�0��w!P-.�*�.�W������H�v*�B�+4m��	�H�z�*6�!��'��GqL2��>V���!��6AV�9e��-A�mC���,���c�i����e(5n �<���+�h��"��D��Va�] ����	�1�P@qP��s9.@�D��7�8,����[�d�qh�@�D5" ��b�!_kB�d��X'ls�CCAI%$��QgGMtt�Ţw�C;�%-	��X�p`@-�����f�8�p,�2/]$6�]��#yj��4�?i����7p�O��/�������@�j���ťǎf�qX�T�h2ci&�	ǟ��I�0�'��*��Y
Ɓ0 ^)!��=���H+RhO�d�O֒O˓o$@�smK6d��j��_ m<�Z��U��?���?I.O��@k��|r\M��8	oV�D�E��A�2V�	П$��t�IPy�F�������ܩ�P�?��I$G^0+��	Ο����\�'¶�Yb	=�韶x�X9F	�y�M�%�
���l�џ�'���'#4u���Tㄔ\����0ǟ	P�l���ٗ�M#���?9)OJ��aB�n�S����s��ч�C�6�9S���K~H�SawӲ��?��0���F�t��M��>�L��U��\dzd�*�禥�'��*sNs�Z|�O"��O2� ��Tںsi�}q��!;[8yn�ҟD��(�΄�������'!D�X ��N�n	�"������ߴj�n���i���'R�O�:O���fp��r��B���67�fqo�-@���!�9O2�$77i>Q!�)]�H@%s���m6��lZ蟠��蟴���+���|b��?E��a�v�3ܤ]۬-�P���7F��ɟ���^�c�D��������g��!�H�S�x�ǬOz�4�?y�Bb̉����'�ɧu�@x��)qF((�Hd�Ų��$�L�1O4���O����<	�O�$���h҇p�R���ѧ_?�`P'�x�'���|W��;���E/0h�b��!z�81I�eb���I��Fy�	ӡ$X�3� ��%� OG<�ca^6'�R���[�p�	۟4%�t�'�$�Od�ps��)�bq����
�,��Z���Iןx�	wy�����T��\�EG�/�@E�FK���넭��	��h�	Yy#^4��O���r�*�"[���2װe���ܴ�?���$˙Pb�4%>	�I�?�X-t�L�O�����ҡ�nO
˓�NE�$ܟ�3�Ø�^�f�3�Þ������i��I?b�f̀�4��S�Ӷ��䄁~j��Ж�F�\+��ce��/����'�bA�j��i>e���?O�6�ԉW��U;�d�#��	趷i=��3��'2�'���O��i>q�	�qal����@>| �\�td7�۴s`N�1p�_h�S�O����Nht����Lm�� A�&Ê6��O����O@a��D�<�'�?	��~҇�$�I��N�%��]y��ܺ|�b�PzD��ħ�?��~roQ&)͐L�F �Dz$���M���%�h��,O��OT�$0&��hA��m�Q1��#=����4��aMw~2�'�X���I�=x�z?�ĨP�Yv%ᄥ�ky��'a��'��OR�DJ<�:���y�~�e�ʼ�ԝҦ�<5�Iޟ��IDy��'����ޟ@1�2ȤqV8)!t�Nd��-zװiSr�'�����ONad��/�!�P��̘���h�v������t�O�˓�?jN����O~�Z�a�
M� �I�L+���穂ʦ��	D���?��a�-LRʩ%�����/��!��;0�4�0�b�v��<��v��x�/�2���O������CAk�!�V@ڄE� 0ޭ�>���v����R�S����25q� �oW�?\���O�7��$�O"H��O��D�O��$��Z�Ӻ�ŝ(Y��	�l4L�:��`FQ}��'D�՘%[�̘��O��D" "}�p�!��J�Y�i&�P�'@��'/r�O��i>���1A�"Q�����L(j�36e+f�f��ٴ]i���e�R�S�O"`ڂw�P��tL���L� F[	�26�O����O$�3`�<��ݴ�?��'Q�U�ċ˿t��$��}�y��J%��oh�M|z���?9�'�t��%�~�Ģ��v,��۴�?Q׮Y���O|�d�O`�d���� ?.i�2��40[�*�>!6iX7*P�'�B�'&�I�$e��0%���Rq�ʢ�>�ٗŗ5\�L�'�r�'�2���O��0��	J�$!�h�{�QqP�݄�te[�����I�@�'�B���V'wE���V�B�TX�"��v�'�R�'L�O�˓|���mZ=g'TT��A��$g�y)�Cϕ|4�ꓚ?Y������OFmh�Ĭ|��*�,��$J�\�yp�,l�<)Գiy���<��\S�I�2S�+�"ٌvJy���}S�6M�O
ʓ�?�V�Q��	�On��㟆��]�Z���S+�&g�f1� @|����=%^�֝�gLu �i�/;������	����?i1��?a���?����z,O�Ο��ɧ"ha�JFf8�	��PR�͂%!�)���58\-�G�>Z�3�'��:m*7��h�
���O����O����<�'�?����8���E^,/O(��U�&F����νiB5p�y��i�O\ �⅄?`�x�a�y������ܦA�IΟ0�I��������'���Oh����\�a�&{�fU��a�i	S̓N�l։X�ȟ���Y?a��H�4ēsbP<>���viӦ���!(LH�'�R�'�"�dӐs��MӇ�ȞJ���������+��:?A��?.O>��F���y�4G�m�����;d�΄*���<i���?1���'�M�0|���c�l�|��%
�G�\v�]2��և��D�O����<I��V@��O|�h�&%o��w�
�fbF$8ߴ�?I���?!�b�'Ջ�{�n��I(�u��m\@����P�L73�x��?A����$�O�8�Ȱ|����P J5Ñ;#�h��+�9:H저�i�b�$�OF��tc�O�'$L�`�j�=�,�E#��	�F��ش�?�)O~��B�'x�'�?����j���1�2qq�&�A��B���*\	�O��:Q03�T?��PÁf�8��O��'�u��>���3R8���?����?��������U�͝f>�-��B�?�~� #_�0�	"R�9�)��p\�T��m	�SH��81�N?�7M��E����O����O$���<�'�?��僞B�p���J��|��3Ƈ��̛����E��4J�y��I�Ob�r�&�6cM��C���Tz��j��립�I֟���;�2Е����'�B�O&%��H� 0*� �%(��ᑋ�M̓I0@f����'�R�O���/G�_9��3X�+�i_��V�g��	ӟt��۟��=!P��k�@DQ���h�I�PI�c}��fz����O����Oxʓ�?i���R>�j �̈1��Q��8RpjT�-O����O���4�	�P�%o��O���J�H��o?�#�d63/�D #�7?��?�*O���J5	�����x�T�z�*�/y�rIr�˔0 �6��OL�d�OV�H�	*CChܳ��a��4a4��[�p`c�j3��`[&U�d������'�b憘l���,�%@� &�^S��<MJ�mp�)��M���'��oA ��rH<A1�Q�Z;��e)�>�PT�!�ߦ1�Igy��'�ɑ�X>��IȟD����� �@3En��R���b��ԘK�f�+c���OH��p(�:�1O��y�T}c��s]�@�cC��`�Z듻?Y&�A��?���?�����(O��Y��kR�D�@�0$P�$D��	ӟB��GW�b�b?����F�b��H���l5��!3n�N�""�O^���O����@��|��{6J�%	�b�h����\=W&��z&�i��B���2�����瓤M�H�G]5v0���I){�^8m�����Iϟ���ʚOy�O:��'.��Q�I�����Ҥ����JG�(���<i��KW5�Or�'����	�.`���Ra�
�I��_!���'8��D[����ğd�	i�_S���dY=vI�D-<8F���'y
�{ѧ�����OV�d�<��$.�R�A�*�M�߶�$dh�
����d�O6���O⟴�I5N��=�Ƣ�q�%#��R��UA�z�0M!?���?1+O����7��S�.j�y��%�<PU� ��iq$6m�O��D�O 㟬�I5]��9j�Ot�Z�iU�8eg������]5�k�_���	ޟ��'�"�5Q�ɟ�*��.&*&xZ%E�4�(x1-�*�M����'���<_K�-{L<y��O��C�)V��9f�ЦU�I����'R��Qaɥ~����?��'7-R��@˛�Z��Ya�`̍Ǌ�`�\���I�p�	��v#<y�O�1��%G�k�B8a�`�DT�ܴ��D��u�o�ϟ�	�h�Ӏ�������G�)��i�qB�����sw�i�2�'��X�'�n��<������,jm��GdE�{���4+���M��}��f�'���'��4��>�-OQ;��I�H����: ���7��U�5�s����{yr���O���H5Q�
̸4��w� �3э��IßX�	6k�QíO
ʓ�?9�'�8����*k �e�@#ꔩy�}b���ژ'9�'L�̈u� ��x0�S��5m�6��O49�eC}RV����dyB��5F�Q�zcr��0�ʙv�`i��T&��וgT���O6��O>�D�O�ʓl|v�Q�'�/�49bv�R�r�&�p"�)|�	qy��'A�I���˟H(櫕"q��3ց7���"�n��bݒ��?9���?a�����R�R�Dϧ����,Вz��P2䀯2}��m�Cy�'��ß �	ȟ�C�>a%�U/7�h��Sa]%r$d�5�ꦹ�Iß���p�'R̠0��~����IR�}`b��㔋��H�T�O����Hy��'~"�'��y��'a剫68��)�͜�Bb�
Q ׿vj�=I�4�?������:[��O���'�d�\6&���p����t �##��;
���?����?qD^�<aO>I�O�<E�"J�9.$ pCq+�!D\ y�4��Y(}@�,nZٟ`������,����j|����bp�!�K�X�Ε�i�B�'5\\�'��':q��8�$.ę�� �Ai���`�iV�)(S�e�$�D�O*�����i�O����O�����;��3`�˖@#����Cͦ� ��\ܟ|�	Cy�Oq�O&�� ^�@��Sbz�!˖�# �H6��O��d�Ob�$�I}�V�@��@?QTM�7�\����߳aL�i�#����'����yʟ����O\�d1�ki�C��������l��lz�l����<�����$�Ok��"S��ׅ�/ �v���,F�V��ɏbE��I쟰��ߟ0�	П��'������8d�bo�S H��W́I�:����O���?	���?ɐ���y��I󬏞)����`U1&aD4ϓ���O��D�O�ʓ:��#%6�ȑX�
�K������p����i#��ȗ'"b�'�2ŕ��yR"^� )�G@$�ĩ��٠t&��?����?�+O�,"��Fx���'_���Ƨ�LwdHjŧ�!�by��q�:���<���?��&%
����	�j{oQ
NA�%q2 T �@6m�O���<ٕ�F2��ҟ���?q�eᇃn�ęh��ǰd �Ł�(;����O���O�3��?�'��Ɍ�4+`q�t�F:��H�2�> ��V��a�b&�M���?����3W�֝�AŐ�@�.ܭ4��-Ϟrm27��O����+%��Mf��'�q��d��lPF��8r���9æ�I��i&�8�dv�R��O����r��'8��d���µ�ǋLa���I��^�ƭJ�4"g��͓�?*Od�?E��%\֒=���5Ҋ������ߴ�?����?q�
�+���Ey��'D��^�y�տn���#H>��IKyB�6��4���d�O^�dǃ�U����.��A�V��"���� �i�R! �(,l����O~ʓ�?��<������վ!@��fO:'�6hmƟL@C�c����Ɵ��	ϟ�	\y�f8md�	���m�XuK����'ҵ�W)�>-O��İ<��?1��Qg�m�פ"�(y���%�0��GD�<	*O��$�O���<CA�~�!���`�P�/���#_n�fQ����Myr�'��'0 $�'J1iƠ�oY^�Ru�һ^ �����>��?���$�)x�Y�O�Ҡ�<�N\2�h�l<��Q�Ř�j��6��O2˓�?����?�E�<�*���ǘc� �ه��.��h�����MC���?�*O�9�cq���'��Os�i�&B��R!"�
=݄�rЁ�>Y���?���4�N����ģ?��WL��z�5S��Ip*
�j3�`ӈ�Ǡ�Cd�i���'"�Op
�Ӻ����/#�p��o8���LW���	�(r��k��J���9��.l�hIAUkU�����šΚw�7�Y��.�nZ�P��ݟ�ӻ����<1G� <����)<+����<]h�M8$�i�:���'J��'�����O$!�oϟ$bL�D�O�m3d�¦��IΟl��&)/��H�Ob��?�'vL[�#��Ȑi2�B�0;�4�ڴ�?���?	��Z�<�OaR�'"m~��4��CM�WS~���$7b6��O$�#�jO��?�M>�1);��Ӂl�p�l0���$Ƅ��'#T�c�'����������'>�6J_b�,eC��Z�VDLa���l[�c���R�����I�X�LkT�G#�E�śs� S�ǻ._1O�d�O���<!��	j��IԠX���b��*K̉G���,���՟��	x�՟��IX�a��,v�ݸSCׁ�P$	���h_�L �O�D�O��D�<y��R�PB�O6�؁q�H17�1a��'6.�Xq�y���$���O��ЇLh�d&}LF[�Hʑh����iT���Ms��?�+OtE	���c�ߟH�	FǄbT�:y��c�AӴ�H�O����O���;
�*��?�c�@E�8d Qd�� � `�Ax��F� q1�i"�맲?!�'k��*[� )�C(S-|)�rć_�->7�O
�B J����}���_��T�s`�ҕ6e���e�7e]��M3��?�����g�x��'�rͳb��I�����.�T�[�r�t(�C�/��u���?Aƌ��j���񵫙���3'�'gx���'���'�b��dc/�����f��Ev+ɬV�����#J�2�H�m�p�	�~�)R���?��OVV�6��!VJ�������Y�4�?9��D��'rb�'�ɧ5F�ŗV�n8��������a :���i��<����?QM~��N��Z�:]��
؜Oi����c��x��mi��O��O��$�O�帱�	uDl��k	W����";�h��<Q���?�����d�>%�'
0���r�L>H���`����d�]�	ʟ &���Iʟ�`f	O?QS�M; DkT&^�c�I��~}r�'���'y�	:��dPI|�c�*}��`"� �Ss�aJg���8ߛ��']�'p��'\�X��'��HQ��ʒϛ$"��+e��l���	Dy��P$(=~�Z����k̅
NY��z�^z�����@/%��O��d�-l����Oz�S���Vo�i����'� �:gC��M����?��T��?����?���J,Ok��Cfl�C��y?�)���<s˛f�'{"�ɟ�O��>yq��[)�29����1��a���i�^I�7C�O��D�O����p��O�'#�l�k�@_�E�V ����9����"�i><2E�������䛃lGL�s�!��8Q0�E��h���l�៸�	�۴�
���|���?1D/�9n)��J<A��L{�EbC�OTBrf9�d�O��D�O�LptiG,�h���NM�ucցPR}2�&��	`y"�'��':�x�,�� �a�ï8z��r�)�>�K�\�8�'���'���'���D7uj��s�H�3n�:PHZ9�� �qV���	��t��]�I��p���DT��iҬү˾��u�h�"��d�G Y2���?���?�-O�P��
�|�S�:x(�a8'$AH�!���ߦQ�	�������?�+�!�~��ק{��Ls�;��R�����D�O���O,���Ov�*���Ox�d�O8�k�e�pǨ!��HL�������	q��ן���*DD���w�6��?}n&)�f�{�TĪ��x����'��	՟��p�~���'S2�O��D���;V� ���3 ��EP��/�d�Ox�D$�ƅؔ�T?�Z��ʩl��ӡ��,\��I{�/`�:�N��R��i�꧶?��'i��	�2�*%R�
��X��,vֶ7�O"����4�b?M��A��W��p�ܕ1Q�d� A��O_����	��D�	�?	0H<����1` ʘ�*�I���U�J��iɈp*���!���p5L�+F��U)�*�J�F�������MC��?����jU�e�x��'F�O�y𠇒�G�&e���D!v�B�1}91O��$�O��<讜u��5o�. !	)n`&�oZԟP��\� �I�����O,�O��J��B8=~�*Bb[�b��CF�u}B뚌��'?y֪�WUx�!@�AE�����U_�I C�ɀ~΄��u��y���=�4���FqsT1C�k[#��O�����:\�|�A��T0C��q��GE�6��\����g8P�џ{~�-x��[�d�K �ŇҘub�X�'�ţ#"n-���e �]�da��O�vl��+;LN���F��˗��aF�f$@�h��7_�TY(��!���%�
:TH�"6�ښ-}p�cA Q�e�:(˒+5rYy5�V= ��!Y�'�R�'��Q:щ�L}x�;��	;�Y٦j�fz@��MV��9$FD�,�0� �d�'�<�3s��3z54�7�	����s�Q<6�J�;�2i���W�Q<]R��g-ɦ 
�
՘|�ɦ�O�>?�̝X�e_�t�t8����|�<B�	�6߬\UK��c�*T�������^��<[~D!,�Bh�t#�:X�g|��l�'����Ol�'A ������?���d���vF�,���開Ի7%����e@[�Mr��^׊� ���%��O��1���F����E�!3�ȘsdF�D�R����'if�; NA��"~�I�|N�2�J��@��
Ƃ2Od�T���D�p��b~J~�M>��K�"!J�س��)��g�B�<� J%��Α
,蔂��"��d ��I&�HO��=��E��c�2,X��1(�:�����1���<".Q�Iݟ��	ٟLZw�R�'r� ���^_�|�+�,G�w��(iÁ�OJ9Pf+��B���9uh�	����d�_SP��p��:y��AWlN�Z!*��I.=�n-ِ�d�,�ʆԟўH� A]�wؔT��	�p����K���ۦ��Ol��*ړ��.u�v��E��#(̑�DC�wL!��_��܂3 Z=li����A�+�.@Fzʟ�˓�,hj��iM.���>=���B(�G�V����'���'��散<L��'��)П}���""�E��6�Q��|����W���(�T�����,>j	���p|��E��,�Z1��&"an�ۆ��lj��i؈!�����$̾A��'Y\�jb��!h`q�������*���Z�'=BU��X�e�T�XƋ�M�0�'@*�آ@V��́��_ ��J�'�����$^�:[�5�'."\>�{����OA洪��>���9�KI��h��I���K�|� �B�|av`�w����?�OW�˳��O��8�h�ٮ�:���е>v��BG�kJqQ��;�r}���OC֙x$��;Z�ՠ���v��T�����c�'<�(��0�C��X�L�q88���6O>��$@)K��`���Z��,�d��Nda|r�6��I*�|�to����`�`��D��.Ռ��'�V>mSGSٟ���˟D07CV3]��-��e�?E��Ð)W [\�����^)n|�}"'V��'��?���PيHs�.�j;���Z�T�ㅎG2[+�kOG�*�)���iw��
�3�Ś�U�<��k�uZ�������'���vL[B
*"p��T�N�(�D��Ȫ���@�(�r��J��)*�Exª:�S���#1��Y���k�h�V�Y�r�'׸��mT�o,��'�r�'��ȟ��I1�2�	��3�9���/Ap���1�,(�����ؓ(Z�iP��ș�i��I�r�hd��ɮO����wA�+���(f��	J���� �M�����,O*�D�<�$�VX���^f���m�b�<1�,�9t6,�Z��T;}G�I��K�3����OC�ɂrB�k޴æ���
O�1!e�<���?���?ѱ���|�����Z�!6�����/X%�� ��Bx]����\���<T'��	E�O��0��C2[^�X�d	AT�ȝ��'LR}+�0�6�>ov�B�ܪA�����'�<|6��O8��?)�ʟ�[k�'�Щ
���<A�Q��"O�U�bM�RXl�"u
�3l���5On��'}削u�t��4�?����iʍ@�\@����t�0T�$�	/�(�(�?��?qt�Eo�6�T>	��O5��8kF˖k���C"�@T��؎�	H����P�40���AU�j�Q��F��O��5���O�=+/X�un�E:@�#4�Y���O��"~�H��%����<GsT0Ȑ��+3�z���9�ēd�r�B�|L���ǜ|�b�͓e9~���i��'��S*B�He�	����D!
$��U�	µ`�$$��0"�ٻP�v��<�OZ�OQ� k�8>R88�f� hc�`:e$�<ޘ���+�)�矜b�?6NZM�QkX�o�,�%��)!wni�I��\��ҟ�F���<����f�l�v�0��\͓�?q�e��2`ɓ�h���A��7��%Ex�-.ғ��%���~j`�e��5q��4s�)�W�
ј��?i��ṟy��O����O:��P�c���?�gD��1����V�C�v� n�m?�6���h?���@0�����a�P��G"�i2X���6,"���Hס��=��⚫��Y1���6;�9
e� �?`�N�?)��iI
7ݟ�	��'=�s������UN݂;I�h��'@:%�4�׾(`��\ji��K,���i�<����$����L0M�����IޮHE�@h��֓$r�'�R�'-Z�J��'�;�.��E�2��&�:6-��*G�sI��@�f�f!�@F.lĮ�?�@�~g�䱆抿Cʌ3iD�Qa��IA�S�:�DD23�@�'┘h��dEO8��lӸ7�[�_|ԡ�K�:�1����M������OR��'7#� �%��!v��X�sN�+N^���d�>,��PSޙ��)L8ib\̓b>����ɱ+ �����?�����i�dJPZ�^��q.��6n�Q�e�32)��'�`��e/�����ZD��S���R�'(�w�A��s�o�!�(O^�����*�$x��#�S�=BBAs�I��}S�I�@��<DO�˟�{۴"6�O��/S.!��U�]6���HX������������(F����>���j���uXa|)�� ��w�U$o�}A���W������O����F:h �cl�5�8�G���K4!��#e�z]��IL�'�	+vmŵ !��L�PtB,X$��?t�}cW1p�!򤎬�$�xQQ�|�Z�S� �!�_\�@(@tጸS����`^�5�!�	SHt�ٱ��;o�up����!��G� �;R��:Aĵ��
\""�!򄅦j�xy6MQ\V�4!��1!��39����7�Հ�N_�H!�$�g,������x���k�''�A�ė�"Ф���qUx�"	�'�L�U�ɋF�h��BUjAR!��'t�RS,�$6w�҂�Ǎ9�s�'p���"O�'�N�؁�\�_bL�'ڼd�-޲wdu�VA�U���A�'�)�	rZ��E�~����'?�I� %"l���U��'K4�S�'�>,jf�H�Wq�`p@*T,���'*�\�s�N)H<�90���Ԅ��'S��D/�]��qZg�]��I`�'I`�K&e��*E�$C��P�� �	�'� �	sD15�D��K�6z���y�'0V!;�+�#}\rY�6�;v�`3	�'��;s�ߧjD(Er�
F�PZ�+	�'ʤ��)�
y���x���b���'b���T6�@%��/F����'�D��N�j�޼�g����ɀ�'jD� �˩x2r��f�^�,��u��'Y M�A
E:w��]�֫X�&�tC�'��YSagM?,�L�����5/�"���'�DI:�B�9�戳�
D9 ڶX�'�-� #�)A0�Q�E!f�PB�'谥�J�e�,����7����
�'���`G�.���㵅�8���'W�� ��Ǧr�T�G��b��_ʌ�Vɗ>)�M�U�õ'�� bu+0A����M�E:��!7� �[�^Z���$�	0�@�UG�l���I�'���c�8@������$X� ���{�'b<�|q��%�(�b�\�K����x�P�F�é8?�ĸQ쐖�F}��i/�>����Yl�S�t��m�����w����*w
��%�f�� ��'������Eh�x['��S6���*���0扵q��A:1hÏ,. �u����Y���U�&��E�c�M7u
����̶~|ax2%<{䪈�o�d���g�\1 9�(��p��ٺF���c����ѳ��H����+$�{� 4J� ����"R	b"�ڭ������*�P@L����BA �y�äB(ED$Q��������o�,P�'��'mb�@��"O�li&o�\�@p�げ'��8�e۶"z�����<8X���^�ڦmk"g�|��҉�^H�;���@RK+�Ʃ	ց��'&Ȅ�EF����-�D���C�\�n��!���Zҡ	�)A�:�ܔ��� L���'%� �����h�ra�bL�W����0<�5#�ص�F$�- �	�T�K�=?P0��N�YΘ'c�XjnT�s!��t�q�	�y��V�y�@P5�?�T>�1�iV�S�My�A�5i��i�'"?���&+R
d�,_�z�0�(�bK�-G.H�Qt?�ӛz�j�R�&M8u�Ĉ�G�C������U�҅�W�>E��'� d�$`� &��
��5d�BibR6��b�i�1<p�$��~*�rX��dH-���e�ޥZuMU�!z�P����j���M�WTt���?0ax⁜����hp�ʳf�����a��"P�I�D�L��~2��K�4�2O�'nj5�s�I��?�0AP3ls�}��z�Z��C�B8��.N�v��H�2O�����*�Q�Lڐ=�(i�KA�Sb�1g�ٷqNT�`"�MUi4-�:3�|�L�O���@I@�B�r�'������
�
U�q��B+N�hH�'��9��E��В���51�\�Y�{��d���Z��=LȐ��'t�ȅK��ڊQ�>���x��9Obij 9�UZ�Ak�H+��v� �E�@�U�qO��O�zp+M̼�/�xL��D��v-,��@���<����?F��(W�'��d"�dZ8V���0�\�;��2V����	�@���dS°��O����+t�mm�U�d�	�@%ֹХႩB���$۠lȈ(�ƕM�LhTg�
B�� ��h��
.$0�q�Cݹ'j�Y���'ܬ�@�N�Ԝ�'�`��&�D�5/���j�MI#s��0��߆���r$c��}��	�M��l��@�{{x(�I<F"��40�m�s:Q,�&d� E�����K�W͂H&�l�eƍ��q��$ɫuMZ���N�\�����I풽XӬ�O�U�q�����$ܟg��]j�������g�����šF�t�	!)�\�;6o�(Ͱ<�EE�5�0�
�#Ԯ7VܪD-�*"��O6��)O�X��)E\!v��O:T���Io�z�x"�-[7�p EH��=��A��'6lܲ�	}.�=Γ����ȕ9N#� 8@��<q>��-L����0*�C���!��<YU��
��'����3�a������ 2$/(�X�CB��0<��i�x@�O]��I�X#L*⠁�Hҭ
6�ا]�a_t|�<4�!�x�AU<t�H�}ΓJ��ꑉK팍�[�Tq���\hcd=|��0��nSLwڄq��4�i��!����eÃ�\�s�i�Da�̲d�N8p�%z�
���8"ꑒ*�Pۡ����|��ȫc"({��U�S�Ʉ�}8\��B�\��G��5,���K�i}��.T��FF	AFYCE㖧9�X�ŋ-扇y	���k5x�c����a&�D�^ar���)k�R0��I>dV��b�i��}������FO"P�gFސN�J�Fxҡ�Od�qA�ۭF��E��ǜ���X&h��fS=���򲬁��#=��GS�4�B���)�Xx[��So}�
��F��bi�'z��H�ƅ�s(ːm6y�#�(�h���gZ�C � �1a��ʁ�Z�h���\�1���3.����Q����Mk3y��ܴ|�(�5��vO�m�N���c����(Q�&(���R��:��d0b�ԸF>��%ٌn�
��4"O��ɇDs�Ic6J�9d�aߒ�]�HP¡q4g!P�T\r%SRC�I���h��&R)�8��ݢ:�.	9�@�&Q^`#�J�3-��,��犰��h��F�'4`A�
�$a����f���X}s�k@��듂��a�^5a�ŝ0m�����^'�������2�R j�(�J9��s���Ox���q��Cv�h�FhO�55>�b�C7O��I[�ʭ��l�<i�d�'�r�Eo	&�� �fÂq8�|YH�-KF$���� ,�6� �iq�:�C�ī\
n�`S,fa���to��ɣ�<E�t�q�望���98��IhG>�O���+rb"�;3�ӿ3�.ٗ$�|����'!�!Q7@�vUKr%Z(,��{,O��:R!Ч,�1�1O*Q�1�ȍp
x���^�&�:���Zc�݊��'kX�P�g������U�J��D��'��koи9pN����3%�>Q�w�'�"M`f�!T�]b"�V/x`�Dc�$�$�OD��*Ēc���F@Q�~����:�^l@bB�gg�ǽ0 ��W�a|Z�`���	�&)bE͏�"�f�2�G
((��������j2o<9$�� &R�{�0@�ɞ�f3f�0�O.h������3D\�oP.�d�zFf	?a�J���ꚍ�O\\�U�΢X0p��u��zʔ���;O�ȁ�[����l�%p���
'D�8Y��P���m@�X�E��D����5)��=�Nj#�a���՞�&c`��b�)�Z��� �V`�*��`���NU��"o6@AnR6�=���v�f ˣ`,���҅�A��t1�J�U�# ��I�AG�R�Lx��'
��#��ɒ �d�h�'i*�S��Gϖ� �U뼻Q�CN�JE��+�0.^&��V,�e�p�6!��f�>�jC)'(�����Ί>D����Q�g��/����s@%K��C�}cG�kz�O>͡���m���љB�eH��	�L)�]�ï�)x�\(��a��sX�ɇyt��qeN��RE�1L̴m�R�sl�;f4�95&E_C�M��I�Zo��ʖ�Ɣ]`����ƫK�t���h�|m��n	l�|�� Gw��Ȓ�ִ�����̶���I�Pܴ(�F�(S���`BMϒP6!��ܻ'N�[D��6 �T䔏�μyt:O:�#�0NM^ٸ7�O�,��a�H��ph��֝�yB����#nI�?/ҼS7DΥ�0>y�ez>5A%��U�T�kѫ�Ij�ː�<jXQ�I�X?IV#L�t/�P�6��"ĵ�Q�j�R���E�h	 A�K.��P2�U��A`!/����x��O�L�Z��z��ر�Y����<�R�#gC�]����@9}�X��p�zy#�e������ʰ�f����6Rvp4�ߒOt�,[�b��<!�m�E{������<�;NZ�p�B���D.V��gN:���'�L�j�ϝ:�0=9����H�Ԋ��
O\�Y�d�#{Z����^�|eN��w�T�G��ϧ���|z6���s⍸r	��W��@䅕
.��I b��U�taЙEqF�0�@4�*��aB��V����M�
E��h�	�I�eA5�3�i>i3�KB���2#2<da�h9l�,�$n�1B��T�!%�dy�.��	��k_�r��g@P�:O�a�-��z�1O?��0K�(�48��l�iX�ƨ�+I3Ta��G��/I� ��)�/*�F��w��ő�/��=��da��W�r�P��O�ىBn���az��I�<�H��0OE�-1j�j��6Q���ʇ��;JsT���Ƌv m�Oh�'(MQ�H�8� �� �	ڐ��eE�{�}I�:�V���G��D��!��Nċ�����dE>w48�7���wiD�
� N�̘'aT�JU O���� �{qc	�-}:���L�/,�\�s��W�]9��խe���t�)?��O�*Th �"/&6�I�F.A�6H��'�� ��bB������f$C�ͅ�;a�)&�)ij��3`Vt\\)�.��"������>��>���V�nD�в�����Y=�P�'\�a�#���0=!�\�Z�l�ˀIؔֈaS��O92ȵ�!��L�L�d�uY���;��'��k���8�,QRG_/T�p�rv朄Mv��C	ۓNΝ����4�p�[�̝�}�f��кt�=Ô.��{�h�cf�.�p?��ʐ�\O�ͻ1(�H�`�B�X�X`��!.�Rr<3�ր`�"ԀM?Q���l���@�n���x�m<D���Ԓ-L020��g��c!]VZ���G�,�;�B�V�#}��'#�ۥE�_wb���xȞ�y�'ج�����yr��330��Z�z��U���cO�x�  �u��I-$H��!ݝ~��q�u3= @����>�@!"��:i�蕣J��£ݭ�.욒͜)*^88��+�OPD�)֝\�x#b��4DȢ���%E2� �mY��b|0d���bS�O��	ɔ
4y9N!��e�6	�68�'^Ys �C���-#��-L�b��C(e�d�����Ì� �H��Ƀw�B�)��F*|��p���qt*C�C6SkL17Lh����H("H3p`�59�51G�G�?D`M*r�F}rɊVhA�3�:����N���=a��G�������Q��x��& i��ڄDY-C��q�A��)�� �
��J8��E�"1���pqbȟ���>��S�fr:�rD�/ �=�W�թ��S�B1���$C�Q�`b�LVb�C䉢D'��@GIB�24�@(@l�S�(Hpj,4$%*G��BD��:A�<�'�~��S�}���x���$8���创(�y��޶�`D���KI� � J\�*qx���e�*4����,�M"��^wpQ����G��Y��
�(�/A;�$�2:lO��!`�$��AA���"c�Ty`%΁dJ���w�[�j~��2�A��A������#A([bG��-��F�I��Oj��j�~�s\c�v��(˲���00��CK[�>�*Zb��94�LC�2UX���F#!p��Y�Eo�S��(Q�M�/� �&��t�H3�)8�g?��Ʌ8v�`0ȁkR���1+���c�<� -] �RѸgH6P��hT��_�<9c�ʪb�]뗯��K�Z���d�<�%쏺�p@�iބWc�X�DAe�<��&�ae4q"A�|�h��Nj�<AA�N>V$8����c�&��Ig�<�QkTv}Pp��F������x�<�뉥b��C�c�sC�(C-u�<���7�J=j�4D� �5Nq�<y�gJXB�cDb�`:I!��e�<	���<���"�!@�r��O�_�<Ai�%i�t1PgF�}���XWʐZ�<A���
Q�:��-����VZ�<e��
{� ��� ���d��U�<Y�
݌A� u���Ϻ�� A U�<)5o�!\ ^�0���8�B,���P�<�ҩV�<��4q�ˁ8O��	S��O�<�ȑ W���a@�l"
 +��K�<Q��Lj1ҕ�Ҫ�1bV.TR	YP�<�ť��0��S��-RE"�K�M�<����;42��y�`ذT;�y�c��}�<9ajYa+U(�"�8���;E-�|�<��bO�W���:%e�	��	�f���<A����c< ��t04���QU�<�bˁ��*h0�
�=��� R�<qp�p�$����+v�A�&S�<��/�|4�l@7!��T�����u�<q�,R'#����tř�@�zH ',u�<1W*�C�h���� ��R2�XF�<���!Ne�ױY;�Qra�[G�<Q0��'�Xy�hT�#u"�	��~�<�TU1�֭#��YfN����v�<B������ ˨6( uf�v�<� 
P�2��;or����"a�Z}�R"O�5�ă�?ެ�����p�.�(�"OR�㲨=���+�o�*|�lK�"O�L�Ć�+#<�bt@K҈�YU"OЫ��ـ7(,�ȑ��Q�bT:""O ��1��E�<h��ꄱ�l�y7"O�����I�]Y�h�Z0����"O,H�4L�5�x��%΀�'�(xV"O��BEFd2�Y`�LK_�XM��"O��G��yf�`	���=V4F"OdUc'ܡK"�� ၚ�Gh���"OpIQ���{�X��`NZ���"@"O|�!5h!!��9H�፜H�d-"�"Ob!Љߩ'�L2`�L0d<f�J�"O��8DAJ�Z��8��O���Z��"O4D"D@S�0��Sqm�9J"O�4��a�x ��x�·&bv�h�"O��u��5s�^�K���b�����"Oְ�EQ�Dk��w�]�e��k�"O~ai&ƺ"_TA�Ņ�%=�����"Oq뙝B�
�Sq��7<���	�"O6Uq�mU� t�qR��7e����"O��h�(R���06�ՍU�h
�"O֔j +�\���+�$
�m��<(B"OHq��aG E��U:�bP,�`@�"OX���G���P��!@xNIw"O��c-�X�6A�"g�Xs"OyX�$
He$X����,����"O��A�l���p���%*kK��y�"O�xZ�]�����%v7� "O@Ax��C�C���䒾h�E"O��� -'C{���ad]�2e���"O")Q�V�y	�pr�ͷF_\���"OD�(b����	P�8f��Ā�"O�HX�� � �p�U� �"O���MҬ=�V@��E�c�2Is "Odm!�����pya��5t0�"O����Q#���c�ʺS�n��"OP Z3���},H��n��lY�"Oj���;BŲ��0HJ�/��;@"O:ш�+��K||��WaQ�OV�X@�"O�`^�K���i�O�+�ã"O�Uqq@()�����n�.+<DKR"O"���R�]
����H#Ä5+�"OJ@��g�-	��v&K�y����C"O�U�S+FJ�Z��Ed�k�4�"O.�:����{����p�t ��"On����h��I��@��J�5p�"Oʥ�fJ��&���w�W� �EW"O����*�8v�T���]�!.��"O*�0��-���C�*e�Z�Õ"Od����)}���X��� ~��"O��ٕGͤ$�rr�oT!�l�3"O��a,�6%� ��+?���y�"O�D���J#<����Ԑ�J]�5"OR�Yv�"1��t�����`C"O^�)f���k��a#�l��0"O��6�3���w�Su��$i!"O���4.��F�"L��Ѡ�J���"OZ�X���.�}��a�!;��0w"O��!��=]
6m��A�39��r�"O�))���+�f-�oS�h}p�ɑ"O�|z��Z^�B�	I��IC"OKŐJ�
q্[?p.�X2璂�y
� ��PG&��oB�h�!gG�M��CҞx��)�S�k�����\=)�dX�@ބH�C�IgP6<(g&`WLj�Kߣ��C�ɄZ ��B�56�1F��f�jC�I�D�Nm@���J���f�X6S�>e��U��(8�ȝ*�č�"N�/}�()�����v��RxK�]�E=�ȓb�`-�p�QT��y��\&w��=�ȓ9�����-Z?b�
\�sg�"hhІȓoO�(��ժ"r�)3ßA��5�ȓͤ$�7C�i�� ��/#~9��^�xṶ$EKl �p�I<7P��ȓ ��p��4r� ���C^��10�����~��I	�l�Q�Z�ȓ$���;F`H'��}X�"�**�U��V����.��X= �xb���2��ʓ%)�����S pҀ��C�ٴ2��B�I [��8�5 �6�p�#!�t�B��+_�0����4�j�
ɀUz�	j��h���ؓ��! &jP�"��5�T��"O�9� ��%u�T��#ѭ0�����if��>�p>A5G�;=��[
��(L�Q�C�_��$�p�9~U⧆�h��i	�b�Q�<4��n�(��1EO�>I,�C�O�<��ѻ�h�q�o�*�����V@�<�ħ ��F9���?G1z@�`�~}��)�'{�ЕX���f0� 3�K;x���O|��K�E�4�VA���0rT�ȓ
�.`#���)S&������	C<Bȅ�~_X0��˒�78y�C<��ȓibW�\� #���A� "OT���K��J����'s���"Od�C'Ԉy��d ��*,�(�j�"O�uB�璲m��h�4o�8/��[�"O�a!�h7(�+R�_���"O����� ����!ǇR�,�W"O~)��/n���kցe��p�"O��Q�
'���`G�!a� �"��'(ў,!GeT�dP>�ӷ��4=�MY'"&D��"�D�q�)��*թ_��U��'D�l�C �z����D�3T���q$%�O��I3�\�91@�J�}H���XvC�	8O��}�hX�t��u��D `NC��;1�h�Sߜ)�f8�S�F8BC��8]��Y����@0T��Ua�[l$C��4rP� aǟ�Ћ���0CTC�I%o����ȗ<����X�{�0C䉀$rN]s��ܝvl�3�
���B�dҚ�HQ�K�~��`��m�$r�zC䉋\��2�,�~L!�'�^�<C�����◆�}�^x���/"�C�ɢP������-{�0P�G$��8�C�	V��)�G��Eb�}Q����Sc�C�I�4x�B�րj��ͫ�����C�"M�t�A&�OY���A�YdbC�	 �9��C�%{�x(�3��2W;
C�I�	V�jR��"�^;f����B䉑c�nM��(3�*HB�3�B�I�*`:��"��0�����P�<N�B�	86�~�jNީW���� 9�^B�	F�XzT�^o~D��J�6�
B�Ij>T�b���ٶN�86o:#>щ��+X�<�J .�;�z�rPdU��!���>q��f�0�PAA�=|!�� v�9@f�<��)��2O�\��6"OԈb�J���$�qeݙf�p��"O�xw�K Hbȭuu�A""O��	�N�8�N$�U���ha��"O
8���)T䈓�.'"�\�"O���6\׈1�4��>����"O؝8B������2��5�V��"O���JIi$�Y}�&}Ї"O��6R����}�^���"O�)��
�T5���$�8H�"O~�ⴉU�8X�� 	ͯ?�h�q�"O���5Ȍ$96mcr���H�jT"O<}0Q�:1Dd@�Ԣ^�Jm����"O"�B؎Td&=�r��	R^���"Op���D*��xt�]�@<1�G"O.� ��*������q�Tt�<AǩN"
�3JSl�b�!�Uw�E�ȓr6`�
��0�N<��O��.�L4��x9z��%J1�*ܸ��ĭJB�ЇȓB�
��%�5L�,�0���(\@��fߜ=�0�X�j��xU��3��݊2f�&{P
`Z��z�؄�_(����<p�艖`�T�&���Ov"�	f��2pm	V(�*n^���<�:p�N�	�!�t�>E!�q��K2���b&�A��`a��6����"ʓl�	��b�,G�5�@	Fod4��������KR�X�C��<2(1��L�FhI���
8�%cP�|-.��ȓj�=��,8	
��B�RjY��ƓXe�eJV�OjXx �${X����'):����O0VQs���-u�� 1�'Ǽ9�V��)xx�<��gܖoR Y
�'Mm���̽�|��s�Q<mJ���	�'h� ��-�<a������Έk?ȀR	�'������uT���1I��gvL���'�ސ��N8�J�j!e�N�����'�.�����|�! G?K�l�y�',��!L�NʑQլWJ��a�'�D`Q���s�:��C��*�xz�'�|!J��I�oLe��癰rs\��'�̨ۦƬK.m8��T���'�b�ӓDP�N4`D�q
�3����'>���֭����N�	j�`��'����)�TWQ�ˆ����'�Ft#��>:��H��[/N2v3�'�����*]�1ϴ�0VƖ?>+���'�]�byX��ƌbצ���'�,e ���33l� �"b�
A9	�'ވ<3��E�r(��RÆY��S�'N�	�V��]Azyc"	�R@��2�'�:ȊUm��Tx#
�L��ՠ�'f�]�&�K�Wp�9gTW͚���'[�ea%��8�`Đ��@"Mc��`�'�&���\�8=���T�R��hx�'"��3"��
#��m�E΢C�r4R�'(��3r�����\)A��
�'$$"�o�<��2І�gkv$�
�'����ȇ</=ܹ�qO�qQ
�'��a�Յ�gS���Ԣ��e�t��'�Av��#!��@�Y<S�!	�'n��"�Ɂ!]�>U��!J�Hұ��'�0u�d
"G�Ɛ볌�;��p�
�'�2�(�Q-4�
�x@�Ͳ~��I��� �E�� �Sf��W%�w��Y��"O��Q��PZ�<��CˠB�:���"ODbw�]p���፴A���C"O�d�����U�%�JVP���"O�ě��=\�����N"1�"O<��O�0�|�ZgW7,Q0d�g"O|�Y�&s|��ؔHAL@Q�"Ol��욪P�����B,�p��"O$i0*M�2�t��V�Bp@�"O�7Þ�H��KC�K�.O�9��"OM[F�X,�d�mV�<�J���"OAr3�ͱ[�2���["����"OD�ڕ)ֈn��I��K͝�ĂA"Of\�G�� 6k�J�Va��"Ot}2�h�<b$X�e)ޟ;"n�""O2M#@�	:˲|q0���s���"O��@�F��,�R!K<i�7�0D�(�$/�7Mj���� ��H.l�`R/D�p��I.x��j�����;f�)D��QwkG�W�x �4���y��\)$�(D��⡎�X�6�[���|�%+D�l��S)/���D�z��(��@(D���'�E�M����M[�e�� ���2D�t����6Q���:�+Q�/D�  ��49�8ˡ�U:EV�<"�(.D��s�HTM�>��V◧7���"�!D��
�oٔX��� S#G���%j>D�H���L�-���$��&
�%y�o?D���r`�4"�-��b��x4���0D��ӇO&2��r�C/-)B����0D�Ȣ2a�!H�`�P��<	�+�g<D�\[��\}վ-Y�獄V/�$2�+;D����ę7V0a����;!��\)�E8D�`�Sf�^��A��=#ϺP�"� D�l:q���Q�H�
D�Q�ʜ��)D�X�Ԇ�v"�]P�e����P�R�'D�\��X�)b����(x���1&D:D��[S)�<���Q
Ќ�B�<D���!�3X���rw'ğ'I���8D�49��īhpZ�C�n��\dV��y�K�M�`��Q:X��@�"�9�y���T)>(y�N�
S�������y"L:q>T˶b�6����D�y£�0)�h@�F���Ǆ��yrF���tT ��)k��Lx��M��y��9����d��.����yb#Q�@�hk�؈7F��a��y�	�5��I��/T�C"y�@���y�P;\��6*+;���pe$R��y�f�n�j�A��	�,�:m�T+Ԇ�y��R�	Vl�h$�&�T�3̎��yb������A��*٘�e�
�y�# 3���d�L�CB�S����yb�цp�1#��%�>��E�-�yZ��Q�͙�l�2�p�����I	�'�����e�}���E�~�|��'�M+".M�f*v�6r�^` 	�'< (z��Z�L�e��kH&���'����擢#��@Z1��ip���'���S
	�pO�8S/R���
�'!JX;�+��JeRA!��>XĎ��	�'/�]�uޠ(\D�&��fe�	��'55����=>��0�k�+1��1�'2�P6���} �����.���Q��� ����^�,I����WcV���U"Ov$14�@m$�7
W�K(%��"O���U�X�	a�)�(�԰�B"O����M^7�AF�A�6䪕��"Oҙ�V+D�33iJ�[;E�>��"OD���옱w&�=���ڀ-�,��"O*)0t��/V
T!Ш�F;�A�p"O�=�0k��G���+ �"OP��W�FWڬ3A$Cvb l��"Oi��$<��&Ը,dV}0"9�y��Jh����.Y*;�H���y2N7T� # �C�,fh���A�yb�N@e�"FH��"5j��Z��y�N��x�p썞L���y�+@�55����C��@ä-A��y�l��s��9&��<c�%y��T-�y2ؿ-�$(��ɑ�:m�tP!���y�k
�.` )`�c�."����
V=�yr�� zͼ(8�a$��9��&���yblK!�`F��%��u��I��y�F��,r� �T
��%�ݳ�y�
(V��0�B�$^l�*�+�y����]�t��SJ��"�$x3�����yr`۰ ��kfkH��J�c�]��ybU�ي׬����bS"΄�y���2�2pQ1����Ԁ"�ڱ�y�&B'=�,�YrJ��~�V�3��ֱ�y���I/ pނ*�09�c�-�y�+�]���`���J�0�,�ȓX��غe�N�L��,�e΅>�ń�N�~ٛ�Q�2*��30B�20��\��^�����Z��R�@�t�Y�ȓ0]H�J"��s=�C�*N���ȓ+�@9+!(r��A�v.�(W���l9���}�����%"��A�ȓQ���e� r�!�&q.@��	�XZ#WHL�!��U�Z�Y��;��EC�*�}���̸G�	��5
�����/cTd�7���p����@Cx�!��B1y�I�g��)��4��s~t�j^=_RXYQ�'��2�ȓL�p\�Ӥ��d�fаc�*�d���7
� �1 �0z3�iHA+�*BDD�ȓm`A�.�X+��"�H�Ht�ȓz�PH�Aא\�����EQ!����p.v�Ӄ��k����`�2tU��^r�Swe�1��Y	�IO	!�䌆�cQ����$��:$Q�ڄx�f��ȓ=���O�5Rv%�7)s�6D��@U\�7hZ1
���QŠ�	 &6��ȓHG��kA�m؁��O�ސ��>� �v��:&�zl	�d�_�U�ȓ:X��G�I'Ur���5El��h��5�2MЛn���H��Иm��Y��W��]b��ہ
0���&�@6�@��b+�И����4a�̂�]?�}��(azUqc��#/PD8{ j
v�p�ȓ�rQ�5�����a��6�`�ȓ'@�U�r� �
v0���#B��2}��$pH���酢/ٰO�����h���Qg��>��� ��W�G�e��r�\�yf�ӋI(��֡Ǝ,��U�ȓO�BQ u_�;7*�R3a�&l-
���F%ni�3�m���Bң&+���S�? hY��_
T�`pԪ�����$"O6`�gK�X/��
��s��!�"Olh !�Nn��E��)<yQz�"O�M0v��$:m2��U@1^�
p"O��0B��2��#0�1_���"O�T	��6^�
4R� ���i�"OL� #�\3gC"���b�4`qe��"O�y���H^vq����5��(ѥ"O� cb�/w�4�I2�؞�<Q�"OV@��Ҿ>��}�%h{By�"O�����Z�i��y��)�2� "O���Ɖf�&Q{aƇ�2j�LZU"OV&�;r(��O�a��!�"Oq�1��z�)pU��*d1�}��"O���.�`9�$p7�^�23t�SE"O��2 ��
'̜�S�	��@a6"OV�.QC<F(�� c��)�5"O���KR�XLbp���"w�A2"Ofx%荺�8S����!�Viq�"O*���)8(��A��-���"OF�0cȋc��c��Aj4%�"O4X���ȁe^���ƟX���"O��j�o¶�-	��lاI0h�t"OZm���T*?�(�	��N,2�D�t"OX`�bo�vs\u����c/b��"O��;�:SRQ��-�/�M��"O��E���	~9h���?%���"O&�����'�����i<'���"O|���+�.2]� .5$Qj6"O~Is��TH�����B"2 ��"O�ʶC�0Jᨱ��������"Oځg�K�-�h(1��܅5��U��"O�!�bF8,ڦ0��BO�G|j�A"OT�b��4J. �e�[�Z]l8�*ONHA察�v)�����P�'1��;@;I���7�����'�@�[�^2D��5��߉l���2�'��p��B���ȡ���bcV@��'{�P���؉,��ĉ7jپ��)	�'øMr��L�i�F+� ���H�'������� ��X熟s	����'_��r��"a���$�����	�'U@�iRElo����F:�x��	�'�xXr�J��0s�b��P?Ք�Z�'��H��l(���֤z���Y�'����&���ڱ�@�E��:���'\�lk��U, ���i'�5z-��'������\��2UY����b@B�'ր�b&k�$) �T�@�JHX�'Rޑ���T���k�k��O9�'�F9
�/A0T�6��*ëB� 	�'�:ɚ��O�jGBY%�I�-X�r�'S��@uʜ�H1FM�D�H*E.�2�'6l	"cd�4{�<a�P�M�x��
�' ����nB�n8ސ��
��;��� �'���CCN�l��4��O�(3��(��'	�����P�«��6<\��'y@y��OP�S������YԶ� �'�xh�.Ո\�a��9I�,P�'�����15��J A;��
�'�Z8�g��cM�tK
�'��\*�le4"eA�8�9	�'�`kOW,� �۷
�6,�>�	�'@1q��U�:�Th{�@�[���[	��� ��#�������Z���"�'�B�'�D��~�M��cZ,�|�rgGP(	y!�$HRU�� F&Pҡ%M�iX!��ɮ{���P���Ԩ,��jڏ#0!��S�(5��>b���*�(�Py2A�S�~��h١W%��˶�#�y2h��Ḧqq2KO�s&"���y2É�,Ϣz���2*�Y�%Oը��=	(ON�	�!O�8�0M<>���ip�	3t{zB䉼k)8L��դM(䙲bI2lB�	>��A�]Mj D��o�*B�I�w�Lq�b�ږ6@M*��ďr�.C�I0Ij�B�$!�i0R����B�	'xr�E�-�P������!�B�ɵQZ�C҉�@o\��g'����$�O��d�8���B&(�hf�Ӷh��-��o:D��A7�AP�Z��#��%�Q��8D�̡a�W�
��cG��+��y�� ;D�H �"����dl���x5.%D��[� ����$�v�3L@���&D��a��P1I�M:�O[l��h�� D�|Iwe|��j؛{��r��0D�$QƦdP�飀ՑLp��c�/D�`)TfҦ+z(v�S(]ʦ�#h;D��)�k�;���B$F�-�p�ȣJ,D�`�C�٬��)�E�t=��q�?D� '`�>
j�y�ʁ�~$���<D�H��nO�Z�����>( ���j<D�$I�_+=厽��.]rX Lp!�?D� CF���W���ђa�#w �C=D�L�t�@�D",� �>"�q�ŏ9D� !�J��r�
��E��KތAQ��8D�|x�m]����𐥉H��8g�(D�dSં�N�$Mj!��˄ͨ!�%D�0*��Y�l�D+F�[&"}Ia#%D�L�NK%g{����E':*��1�5D�Ѐ���4��d"�l�.���T� D�H
"��IPty�b@���iRL2D��CF�ɬ�r��2�݌� �7�;D��!���>'�u�rEI"�$�5I;D�L
�,�ʲ�SE
r )ǎ>D�(�V��|F�T��ē�g�Xx�ǯ/D�t�b��� "��`n#B$�6�?D��R+Ȩ[���)2�V�fN ��c�!D��c���3��  �׍RGH�KU�5D�tQb��g���� �C,4�1D��bn��J������g`T� �/D�0*"
��z�.)��,���&D�U�2D�t!�� 4,����E�RBRu��2D��c�L`� ���q u��2D�@)EOB0+��Yrק�O��XS�@1D��;&iN�0�,Q�a�G����3D���B�Pf
 0;�Q�$^6���%D�ʣ͇0t� d�c�� 6X���t #D�l�S�\�+nM�!�K�f@�����,D�l�
��*��vG��b3t1�2�*D�h�'CԄX���򇉲od:��@)6D�㤦ƚt������Ďg�U��N>D�Ыd�)l�j�&(C�#���Ո<D� � �>�ؒ���T8|��;D�p��WuBšF'_�;7�fA-D���iNI���8g��(3�	JT�)D�t�/jy
����ƺte���l)D����I	8��PG$�-B�P:F&%D�� �8!눹LC��Y�>� �9 "O�љ�T�b������l�:带��S>űG���s\as6����f5�2!>D����)OTA�TMN���'D�4�T��d�Ѩp_o�%9E:D��(���o���!��6J��\ړC3D���ږ>��m
c��T+�a&D�� %M.m���v�#\��H�C�#D��0��'C�4�X��@�C�p�b-%D�HZ�`�5$���+\k+2@�Q�$�ON�b����4�^��
�Aa��Kr��ȓAپ`Xd�V�r@m�5��6*7B��k�AF��U���Aj�'n*���ȓv�ve� �ίP�8mB0%��~�؆�kn\�2d���8a���.`^�)�ȓ����@,,o�bH�E
� �HU��/�`�T�$h+&D����x�������o�6���9'���5��|����|�3ʍd*Ta)���\����ȓ��t�%�#V�*��%�J0���ȓ	�.xɀ
Z@u���]�ư���~���
K�< �K�5��1�ȓR�>]�a�{���ʙ�{���k���{�O��!6�2٪���mU�m�V�c�'u	W��r� iq��١a�>l��'��� �	|�x�[�-��W�j�'@H:U��$hQh�k�ƖGy&���'��$��&28�́�K��n�X�*�'��2��:
!����Ԟi�T��'�8���V]��y�$^�/�J 3�'2V�C'O�;+6��O	䞤����)��U�I|�$�����5�0�ӷ�yA�>��|�Cc#V�zXʆ���y�L���KA�E�U a 5�y��B�r ݂�jĦq��dEש�yrNu�QY�F�_t�IT�Ψ�yB�Ё4y�ʄ+X��	w �y���*$oF��2&�&}�5�6���?����0|zw��V,dR&��~��Щ�M�V�<у�ߦ>>�,�W���(�@�T�<!�'W Y'mkdG��8r�a�a�AG�<�C\�LZ&*��=�P!��g7!��l
��2�ͧ>�YD�(H'!��O��P��E�:
r��ć��	%!�/2���"N!�輫0��6k��'�b���\�C�(��j�`ݼ{�Dx�!��fh�EB��H�&׊ͱ��%�!�DP36@R9aA�;��i��� q!��R��p�&��1vĪ""�K�5p!���\���a�GƝQ㜵+�C/z�!�M����ê9�-y�Y:A�!��ٶr�1fF�x�4����_��'pc� ���p��<q�X�u�a�P}�4��iB��@ �R/C���r������>|��ҵ���p3�H�Z2h��e�l��vj�a�챕�G<r��ȓ7(�*� �^֢��k�S�4���w,x4T�a���<N,��ȓ1�ڔ�4 P�
�Q1�O�  �"e'���	�����e�Ou�9�'E��D!7�K<?� P��'�$8{�@U� 	�CgR�5�D)�'�> ���^&�Xya�R�1=H
�'��Y��� �8(���.�ʱ�	�'\��j�掍\�uh ��Nx�E���� �X��G}4�P��£a!N��Q"OTH����
�ģ�>`�Vi#�"OD���v8k��C��4�J�'��G
�44QB}Iሕ!U<B�8
�'p�y[��
@�
���I6�h��	�'�8l�2e63���JAH��,�.��'\�\�ֆKV��@k�.K�ӀtZ�';D��%�7b�!�Wc9GXٲ	�'J�@����3l�h��B^¥��y��"�0=�Ui7(�����5	}��f	J�<s��	7���ڲ&�H�Zpq�J�G�<���+l`��B X��<�t��{�<Q$�΃GB���4E۟OH�M��{�<ɲDH�`|ї!�w��Dі��u�<��m�)o���wdb֚q���n�<AeԻ��0�G�
&L���O�g��0=y3��=R���K��K !���{gΓK�<a���_�X({r� �\�詢UD�<QvOY	5�`�(��A�HXC���<A��Z��d̩�)� -���!"s�<�+ǐL*�#�Ѳ>S�D�r�m�<)���O	 lYE�H-L���c�J
h�<y0`�" ���SF�aO�ؒ�I�Z�'-��QÓS�������a9LQ
Q$D/!������ ����#U����b��B�
B��=D���p�[�&*"�y�Z��C�IJ����%%��k���qe� �C�ɇdu I�����d��H�G�X$�B�ɈLSּ�Q+�<[ d|�����B�I)k��p��cDY�b��DL�&�R�`��U���e��������C�0�+��(T� �@�3rb���@��^�lI:"OR���D�}�x=�0���h��"O ����%4T��*Ⱥ&hfAb&"O"9iT�/,{�D��-J��s�"O����6X�0�-�#kt�w"O��j�K%���m��ȓ�<ON��V�'�d�8���{�6p�ՏŮs����'��T@n��d�-���D��'ʦ�ф �D�y���ɞk�l���'A`����*H@Tc�cIa�^�
�'~�1�gKOYT�[w�җm���(
�'ռh(ŏYpP�S��_f�h�':�tp��^!���\�(�:���OZ˓����&qF����ドf�D%y��Z���[�f#D��zD�S�l2��Ҝ&R�U�se/D���abM�Vrj�I�&қJ&�U�@`(D�PƠT���P���!-n��%D� :f���!2
/P��lѸ"`#D�d�s��:��)D�"T�G'D�\�ц6^�hM���@V=�B��b���YS�Pr�H����g�;M�]�6�ޔ:���#D��Q�'\q�9 j�)n7�R�I"D�t��
�x�p2��-aŸg�$D���vM�`��D�ũZ/Kv��2Ve?D��c�F?f�t�ٴ(Dj�~yi��<D����L(R.��2!��G��k�*O�̒A�ǲb�@:ō�8.���E�'9�D��a|����=а�1�Ծ5�(9Q!ӄ�y"e�$n����� �-�ډ{ +̫�yb'�" v�Z���;:�H����ܽ�y��ҵ9'.��FF�-��A�h��yR���6�n�X���'[W 9��KǸ�y��Р"U�U˙���H���xBC�̀ Y���*s�%I��JP��Lp4�'p!�N�8�.1j��{ۢ�x��ӥav!�^%4�<�	�ɍ=�0DRr�P�u!�Ğ�u ��đ:�6Ē��*F!�dW/k�����kK�AL�JJR�7.!�D"C� i�-,�2�"��M!�$��8���D��=�d�'�R>!�DU�U���#��H�J�yF��,!��QU���'Bn�Xi0�B�>!���O�iɔ�;Pxx���"}!�:O����� O� �5�G�!�d	�A." #��� W4�q�D�<}�!��+�ό=h
D��@�J�l��&#�Ђ�`��!�HcB�I��]�ȓC���W�۱L��1��=N���0qxP���ޠƎlP�/E\���W��0C�@5��1H֯]?�,�ȓO��
�#�(��d��F��ȓNJ�I�J�,c>�� ��A���O���Rvh�1@|�x7b΂!~�݆ȓ_K�9yW�� v�H�����;HR2ц���Y;�� ?�l�)flA:WC=�ȓsn��I���4�Ā���
im�ȓB��C�ƍ.7%�8A�/W��d��o��+U
�-g�ðၬV7��ȓ%��D��m0���M+.�
L�ȓ
|��Z��2n�r�R'��'�&9�ȓ��bCZt�$p"�HL�(��5�� 7�0u��:[�Dm:d��r}�ȓ]��
%��X�faʣ��Y��)�ȓ�0XV�'(N�XF���N���ȓ٨x�q!�$ZH�P3�+�d��:i"��!˭OJx��!��Z�X%��F{�O}�ɹ^�J�Q"�Ā``��pG߯U}pB䉵NG��i �m����@�אCA�B䉐*�^L��Z�	� ���+g�\C�ɱHݘ�BdE�::����"ӱK��B�I�=��aHnΑ=Pԕ���ܑi.B�ɞ� '�S mj�S����%�B�I9��H�ua��^BD���U���B��0-�H�yW�C!_D��eƪ,�nC䉻t�4��So�"l���q���,O@C�I%%J5��͊�Y�>Q;7
ģ)<�O�����q�$���� ����u!�{m!�$Z�RJ����g֘W�0���9!�do���׬
1Ѣ��ԏ��X!��&vzk�B��|�r����<ig!��Ê/������x�iQE$3T!��)]t
U)$�@�KW��萪�v>!�D(	�z��!̀S9 �1�hԩ!���:G�г0��%p�Kq(>�!��1ر�5inb�<��@%=�!�D�n�H���JX( �r�팂z�!�F@\����$
�Nl�2��*f�!�$V����1,��!��|XІE�{w!�dͦʀ�wCF'3� ,�P�S�8[!�d[�H�����`�'�֥Y�	6!�Dؕ ���z����t0ר�u�!�� "L&9 g����@�͖*�!�dG�'�(�GI�z@�uygʈ�!�_*2��x��C)�L�@�0W\�'R��i�<s�(�(#��'�C�(1F��)�'o<$�ۤ-ա$�� �v8MC�'���C-c�J���H0lX!��� &�	ahC�,�|��sg��0!w"O��[�IJ�3����,`T�x�"O��)�L�X�+�HC�T `"O��s�N�
4KԬ58�%���yR ��p���c��12����d���'�ў�OF`3qh
�e"��	��#��`�'�P�öN�|�$Qd�ג�A�'�D��D��S)����A[�D��'e�H1�n�  B}`�&�2�||��'"P�k6�O(1�����.4��<��']�D��+�f8�3jI 7$5B�'��I�C'J�=ti˒ �t��Ub�';v(�AJ�,;�<��D�|	�'p2 H��_=2[jt��B�'}]��z�'
^�s&�X�@M�d�*ĘZ�'��H��ڛDF�1���*��� �'l�\�"�W0��k0��-��t��'^T��"n�.i�TQ�W�)|�Τ��'_�A���|B e�I�!I.����'��l;���D���z�(�3c(�q�'n���lG?�����K��y�n��M>i����^\`XU�dF�:p��ل�V�S�!��"Bp���^-F�	���� a�!�d
���rǝ9B� ��%��t�!�ĒRu�i0e	!FW� 0Ҧ�'�'�ў�>���ό�,��c�G�Y��0�!D�4ۗ�0R�����D)&�Ф�e�=D�l���ر7�ԩ���'�<�@�<D�����RbBM�FKσ���z�m:D��j� �o���f㟹z�x�`&9D�t�c�]�Q�R���?=�J�P�L1D��Y�mU>�9@��ϙ,XDrD0�Ijy��Ӿe��ʵ��C�����E�d��$/���ቂ�J�L�SA����}���8D��
�(�-v}f��'��<Z�0��+��Œ&eK�*Vp�j��Y"�*i(�"O9`�Y�&�(�1���3���r"O��C���q�ju����	�U��"O8ݺd*���\�JW�۩)����f"O����)��z��J��"}bw"Op��s|�ݑ5	�,=��q�"O:���MܸC�L0q*ܮo�.f���O>�$*�w@�h���;3��a�R�H 8f:���%�ڄ����]Ӯ<
g,�Y&���pb�d��@r9.Y6��8T�μ�ȓn��st%�_B�qH32o����#�C�g�	G�$���y�0��ȓ/��q�JO�0}I�Q*�@�ȓoĔ�S��	5D�jL�Q����G�S{b�yg�ģ:�&��ԃޅgB�	��dY�ȫA����t*���B�	lL�dY��9��Xj�À�*C�	�R+���%�f	ܴ�6��>P��B��&{��&��QܰP���b��B�	 ��P/Mx��H�iZ�8�C�If�v4�Ca�{���K�EԦ[��㟸�	؟�F���!A��9!匏� Hu�Q��y��ϲ/�e��� �d�@�Ǜ�y�&�,$�<p3so�F�L�rq����yr+ڋ �J�1�<I�Q9R��y�k<NTD0ӵ�ԙ8����Z��y�⛈��(��	3�h�[a�R���'��OLl HC˭x^tXA�W_"��'��� �C��c��� �_�
 x��	��� ���0e9�ܸ��m�=k	:x�"Oyui�(	�;`�п��Ae"O
L��+��fXi�r���M�B"O �b�E�� ���C�UH�"O�5�e	X�����K[8@>	�g���O��ɏ�v��tk!�9I�PubG�7(!�䊦@O�r���8���3#��:"!�fg���sOǶ�|��ƪ9!!�D�m����cjF�PJN���j $sy!�D�%Y������-�5�2`� v?!��,P���3W	 �1J�!�D
�dr�	�0� I١)U �!�� 0U��r3l%�Б����A�!��K��&i�&ȥ�{�Ԯa�!��K�Y�	���4�4D�MO!�$Q�B	~�ꅂz�(��$�؇V!��E�(kƋ��X2�ا���g�!�Ą�kƚ����vA�蠋D%C�!�D��V�Z\���=�m{�+B�k١񤓭�$��1Mn�R`AF@Q�BC�I�1��E ("YQ+Q�u�C�	78r�� �J-:lX2
N�}� B��,�R��`l�H4|�E��5rxB�ɶN�xP! '�>!6Y1�#_"B�I�@e�	ᵢ��Z=d� ��(w��C�I�9�b܋��Y�{��$�1� tp�B�I=�ڐ��C	Wn�Ԛ���;��B�	�%� a���+��7@N$Y��B��%�H��?6T�p��c��B��B�	&j��cCD�3�`�3�޷G�<B�I�9ز����9�*2)Z�T�xC��VOV\�1)ө"�
�J�X5"�,C�	���)�(Y=3�8��&�:"j�C�I"PF��Ɵ;4���D�R;�C�	2*�tq��!V�l�Y��AL�\C�ɴ�"l���n�����@�{�C�I/m"Pه,�@!H�gA�}�B�	�-�*��6͙7UOƑR!�_��B�I�r� 2�eٱW�he��#c�B�	��t%� .QT����`�,VҴB�_
ى@ϛG��`H2+�6]�ޣ=1�'5��@2�@�M$�Q&��7U��5��c�NH�d`Q��x��UAͳ���ȓ)kT�+�i#e��P&�-bD9��}OX�G)�=\+V9b�Mɢ���ȓR�IK4�*�
	�5.�%v�*ȇ�Z�qg(ɿv���v�%^�A��/�Ռ[)Z����(��j��G��'����Js&�36.#~� �2j�0J�!�$�Ct�ʑbڳyl>p@�7�!�$ܿ�Mb�M�0^lJ�C���Q�!�����Њ��8RWƔ[�  e�!�d�>0�p�A�;7ИaFG&�!���7�u�5��*(1�����6jb]���I|�$�G����yB%!I�
,��N���"��bJ���y"BS^+>��iԇm�x�Sg�2�y��AJx@"�N�g��!Bi���y��ʽc�@�� R�]0(jQ,G�y�N0MI6
[�[R.X[t��6�y��Y;@���۱��Z�yz�-(�y�lқ	�P�(�,���ŋ���&�yBfO6�,��dꖈi����!	��yb�Q�2|���F�ڇa�j��j͆�y���,Q��"�1F�"0�@��y
� B�¤ߛq�:��!� ��#�"O Aj��R9.���0  �H��;�"O�S�(�;4*�]ه.�_�8�"O
l���V�)
��*W�I�����"ON�R%��	
U�1�p�65��P)�	K�*-B��s�d��d�/���ґ,�>��I�1D�H��G/Q�&,  Ƹ�5��1D������v��('F,Z��H3@.D��B���2'�@���N��ș�fK8D��R��x���2#�-������6D�\@�A�:�&���M,��Hjp�5D����/S#>�3��,n#�p!�4��҈��	�0�^��ggд5�HC%"Oh��ԋ�/\A���,<�ր�"O:��ҵt/�8�"f�&���
�"O�T�R(\/S����Q�̨%00�B�'4��h� �d��i�Qb���(�'�Z��N�9<%#a�(�(��'^8qᄅ	�|Ls�G��`-�e���D�Of"|�cE�V��-Rb)�+�*f�^�<�a�ê8s����jN�M���I]�<�DK�r?��&���^�a�GUt�<�.Хvdz�� ��
Gd�!��D�m�<1уz���KBl|����a�<Iª��xU��֝�����X^��I���O��E��Q�W�h�'
%�6�"
�'�
��V(��4U�� ���|:	�'j֝2�` �Q>H	rb��*Ț�'~� �G��l$btK1��!^xq	�'��(��A�\4+V�� R���'���K�ʥ1b^II%Iô}v�L��'0 �ɵ#��E�~-�t-��|6j90�'@j�sFkN�)�Ta��q��	�	�'}�(c�̟0�E�Є�yL�%��'j�k�-�r�\<�ƛ�G��3�'�>��Q; ���+�� �Sq�Ղ�'aƘ�B��<KϸiI��5L
|�:�'�&�p`�ǫ�FLr�nЙJL ��'���m^Lh�ty�΂�_!p�"O�[�"��BmM�M�,�k��,F!�䞧k�Lʃ�Ԋ]���O?]&!�d��h����	��Ƞn�/#!�$=A�*|�F�%l�X9"�ǳ}!�0V�{a�!���9��D�~!�D�AU�e2���v� ��X!�d���Q��ƌ#T���	��O\!��Tg`�y�����R���"�_K!�E*��Iv"O��	B�D)�!��&m�бi�I�ʜ�`��((�!򄏼W�H-s��ݮ	�*���CF�!�$u��;��\$(�D(�cH4}�!���I/��P�
��A�Jx"W�N�!�?�6�p���!ʶ�3����g��Ox��?����C��"�r�3�2q�\x�"O�sՁ��Y��Y�)˳O���V"O>�jR��$������э ��IЖ"O@���� �\��9�'̐�4qD�z�"O-;��E<�x3�I�� Q!�"OF�!����?
*-J� @�u�&"O���7L� *���v(�I��.�S�i�!c���#���)�`yb�!���!��]���X0�C�^Ĕ1p�Y<l!�0�P���T��Yxg�J� 8!�$ڑ{��� �Ό�C�!��
�2!�� �h��,g�lѱ䬍�^�`+�"ON�2�@4k����,D*o��!�"O@��إ'���B�(S&���g"Ob!"��
�CWi����,y�q�0"O�p�	X)G����Z20���r"O����ɱ9���2#��P��й�"O^�"��G1�HH	A�\��("O�)�
�.�
ݒ�M�h�|��"O�0�g�P�Ҟ�¥"��^4(1!�@�^Д�s�ڦc��ʦ���V�!�d�8i��°"J�Qjp6c��u�!�$�.v�XA0A�`N�$�<�!�d^b��9!4"_H�ep�	Q�^z!�~=�AqƆ�	('�a�!��<ZmRjZ�}���"猥2�!��<;���h$Qx���i�|h!�dN%U609`M�{�n|уg�k/!�$��0�x�P'O��ax�Yx���?�!�dD�*W�L�T��
M}.й�`��2�!�B3�&���H!P�����σ+b�!���4�tXs�Ǌu����K�o�!�$��0����!�=*h՚Uy�!�HV����&�"[l�Ǚ
j�!�Ď)"B���`�ײv3���
�!��.�H���2����0$-b!�$H\{V ؕk r���w��,{,!�'w�h�PU◬�� �G'�%J&!��Y��8�S����TG�X�!�d�"K��-�F,T*�DCr@��n�!�æXQ���] be��3a�S�	�!���9�v\˒KKY���Dm�0(�!��8 z�Ȱ�)�%�b�%�ћ7�!��If*.���)%��%�a�L3T!�$E�^e�	 D�I�u�$L)��K3!�d .tM�p1'�ǻw���P�w�!�D��^�!���.:�	w���!^!�$��\>ڼ��jކ���F�ƛd_!�$�P�Ƶ`,³z
z!���G!�dŹ'�%a��b˾ ��X(~!��� D�qcrB�̰����3�!�0U��9�0�J���Q�ާ�!��X�jŃ��H9,T| C��R�!�D�4���
�7fh��3�C�i{!��*Z��s�l�25��J4f۶Fg!�$�>!e�Y��)��g�:���#;!�Dǈ$�"H��B��>H�ȩ�80!��Uݼ�YPi01������(|!���D)�!jV�w״y[�ֈ!�d�}�n�s�С0��\��'Q�
!�D kx:,iv-�9����7�C\!�&�Ҍ����#v��9��ƑI!���*��}	gc�{�R�xֆ�
�!�D�^�fP�BJ#�Fa�ƥ�t�!�Dy�*9��
�&	��A�䒔h�!��ւ9PE�hb.M8󢞆/�!�$�:X ����
�:]N��!]�Y�!��C�{�4��k؟M@���vUa�!�X��*e�HP�Jj�	�̖�#�!�D�
_��`�ہ�zaN¤�!���AT�(agڨW��� 0k��t!�dP�})��1��>|�DeHH38�!���D��`��N�3B,P�O!P�!�ցa�(���*>ҡȰaןs�!�$E��̑S��4[�
���?(�!�� ��C��A��� *�`��L�W"O��#��9H7Lt+O�����"O*��%�I�d�D:�����"OBL��I7m6,i@�K�)�h���"Oջ�!G��X9�ڄ��!��"Om��E�#8b�#���|l�&"O ��r��.�-��c�,�yPq"O>U�6��Mv�l�C�A�DZ&"O�xΆ�l�&�+"W�Pũ�"Ont#�c������b/�N�\M@�"O@DǢ� ?p�:��ݴZ�RA"O>�b�g̺8����$�s[�h�v"O2AQ�oI�[$t00ᅧN^��"O�� Df�=/�z�{"�ř|C���$"O���F��q�*	Y���9�\z�"Od jwO[�{��]c���� .���d"OV\Rv.$)�8C�f�xf�S�"O��8�A;e�5�����/��p��"OdԢ���4L'�= A� �X���:�"O�qڂm�%g��E���g-�h�b"O�2��]w|�q�ԗ3fp��"O���I��_-����#X~�tpq"O8����S�3�\P��
�B�����"O�A���>��ԩ���(+�"O.�p�(�1�pd(�Ȅ�a�����"O��W�މIsD���`I1`�Rt"O��Zǫ�q�e:� K�bY\���"O�=��
�(6�e��/�C����"Oha�Q&��0�^D�A�J�b��x:"O\q��ʴ9�l-�P�3,ѢaS"O��6�ĐF�`t���2ʾ�zB"O�i���W�4A8�\(h��ty�"OTp��M֒7�U��*l�����"O���+Ȉ'�QT���a��=��"O4M1��-8j�p��J��}���Q"O�|B%�/"~	ZEl��qeX�J"O��@V��)ɢ0q�J�(Q<�"O^us�'�7�������)>�"OV����ϕ �a��i�5~)R��"O������.=�}��B#t��8�"O�	d��
* ���v䋴
TEp�"O*��U�ԜW��S�� 5c�ƴ��"O\��S��f�V�E	�}2��"O�HSˁO9���n�!hj���7"O�X��F��كe��-2bf��"O��'�H-U�R!j�~�4��"Ot{u���#Și���5~���u"O�05I�.U�"�A��_���	�U"Ol�d
�=^�,�V!�#$U(���"O�����\:)��]����FH�Y�U"O�i9թ&1����1�Q0FO|�+a"O\u�D	��z���eG4U=��[�"OdSw�W7_���ݠv��H�"OW��*Lن4���	7/F���"O�(q!mH��ָ���A����2"O�i�c� �h�N�t慹�����"Ot`KV��H��,
"E��\p�0 "O�P:@쀛-Q�}�B�	����"O����ª.�`0c���=����f"O�l
F���_�JU�7琋l^��ӷ"O���Q��6>�A��ENPM�x""OȔ�1�Ob��s�"YN,3�"O�� B�,s���.;<@���"O�Pb�b��`�AL۞:��"O� ���a�8 ̨u� j-J
(�$"Or|y������c�T�\�n��"O��r��d+�x���\�ri�"O��S��r�TX#CT"��a�"O�)"E��⌝��bޙk� "O���GR(��CEB͖9�( �p"O�#�*�:#�����cw�鲶"O^!X�D�\q2�@S�eτE��"O\�2&���T1ֹq���0U&�JR"OB�Q%�©F��/%�ơ��N��y�L^�U��{s� .�]���y��u�V}�!*M�s
8��ď�y���;�Z笉�d̘����y2N>~gDd P���BF_�l���	�'W�(p�K0-�u��c���	�'��!��kL�(�F�)T+��S}x�C�'U 5���,���"ÊH�H��PX�'���C�~�������:�����'|�Z� V(8�����.f��
�'��=:My:��Aw�؜R�
�'@���w������;w���	�'��S��i��y��H�b�,�C	�'�ye����"�L�Q �b�'����Py"�4Z��R�H�r�q�'�u{F!8Z[L�Zem]�u E��'R��Ӄgr%X�k�k>r�'�%��Տ;�x�Z��z���1�'����BC	 E^m�k�.��
�'�~�2G��`��I������QG�<AR������������pГ�l�K�<�EC©�dh�ʅ�#���c�J�<�!,J10��ii�������祚E�<�cႴp����t�w&�`�K�~�<�f�p�|hӓa�`��h2C�o�<i�M��Ͱ	�u��\�`@���h�<� �y2X	1��KIbt���gf�<�.0�������N5��-�w�<��&I+J�6d���?@!��Ry�<� L�],����� < �V�0G�HZ�<��D٢V��k$�40�8XD$VW�<ѡQ*����2�'w�<����~�<W��?-=$�iU&-��w�<��Oə1 �͉E!�D��U����r�<�/�0l�B�ңo�xQS0�JI�<i�
��\�qq�A|h�x�n�C�<�S�+z�w�!v�8�Hk�<���փ�PBXg7�,��"
o�<��k̀�@t���~���l�<�D�κ,N����*|,���b�<����k��\�_�0�ZG�3y�B��&��AT$J,C�$D��� ���B�I�cJlt��&�>q�Ļ��w�B�6��u@o�T�˦�ېCSJC�'0{�X)��]ux����t��C�	t��!{E��4g3ȹ�S흴��C��$���)��1��qi��Τq��B�	&Orf���B��d����|��B�	�S��Y���2�dr�	��G�B�BFFM�2AD��N���2q�B�	ix�Dvˊ	a.t����!ny�B��i	��#�CՀ?Ʈ��g��\̜��(:D�L@��t�Rt�O�:��|�S�*D�����<m�	82� "@j�� �=D�4��j[
T��8hqO �1��9p��<D�� �Xf����0��!UE[�9c0"OlXs��\y���r�+M�C�"Od}�2�[9C��E�aڴ���"OFպ�.K	,f�P[� ��]����"OV�E؅5���&�ͩg��	Y"O�iQp���,���d����4�Q"O$�W.uS
8�hW�u�2Ր��d9|OD�� (N!NL���kem�+�^�<��G~E��q@ё1��a�kr���0=YF��^�챀N<SvA�3�w��E{��'k�Qp��=)�6���0=y��)L�lX�P���)�~C�K1�yR���YGv���l\m=p�m����yr(7{�U(S���e0n��	Y�?����=}�r�;�C�+���ZP��!����<�	����TL�.+^8��p���A ���ȓZ�$�X2�HZ���Q��z��)���<����=H`c�@�#�mlZ\?))�!����x����_�][�G�3�&T
��'%�I5���q`���e���sQ����	�K�Q��}zs劒j���+� u���%Bx�'�a�T�@L��m�V
s�EI@�2��C�I��j�b��{�6�.�J��1�S�O����&8"�J��NEQ@��
O�I�'�'m8@���	�8R.�����MK�O4�Ia?ͧ���M�H�0w`��1�]Jk�@�c��8�Ѐ�#/��m�x���va��'3Z� J'!=D�x�T�,"(By�ti� .�x�a�6}�[s���OD� �U�8X^�9t��eF��'�铉p=�0�L:d�y���F��B��d�gD���$�#	�nu:��
�Fb�4� �Ða�!�$�6�h�!�F���p�����g���{��'-赢P ��+�.�	!�ɀ����'���A�@���P�']�|�r�'52���H�j�h4��&L0	p��a��퉄��_)CV!+B/Q3L6�X�̓��O��$Ƀ���W��}Iй�2o�('����Sb�4�v�`ɀPLܺ t��ȓ%$��B򇃠P���!(B�_��%� ��'��>���$lb�� �
̌d_Ό(�-D��q!�e�n���]���'1D��#K
�p���/<�B����*D�TӁ�H�d8��B��B�`��*D��ړ� !*X:0K5��T����)D�LC�.�,.9c�
�g�����(D���ʏ�3��ѻD݉.����%D�(HD��!DE�	[ #Fh�)�j%D�8)n^d`�՘�&�5�:�"�%D�8ʰ��[���Z$oH�+*"8��/D��
�fטk��	X6K
�'$��s���O"C�	�h�}j1/
)$Mp� ��<2/�C�ɘLx9PQM��c�"E�6JZ#.V����w2���/r�J]c"�ļ:������2Q���'z�~R��*A~0r�Y�l�A���y��H�3z!*d#�	P�<!e�֠�y�m��J넡� ��"�p�e����=�{���2mk k$m��{�\5m	-��:�O��(�Nr�f=�N�$r\T�@"O
5(I˝!�F!!S*��om���U"O41�J'2[��#i�DN��96"O���P
۬W�2��b�������	�]�qO���Q�D�C�ǥM2�{6.�t�:C䉎4B�sJJ3"}Z��'ē�<�C䉢R^КQ:<puȲ��#���s���  ����:A0��sLZ$;y��7"O����˨l��D�ŨL�=QH���"OF)�E��Jknt���>�<�7��@�'dў�g�5�@a��L72���͏'2$��ȓRW��(#K��ʹ6�j��+Ϸ�!���d�q$�ϊQ�$W#!8aDx�S��D��
��gH�f\�i��M������'OȽ�Ag��`+ʽ��,' RZ$,�(OX�=�O΀e���JM&�v�P�i`���'(��S���ot<��-ȱWX��O>�F�@����7t�RD��	rJt���	V��*<u(�<2���V�呁E[��yB�'�T���`�p@��յ	�P5�'�|�{p��`�R�O��L���'�/X�
�*�t{Ҁ�S���?Y�'��	�L�|N�Lȁ�Ʈ2t(u�'�6!�C!�3R���.��1Dv����#��<��p�L��5G�	V�T�he(@Z$2B�I�	� ӖC�e,�@Sd� 2�Ƒ�"}�k�8�r)���˚���Yg�T^�h�O�� 1.���c�Z�!�z��"O��zBH����0�(ɻp��[��'�󤘓r�>�T��:$�J�Ж�+K�!�ٮhĸ���Z
fV����ʾ.w�O�}����@��"�\u����"L��isF��yB�T�Y�LG3�Ԉ�R	���$)�$ڼ�0<�1p�`K��3]x�g�R�<Q��D�H"�[���$B���qJ�'$�x�c�*�5��3Z�X�{"�ê�y�.�+Dȳ�*$��}�����y2D�9h�]�?a��b�ٖ��Od�~
��O�n��2"چ(B��I6��`�<�q�����Ļ唄O�.�q�)�X�<����P$�e2��ѦvX�
�WX�l�	{?�g"�b�� �-�ؑ�D��<)r�Ãc$�!heˌf�yjr'Uy�<9�d׏A4��S��]-GG��e�]`�<q2+�-*��-'C�Q�B ��hOp�ڏ�4�~42a�*���gH�v�%���Ie�O��СG#�Q�\iD�
��T��'�����Q�'u��FLV�}���'��H6��?m^=���V�ru����>��SDȳ�����AIDB���o���7L����Pv㞀+nP���w�Q�@���ħR#�Aa�3T�J]�<���ɂ&7��L�dn,R4Z�Lߟi�!�Dɂ#&���Q���.�t�!��'�!��O�����S	k�0�x!��-)a�I{���x,�n	�)��`��D�:+�X��xr[�`��ɘU \�@�<SS~h�u��`VC�	#g��rB[u�Fi��JXM�B�"�c1#-��T�4��"U.��(���O%����+�+
�CݼeCA��z����?!f-Mb`����,^��i2�|�<�F�C5u�`б(H�>��X���z�<�$��*BYF��"2�a��L�<	��A�)@ +���+��=J@��D�<13�/��A�/���$*&iLB�<�f]�:(L�E�=;�"���z�<�4�Z���wH��&�p@���x�<ir*^�!o�����j%�,���O\�<ٳ'�>_ɰ@jQk���4�S%�[�<yt�'�U��Un;���#˛V�<���Z ]j����1oV�a{p#�N�<� ���-�S�	���ӁWp�v"O*���T1Wܰ�Ĉ@�B���r"O�9p��8[������C<0�����"Oj���T-.���i��z`ƈ"OyA]!KJ��@)�R8��0"Oڌr1��Y'�l�u� �},����"O����&Pw�����1|i�F"O���D-~�ԍ�gŅ�l��u��"OL< P�[C9����҂>����"O.m0�P>P�Y�u��jk���u"O>�7e�-^����u�3.Ljy�A"O�dh��b����B"��&�����"O��CH�t?TL�ĀF�O�P��U"OX�*F%(���z�l��
� ���"OPP(�ria&!Ș+������y��A�I9�)��C�$�b�Q���y�'�5i2��{d"��dht��+�yҢX�Orl��V�eQ�p�g��y �-fd�qa��;4˺`��n��y2�<Az"���0^n`A¯��y2d%-�@ j��� �@2���y᚝�J�."x�B����y�
�nt��6�����[��Y��y�
� 8�V�a%#��S���y��Z��v�9G$L{
��8��R��yr�ۍZm"���Bp��ҏ��yf��/�L}K�	�AHz��G���yBK1F
���%E=���p�@��yf�h�l9�g�G`��0k��J��y*W zbXy��0a �؀�E��O�\"�J��{,Tq��S4�X��2"OhI�
�/e�\�%%M5Q4���"O M�&ݘ~�:�E�?`W�Q�"O�yk7��H
������&�>!�"O�b�>*X��ڷ#M���z�"O⬡�i�Fw�D��%�
�hXp"O�A�>c��xx!��z��x�"O��r�F�
Cc��Ղ��=�*�q@"O*�b1�J�V �U�j*,�X$"Ov0ee+M
"����8��2�"Op`+�G�Z������5k�n�)S"OB�{�A�E "��̊'(��pP�"O���wMѐ;A���ak�(_qP�SF"O~%�X�1�8B�˩wlx�9b"O.�����ѳԁH/P��8W"O詊���3m�
"� �:`Ђ��#"O.J+�B<�=�o�'�>��B"OLdq�`�]!b�� �V�1�\��"O�S�荪���qʝ�J�����"O(�!cI<h(U���˼f����4"On`��(M��d��鐳)�H4h��'�9���#le@Q��`[!wB�QgC�:�n��FO��{�Aޚf����eI%Ti����	�~��d���Y.��p�|r�H0�j�޿q����%�_�<iD�ǩE��k`�2 �Z\3�����(E!Hw�iV���j���sӆ�r��ɿ:.X�BuhB�A��4��"O"m1�l��[�\����S�`�c&g�֟<[���-)��	�F9dq��	�6�AǏO�5���"v��Z�6���&xd��D�L8aE��lQg���sM�/��HP��ѕy����G�%�r�	�WG��+&E�Z{���O�:B��@�$R<��tG�~���\� M���U쓚Oւ0�u�M�<p���	լ颕�B�8�������[,\#Da�`�	qΎटP�@b�� ���'�h�H�n�|�A�Zd@` J	�dBdR���0�΅!ƶ�"m�ge,8�8��Y�1�܌(�.S{[����L �������V��J4�͔/I�퀂�
� d�� 1c�M*I�R1:�&��$�pTy�EG�4�Ό�� ~�Be�a�>esb�{�pl(P!���0h��=9�y2N@�v
4�t�@�dC��ˢ�H��2!�2N��`v�Y>,���ٰ�/{ �ĎA
gF���g�.&'�lZ�	ӥ@!�T�������D�'M��0b��"��)ʧB�\H(�$̂y��i��A>��"�n�FD��gN��g�����
kj"�A�v^��u/!T���Gz�����3��(�M�j��s,O��:�d4��&>7��_)�@��J3Cr�yp��,���$%Ny$���i^��x���)IX���`��8��m#�}�bN�y�H�c��
_��2c��?N��{�N>�0ċ�e�n~�S�;t�I���JYn� �׉؁z�2��C'�|��q��Z$>(T`���7/,0e���%_�A��&�~�zh�d����v����+��OO����s@#Hl���^����)J����p�dV
 �\}ѥ�����C��"I�s�5p3�C�
�m���DQ:RS�Nh����:7\PXCD�V�0�Oڲ��A�C�*��Z74��h `�;6и8�� �4a�c���c#-J��y1a�':�)�4ר�0���"m��� f�p�V<���5�[�Io�'�D��$�\��q�D�ykl�h4�<����DF��q�P&���%NХW&�jb�H�$����P+�M�Ԣ
XN
��=`=��\�H+�P�ń`Ӑ���G�/Ai̱���MThZ��R�@ybg]�\d@���<�2EI�q�j�y�dR�\�j�OQ��I7j��x��c�^2"qp����MMȰ�y �9?A�c�F*��J�IY�4��:�	>bK��X�44.0��S�I�=|����_�RY�-tL��c�;��Ƞ�U��?E��'��P�Pi�;w��4�sa���7ɥ�x�c�m�:����ΰ{��D)׺u����!^���w��@:�{�-Y�6aN̛��0�?a0S�׆�
����=?+H>��96 )K�.��0��B�ţT'����K�!d�Y���/qR$rک]w�{򦟚 ��*OtՑr�z`�cāZ�� ��:���ca�$PUHh�%:�$G�RRX 0P�[�$}�೪� 9b`R�ŅR�@���E�h�.،o�`���6u� %�p$)?�Эښn��a
�� �c>-c��6
��l�A)[�{��}Ae[�W,�A��������ߕ\�Ub5��L���ۨy���s�]����
9�d�)f� \D����O*����Va�d��A��"~�ɬ|�&-{��3 RE2A��2>dZ�-S�a9�,��U������d>%cV�1%HqZ�
X0;mN�I�+~\�p��X�V�Jȝ�B���k�����
�B�B��{� v)U�����0xӁm׍v�J���6n���I�+B��`�8(Uy�V]��˚�G�$P�<���ZF�"\��8owl��O*{=Xq�-�2��㞼�r��Q��K3!uD�	)j#L�A7�ݴN��e�3��tH�5iB!q-��4럇8pdb����a��C>�s����'>��b�^�@��e���_:UM@bc�?'���i4�5}��K�!1��C�MA����I���xK@e��k�$5��
�o=T�@�-b1����+[�{��x�2.��x<�Rƃ�z��a����)�(ҷ��,a6���wk�}��T��'E(���W>G̐x�ƃE��pi�2'V��q`P�7TJ1����.>��r��1Sј�b�`x������(;�[��C�����W���O��S���#PP�F�6k\��q�d6	nR���G�(:�
���B��Kd�]�Ɣ�≺��3$���sgCV&�`�eEҫt��{
X�v4f��� W� �0�8��ɲ"��( j�eI�QJS�ʱUV�S�	KS�a�DY�iAV�Kd@,�~ T�����{�:�1Şp�B䉚]:���J��5 �8��oܮfþ��eA�|���[cbN����,��\4��w��>3+�����bʪ��ݴA8PP�@�d��(�[(��E�鉲M_��"ȗxö-��BZ"j`���m�l挝���Cn�� �6�W�O�$���ٚ� ��f�M�nv���Ď�Z.� ��.�;�N���⍕V21OJ���S?���Eb�9��h��M�$�D)���\#�A�	�0J���x��%p4�a)t@��,��OZH�'9>Yg#��C��9a��/Q�Lz�nR%= ؀�� o��BEn��S�4I�s��HF8�֬.U�Z9
�Ӧ;,̠�T�E�m�
��ҤIzm�@�N'��#$kN�-kqO��G4� A:�[A�x*�$ݡXp�eQ�O�2��#�I�tB4��n�+Tt��B��B�:�\Y� ��Xᶜ"eǋ+P�2��S��qV��Ί�W|��*ehc�^�� ���5�,�)c'�:E���H�Lկ7`�q�m0s�K$�^�G�T�� �v�q�pƌ��y�CP�T�6��'�P�R̐Y��A�;�R$������}ReL��QM��� jc\������T�Q�l
fJ�	<@Bɱ�؜S��B��b�b��#D��Y8��U,)e^N�"&
�	=DD��c��U��J�O�V�C�@�<������,E�͂�L�<a�۱��(O����.A���4L�>e\)u��]��p!�]F:��a̚SĞ���`��8�$B/˨e9U�Y�Z��.p9L�pKǰi_DS�C3q8L��EթY|�xȵ�O���S��(�KT�_�b 3�.��l�����N
�Dݑe�G0d�B�����X-�A&�N,nG�y��O:�����5b����|]H(31b�3Myj��6-X<8������?��)�Qo6���a�E��i�b�H�zMzE�K��T�$k,�D)�'Sk:�Ta
�A��u�V"��O�n}J���$9٠���DK/=Z�V(DR��qO��hX��	�e��,R���U��6#=��)�]�ERsG��JD�����[>5v�X��`��7}T����8+���+�OX�i#�D-IC��o�7}j���+��w�9��ň\JL��P/1�@A�#y�ў�ra����S$�ͫ\^�Q��ˏB$�Hr,#~��h�$�.	n��X���� �h�
-,�<��ī�/>J Ѥ�H�X����"��I�2��r�E��q�$E�[��m����rq��M<�6��,��8Zu�\<[Î�����i���ځNO"W���E��h���{p�X�A��@Mų2�ȑmZ{�A��6F���FԻ7�p��w 0��c�<y�"��"���ÇF�p�]��'Rr'��pIJ�yd�Q��'6N}&17��!����w�y�]�T��s!��k���;Nz��g�%j�\�aAS;P��q�3D�=x||L���5,OF�[R�ͼ,�^�c [�GT��0� #���˂M�����p4e�	�=R2ʍ�+�^�S`�[�DU�V�0@HJ���@�Y���@C���ٕbd�#e���D�Dhy��dJ%i��@0j��vfl��wB��1�p���7+�847��[��y���x�J���K�c=������p�|���L�:01� ^���m*����I1?��u��|�1=��i�v�ԛ�h���A�Mu���m�V����0*���E_yb��r�F"+������Y��g�\�/�z҂�	5 ��*�ş{g1OИ�!'��j:�JեXl��z�͘ul�f�@�QZ���vJ�4_ڈ�G��i= �
U��o����7al�q3�T�(�:`�Gk�c�x�gD&2X��r��|���V�7\O����P�\
pL�dRP�ХIP���:ՍD���L86EU�^��pL�/Q�^�)Ǧ��' ��3&���l"B�Y�AԀ%�d�X0=|OF	H���ީF-��!f�Y�`��r �բv�P+��\)&ޔ	ƈl gB/o���A�L�#b�U�P�H�s!�ѲF���@b�^1�q[����!���dd��d#=1+C�9���1��iI���V>����͐b�����E�Bw&�;�C�ئ�#�9�0�h�~�r�c� ;�!��O~�f�h��r��Ȓ'.}Zw�'G�ِ��*��׈6�Z"@�DzĈ	F���E@ڐ
��(4�ŵe�Zҁ+�&�~��P� @fPLCf���ȕBBL���>�"��m�|��P��Y�QJ6Eğ��F�9֦�ѥn٧bX�e�B-��?� 
�Z�Ej�+�t�y�	 �,���ӄ���@4J#H*�D�B�X����#���BT>�Tg�W��	�LM�8i��C�Is�1`�J������FAA]*�Ʉ'�W��Yq�l���E�߯"1�͑�͇lQ�l� )�O�M9���'�r�G#)raƨ�GFC=.fʀ�e⋄6r�
�f͘|k*��M[&�|8�c�tnܘ�Ǧ�/dΐ��ʆ<�!I5bt�H�OՀs� r��X�(O��P��I7fd�fu�:="%
�E�@�c <T�9�5��&m ^� ���;'<=��E[��u����!ʔ;BC��9Xў�0J���2��*۵#��ɲ�	��N�k�n�m��ys�,�)1�0�@�8�<��V��6%�����^j�%U6a�)��f];{2��%�# VFE{A�rx�,1b��4Mi|�g%�^z���G�&�,d�DF��|Y�Y�`� _jza�*·I``��Xj8�e�f�1�fh��J�L��E��)t����$�OJ� ���B)�u[d����0�6Μ$d������m 1P ΢j��IZ���	Z l�6�A����&`����'h ��Ҩ/ۢ<%�;P�j��� S�C �h2!耧TS�y�K/r����A ��L����)W�#����5R�Eu�߁�4)ゅ\�7�H�
�%\�T��- �h�0-]�1G{���R_,�
GkXYμ�p���Tu�-v��%�%�͹
���!� QZ*�2�+܃^TԐ����dxMM!x��у��YV�I"ЏZ;a��0J<��}�D���Hq���W�ꩃ���,cBR	A��W7z����:6�*D���|�#�Q�����Ү�ywK�43���`G��<�D��A�
�0>y����D���G�q2ş�r.�1`#G�| y ��Q~r���5�`"�I�&G���N7 f�,Mj4͓!��	S�׉��!a� O.�iGy�B��"��)֋��=!$ K&�I[m�K��A*B�)�
�0p�ހ ����hܦ4+�l�/��� 2�ʩO�ģ>�Tց,��KƦ
w�h!H2�L�d�RO�>gk��@�L�'$BI��KW(���sF��	r�z	�b�%I�pPt�Vx��a�!K�Gs $���G�j푷�I&���#��MڦerDB֛F{~!3䝖�J��$m$B/~�!dG�3A�]��K׸Q�b��E|p	cDݗ�Z�ͻ�b�;�%V� 
�	�^��d��O�1"��<k&���D�ĠXbL��E�?7p����a=HI�B�^�(n-�s#�9p59vC�&(����&�;=d��@c֑g0^a�J�������5�Ah���`j��*��u�'4x�q*�(7#����F�s�r�)��Fb�(��b˹~�$�g��_*l �����Xx8�y���SƬ���O�Xٻ��S7푞�y�`��pr�S�S0
A�I�휇Gel�:W�>vd4	�0�[$��M��/vf�;��H�])��Bhv�b��ƿq���n˰%� 剡ה%��h3���0�"<��bC�!�����+H`�j㨅@w��c�(%� �m�9���
q��<i�0X���KQ�l ׍�a�"1� E�i�ϻ لh�`'Q|����@����'��ؠ��Ԝ"�$�TV�mC�v�i0��`͟�r�[<u���g�-h^"�	�#�R�;��	y�P؂ƅ�2�xY�>p���׮D/mT6�aQ�ʖ\��	7�h=�V+�|�(�G��s�6y8�L�o�P�� @rb�h�
r>9��x�,@�Gr�4a�,W=x�.��M���L��D��פ�;t���_&=!�,saI�xE*Հ'�jܓ#�`������'c�R2��$H���G7N!:e�@-!$"z�D�4nH��"%d�z�bC�!M��a���I/.MQr��^H�s�Q? $�
��V�{^ѰE @�9���<�u���=��{�"��Lf�ڀgUX����+�2n8f�����3=Ըr��8{�<�#W��LA 6?Ҽr�X8y� �6��L# ��*3Ǟ��ós@D���%ZF ��V��P����/ԤR�7$}��Ձ9"$�࣒���|@;�O�����ޝ\X�$9t
�v�]�AHԐ���%�MD��lz���?��*__�0$�$|�u������$��=H��+KN�5�H��h�.J�y��$�=����k��I���ԟ䝘e']�[>}�$�����e��� �+�YiҶ�O�J�`&�^���5�N��@��5Q6��<�`��R>�0�e�M�(�C2c2�bl�d�A�T�I�T	Ҹ&4��-�|L��� R�U�$ɒ�$6��1#�F�O"��D��$3�����x6�:K��!�0f`�9��س ��<�1Z��U�&#Ek�q���t,#�����ܹ�"�τ>�4�Ю�p�"l��
/[�l����	�fC'�Õ�ֵ�2�O�?�Pqti�	[@��� 7HU�e9�ç<	n� �.I��E@�VI"u ÕV��q@��k[��;;�Y�D�N��19�兆cA���ާd\�4+Y'QJDV��%���.`O�la���yW�^��0�0t�Z%Qe�H�S�D�D��	)!m��@��yz�Ƌ6=xH�yt��DfJ48pF�iD�ސm����M�J�bD�GA�<��$#�F]88�\��/G�y*<�iI06l����I�!q��4�����I���.yv,�{A,1�-�!hQ�4$_v`�wd������X��pX��>!����"�ɏRmh�d+N	+\�5��ɉ)Œ���F[�'7��5��զ1�RK	�-̆ �e�ϷQ��b4��H޸1�,��\�`3en�lyҠ���xi��M�8��Hcc���i,C��h�|>^=�3��b�Q�(�r$�>�a��#Ղ:a�3� 2��O�l��|CGԬPt�,9��=іKN7u�F�����>�Q?�dڳ#�TԀ#�W�����A�k�����p �� D~
�Uç�`�vo�/�@�p�:J�T��O|m8$��K�Yr�B�O�'�^���ʁ$I�F� ��@�R%�+���ly�B� T@�H�.8��D;��M����( ̴Y�Ӈ]�����:������L���fg�&Iq�y`�
������ɳ"����em�/�<�#�K	05���ֵ �4���y�*�\+2/�.Q�2��Kۡ�y�-�{2\�1�']��E.ʆ�y2�ٝ)%�%���!��-�e���y�
	��KTn�(,����уԡ�y"�r��Ԛ���|�y���y��N�"	╌�XQxd�����y�b̓. R͋���E��x����y2g�4S��쐤7<c(�ho�?�y��H�~!���%�2Mc������yҥ�C�t(�f+I�3���[�A�#�yBG�<V���3��@'��MC�`	(�y��;�pc�Eف*�Qy��X��y�,L5њl13��$V
�P�@� �y�D�~���bv�ѡ�JU8dԾ�y����lX�A	r�^)!b��ybKYRh�WD2cY�!�����y��SU��!��X�.h�u��y��,Z��y�
D�]0 ����J�y�!��t�TWvt�HU���y⋏�';TEz1�N����d ��y�� 6H���)Q�1v�81H2�y�,���U
s#ϡ��k�"��yb��b��a�teU�c�<y���L��y���aDm@���)+�r�ib �y"��0�� ��AB(U�؈!�˻�y�%IDӠ���\�ĀJ�M�'�y���j��՚�D9@ CiU3�yR���Tp°�@)���Q�%���y��,����7�(��w����yr�ժ+� p���Q�6l �y��]iڙ��C�I0pH�DB��y��-Y�����@�Ii�g�2�y�+��@ҦL	A�4�s�iҫ�y��?1d�l�5I�)�p�($�̓�y2��]�J%xDgI�$��a�휝�y���^qz�&L�I�|�ڃ�
"�yB[��Xe:���M��u:�LV��yW�A*��t�jQ MpP��y��c��d�W��:����G�ȍ�y2nߙ1�2�A�J
E������y��q3�%�5��Wav�� c�'�yb��?I	� ׏L2E��YSlC.�y�&� =|�B+J4:�ĉ�EO�	�yb�s�Μ��jپyT������y�+
n'��x��׆h�����KB��y�Ip�JFÅcC�-!�����y2��6`����	�]�&���lЊ�p?��J�/|ܔQg"!�X6�գC9�!�A�	���x�7v+A�kH�O�H��ckX�hOf�0���G��
��3��*?���� 2@�avƍ�?jB�I�X��,�t��c3�,`vH�!dH6M�d�d-�!̆��1질���7`a�d��-O-��`2̎��yB.�D�����*����6�0�䐜^�V���ρ�J�*p���hO��"�� ^�	J!dZ"A�n(�G�'�e��$F���cTg�\m�Y��'٦b���zg��BrZ����'#B�!�h �
1"�a�p�R������
p0H��PE�5.�e���P�gN���s��������"O� �ꗭJ��0s�_�`�p��q���n��4�߈5��)@��9;N�O(���7 ��|ΓTd�pÈW&&Jp�Y[����XY��Q!�@�����6�<陖*�m�X4Y�MT�O�f�+S��o��Y�&���@�>�t�NFy����Z�@AcN�'�tdK">���wLs�@��q�F%Uz�P	� �%���	�	~� �B��5�L�P�B_��b��G�q�	y���..�N�*�n�~�I Gߑ4R�ҒlD /�4�&�� |�=c�D,*�D6]?��� ~�)�&jJ2RHR��G�W;D��ɨ(�N-QB��_��S�Ov�1�`'�I������B���wGX~d��,���|�!D�Q;���k֥fb���w��h�����,��`�N"P��i2F�xW��آP����IXh	�I9J|n&`U�9跥	�)�Q�#ںi, ��ÂC��Y�7CԵ>Ǥ��& $*h$��'y4NM�c�d�R�� �VꂦB�*E;�H�22izP��� pD��4�����'4Te��_�l"��cƦL�)�CJ�,*gaG3KNI����.���A �qp8�Ġ�()<(�'��Y��̓�W������`��P�.	%ޏ�^��Ϟ=T���S�JU���S	����U���R�O^���ε~λ Vf#n��'�^(6EޝO���ϓr㮩Q��� eZ���t	�8���Mh, ��'IT���c�V��0iM |�6���+gd��9�)ū
��0��h�3<fޜJfz>��`�M"y�,,�C�M�fd����E�KM��Xf�wF��1�U�������yb��z�p$8�a &99�R�$�� T-m�5�T�YzSj��oJ�jzb�s4�=��E�g�VڦI�r-��v� 9z�U�
���rS�^�(���xǸiM��
�!_�]�X���g�RQ���O0`�~�b�M'��4bZ���jY�2�
 ��*W�e�'_��Mh�IA@�&=r*F.�� #+�	gRa��R�"�2Q!d���1�zA�`f�A�(C��Ӕ@"�7햮����xh�H�X(b|ځ�� w�F�JG�W��Y�U��$�X7)�O?牰S#�e��Q�+��E���R��X#"]�>O��R�5x�.�Q`I�?a����/��m����R��1*�tz�§8N�8�K����	'v%$\�!����(�N�q�I����`.Ȳ/
�԰tj	� �b-�gRDZ �X6�ˍL�� "���_w(�	eQ`I�����IbyfG>��R���"D��u�,\���G8�X!�T�X��':�L:���9^���� ��)B�;$c	'^��5�'B������
�92-�2	�/!�t\b$��9k��"^F��DH7t�LY�	+#ŦA�u�i�AA�J� �Cܫ!¶i��f��[�Y� D�7؁R�웆Yo��5�H�9�X���b�/ԕ�� ��	I���UY)5ʒ���	p���O?����.%
�Ж���D�Va�W��H�^��b��i���A��U}=�i�d;����A�LU��^�L��$PX��L)c�؉8���+����r��	r�F���OoWp��=����/�ܱjd���0�L��1���o?d���#:s���yC�՟(^��6�GN7ʍc�o�5�Xc��s�Y�4�^����r P�aoZ�a�Q+4��7=�qO�
D[y!d�[QJO0}� 8��ۣO�ŹW�V Y�E1��ވ�PS�V�?P(�u��rZ�OrY�g�ܖ��>�(��(=�v8h�ۼW�})偓 �&��3*� 0`��+�e�T.�h�+ë:�n(����"�1��J������VŔ�cZu8�"O����m�H���Y�{UM��;�hq��� �]����Eц%�1�זn�T�%��}XaH�'4����낡
���S�3&��I��:��L�g��.ڼ���.ۦ??l��B-p�h=��j��KD�U�C�(X&��:7�W��0�����:3v#>i4�V$܄�7�W�v�J�Z!DM^�v�B�b�d̜C9ze�PI�in!��ŭE��!��צK>Y#3-�/+�̀��ۤm}��� �0�t��
�w�����?��ȠfS�<���8��[3�N4�p�I�c"	��H��s��=�A)ģ6���'Ez[�w��퓃�G�nl���ɒ�mmZ)��'�x�i��C�8ؘ���� 1VZ)Y �Va"�#��K� 8b�E���|�Q��>	´�N�2QJ	��w�ذAeL&1�"� 'O?K�
����'�h�+瞦`
��GfM+0�P[(Y�D��&@��W�&=�5 �i�O�MR$�Z�w��D��Ђ0�T"=�.7��s,ɤ(�f����T̓)�l��S!�����>˄x�W:�dI�O-M
��RAà{x!�q%ې�D@�t`,:R��I"U�Ia�K�)�$��3>P	�"L��a���M��UYsT�'�́$�A>��D�ٕ67L1��I ��q�a��I��yo�=B��2���@�2��'��E�y~�W�By�~�	bLW�,������=p$,擽)���y ��&Қx�A-[����* .Lk�	�Dg ܢ�� �)���9�ჶ#ۊd �fA/^�܋ڴzb����KT?Q��E*w�d4��3Ut��w�
LP�R���2x��(ke����b�Ó�̝�aL�<3�Rm��d��MWD}A6���=:l�9���<B�U��e�g��3�ǟ%{�L�C�5�(O�%ce�Ň_�
Ac��޺~l�y&�]3TZ|�*P5e_���@�gp�1CE�E�]�AF%�9xr��'#H�8b		f�,}��΁�D�L�Y�̕�&���H&��g�'�.i҃΀�@�\� ̔�"�� �Jq��T�snǖs� �pk߹ ��@y�	$<�|xaw����0)˔�u�iκ_�q�@�,�\r�c�)]�ݑ&ǝ<d�D=*p�u��;x�z�:Ġ�'o$f� ��J�>����L�B^L��Bǋ�F�So�O{>��Gl���iZ�'��ɴz�
�� �'g�H�3�ϚNx8��gL <�qbv�'�n��t�_�%G��V΂Jh�e���Ik�e�DЉh���tFA�P�|��$�4&O����In�Z]c�4�!s"��1􇙬K�"�b���1 Yc! 3Dx�٢ĈB��%���`��Y���	%��3q��D�ςDF�Q����U�
;W���}3�0����iՌ�1t��6ƞ��8���V U*@`CK��2����ЮεY�j	H�B���hO��zT���9�(�ӣ�W�\L��$'�!!� ��W��^���B��Iq�(Z���~X�%M\���l�$m9���Կ���F.��ql.e��Q*'��a�B�œi��p��[� ��O�-�B�H5%L��!5d�	Wr� ����+.�HS�dVI,���F_�E&�w)�
���ҵB�Yi��C$Z�"!���^�\t9�K�=~�&l�U��2�'� ��V�Bt <[F/J<?��1o�k�8$x�g�0`���S���2��Bx 3�o>=�)��;� ��h$n���v�r��(op����E�"� ��*RF.��&�'��M�3�
,������c!�<8�`�غY��dP��P=�0H�c�R&���%H�M����wPt�X(%�6qB�

&��ə�śEx�xZD)�"����E��G;��*c����� C�Ni`q.�3Ҵ�1j��<`x��І�]0� ͸����IHM0��ۆ6¬�t8[�ި��� Mr�\8�g�B�I Lq�H��J�L�^���L�
��T�	� x�$�$��X�T��/ߌS}�����i�t�u�i��ًaj���?���m����W�?��0�y�O�-+`��8#�6w��R�����1+�t7�x�"m�+��t���?������+������#ۆ�!���t�K"d@�7��d� X�vÁ�
:0
ד2Zx�k�K4\pX��.��Jψ�2���V�X���F*��\��l�,3Y~�s%A˵Xb`��i������`�M����{��R!^���I9g�(�eA����Q�E�Q������:Y}��ɛ�]h�8���-�6�ϗB�6uc��-���;��Cu��t1���(��Q�]$���
�j��]�BM����HO��I�_ldi����	��B$��Ic$�Sm��k�f�	ov���O�5E@��#��;Gm��V�J ��QC4d蟚�{�O��6lB7"+p�tͅ6�EH��'�"|3�BǰMF�q߂7��� 5Ӂ�.B �#�i ���֟{��d�@N�/B<3��\;b陗(���rd�0#�G}RL���A&O�'�h�
�K������.`��c��$��Jb��8����c�=!�D�!�P�#n`���/�PQ�g��n�nXb  Jt��#镤#�����څX�jP�'Jz�P��B�Oc��Y�܊Q��s�d�D�4��FI �ܕh�J�>"F`�H�+�Ki�u�X (�"Fw��r+[3B��p��-�O
�b`I42a�ۜ)h� 
&nU�Y��02c���)t�ٱ�O g�H�E�K�5v�����/g�Z��3X�� ���,~�錹��t�6O�	/��I��%�(O�PR�	����T���)���-M$5�Ȍ+��NE ���5P���ֆO�!Ll��ՆT0b�eM�ka�SB$�ў�S�F�_4�tI�PT*ܐ�'E0�fx�e ��M̈́�@��Î\rF�Q#lF^

�ĬV_>���47h��g��:�Z %R�X,xtPޞw�L��� ��>13H$��]z �R�:=�T����6��m:I�%�4��#�i��mq�����qB@h�81�t�f�ZԼ36#�e�2��q��B	n1𐁑]�R k��	��,��!О	N8�t,ův��Q�ݶ~�p�Q��D#O�V�j�f��m��Ζ�Z����s��E�lݴ{�j���|(�	�&�h��zA�>Cu"<�WN�'�H�k�1j%��s%b z��4������$ ɍ8G��э7�*V�{p4�Df�!D��fk�e�WG S�'V���$/ϰ("�y���	Lȭ�>9:雃��yS�,8�쇀�u�C��==Ƭ��W�K`�~p��;5 �	�1)rzIcbD	���Cql��%��b��tx�4��?b�|a��(!�"���A�5b��sV�W��Jp�®.rHc��=`�`a�𨄄&�0Ђbaf��q/&ed���ul��#�����'1�O>)d��8�h�跉[bCV�8��Y��.Uh�m]KD�1A��X����9<��T2l���+W$H����)i��;v�܁i��CFǐk^���J'�!�|���݃m��{&'�oV��CRJF;`��Q�0�B�c9BɚaJ�4��x��Nė(>`6.��d���I�Lp����Z)}Ӥ@�(ʖ�DtO���BѶOz\�ҌI�]N�|y���_#Y���ǵ,Â4�ΔrB ���хf���lX�T��&�~ڸHp�ۿ��O$X�E��ēd󀉻�͙G�60���JY�4	�ٺ�¸1���B[0��d�ɓb���۱���D�8�R�I^�ͻe��-��އe�zYC�ÃHa��Oh����G��ư��\ �i7�*k�fqђ�J'hZIr�i�/p" j5m֔-��hR�U�E���R��B�U�hQ�2�˥bL}	I-����p���\���b �J��!kpb:�C�L��(�-5ĉ�Iٸd$��QT`M,�|��c�z�n5�A�߽s�J���%�e��(����k�.E�Db*�xk��HO2�kT��l�̛��^�M�̍J�`D�hTv ɰ�H=+I�U�.ܪ \���%�
f���2�I�ƙr1 �-nYl�0>R~�(@�m��ii�%@A*¹_7��;�u��hY��;��L�BTr���-_t��(V<X�l���K�"嚅G�g�F�ە�W=U=.��͒�Y{��x��E�Z�f�u�N�8�]���*���rv\����A�W}&�� ��c���2���c���M#�4C���OK4�k�-Q�� ��� @M�7�C&}�i�� >s�j��~�&H�Wm���[��"EF�Ї�B�~�r��6/���7ΔO�P���H�[]9Y��I(|�D�t��7ls���O.����!�K�X���H,[[
%l��_��`�@� E�.5��	�;[ˎ9ـ�ތ=4�S�+�����,�ZqO��JfL�\��(�	�︝*!lK5K�H\�������N�ήh�T�&Z��(��欉1,6M�Vd�E/Q0fh�pvNV&��@E��fM�R��c��4qu�Ǎa����
^�A��� 7ip�X��Y�� R���y2T���%!RE�]y`  `v�$ȗ#�	9X�2e�ؖ	�
g}8^���%#VM�AI��x(��0S���`��Q@}b� z
�Z�G�	2�0�B���LT؇A(asJ�Ӗ#6$B4�\�U�E#�iU&1*ͩ�@�"C�} ����d�^y*���O88rD@��V��Q&I�$48푤��e:&�ՋZ���0��#���2��$g:T���O�g�LuP�*��-�^`��~�vk�JBQ�hɤ"�3��Ă�!��Ay�Rr(A5?�������8�lX4�@�"�
|�cN9'�ز�LF̓'�̊s���Z�z�,����	v��d�8����.T�*DX@)�d�����B��D�z�l���fJH�g�>��8 �|4�CLG��\Z��$t��k�o��8̚�ht���d�t����(L�,�gFX�y8�{7����
�t/�2H�6yaq��9p9���I�>C�8=�4Ӗ~��KG����{�orS�y����1r�p��с:�F�9�xm�	���ny�h���f\!OV���!�;�^�A��|j�)�&���Y𜳒mC��8Pk��8}L��%!�;.�$���B4�"��O�l� 
E���λ.���󱃀�u��� �G	�ؘ�2h88����*
h�������~���)�.���`�	�\����hK�X{��Q菚�¥/��u������[����p�� �O�9� ����9R q���d��-���� �L�3e �7߼&K�nB��7�>�ƭ��[�i+��R�)��U� p����e"%":U����!MP��8�R��"�i#>E)��О$��8�#mK
y�� V&p�%1���=ռ���Y��a_M���MK�z�� @o֟��IF#aɀ��t�jU�bb�K}Q�(R���~< 7oV�,$���s,�6��&�,kc�E�?1vY1���l��M{��B17eZ,�c7��0"�F '8���W�� e���<��@��v��xĀH(a�t�'��lh�!�&��Ր�JӉ f�	�[�8�U��U�J 8��d��#�
5:�ĪI�j��ą�>[p`3*O$1�!�S�T)�|%>c����@�ܪ�S���>��x0�&�Ob� �dBT��D"S�V�&�ñC�a<�S��ΰ?	�X0�Ҥ�E	IV��� ��
|8�C�n��$1O���Ӯ�5;�(�;�F@��(s"O8�����|Xn�D�Z�46���"O^��V�Z�$��<�$X�n�1%"O2 V"��w�"
礖;'��j�"O�Q����69�~�q��	� $"O�Jƪ\A�@X�^�4��R�"O�u-����9k�ӆ>�rb"O��[ �	={�����{�"��"O ���{$t�7��-'�pR�"Ox��c�פS�zx[!F�#>�p�"OT����-^P��K�Gې5�l�"O:�:�]9o���s�S�c)�1	"OX"�ꑌ��i�EPC8"O8BE�6~|4#��~�)K�"O�h�3j�[�d����M��RG"O�qK1g]�Q`�(�W	L�XV"Oeh#��0Rnh�QP�4& ���"O����G�^P��RF�F�hL�s"O�h F�J��U�%)#$5Ɣa"O�Y�`�M'��+�;6���"O��c@l� 8!vƎ�d�$\R�"O���
M`\:h$�<�ܕ��"O2�����#d��q�b�9b���"Ohib�`�;�֍�����Vm(���"O�-a��yGv��!�$J��Ї"Od��$I�'fؔ��1f,<V�%�?O*@v�l����%�{�z���cx�u�O:^?���K�U/��!���Q&����#�?1.��P�B>�zM)0N V��u�f�_�C=������B� h��oW��3ܴ4������u�`�c�2!T Re,�5�<��A�I&8G�-ڴ@��A������w��Tz� E�'��B�
��غ�l%
P@l�!qBjP��r�l��)��"H$E��B�0W`ʼo�p�yش ���F�hy�'R��N|��mv>���(-cJ���#�A���7���"�T�<�i��yR���IN/��qWb�o�%��.��� �R j����2\����O#(�ू�� ����O7%�\�+#2O�� �����&u[��U<2"�>�݂\�D�)�*�)Pt`�q���Sغ,�uk��Д�eGL�O�O��qQ��i�I+�Mм~E�;���'*����ݴi��Ǐ�4`����T��<E��lA���)��Q7`���RD�R� ဟ��#ÅȊF�a���J�M2U��!��Q�dy�	��v*�	��t�"��S�m�a��(�G��f�@�4?�49�����~%����a����y�iF�"}��*F0�hr5�*1�lБR-;-o�j�˦W�۴:S�i�''8=ꆇO�V������A0Zz���#nyZu��4^6ܘ#+�0|��LY�q~D�#�j�	g�٘	[�o͖�ߴx�Ti�I�R e#L?��f"��?�eI��N	�_����	�&TzDY���a���5L]����O�&X�HR�D��͙��_� ���K¥�&�@TX��c@D3����d�
���Z�&��P& �<�(P��H2�'!L���i_|<0�,O1l��$j��4:?�	b�8�AĮM�iu|��i�tl�\� jF";�60r�<-��d ��HC�g��)� x��*�]���HCU�P����-QR�����I~
�'B�M;�iͰ+���/A�C�)t@�4���'�0-8
�'z�d�j���>~�c����,��p��x��]$3}�lKDgZKR��i���eI�.��C)_�{�؅ȓ$T��N�rB��ڠ���1%ƽ��S�? �xpY�Z��qk0@�:B A�"O��&l�-�DL� @�fP��AU"O�ja�I,O��qk�jZ�wMre�V"O��u,D�����
��J�R"O��[�b�/����uOҊ/R���"O�L��A�t� ��aO@;<Z��Q"O��SSO��
ԔX㮗�D���"O(V�O�v=jA)8�l��!J~�<��Ƹ۲\�1�[m��'�w�<�Dm�Bd�"�ҕD`�����N�<�a��G�*i뀥��"��x�BVJ�<ic�DN[���/×N
Z��E�<)p$�c�^����)B���ŋ~�<����S��HK��91�N�>�C�I�~�Mr��	tj�R_�]��C��5K��t���Z.5��ܰ�aޢ>��C�I>x�&�����Pς����P-'.�C��O�H�@�
�tF%��g�#[تC�c�,P] u���"��f��C�I�u��tK�$�9�&d]�Q=�C�I��jH����0@�Q{�� îB�I�CM=r�iP
P��x���ǤmӰB��-�bc�L�B`R��O:ZO�B�ə8��0���k�X��	���B��	bq����,~����e*L
�C�[gf�q���_oh�P��b�C�;fi��Ǯy!h= �F̀']C�	����*R�TI�0Y�E�J�/=C�ɑ!uB����	����V`@C�	���p�7dҎi�H��r ҡ�"C�I��RqhdkH|�f��U@��e� C䉪-��	a@�s����j޷.�C䉦~v�E1eeدAl�3'�>,��C�b���qE�u�Eb��ܔ8��C�I>$ �3���7�ԑC�ڼ	�B�ɹ!HX�5c���:Ø�<�tB�S���L "`|%���T�VdB�	+{��YǬ�y���rKҋ)�2B�	"L���ӕ��EӜr�,͐e`(B�ɮ/�T41@�S��<��
�=a�B�	�S�f��F��rQ���A ��B�ɰ]e����^H����C� :P�C䉅a|�;�)X�n������\x��C�I�0-��xs��	^zn�S���,�hC�I�r�b)#�c�%4T|a䙅b<C�ɬ-�0��lQ.���"6&
�Mt
C�	�ε��D�w�����ɋj��B�`��hѫ��r�  	՛ue�B�I,�j��ֈ"D�b�C2AEc��B� �n%���Һ�D̺��aF�B��/��l�׭F�<�(X�4AbyB�	.)N��[�m�0O$` �f�T�|�C��{��H�E��k�4$����-OrC�	�K4���ׂ@� �J�Q�)z�B䉮��ю�>�v\Z��$l�B䉜J;~`i��BtlH���Y]�B�I�	���	�&B��>�r� '%�C�	R��0��m��p�/#�C�4|΁y��	��@ZJ&@zB��roj�H�`ѨZDҙ ���'��B�ɴb��,��C���L�f�
_TVB�ɖd�^lwɄ[�$E�
�'�C�� glа�RK�-7>�pD��#˒C�����f�
!���b��\B�)� *�s�h�8��I	�.�2� "Oh�"M�5���G���s�-�"O,��3oQ2X��+�Ο�&@�t��"O�
q ���l��>T쀹�"Ohm� Κ>{��}*�m�ETz�Rc"O��{���g��@���0:��2"O�+P�9G�R�XT�D�w/4I�v"O�m*FK��E0!�(�.x���"O�`YQ9���I���#f��Ej`"O�u
�)�;�`E�E�Ky�A#"O����-h����e�'x�Q��"O
da��Vf�k��ȴH;�U�d"O�A�l�mIy��D��
�FY "O�pQ�I��.��0����2�jqP�"O\�����Bm�e<�t��"O����k���9@�F	 o��2W"O�D�T�@bE��M���"O�R�l�tg~�12K�'&��Y��"O�آ�+�{�|\�e����r"OJ��!k%n���Q\&T�#"OHـҤG�~��@��O�Q&�	�'"O���3�\�+s���(�0e���E"O&-ceG�,R	i硎/D��y�C"O&�	��;��PgA�XI�R"Ot%���]�~5���fS�Re�qc�"O���TH��Zr��2Ƈ�]2��q"Oh���2swT��p�U$3!
�AP"O��BD�C���W��C��r"O��Ȍ�6��"��g�l�"O\=;���#+�Xk��q�L`k%"Ol��� HTT�e���_;��a`"O����c?ܶ�E�I
ܝ�w"O��	�K0S .\[�~����1"O�!��![�
�x�a�M9v���"O�]Q�F�(�`�yK��p	�(�"OV����5L�P�)9#�҅��"O"�y��N/�e3��Ƌn��H�d"O�t��H�8|��٩��9q���"O���ë��Y�=Yr-�ynI�"O�����U,�	Ь+3bD)�"OpT���;
�*�A@kؓDL~�#"O��3Ӫ@������\:6<�� "O���w��m�ncAӧ{x�Yb"O�\;�g^7��k7kZ*:��"O����*�,
���!��+�\��"O8��V:G�6yk���>O��E(�"O� ��(1+j��ѧζ
����"O�1(�U.it �$P�hd9+�"O"9����z��M�r�ƺD���V"O�`&�ڟ@x���_��$��f"OƔ��$s�q���%�2@��"O��
&M�9�6D��M�<W����"O8ek� �2Y\A`1,E*���:�"O��I��ȱ�P�ԁܗE�&�"�"O�E0�C�w��̺��M�K�
 A�"O)(�dS>:��A�a �j�{"Oҽs6�Q/ܐ��'�2�� ("O0E@e�
��l�$@�k�,a*�"O�Z	E 鈁��;~M~#Fgi�<i�ϙju̽	#o��B_h�<��� Nr����L|��� Wg�<��"��D���1�E�M����e�<w�
�D9L�1�C�r��X16'b�<��)�h�>��6,��#|x`���Mr�<� ~0Y���W!v%(�aB!S�S�"O�b�@VF� x"�/׽aD���"O(�k4��$4P���A�5�c"O�:�iW:8E����:I����"O�e3�N�.B#��Xtߋ:� aSB"O^�Xv�R"4f���"K�uE�8��"OD�Ђn��m}�0�7K�>:,*"ORdKG�i��[e�N�;Y�ʡ"O.r��.A�\�AO�Fd� "OZ��E��_��m��˻h4�]i�"O.�bǫڻO��2�O�0M1N9�"OV�e�Z�t��.�3v��$�5"O��BF��N�.��L�O�P"O��	O�h3�# LM�?��	H4"OF��s�"`��Z�ͻQ�F��D"O�D`R��+_��=�cC�7@��`�u"O<m��k�P��H���0��"Ox�{D��.U�̕������@"Ol])2�,"3$Ěg�T�b��"O�A��DE�dd�C�M�>S��:t"O,e�'�c�d��D�/Q��Rb"O�	j�E�t�@��f�d_&�Kb"O�i8��B�p�~�f_�zB�q�G"O���H�f��b�B��.U8E"O�A�!J�^��X��4nq����"Otx��-��.�t8(��]0Dp�Q"O���Fɲ���"5�i(-9d"O�I�h�5_�(���<s��"O(��h���
�*�&<��Xp"O ph� �((��d+`�52�e� "O�kD��#�VQsdp��aZ��!��	$z��b�Z�1�6��@�C�!�ą�it��bU�����Pr��=�!�d[�*��$��N�w)��C��/<�!��؅Z������Y+2�3�o�r�!�d�	��I�`̛�$%4l�Xh��"O����+JSp�x��	OԔY�"Ohe!�e 
*Ё�� 5V���u"O��@A��;���8�Aă(��8��"O��.���}����A�Z$s"O\A��Bǀ |��NK�NIr�{�"O:�ì@��p�y�'�_D6Bw"O��B��\F�.�aχ$	��ؗ"OX@h��ڃSu`�B�����v%�C"O�`�ʅ>`�@���e�^�i�"O�ݫ�Ǐ3��QФ�1~�4P"Oȑ�hϬ1�T�caC75xR��S"O�����׎8�^9[&K8!p$�8�"O,0
 ��"�+ �C����@��y"kP�l���J��9lM"e��yr� +)B��d�6 �ʭ�QD��yB���Rh�л!�Q6}2`91&n֫�y2o��+h��	�p�T���c��yD8&h���A��b�f��%�&�yb�V�H'�H9��7(̜92́��y2��rN��t��	�B��c�"�y�D�c���p�ފ,qԽB1���y�.�5� �D�ߜ!*ѡ�$�y"Ə�/RT��s�Ս
��@�]��y�G.Gݜ5�Ɔ������y���w˲�ك�K-1zxa�@,��y��=y�6�9w�d��M0�y�݁*{�h+&#��� ��N��ybC�&���S���s' �Gs�C�)� �m��¨]����M/i�p5��"O$E�
�	s���t�~��R"O<l��   ��   �  ?  �  �  �*  �6  �B  �N  �Z  �f  r  �}  �  $�  Ϙ  �  2�  |�  ²  �  I�  ��  �  ��   �  h�  ��  4�  ��  ��  =�  } - � � =( �7 �> M �\ �d �j /q pw �x  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&"O@%����-Zw*�`C�#���"O01#�m�{�0Rda�#�"O� �	�e���Z� TX�؉B'"Ot�[��*Y�~����4[�h�1P"O��@�K�4Xպs-َbF�ģ"O�-��H�l붼�t,�0F(���!"O�����G>�`R+�0Zy�6"O�eXu럋>���i��wf�%�Q"O����d"�9c*��h>�`;�"O.T���T�`~fM����q)X�h�"O,�YD�#H��k\��t��"O�ɢ%b��/�P5P!m��hb5�%"O���0�φO�Z��k͡1���k�"O�``I�4g$�1шىK�yR�"O6|�D(
46�jf��\��A8�"O�ukg��<Pz�Aa`�#�h��"O@PQ%ƃ^R��p� �p���"O�xjd�j���a�ݾ
L�t�V"O�(Z�[�3p�����CE���r"O.��E�	Sn���
W)^?n��D"O����)�e=!쎷E+���"O����!,\�| �-Z�6xtb�"O ��.X������.��K
�!	�"O���*� �|�S��N ��irU"Ofl0��h=��@�D 5K��� �"O�<kqO�D�
�AۣFj�@2�"O�2���w��"��QL�.a��"ORp�2H��X��a�Ԇ	���A"O�u3o�A�dr�R3�Vy�!"Oؔ�sO]�:��@��z���U"O4�k�a].����E�j	�p"O�1`�	
 ��x1�F�C���XP"O�𪰇O�<�D�8��$m�p��"O����Ȃ0z�L	���K�(��	ˆ"O0���<�*��4bڥ�V<(�"O�m��OE SX�7$�f�31"O�x��R�8�k�]8�U��"O���/�4Q����TdN�lЌ�Qc"Ov���j�3����cč�Dm��"O��ۗ@^�?1�H��ի:�晀0"O8��M�T#Z�h����B0p�r�"OR|q5��*?��ATn�(Ta+�"O��zc��n��w-ݏ���v"O|��u�&�j���?$��q"O~4���7,��)q�V3h���s"OJ�r3M�i�[��V�ZY�u��"Oҍ�dD 0��ER�<hbv�A%"Ohx�  >,jȁ��"){�M{�"O�(�b�Aq�tQR����]���
�')\5fŋQk���M�r���b�'�~-2�+��'4���Ůe9����'��1gOJ)'}.��a��^�F�'W�1�( a��IJ�s�ź�'"D8"�J�,�^P�"�ب@	�'�ʀ�F�9Q�  �����X��'�p�Z�-3�����5{?���'���-c9@yq�U�i���s�'�5��A�g*f�)A��$u���*�'В}�%�G(}b`�e!Эe���Q�'�Xi���2���@�T�^x�a
�'�^dk�D��h�J�Q��B�d�H��	�'o���� ̗Q�l��@R�]� ���'ƶ�3�ʑ�����F`[�J���'��� !L�,Dl�F��6}� ���'�8#R�F!*(@��5CA	z�����'Ϙ�q� ]�h�P�g�fMT���� �ኃ)4�J&ךF�0�x�"O�\��]-|�9���G��0��"OTE�2cQ~B(�b��)��"OD)@p�1�uKЧ{�a� "O؈+q��6$\�s
�<4�d5h��'��I����I���˟��	���ɮvZ�Bȅ*F��S��JR�T����(�I���ğ��I������|�I�RƄQ�h�,1QǙ,�M�	ߟ��ݟ|�	�����ҟ��	ԟd���wMBI���ƙ_�4��ƛ1<�-�I����ǟ��	� �IܟH�Iٟ�� F*������\���XQ���l��H��؟�I�����՟��Iҟ��I�p�A	�$%
eq��kgH�d�	�������	ǟ|��ҟ����\X��X:̔hӎ�L�h�cŅ}����ϟ �I��@��̟��I����Iǟ�p!�B�U`�K߃[I�P�*���	ɟP�Iԟ�������IƟx�	� �p�H2gU����\D�d���g�П���ß�I���̟�����	ҟ��%,�`h2��M�7&<躅��Ο�I�X�����	��H������I̟< �H[��hw	Rɐ�����O���O��OT�D�O:���O
�$Dc�.@���*npja����&�j��OR���O��D�O�D�OF���O~�Ā�uC����Sq�bQ�ŁqI���'2�'���'�r�'#�bӘ�D�O�"��.��0
⩟7(9�YBCE�Jy��'��)�3?���iP�����o*�:#Х{�����F3���R�A�?��<��%@���`�?\c��� �J/@!r�Q��?���+�MK�O����J?!J'iX�ZSX�� �9\�*Y�2�/����\�'��>A("��1���yd�%H!ڵ�.��M�*R|̓��OJ�6=�F�ƣ�$A(̭���͝4�y�6m�Oj�d~��է�O/��տi��$N2&l��f��j�60d �f��Dg����A��=�'�?�0��SW�h��ȝ� ��u�Q�<9-O��Oz9m�&�.c�hr�HO/Ve����@0��%qCd�f�wj�I����I�<A�O��8�(��_�DK��[��� �	�����%� ��2�@ߟ��&�\�*�xElǞm�eR��qy�S�`�)��<�I�<T�9Â�ʄq�ƬX���<�дi0Tm��O�yn�G��|� _y|�� �<1KHq���<����?���L�����4��do>�q�� ^���b�n^d]��śy
��6�5�D�<�'�?����?���?�Ix�%��aA5o$e E �������0	c�T�I���$?�	�8���
#��dt��8�M���]��OԱo7�MCI>�'�R�����A�]-�^���l�8u�b�3���.�����H�Ĉ3ׯ��b�A����>i�Ρ<�t!�2(���4Z�F8iԯ�-�?	��?1��?ͧ���)0e�v��)��صt!F%�'�g�HzA"i��i�4��'���A&ed���d!| ����	�<�t)���>;Ġ!�%i���	.�4�G�0@�r֝�G���ON�I���w5��12�J�_D��{���$��'�r�'`��'�'n�����2b��q�I�y]�h`�@��<����?G�i|�:�O2lZz�Ii�Ȑ����a���˧i�
�%�`�ش2ݛ6�'mX A�i����O�HC�gP#AfR�IT���c�10��'_^%r��i�
<�'.6m�<q���?q���yr�ׂ!���1KR�Uy�0��M��?�����K�j�K!?1�����`Y\4��O�x�a�B�.S��'��n^��j��O������Cς�T%�ؚ6�F��,5�Eĝ(����g��f�h˓p�뮊�Kh�6�XMyR�wcn�a�c@	A�hvo��L�L� �'��'�����O��I�M[4H�/	�fT[�,l�\�ᓆÃ9�R��'rL7M/�I5��d����Ƈ�}�^����T"R$�hCj���M��	m�T�ݴ�y��'%��cu(��u�c�Vy2�$Vd ��M<x]�uKf��vW�6-�<���?����?���?a-�|'�	A��X�Ĕg�`�P��-0h���IП0$?��:�M�;.��p�Ҫi6���d��vPC1�'Z�v��O%�D�'Z��a�i��Ƿj��� g�/n���I���%6��P</q�킶�i7�<�'��7m�<q���?��,��s�|�t�M9xla�0��?���?����ąڦI�Ն|����ş�p�f�`J&Xj����Vq�a#UM��R=����M�&�i"�'ׂ�*D�ș�T,Եj�'�2�:J GL�&W�	��u�bТ�M#���O4�ȱm��S���z�h]�fᜉ���O����O���O`�}��^|D���?-(�\kf��8
$���	�����$�֦e�?ͻ]�TmRc� �Ȃ�څ$�8Rw����M#q�i��-�l���>Or�����9��hm�ӣ�]' ��R�sʲ�����
ͦ��'�R�'x��'l��'�pmC���G�6h��Ƒ���z�^��ش[k����?������<	&	��Z���-�"F�dؐ!ĝ3�����n�I��?E�S�@v�H38��	3�<G�)C��c�F0���zyR,4�%��4
��ʓ`h�fS��6f��x�(�,Zy0CdCʟT�	ğd�	��_y2�u���J��O�!����n�g6Af=�'@�O�AoZ@�<����g˛�li��Hk���+�=�坵?A)ʡ@G�0b�7M6?�(�$��)�1��'��� ���
�*G�Ԝl�zpA35O��d�O�$�O���O��?5H�(�3f$U�d��G����ß6�iY��r����1���DѦ�'�8٥�ѝ	e|q����e���m���Lϛ�t���/�>6M2?1�K
�Q�Ej��*)k�uk�,N5~V��@E�O䨒H>�(O&��O��d�O6Ѐ��K@�X�f�Bق����O�D�<�f�i��]I��'���'���_�ܸ�3,� ����+VM��Z�I��n����S�d#H�,NP� �.����*GM�*l>����bL/���X"^��S3��b�h�>�X���k�{1��kwj8J{<��I��d����<XC(�<Ac��'�?��'
d�[}(� � i�p�cL�l�0$�Ɨ�P�ܴ��'s8�\K�v�ԝ���FGN�3��I��)[<�H7�^��	S����!�'���f�N�?���[�p���Ҍ&��Ճ�%�0>��U�m���'�r�'���'���'l�ӂKk^��S�Z<?��I��۔`7�Dp�4W,p]��?����Z+��^��]L�n�IaE�G�ʅ�3�^YGBD�ܴ&-�f��O���|��'���b��M��'}��%Έe�����'[qf^� �'\�S��j�MS#�(�d�<9���?�� ̀31P�{�`EY� 0#�G�#�?���?q����$ʦA�bk�L�Iҟ<��i�;�����ʷ��aӍ�r��ch��%�M;2�i�d�$�>����@���Z�\n���G~2# �0��+5��O�8P��#5����.]���X��J�Њu�'2�'��'��>i��	?Ԑ�O�C���a�L��B�<��ɭ�M����W~Ho�|��]0�HJ�KsC�@�c.�-�牌�M�E�i��6��q��6-o�����?& ��O��:��U=K��p�CB�Y�W��m��'H�	��8������Ɵ���w̸<����9%.��3n�{?b����4`m���IΟx����M��y�i�'��1��c	P�F-ǞV>�?o�AzӾ���c��?���xL�H0�jK�+�H��� ���P�'��s�^��'�.pYB�䟸z��|b^�t���<\�}h��J����"�o��d�I͟X�����my��|�����O�$fg25*L!K���+`l8%��O�0o�j�����)�M��iK6-�3{x���}fN K��&^�$�Y��~Ӫ�	Ɵt�Di�e���+TyyR�O3���J��L'�J�)X�XC`��)�y��'f"�'�2�'���I@�Eh�YsGR�HbA���E�v� ���O<�DR⦙��r>��I��M�L>S�� ��!�9���򆒤3��'�|7��ڦ=���yb�m��<��5�p��7��E�~eɕ��9`L݀:k�$T������On�$�O �D���xP��;?���`f��I���$�O�˓S7�6�ё{���'n�[>��҄חa,��/K F�r�j/?�d\�DP�4fR��8�4�X�	Ā
�l�#,]�SKj�9�A�l���@I:r�J����n���h��ְ[��S?hҧ5��^�f&�p���f}�F��;���'�2�'����T��sߴ�f=p��I�>@S�W�B�ҩIS���?���a���LE}��b�f@ѧC̿廅l	�]�"pӅ�Ԧ5�ߴ��)3�4�y2�'n��Ȱ��?�R]�� '�T�Z��`p��{T��:A#j�l�'=��'��'p��'��/����DΟ~��bK"���9ڴP� ����?	����Oʀ6=�. j���L��(��ުK��u�w���][۴9ɉ�����5ش?�|��ݴ�yB��}ɬ�R� D1O�������y̊'4*J�Iq��'/�㟬�I�'!L\*�"�ʜB��/�8�	��L�	ڟ|�'�x7mċUd����O<�$��	�0+lpL %���\����O�%oږ�M���i��+t�=�FcH�>�d��n��/�dT��?����S�)���E8��d����Db݅���<ؾm�P�E3��(j��-Fv	���?9���?���?9�rE�i-B��?�;0��XXrh�+(��-ĢP��h�B�*����"�y�'y�'��ɂ�MG&P:g�P���iJ�\��.���R��m�&�i�p�oڧm�inX~2C��!6@��
lا����d���������|�T�`��͟������Iş<�̱W^����A5&5��dy2*o��a�!9O,�D�Ot���)����g*]zL�M�7�/��8�'��6mQ�m$�b>�1kT;/ք�Q��(@�!��$k��d6�ʓ3�
�b3,\��Y�Q�|�V�����������hkl��|����P������]y�`e�L�$O�O.M��O��Ů�����#ec�}!��O��o�t�3����M㣱i�ل{��pl�+lR�qc���s���4�im�I5�̉x��O�q�",�1���1�]�B�;t�Y�_^�Γ�?���?����?���O�����Z>dt0�RE��y��8��'
��'EV7-L%1f�i�O��l�S�	.>޼1�G�/����e��7;C��Γ������4�?!��ǎ�M��'����/Ů�Q�Q$D��+ � 7Af(a`o۟�B�|r_��Sџ���� ��#�� T��qa��B/
H���O���� �4n�	��H�O~����k��aY���� c�O���'�6M��u��ħ�*�LВ(���æ�A�\���@��B4?Ȝ(��.0F�H��'v�����0���|r(R6b��@!��ӪJ������ 4��''b�'���t]�tBܴ[�B��H��;¯�({x8ዔ�R��?Q�v��F�d	}�g����R	��u��=k�-*V<��sC�A���ܴ}}ꈣ�4�y�#�J�:�4M��?��18O�� ��#Q�T8OO��ǯٕ8#X\T�i,���'���'��'A��'�S�\ ��4-Ǧ��=�7��uPM�ش[�|��'I���\Ȧ�ݺ�\��@\�M��A�qO��%�V�Rٴ+ћ��O`��|"���b&J�M��'��B���I	
dj���B�Ԃ�'��	��#@�L*��|�S����Ο���L��`zP�ITg�mj ��Qd��h�Iҟ��IGy{�J@à3O0���O���U<�DP"�~r@�-��'������ѓشz�RY���b�"C����g'_�r�.�RՅ#?	���Xz|1�����'\Z����?�(�VxΑJ0����,ɷ o!���?��?���h�v��.`�\�g@!=�T��c���z��æ��vA2?���iJ�O�N��M���P�M�;6�~%#��\�=��̦	j�4Zʛ���$қ����RF �5Zk���߳3pv�x��&H��hR�d�{:�'�d�'���'��':b�'�����b޴ �:��BQ��n	0Z��#�4�h���?)�����<1�hU8.l�yXc�[���çU�0��ɂ�M�ֹik���1ҧj�r�)_s�pL�W@��kMZmBp�k��58.O�5i���8�?���<�D�<a�A5'2���I���L*�����?A��?���?ͧ��E��1��aq�t���h��h�)$ZG�С�n��޴��'!��8��Fi~Ӝ����D9�wf�w�4��[�5g^Z7	�&�j�J�)!����;wf1�)��諱nSPO�@q4�G' zl8:�5O4���O��O����O��?Z ň�Lƞ��hQ�G�I[�-k���̱۟�4{׼a�'��6�/�$؄c�u �$�;ṯ�U(�kM��O�mZ��Mϧ#��P�4��DلDfx���La���gf.y�(��6/śƭ�R��Fy��'���'b�V?mT��f�<-'6�p�%m��'Y�I�M�����<���?�*��hx�g��>d��43]2"W����Orn�9�M�L>ͧ����0c2ْ�bؐ^0I�4�'h�3�/I#G-���)O��I�"��6�o�	�]�J݋@וa����`BD8U�@��I�,�	ğl�)�Jy�Kt�){�M=�ʸ�@�C@�}�v$F��	7�M���<�ܴ B�S�[<��1�f�+���Q�iR�lY�
[�F7O�DN�HB��jµ���.O�9�Vƞ"!���]��W�Ȝ�y"_�p��ߟ��I�������|�Oxڠ!FA�Z­�����s���B&�n� L1OP�d�O����$D���]bW�8Re�Z�$ƌ+kߨWi�ua��M��y���J�� �m��4�y2ϙ���!AF�"�R�����y�	��M�:�4|�ВO�ʓ�?���|����l����"�"�jzzZ��?���?9/Odo�[>v)������~s�CÈH4f
q��Ě�8`�?i�S�X۴ϛ�9Or�u�HAc����]�r��E�$-f-Γ�?�$�N�xK��:�b�~r�OǞ$�ɬ���V14 4����BJ���	h��'"�'��S˟��'�T(��bN "а�3lßtyٴs�Z��'�r6��O̓O�΅P>��cJ�H��pe�������=�ش�?���6�M��'R�S)��8]w�� C��#Uv�{��!v ��n�l�]y2�'���'3R�'���\K�*�C��#=��cqd�<�����@O�0�Z�	��`��}�S�����C=^�$����)�|��Ǣ��������ڴ�y�����Osb��7��%���Z�7����ug�?D:���s�\����Ϯ�$I��$�t�O�),�r�j���j�҇	�	�:ȱ���?����?1��|B+O�m�9EL�@��?F>D��0�J�a��#$r��	��M���n�>)C�i$�6�Ov��"c4���  �����I� 4�6�r���I#It�$�W�O����a�ƪ�d畘q=X��=O�~Y�G>O\��OF���O����O:#|�g�6"�cUA;U����)�8�I����4~V�aϧ�?��i��'Y$]��ִoڑQ�N�2�`)��5Oh�Jr��v��䅗G6�j�`�IIۤ��T���u�ᮀ�5ʘ�2�ز2+r�g��sy�ON��'���@��3�V}��\ze�_.T^B�'
�	�M����<a��?*�T�2!U��ؔB�@ʌ57�<Pџ�,�O� l�
�M�M>ͧ�
v�M�a��pjc�C"����l߽NF��A��� �3,O,�)�W����A�	`����)D�q�I*�������ğP���\�)�Sjyb"{�y����^�F��H�F����G���ɺ�M;��$�>QP�i�NeYd�z¸
���g\��b�t�: n����n��<���#��]@B���X8�+Oh,{���dVMB���1�`�h�;O���?I���?��?�-O��l��XN�>~g�X{�c�4 J�tm�����"0 Sӟ����?]���0�I�M�; �A�%�I�\�8!�B��Kp��i.6�V�]��O�����鏍-��6-f�lx�F� Q���v�V�H�iWb�8`��j�Ҍ�J�Iey��' rN 8�xc���;�-�Q�v���'��'��I��Ms���?���?����%LƤcV��5�N�7ƙ�䓴?!vV�`�4&!�fFtӊ��'@0qAKǫM�>���6cl���'�B퓥|DRB��0T���?QqE�'d�P�ɽ}�r�4l�5����6	)�4�	ߟH����s��A�4�'��УeCյ4�j�Q��rp�����'#f7��&'k^�d�OH�mK�i>�3+�ɋ�n�~��ZR��5�t��Ŧy��4sI����&���;O��DW!��� ��� ���W�K2q�\��6����0����6��<���?����?y��?�+Q)��-ˤ#LKG��2�`U���d�ȦI�L�zT,���Пp���?��ڟ$���?@��`�L�� �����F���$��*ش8���2�'@�xE� -X�$S�Uť�Ɛ� a� <о�@(OV4 v&���?	�)���<qHN!H@��gŖ�\�%O?�?y��?	��?q�,��dGѦ�6��?��f��rm�����nq�A̸+��	���$������Z�	2ߴPۛV�֚h��H ��3itU���&Y��=KG�i}�d�O:�+���r� �<��'h�k,�<���k��A�Y[���M	���D�O����O��O:��&��{pp�,�#B7�,���Z�B�:�	Ɵ��$�M�Mg~�p�"�O���F)C	is�-��B5��q�r�-�D�����޴�?y/��M˚'�b�ϦK�H�UiN���R�#��h����ʁ'�M��O+�D�<���?9��?��F�@�����`Ʌ4uޜ���Ñ�?������Tͦ�4�v��	ٟ���?-#`,L�B"�D�S�8�L8T�3?��W�� ܴu�&�|�O��Ԩ�F���v�6VHtz@h�O�
�yT�ڲX�XCc]���S2i�P7���o��mJ$捗W$��!C��[�H���?q��?1�Ş����Y  ��u,��v���TÎ�-z�w�6�$	{}b�k�$�&AR�a���� ���_e�����+%To��<��E���B�%��<��n7e�R�
��&OE���n��<y.O>�d�O�$�O8�$�O�˧f,d�{���+9W`�xc�˥r�,�V�i���r�'mR�'��Ol"$a���@�+� ��/W�Ҭ�����,9N�oZ��M���i�|�S�'d ��ٴ�y�j� �$䒷�;[M���c���y�O��xE����)<f�'F��ٟd�������X9
^TœDmHw�<��ן�	😕'D26MP���D�O������"���
.
UʵBZ6)����O��nZ��Msd�'����<��b�O0��Vc��@�d�n��e�u��z���I~b4��O����]��A2+�4`�G��DD�0����?���?y��h�x�$�&}�ݱo��w 	�M'2�����ۦs&H#?��i��O�n_? ���9u�W=bd��8.A�r��Kަ��4)5��l�)~�����|�q(�b��4�'@�=@BgW$��vf� M�|�&�Ԗ'��'\��'G"�'m�k񫐬{ �c��K&f�T���R��I�4as`5���?y�������?Q�!���gCס,��B�1$6�#*O2�o�M;B�iE��������ɝ�V��J��y~%R�Jū�>9�%��<����+�n�����䓃�H),�Q�1��o �Ms�i�+����O����O��4���[ʛ�A���ybIǅ?��x�mJ�4DJ�G��y�Ԟ��'���
��g�:�l��k��)+�c�@�$��& ��#��YͦU�'3� #�BZ�?I
U����z��I�Χ@)"D�p�B���ҕmu�x�����I��d�	����I6w�\e)b�j>9A�-�\:��s&�~�l���s�����(�4"N�|�'e�6�%����@�� l`H��NC-&�����͟�'�,6 ڦ��S!�\m�<��y4�Ւeo^�_v�"GT�|�QP�A���+�����O��D�O��dW8I���"U��W�t I!�)� ���O�M{�׿�y��'3RX>!��(���fn��I^Ne��3?�F\�d�شa�6`�O����)�yZ��bۍ��P�� (�Ȝ���E(X^ݰ@(�<I�'������|f8�
��`��t��͍�(���?)���?��S�'��d�¦-yD�ɝ'Ӕ(�3J2E+�0��bըk���3����$�b}2�z�8�Q��4h�!�c�JB+%��ܦ�ٴ��Ѱ�4��D�v5���'J �^�\@�&H�+`���\ $b��'��	ß��	�|�	��$�	B���Y!v˲d Q�K�m~⎉������= @�d���	ڟ�%?�1�Mϻb|��W�K�.�z����ΰ �����'V�fE�OR�S�S/���mZ�<Q4,�)�r�@�B;e�^�<�*O� � ��U�������O�����b�(2S� �LD�� �k��D�O����OV���[����O�a�$�Y�Sy ��ϭ5���xe;��������Sڴ9��R���Y�X���j�
�����'?�ժM����wi	��� �����?�$�fF���)ߓ-�v���]��?����?a��?���)�OddSү��K�\[��Cg�F�9���O<�l�7 ��q���T�޴���y��Ԥ:3A�JհH��k�ڛ�y2-qӀ�n�M۔i���M�O�P�,K5�jT�$+DZ9ĮN��@��'gK��O���?����?9���?y��"��pk��	�P�
a�QN��f�h)(Ov�oZ�^_���������?��y�Ƥ?�<����ֲt��p�1�-(y`�E���l���IL�O���#��ٳI����̝8̘��Ѯ�2MG��;_�cҫ����t��wybm�)]��0��@1+��P���<@���'?��'2�On�	��M3Q�S�<�D�A&�+���;\Dq���Y�<i!�i�b�|�Ȥ<���M�5�i��lkS�
@;�i�%����	���-ϛF?O��B`��Y���4ʓ���rB�X9�<a�!ƕ�x����5O��$�O����O��D�O��?9a�aO���A�bh&�kኑ-P�d�O��A��Qx�&*?I�i	�'}�E�I�D��-�KTX"ƴ�a��O�����)l�n�		���7-y��	{ц� .p�mF�d�i�씣��A����?�QA2���<����?����?�q
�
;��h��(/�����A��?!����$ ����Wje����՟|�O��X`�Iɳz1((�ÈaL����O,-�'�6-ئIJ���'�R�.޼g���DGI�X r�jp�K�&�b���\�utҴ�,O��I^�?Q�6�$�5^��K� @0s���V霫t�$�O^���OF��)�<��i�Y ߖ ���SF��w��bw`ھ��DY�E�?i�\���޴+�шt'��Nw����g�aD�����i��6��jۄ7mg���i��h�+9p����xy��L�@;"����_*#�6��n��y�S�h������ٟ�����O<����&�K��y���)W��+cyӈ�Hs9O2�D�On���զ��r� Hx4�'(v��j&3d"İ�4i��֘|�����.��f1Oʑ�.�-!�4Aӏ�Jie�u2O��bpAO2䛦(MA�I^yB�'�R��;4�Z����b;��`�!��"�'���'Y�	6�M��-	q~��'���{�@�.���h����WU���'�'��V@�k����Ic}b�Z�^l�W��PE>����Ё�yR�'��lI~cK[���D�Fyc���N��!dɘ���F�E�8(�n �W�b�d�O��d�O���/ڧ�?`Nؚ`Z�PwM�AB�����)�?���iBv��'�rJ|Ӷ��ݩRH(��	H�:�����,Z6�v��3�M��i�Bi�5g'�6Ob�d^��F��'0�<!Ywx=���8	����v�\��䓉�4�����Ot�d�O����<�"�2f��D8Hr�X����[���E{��Iǟ�&?E�ɴ�~�-C>k�Tx�W�ҏ=Q��	�OrMo���M˙'"�>a�gGG41@$ҁ'��:o��T`�,
�v@��/?��)� @ ������$QSx`��E�ҞN�x�V�ĕd:F�d�On���O�4�4˓3ǛFg��M**�ώ|N2��d�$��J`�(�$0�O�pn�M��K�X �a��* f�[��	N�U&�M��ODpXS��:���t�}�i��JE(%�����=HN*�Z2�e�0�	�\�����Iٟ�����~)�tZ7a�/_� e����?����?qU�i�h��O���b�H�O8T�e���\�!��c	޹��Ac�ܔ'�����A�c՛f��P��� �N찅ۄ̘l� s����m�d�'��M$�h���4�'{�'��Y�\�7X	J/ٺPϴ|K��'�rQ�Tڴ`t����?������%;�Ta� !?Ѩ!r���`�������Ц9��4�y�����O��h�G��6�Be DR��R7K :��&�P"��d���`��P�N�O yRD�Th�rB�fZ&7�nh��O����O����O1��M��-ө~/�$��Ⴆw��E2�͍�l|����O�o�v�P��	��M�#Î,H��%ȅ��h�
WZ�ٴ�?9b���M��'��w��X[w���'.�a;�˞:�҄Cb�D����'��Iɟ,�Iޟ��	����p�$E���+��+,r��HF7�T'U�X�$�O��$+�	�O�!oz����"C3ތ�*�e�S� P��C�Mk��i��O����i�BR7Mm�(H�!ύ/ڔ;�I��R���B��a���B��1Q�®�|�qy"�'?R�n%&�0�����F�٧O��'�"�'���M��'��?	���?�'��M��ݝ�H�d$���$�dP|}�ArӶ�m��<��Op�8A���Kg��&�,ݢ|pw>OZ����D�I���c��	�?E�3�'�&���5b	9�w�K�[\�x5��p��Iǟ��	ܟ`�Ia�O�b����д�D��J�&�j�#Ѿ=Z�)nӘ��CI�Ox�$�i�?ͻ9�B+�M�}���5mD!�܅͓ۛ�-o��\'�7�v�����i��F�O	���� �O��젦D j$��r#	Z�	`y�Oy��'�"�'\߃_�\����sq��sD�8*�創�MKd���?���?I�'��i�Oz�6b�l󘥩N�\J �P�CCO}ªm��(l��<�I|����?3D��jL)��P�y��X����*R�@�U��I~2ꁚ	f���I���'g�	)P�K���)䜼7�ߟ�d�I⟨������i>m�'��7��p���$�%�,�h�@�<L��s�Z�+Gp���ͦ���]򉆙��������4�?9�bAT��=�2�(uBÊB��q�4�y��'�NXSQ��?	0�O&���k�ٶ&���bwjơ����M
�<a���?����?����?����[� �t�����2�sWoA�nr�'�R�b�
�aƝ?��ܴ��ib��Q ��- '���X�x����'��I��Mc��i�" �?���1Ob�D�iX�@_2`LfLSf�'�8L+RjT�%C�D�OD��?�;����'%"�'���8E�[���kq��<1�f�2,�D�*�'�3&��,>�B1��O�r�'��6M��(�)���>^�,�fCR�M�b�ғ5O��o�5|+�]�I4�M���i�9p�`�E&?%��`���:��0ʈN$n��#� ;� �CÊ��d,���4����|�CϬ$�w��C��� b��':��'���X��۴a6��WA¿b8���r���8��x~"�e���TI�O��mږb����w�6?ޮy�j�qy�m޴=����\�v����w���=���hHOy月��H��
�b/�!�d��,�yRX���	Ɵ���<�	��T�O����c�Ҋ*�����EA�B�SnӼ83B5O����O쓟�D@���%"ې�+��*-�~8�.ϝ;�n\1�4��6*�O�Ş���ߴ�y
� `hP%��	2d�$h��1�x�Z3O�� U�O��?2�3���<����?�$刖����k>-.�9�˞��?!���?)����禵� ??���`��88��B��^�#�
�9�")@�B�>9��i� 7���'�%R���=#�^(B7Aǩa�}r�'k"셒tR�Q�/}����?��?��/�O��6['T�i2��$%8`g��O��d�OJ�d�OR�}:��$H��S�s�)�:%��(��fg c"�'��7+�i�� ��,\�"�J-`��LT�~�X�ڴ
!�6Nx�r�@2�jӘ�ɟ�F�ϟG!�Ĵ�xC�Z�,�8eR�쀽8��g�|�\�\�I����	�������"ܼj2T�%!��k�����[cy2w�d�s�Ž<���'�?�3G7-%p9���d̒��6$պhw��	�MC��i܂6�]��?	�
n I�J�I�p��&��2�$��h�0^�<��'a2T�F�柠�P�'�	Yy2� �Gkl����"5V�(��	�S�R�'@2�'�2 �&8*�I�M#�eɩ�E	�R^�� F"R� ���<��i�'�BK�>!p�i�66͕��:�e�*��X��G�,�8�ӵ�©��n�<	�X�XX��"�&��,Ov������,�	$�N)�֏�\�:!`�K��<I���?���?Q��?)��D�-N"��$��~(ܡ�HEU�R�'Br�~Ӑ!�:�H�$]æ�$���򀚊 �Z%KC�ǜZD�L`���<�O��n���M���c7�-��4�y2�'����
*���AR��$!f�4Hr����$$�'s�i>��Iߟ��I�J��E�%U����ъ�4� e�I��,�'.�6- �}��$�O\���|�)T���q��Φ�|�v
�`~���>�2�i�>7�u�8'>�ӄK2�Y�f�NH>��3.[38�.(��o�1L�~��f=?��z���ɺ��F���WKA:^�����X0e�h9���?���?��Ş����Y��LWM���"�g��H��$��^o�L��ϟ0S�4��'k��7��F1e�� F
J(��4��ڧE3�7��ODA#�h�.�	��4��/��+��Tj,?�uEJ7JF�pBG�#*&�(��<Y(O��D�OT���O��D�Op�'6ؠ"fO&YIjD�N־z!JѲ�i�4-��'��'e񟤔lz��s2T�Z'�3<$TB���X���v�H�IDy�����I^��ܴ�yK��j0^���'։:	E��O���y�㕯/Hj��Ii��'L�i>��	!<�NlP��ԬȆ)Y�h\�������Ɵ��'�6-P�kW�D�O���Q,h��0+T@�CH��$��g$�l�)O���d�n�O�	bAR(,ϐ���H�EU�(s�8OT�$�GlSVC�2H�����`�˦9ڇ�'��-�
�Y�`y��._�6���g�'���'���'��>����}�^�ȥA���ڡ��'䌭���M[P��� ���4�^�ӓB��p�(�R�� �4�b�;OԽn��M��n�i�ݴ�yr�'��A'8�uG&��&�f|в�F>��4e\"x�n%���'F2�'/�'���'�#��ڳ}���
ӎg,8�@uU���ܴD�p8��?9����<)Dk@���`#bj�;��0�E��	!�M�u�i�ɧ��O������� �Kv��Q��	,v��	��52�5hN ��q�x��M>!(Ol�񋁑9��0�R
H�XfG�O����O���O�<1�i�� ��'���Y��� �
,�q���{>D]	�'�7�1�I)���N¦�9�4�?	Q�Z�|���{�
`�@����H�r����4�y��'$�%P� �6�u���Sy��O%'.��%�ҴI�M8?	$�0ծ��y��'���'�r�'���IȴV��t�c጗��A��G2G���ڟhKڴq���'��6��O�˓J�6� ��w�2�Y�*r�2L>Ya�i�:6M�O ����n��	�xRV���g�����X�$�
�I���a���[For�@�M>Q/Or�d�O���ON%���L�E�49��'
�`9��O����<9�i˪tr�'���'t����
`j^=m���^�< �~�I�M#t�i�ɧ�T�O��\�2��Z��P��s���L-3$�F��2pp��?i��LxӨ��O>�VF<pN�Թ���j�*$���W��?Y��?��?�|B/O��m( �X�h=�^��F��z.t�a%�ɟ�����M����fu�	�M�A��Z�B"� 3c6�b�Uq���'ʺ9+��i��d�O.
wKO������B�Z�kʴ����>Liɢ�i���'uR�'���'	��'�S�rN=�� �X ��I�/<2x�ߴٸ����?���䧸?�Ƿ�y�5/�x� ��<|%��Y�oQ�����`��Iy������W��@:۴�y�J�Ą���	(y?bM	v��"�yROL�:����ɞ`��'��i>y��/(:�	9E�j�5�Ma���������'ݼ7�͹e�h�D�O���`=t���L�7N
#*��j�2��<I��M��'�	�u�����N�oL2t�$& ;-2��П8�C"l��Ѣ�2?1�'@��D���?i���-b �&�QT��H����#�?���?!���?	��I�O쨘��^"j�l�#����L���G�O�An�F�|��ɟDsٴ���y'��)P�e�� �4g��8
�ٝ�~��i!H7��O@���BxӨ�ß̫"H�e}��t��p�ì�.O�zLʱ�\7��rI>�)O�I�O���OD���O��;��N��@�E!78�9�i�<���i�`�p��'�"�'k�X��HQ�("6ڪ^j��#��t}B�q��n��<�N|��'�?�bM�? ���-�/H�IsnՌq,���-	��ɨ/Z Qq�':H!'��'<��3���Z0R-�a�:d�S��'���'W����$]�4!�4^R���*m:#�.Ok� ��YW���dV�V�',�'o��	�6ijӦ��Jh"�yQ�J	k]�xõnˇ� �3av�b��ޟp�Џӥ��t�(?��'R/kLG>�r�Ӡ�d�Dx��ܔr��O����O����O �7�ӕZ��*!�ѭC��5#�.��2��T�I������M{���|���v�'�剓X���V��l땃33�� ͓��w��m�ǟ�Z���	��?1 �!.�V =6i2(z�O����P��OB�kK>�(O��O����O�M�m�,N��� g�?u�z��s��O���<9�i�����'���'��T�O��`F��rnYؗ�;=����O���'�6�Mڦ����'��D��7�\.o�Pa�t�ͥkM�#+��20�u�;?Q��pat�D���0�<*ī��X9{Gj�/dW�����?1���?)�S�'��D�����ɭK\����L�;S7��sM�I����۟�4�?)I>gZ���4@�:œ0kđ"˂�S��_���A���i[��7z�:O@��ìwF�0[�'k���Ge��H�ʢ
�	 3H��+/��Oy2�'L��'R�'9�S>��/����hC.ٯ ~� b���M���Z�?���?�����OD��w�
�s�d�5M�)�/ܒS�ZE�p��8nZ�<�O���x��ѵ$�6�v���cN:�\��q�W�,!I�Nx���a��m��RR�IEy�OZ�6R�̫�˃3@�U��
�XR�'���',�ɏ�M� g��?y���?�D��%Ɲ��'M�Y����)�?QJ>��\���ش_z��9O��ct�ȡSi��T��q�`��c�JH�'���
sKU�Y`�50��D��럔0u�'�� JC�ټ3�2y��aݟ"v��K��'�"�'S��'��>���RT��n�H��� ���$+�N=�I�Mկ��?��r&��'�ɧy�U�rF�[��װO�y*���>�~b�'��&�'צ𚗹iq���ER��O�
|z�8fBuქ�IQ(R��g�Iy�O�"�'�R�'��E	4�l�aѣ���gK��2剞�M��<�?���?K~��tw $�"�?�r	£�C6.���z2W����Ϧi��ħ����$5�<�B�[��x�%�ٕ-�xs�G(U/�h�'Z8y�e�͟��r�|�U��9t`@�>�b�#T�H�SgFr�A�ן��I��I����]y��w�RY�	�O`M�7D]��Bp���%.T��'�O�m؟P%���O�o��M��gJ�ؠ )͍Ex�8��
7�2훴�]�M�'�"�V}����S���D%��Y
���Z�em=궄B�WUu��?Y���?y���?����Ok���h\%+.4	�'�j`��P�V���	�MK����|B��D���'��ɴ|(�>Ɛ��� p��R�\�<1)OV6�æy�In�`<mZ�<���m�ȝ��ɕ��l%Ώ�H�|��/�/�H��S��䓂�4�^��Ov��]�{Ƅ	���{���9%'̀S]x���O�đ&,���"�S�����O�$����?!�0ȡg�	xp��ĝA���@���*�M�r�it��>������p����������&W�`��\�n6J��J�����?Y���'��$���cJ�1�x�J2HG8�~�k��Mş@����I�b>Q�'3�6\m(Na!�̎n�)bCP�ub�$X���O����ܦ!�?tW� j�4{$�Lhpb�,n+ �c���4�tM9 �i5��H�H�F:Ol�d��/�ܱ��'S��ɮS�`O��M ¥���&��IIy��'3��'d��'iR>�Agh T[& �����ZX�Ѵ��McEL�����OΒ�N����睷MS�m8I�=r_,����O	b�Ty�ܴMB�?O8��|��'�?�科��M�'K��9��	���Y�- 4����'������ޟp@��|�S���ܟH�C�F&'�|LK�%�'���[�K�ោ���8��ky��j��a ��OP�D�Oh��n��2��͒���m�Dq�&�	���d�󦭺ݴ�ybY�,�gNA�
����)fD�0W�l�D�	��jH�S��q]$��
���O�HP��C^�t����0�2�y1Bߤw��;���?����?y���h��DF37%�8�D�F�$��V��1 �|���妙�A@ԟ��I��M���w#���"ܴ6�M+��ġc%r��'��7����ɠ(AMn��<��{$���c���[����aڴ&�8x9#RHU/�䓝�4�@���O�$�O���9X*�(+a�Hܠ�z�l�z��d�OR=�6�1/ʲ��O�����?Q��}g�}��D���d�� ��6�Iҟ�oZ�<�H|
�'�?���>z��)J�	��}��CR$�.}g��+"��~�H']��0�I;�'��ɗA�@IP'�Q�ȑ�J�*4�����ߟ�	.W���i>��	ß�]wW 
��'�`5C��Eq�|EP`�x̒�'�R6�9�ɐ����O6��O��8%M�Q� ����ɦ!:�8k@��<��7�y���g�JE���O�t���ƞ��wˏ���]rc�^�(�0e��2O����OD���O4�$�O*�d�OĘ`P=��邡(нO@���%R?4d�|�Va�O���O�o�y�(���*ٴ��^��D�c┭l��R�+����۝'%���M���i���hj��=O����/O�mj�H�z��a��#ƴ!d��A�ۧ�?�f�;�$�<�'�?���?!�dƪgE�-�eBV-�x������?���?�ucؐH	>UCB�*�?i��?9�����њd��9��L�W��1��
��$�[}2�w��9nZ�<iK|�g�? B�� �G����-a'6� �ӡj|U+�
� ,%���?1z%/�$|	�hvk
mD�K�� .C�6P�֏ -fΈXjg)�g���E�8w�``'��|�j��V�$W�f0T�;J�8�+�/�S���`^�s�)l�8�� CNT�dXwG4�*�я{2(�
_���F!��~���'
B>2�����n҂7��	��E�7}x^���̀f�N��RI�;Ml)sGf./��\�Fkٔ�\iRC�-I�1Sq�Z� `	��K�Zf���#aӈz2�l2b��n��T�d_�(ג�7���C�ө{r�Pt��}A.Y��/��*-R�Hݛ�ސ�b�@c���v�F�$�%�\�Iܟ$�X�	ܟ4�t��w��=����!7��� @��&�8���?����?���?�*O��s��馉qwe��^|*t�5��7�4�c�����O>�D=�ĳ<��ąI}"�D�q=@ة��ȽN���SaΜ����O��d�O��+�����Dk��t�M�@�8o�X��b�6_�6��O�O�ʓ_F�~�+�C����l��s�*��5�˦E�	���'Z����:��Ot���j�CS�]N���W�h7�8ac�xR��a9§����8YD�sT遌M0��/��M/Or��!���A�����$����'�$�x�HF%$Q<�@]�c�`e{۴��P�A��)�O~nڡ�� з"�*\�j��QKY�G��6�$&��Im���I��S����|2d���I�k��,SA�К��ӻ:X�Ɉ���D�<�H~Γ�?q�d�z@�<a�@P:0�	P�Q9Q����'�R�'a�#�d6�4�B�$��,��Id��P��c����$j`�p���<�r`^d̓�?A��?��+~E�S�ق@��󴌒�D�ҍo�������|z����ӺB��%�l�RR�9rTL�rC
s}��#�':��'rP���#@׆w�LM�`$J5f�R��"�!WNv�cO<����?�O>�/O 	q�"b	8�"6oH&L�x0��e�NA1O.���O2���<ᠫ�U�I�9	@�<X协���p�3)F���I�D�	^�	jy��̆��D)O�Jx�Tċ8S�޵�֪	"m���������l�'�fI��1�*G���v`�.{w��96�(,��anğ�'���'�Xӈ����0���[6�D#e�,���� ��M��?a,O���hEO�S˟��s��xul���6
 g��0�)<�D�<Y�Gl�O����$5�� �F�'Ԍ2��I.Л�V�����MS ]?e�I�?i[�OЄ9宓!Զ��G댮tg�XkC�i��	�cu��S�t���4Z��1�%'ԙ\��B�C�,D�Rao��b����������x�Sky�O�򏉂c�*)���B.�!�D �v�r7�y!�3�����e�9��Q�ե0>e8p���M���?!��'���(O�)�O\�D���˷ǒ
c�������>P��\kp�K��'��$s�i4�I�O��ı�L	� �F�2䄉k8� ��m���_�t����?q���?y�{HW�@��� �	^�f!yҠռ����?oڲA���$����'����"d�� ���$^ː�H���6�|\K�_��������z��?��/ӏfz�)���YA�1I$(�:FI�Q�BM~b�'F�R���I��d��'C��$�0+ƎP'6���L1�J�oٟ�������?��L��p�V!ݦ��A_�A@�p����,�{ �>����?�.O:�$�6/Tʧ�~��3I3� y�엋^�"-�CL֐�Ms���'�r"M&iфqK<	7	B�F���1.A0�� ��/�A�Iyy2�'b��Q>��՟x��`����o�'���I%����<��}�'h��iad� 昧�I�ol�]��F�J�R��T1za����|���V⟨��������?a��u�Ø�"��U#1�Y�1Y��q�f�����O,���PI1O��ب���k���sP�X�$�R�ic:�+��'B��'R��O��i>U���Z���ㅆ2g��rt�0N��uc�4IM���M�S�O�2�����z�LG�*��Ȣ��]~�$7M�O����O��\y�O��'����A����Р(a6l�2��)EmVd�<ٕč�:��O~�'E��ǰ7�̺���&iI.���L $S���'�h	�4\��p�����O��4�Q�X2-6�Q��"N��A`�&�>q��!c1��'j�'��	۟�q���%$�U9%���� �E����'R�'?b���O�0�T �9C^���-G�\<X�JB�Cdn�jě��	ȟ�'db���W��V�*�0e4#�	���b�`N�Qӛ��'�"�'��O����8��Hb�i9�d�@EG�����w� 0a�/�>����?�.O���W"�ʧ�?�6�S	����U$b&"�@�O�� �v�'$�O�˓��X'�H��`����2��/��`�(g�v�$�<���F��]a(��D�O����$MH�R`'X�*b�M`VH��/\R��>�/O"����i��*�'^���A"��8��&ʢ>��i����?��?A�'���Bi�v�ޅ'l��� �<2��$kP�8�'�*`����t�	 ��r�c��TTE�@ �M��J0�?q��?I����/O�)�O a҇s1J��$oH)g��|��f���A��i��)cb�"|:���1I�掻G�V��FO�Im�8�G�i�b�'�2�A�G��i>a�����(�	#��N)`��a� �Q��z��d d-lP%>��IΟ � ј������u�3*p�l���`ƃ^y�'���'jqO� �d:��;P�d�YR��ɤh�D]�$��&-(���?�����O�����P���E	�DL>��'HU�]�˓�?����?����' ���n�;j�M���Y�#S���' �XDX�O��D�O\ʓ�?Y��o�?�q4�#\Q�u�%LY*�h<�U�v�4���OF��?���`ô	��$��6�Ԏ0�$���
k��q#�����ݟ�	Uy�'���[q]>���eg��9�I��)"�k%��r�x�n����?���%Ш�qw@JC≹�	�兎w������ �47��O�ʓ�?��c������Ov�$���%k'�Z^�4%`��N6j����c�n��?�Q�Y>����<�O����*OR~T���0@5��OR�dܜK����O����O��	�<��9A��S���
��h )�Y�:�',�m3S�R5a�y��$�Ϻf8�kgN{�VhI�G�'�M밦"�?����?�����.O���O�5볯�T؝a��y�9S�������J�l�rc�"|
��5L
�9E��R)�u��(ZR94�i���'��a�'��i>��	ޟ��+*$˔Ƃ5fy���D��cB��G��(g�Y'>����`� b� �@]A���X��=��nZ���b��yy��'�2�'�qO�Iե��z8 ��M
`�U�sZ���B�&����?������OQk��ݦ�̤8b-E	J�"��U'����?����?y���'��X����_���f��FU��͔�T��� �O��D�O�˓�?�#`������Rmtؒ�B�w����!�
�M����?����'�Bʟ0~Ԏ���41��J�L��g~�$����+�<�'��'_�I�|�6�OV���O������t�C���$�^���i"��d�O����
�m��'Bz�����#��2��H�Պ��ܴ�?	.O���J�<@ʧ�?q���QcѦ*��C2L>DN ԓA�J3y2�Of�dÖ7�T����T?�3AE�YO�DzF�	�<�
1��>q��r�)���?�(Ot���<��_����ι�n`z�΀u�FU�'vbg\�t��Q�y��$��.;���$ʂ7<xr�B䀏"�M����?q��?y���r+O�i�O(�`6a�'X��b�Hr���JǦ���Ĵo�b�"|���7�tQ�]'ku�ɂ7K�$֘X�չi���'���K�k��i>���ϟ���u�ȸ�vU�3�~�W�^+N���P���^��X&>A��럐�'�4�@��S��\Ab0�Rbq�o�ğ\#Gg�oy��'b�'�qOF�:"j�%Av��VhK�"N$ATS�41�͓	=��?����$�O>���/&Pc���X��E ���J��?����?����'����A�%'3Ȓ��Ivź��$Aa�:���O���Of˓�?鰇����Ԧ��^I���g��Af�U��M���?I����'rK�_nH��4%��\  ��0u \�S	67�i�'p��'�	ןT Q'�k���'_.p���;0Ӿ$�7,��!~A��c�r�d8�	�X�l'��O�|��dG����*�B��Ȓ�i�"�'z�	�H���A������OP��В0�"�aO����|2��}��'���'m��Y�y�]>�^R�b��4m�q��g�t; A禩�'|lb7�{Ӷ�D�O6����6tקug%V���� ��D��&��#�^��M���?)���<���?���6��O2���X�/nB�� �6��ش,!�S��i ��'���OҾꓩ��/J!��K�D֮4��Xx5΂.mVB|mZ3Q���ܟP��7Pk�=�����ΐ9��?�l�z��xu*�i�b�'�ڰt�:��'����8���Y���v|(�W�Mn��X�'�z)����I�O��D�O�Y2��A%��PJQ,���r���5��*3Bɑ�O�ʓ�?	+O�����UZ3���cc&��ҩ�O���Z�l3�"y�t��ןH�	����	gy2OP%�p2��ndN�Fa�*�
��э�>a+OX�Ĺ<i���?i�9�6=0`�Y�B��9�n�J��GP���?���'�F�����?�(Oܹ���L�|�(��X`Y�s%P4��g���Ŗ'�]���I쟄��*{�<��-M���s�m�c*��3�E���HB�4�?)���?����򄀡?����O�����5V�,Q��DN�޼ q�W�-�7��O0��?9��?�Ǚ�<H�(��M�-B����1o ���k�����O^ʓU����V?���۟L���7 �I��K�{j8a���	���ȭO@�$�O���G6s���$�$�?}���D�h��0+�Z�)J#hӜ�	 Z� D�ib�'���Ox��Ӻ�Yح!��SC�ب�eL�	]��l���t�I*��I��9O��>�J�+�wJ
����ΎX������i��bĻt�v�'���'����>�.O%S�֜	��=頯�-%�:���%C٦��x��%����s�	b&��Y ���A�,�"p�i
R�'8ʊA��꓆��O���:U���G�4'lZ|Z���$�6M�O�ʓ���S�T�'U��'T�Z�c� G�Xi!h�� 4��Ie�r��W�,��'������'�Zc���K֡�=�b��;U��<q�46ĩ��S�<!��?���?	����d")�,��b����J �߫�ޔ9P�B}�P�8��cy��'���'?����%4�@��0~8�����yb�'�B�'4��'��/X�X2�O�b��� �1�0���-H4=J�@ٴ����O4��?��?�J�<Y�� ��Ђ���Hi�eC7��f�°iXr� �"�'B剽kUN  ����$�u�J��mW��t��rg[#yhlџ��'�R�'Er��y�]>7���h� D"��_�0�z�SՀÛZ����'�V�P�h\���	�OV�����q��h�pt SD
 �\��3�Qg}��'S��'����'=U�<��{�D�*�,r��h+�"�Gbd1n�hy���6m�OP���O�)\}Zw��p��JWbTrM����	��:ߴ�?��^�>�͓Y��Ӳ��@�}2���;�e��X6)*��P��A�V���M{���?���z��$7��!�%S����:ȅ:�)o��4~`�Iw�`���?��&J�x(�z�6~������q��v�'n��'Q�	�2�	̟,��H�`s��,b�LX��㐋A8�o^�ɻ�H���_y2�'�r��5�)>�b=�l�>�<�I���M���W�FI���x��'�"�|Zcvt	�paL�4¤EP�fG�@*�ݱ�O�(أ�O˓�?��?Y,OexeH��<�\L�bL������̭f�'��	��L&��I��X��""l�(���'d���7K0G�%��Ly��'�2�'3�	
}���h�Og|k&�_5�@ܸ��NJeHL<������?��\"vA��`�R$��%]7�C&K�G�~`�RU���I�����Wy���w b�(h����gflbՂ#���8edO��%��i�ޟ �	G�T��u�0��d�#.L�E0s��%]���'@�S��jw)���ħ�?��'	���Yf+F^��_O1�W�4��ǟ|�D��(��c����T9r5����7A��c�Qͦ��'�����|ӈ��O��O#��o���2W�N�aM\�`���l�՟��I�4�x��IQ�	`ܧY_r����q�>��� ��D]0�lک25@�:ڴ�?���?��' D�'�KM*5�d��WS{�V�r�]�{/>6��n��2�7�SʟH�e��
��%"�[6a��S��9�M[��?��E�p���d�O��r�>�rg6��y�����;]l7�:���5F��&>�������'M���E��4mŸ��ADP2ª}n���֏��ē�?9�����OkLY�L�tM�BS�y��h��M1��ɑ'- �`y��'R�'��I�6�� :��<�`И8�5k�� ����?a���䓳?i�Y���PjW�hS]�`�N�7�����?�.O�d�OH���<�r��+��)S��l���I�����I
�5���E{r�'/�\��')���B�Q�	�M	`9S���I�~���O|��O��;�< K���Ha��¬F����!k�#��6$ړ�?A(��?!L��R�2;P� ��ځ�X�0�l�,�D�O��3w�-2�����'F�\cjptr�*�#�8ؙ��I�p�Qa�}��'����'iɧ�IͰ=��� M�j�� W�ZH��W��a ��M+�T?a���?A`�OX�+S� �&�*�i�D�Pߢ��%]�0�ɡ�r���z�)��<l^�bTÌ�	�`:��ݮV��7MU,h����O����O��I�O�$�|����:=�J�, �4������lW�I�4!h8!b�+HY�S�OJ�c�=51QqLB�:#�c�B�"�4�?���?A6��;���q���'T��P�{ʊ�
Q6��D �o�/_Ťc�Th� 3���P�	��,+��N90.6x������t�s�]��M�Co&XI��?��Q?��IV�	90�Dh� �-h���v��Z����O��`"I�,��������Ο��	�	ԡ�Se`ye�B=V�܋ N�.w�y�'u�Iߟ8&���	ߟTt䟊m������0&̠!c�gB�v��U#�3?���?�����ԙ(��ϧA����1�Pŀ�f@#�Uo��`�	ʟ���w�Y$����'߆e���G(5J�뒈n�P���O��d�O����O��^�3��d�OP��.>)������T�XD;�F�3Ǆ7�O��O��$�O^��Fj�4��'�j}�aE�%0��P����_ `ūݴ�?����?�� +������?�,O0�����u��'��b��U�F��N��&�p���<i�c1+
����jx�� �
{`���KSY�7-�<y���7��V�'n2�'��tJ�>��4�楺ř�P��J���M�A$���U�O���I��X�\6d 6Q�n7sj>i"���왕�OJ��<��'��d�<�V�ŌW�􅩣	EA������>j��mX��\��y���ԟ��b�9�����2�}y�B=D�x��#ζ0Z�����G=n7D���9�OZ j��W�;��d8�D�4u�j�i`g�GL��J�iX��3&- �B~ݑ��5K���GG�:i�:@)�e�Sd��҇�A�E"����ǹ[��ر�D�k*�)��C�� ,�ďh1��D�:���P@�؋K�=B�ŋ2Z��c�@�1�hu�K�?m,��T�T&{FzPH����?���?1��Hxt����?A�O���w�ڙ?��B$E�5p�f�K��C�5J�ePbL�t<�\s�l�" u�"?� �͈lҲE�+�m��Q�Y�JAGꑁl��R��Y-~Q�i1��X�H�́i%mA���K�����XK�͆-y�> 
�ϖ�]�f�c�,�x�'�џ\���|�� �+%tP��E!D�hD܏{�XQ�C��&O$|Թ+`� C�O�BH�@3�X����O�T
�34���J�h�37>-`��'+�\�@�'�r�'0��A-X$�@u"��O�39��T>� )CT���v�4m�D�Y+�:�rf�I�P2ԕ2WH�f��ըG �r��0a+�a��	�%v$H�8�"اҘ�<�����	i�'|�DC�E �h�1]�����?�S�P$E���ǅ�p.I���`�xPO<� ���Eca��&��A�E@��<)D
�(������O�-�$�'�"�'��@B1�#:�H5Sq�&
� ���?.����OX;12�ݻB��O�d��`����8HXh��h�Z�d�;�q0-�g��I��9�6n�%�?E��9�6\ ����p��1y�ȗa��3��?�������Đ|� �:9d4 )��41�V�c��
�y"��0K��2��&�lav�W3�O� Ezʟ� ��O�S�XA�VCK=eO81P%�/4��
s�L r�t�A��ř��	��(<D��ac��U�<`���'T���aB�	?"��u��1�^�cl͸n} C�I�R���ƌE*;��tJ@ �.Ef�B䉈9��+ ,�;�n�SA#Ǒey�C��&vu� ��M&.}��a�DF�nC�	�VaC�� ��}�1M��U DC�I		��I���7Z�6bݞ7��C���@2���e�%��AZ#F\�C�I�f��kT.%�@Ő"	��C�	�����B��m��T,[zlC�I~�ӵb�p�= j� �$B��)k�z�s�\�
Ab­�eM�C�4v�Z���k[=n�XA�EM.@,�B䉿1h=z�Ħ�b7�W�}�C䉾bD�I�D�I2oG1%B a�"O^ukUN-N�#��[�:�h�"O��,�4���D ʚ^��yC"OF��FEŌ.\Ȅ���/`��=��"O�Lʡ��5m�D�B�d�G6^��"O�r2�M2)N,�4���%|`�"OЄ�,�:!��5��.B���"Ol���$0q(�#�\
�,R"OH�1�#wp�\)F`K�J�X�"O��r�H�)6j\��4JDʲ"OfRt��;���2f��y;�,r�*Oh�y�a
�%Tc"�G ^]J�+
�'_t�� ��D$���6P��ܘ	�'�д��#b������$P�Ԡ��'&䈢`�1�8��לB�@Q�'�RA�R���)��`�һ��IS�A�<��L�p�����-l�)k�|�<1tnˋ�BwF%a�b��&LQQ�<�3���dV2Y3ԧ�#:�ɡ DQ�<�b�٤�ni���o�p��GG����Mñ��.i�(�r0�E��c�F@-/v\,[����@(B�	ZEJd24� -BhB0�ďf��S�\#cn�d���kVc �3打M�ά�RÎ�!644������C���-)N��Ηn�� �=H�8�Qk/i|�� �<RP�х�Iz�
(c��� ��1���^�$q���D���;p��5V6�$��*�OL����v��DS��Q]�65� "O���!S��Q3͈�Q}H����ʥj�#+j-� �эA�F�4���VC�I0'��-:B�"�8��D�<�TM��j�]�Щ��9V������ �Tz0��$O$�`����-���I�gc�l��L+�s��p�⅘w���AF$]/J-������M-v�@c�6�O 0
QG#?�(��_�f�p�p!��Y������p~|�h� ��첤��/	���c#E�x�O}P����F
��oK�'W�-x�& ,1Y֤�2�2<��`ً�?14&�>2ƴm�%)97\:��bC��œ�ƙ�i�4%cg�J����s�T���Լ�P
r'���� ���T��Vk��$�(�j}>�D��iN�j�Sv��)?�DD�Ea��d��E^�A�"/k����ɜd�4� gJ�{�ȤC�;$��J�B?�&u�I�Pt>�@D')�s��\2�O�=��I�F�(����I�8"��S�k*�p���	%$�ZE[���1B�AE���0���aoE�e�� �m0$Z(��)� 4;�Y��āR�"�<%�`���'{"�*v!f@+7	��yRE�,g��C�//~^�����<�y�R6s�����r���&ު��	Q$�\P T�5U@�b�So��9Wj��-�� 	 ��C䉨^�a�'f�bҮ��$�� �D���c	�������˛�k���K
�P
(ȱ'�>�y¯I�J���z���K�Ĵ�5F���~2��#T�a}��.���C��,�0T9�O��>�v��̙��KO����/D"RU����9D��i2�؟3'�3�`�!9��Ia��3D�$��%�+�,�Qc�OZ�f�[��1D����0��0�tG�>j"��Zǌ-D��0�ϗ�(=�U�V�W�vĠ+D����@G�l>2�O�C�d��$)D��B��ͬ$<�<g�N+�X4�@�9D��`��իWI8tS�M�?���k��<D�̳C�w�D�b�יsϼ-�t�9D�؁���{^�i���>m��0�,D�T��
D,C�T�� �ē]R	SA%D���`K��
c�Z`�u�'D�����9��XQ &t�(��e'D��*!j�X+$�s���j����a8D�D�sE�.#܎]9�AZ~���0D��y�/��v $|��j�"~�a���-D��� "[�6�{�G
�wm��B֨/D�4����rhR���au����$:D��҆���,"K4S%�%S7�9D��q�T�X12a��El�,�Ӣ3D�K��3��](���2\��e�n6D�l��W ���%6��y� J5O�0@q�!�	Npe䖗oL]q1�ڑ;bC��?g��#pÍ ��Tpؾ>�4�H4����钤*��{vE1Eo
����87!�DJҴ���eUFȓ�!P6�1OV��!1<O��G탠|����ў�CO�����ˋ\�4��ӁljZ���˖	F�B��=mEBi	�D$Az%c��9] n��DJ2p(2�Q��I�r����w��%LOVܸЌ@�?M��� "����x�
4$t�䐘z'l|W�-D��"ФR���s� ��b1Bd#��0扽f9RDcA�/E:P��	ڋ*�qX&�/H�@�ѭ�y$سw�Z��񬉕1��h�(��/I�;ר�8Ǌ�@Q�]E��O�yhG�U�:�ég�x�"O��a$EʛGL�H�Ci�V�8�[��!�E˙CD�h��i�Z؞4BS��7c�&x�S�Tؕh�6LO�����=.�Z����ئ�C��՗s�"����v�ڡL)D�(����1耰B�'��r_�mu�&扬vW�MX��^qX��)óC���p2���Lm �H��E!���&�bQK�&��(N$U�S�U	�LRp+�0`��'��h8�𙟬iEM�s�H��숍/�2m�v�)D��Y�͓�b�B�mm貄ƞ!�,�1 �.�n�	ۓ���FL2C�T�f
�|�Ե��	�%B�EsH�q�J�X�4:��
k�.Wxn�*p-͕Z�� �ȓ(l����LP���h���1����<)U��5����B�Z/iǑ>��u0��q�Q7�\��Qe.D���2់V(�����Г�JC	*�h��C�����R>�0��!%��9�6��IU0#���ȓ4���D)�EY��!0ILJ���C�,D�B��
�a{2nѰ
�����Ϝ5d�������'l�س!����d�;+b�ɺ�Mc��=3����)aD$lӨv�<�sh8�$SV�&mꙀ��^�8�6��'D��s�O$X$>��/z�)�C%I!"zn��'i�>��z�/.D�LI��A8$Q���P, ����ޖp�
��E+�O���t%ҮV���ӕ�
5�敐��'{��
����� ��ӂB�f@lLX��FU�!��"O�)�W���7!�d��G�:��� ��F�>���@�O��0��ER������G�t�	�'�X�xP�Ɖp
��b�?��q����'�5���0H`���h�\����u`�lz7�#D���E&ܭ\���RI��*��H���]l���u(:�O�ePa$ے � ��d��)%t�R��'�@��ǖ��dۢ~��3,��%���a)�!�d��4x��&�N��V�$/!��|9r��6É67pTysu��3& !�Br�x�i"�V6lx�����9X!�< 2�{��9h\T��I�
�!��3l�᪥�	.mf�أ�Z*��'��P1G��<\n;����,��݋ro<.va��O ]�!�DےH��L�a�A�*����H�J������v~R��J�0c?O�\�pD�5K� ���F3il�$C�O8<��`�$N�Ȗ�&7��� ًk=��:�J�Kl�	(
��� ��є{�^t!��Ū=��q��I�-�0�����QsF��\A�P,U�O�	)bJ��K�b ��A�v��QO�e�@�s���o�V�$� ���O3=׆��(4�a~B!&�+�)'�іlB4���%"���B�µ�ul	vN�����-|9��<�`��L<�D�K�_��0�G��h�U�DFH<��G�9��-�)��7���#A��t��� ��y��ɕw�RT���C$	�i+��_Q+d��$F�L&ē�l\����"��mZR��j±�A��N`�B��"EA@��;������K�H��O�+7�ܕ�@�1a�Ӆ|�n�B�a[mN\3T$�;Xv�C�*����W���ؠ *K�|�R����D@0P�Z��~&�`y���|@ޔ�V�_�>��91�C1$���&�r��#�'e��B�cہBd"��,�;z��D�<�T!R�Eɳ�~h%ꑋ& ay"���c1rݐ�J�!��DG�{"�{2H@�Vv��bďs !򄓻Hp�tp��&h66U1G��WI!��_v���s�!�B�a� 55!�D�3� �2(�9l�l2��%!�Ύ^�)�E��+&�BQ�e�2zy!�	mIs��L7\��Ea��N8 !�D�-��ɲ5(�J���:F�	�.!�$B0��H�/�v�u���%�!�_��J�*rd��C@�5�!�č�V=>ق�c�"�v�ч��<P�!�䏅HѲ����%��<kW�$-3�'�ʹJ(��7��� �Oܺ6h�+�'� N�	1w�6� "���""O4�27(�28���L�o~f��"O�Zө@� *��` �ٓHr 9�r"Ot1�䅼cg��@�p�	�$"O��8C+Ѥ}���Ac��mm0��R"O�t� ,��R �ݩ'nC)cm���"O��A�摇4�#��<[fB�8T"O"��l@75�hQ�BR�J�ߚB�	4�JȐ��B2pB��H"ZJB�	#0��3��	_BV|���:�$B�I3K�A�AΏ ��5�u�	L��C�I�R��)�:Fk E������C� ��a�RL5&gp���đh=�C�	�K5��B��F:T��a� �@�A&B��jU�i+�/�.v�5���9/��C��+��)��� ����A�wɌB�ɨRP���W��	$�Q����*]BB�	JP�,Z��@ t�A���e~HB�"y+�X땉�6E+���1�X�4B䉷�nE�%��W <E���NW:B�)� �U��.�j�`�C-P��A"O�U�N��*��s�^�?4(��"O8m��`�f^lc�LZ<��"OrIs#[�Fբ�Q9gE�J�"OX1elV�I���Y0Z��<)z�"O��i��2T��+@,�"OZ�ڣoԯ�n�[�&�f,V�"O�$�P�T��J`��eC�M,^Q�"OB�+�4��(��ͤ4���"O�}���AO�>$PĠ�>O��i��"Oz���8'��(A/�}?���"O��"�s̈ܚ�LƩ60(,�"O��FoC�'C@`�q.O~z���P"Ox�[a��'4�B�C ��(T]�]��"O��'@���
d�yV�I��"OP��JJ�	q��:���s�"O�8��kY $0N�*C�΂��t"O�����9Nm �@\��P�"O���Kӕ�J�� !�&`h�ћ�"Or��` =,�ԉ�MU<L
��$"O����� /�f���Ӓc@��
"OHt��a �c���Sa-*:ъ�"O�E�iמ5���bC��,t���"O ,PE
M�a쒡KW29�D#�"O�5Z�O�M�����*\�&�YD"O�8��͎&?v��%Ɠ0�bѱ"O}�X[x� 
�*�\��q��"Of��&+��P@�k���|���"O&�єDǇ6�@��`�u�`�j�"Op(�%��?�F�ء@~-�(�"O�բ�.Z�inW�"��a"O���5�J�RQ�Mٲ��6Q"��W"O^��eJżh��X�'�
��1+w"O� 2�Ȱv�T�"�.�v>�#0"O����)�"������
���!"O����@�<r�m94No_ %�"Ox5�jE�B��T)dd��F��Z"O�W!�_�tMBT�H'���"O�A 2f{)�3��._��|�d�.�y�Ñ|���S��$��
p����y�ϙ\!^t�f��pw������y�C�Z���d�Y�cԬ�y2�V�m�Y 1���W��jvaʿ�yBDX�S$����B�_��<��Þ�y2�m�X!�>�a�P��yr��7u�x��Vq�^��@���y�ȞV�J6���c<����/��y�"�H��i���D�V��u�1�yrA�0^(�K��S�L7��;vE��y���'	"��C��<�D�Pl���yr��:�FW��<���3q@�3�FC�I�L�6Dx�l�b��"q�� }�XC��6wm�i�Q�X)xt�Ku��k�@C�I�u�t���N��A�(�i��FTVC��&V�a@Reט�8*扗�Vs$C�I�/?n���,QJ��C��0��C�I(����X���	���j�bC䉪\���e��_.����$Z%p�B�I)�q+g)@�R�@�k�@��C�ɯF;
����<~�,%+���5��C�Ii�����	�M
�S�$��x6�B�I�g0��0׉�_>,ٓ�.2�B�	� Ġ�Td��Y�Z��u����C�I���v�S��b,�����C�)� �y+��A�+[�i"a��S���ڷ"O����@�C�`�7{3 u�U"O.�.�4jL��Hs/M(.��Y�"O�d�ϡH=��@b�M\�؃"O�L; e@��|����pQt��7"O�iAD��#2*�E1�"��A=�PR�"OR�I�I�4L��3M3" �E"O*e��@�L�!�c�O"(�"O>@J4O��Eb�y����&r�H��"O,QP�h5@,pi�+��4�b"O��G����9B�l
�{j�� "Ojh`��
���{A�u�j��"O�ic��*X7X���.L6M"dX�"O��!����L�u�2n�"d���"O~)��&P�)W�-HL��"O�1kSF�;�]���;9[H���"O�U93�
�9 ��h�݈
%ʘ�2"O����n�}\l#��]0rԻQ"O����Ʀzf�T��^�VF(���"Om���C�X��* MAB4l�"O�8b0���D���E7^0t*@"O��`��� ^Rla!�a����;�"O`� �ҷD'����N\�{N����"Od	�6B�&9��4d)�U"O��!�� m#D	
�l?B��"O� ���<SVXp�V�X^�`�7"O��B˺r��[���,D��e"O��h��
�<t]z��H�H2+�"O��+Q��3CC�ݘ�L�9�4��"O���6��#ʕ�1AǧDz�`X�"O���6JD)��w�H�
��}�!"O>�#�Kҵ;����(ȊD��	J�"O����4)�z�<S�L �"O�aU����,R�ł7��["O&������6�Ȩde�;T�8 �"O�d'�k�H��"Mɦ��a"O���@:PJ�� �vc�	[�"O�)A�t�t�PϏ�:>��"O�q@E"X%)f��r �-S� ��"O���� J�OƤ��G�?#E�0�"Ot����V�j}�A��%"J��T"O��+�� �V�|�C�ŉ�\%��W"O@��S)���
�#
/C��hH�"Op]��	BV|�`��E搑Y�"O���4�G�h(( �G��?��<��"O���� ��'̉��H83���2`�'���s��hǇ����s!W�S��B��5m|�����1�)Hz��B�#���j�j��e��=bŠC��NB�8Z��<��J
:������/n5�ʓ�0?Yw�M`�r�r�,X0�P��"U�<Y����v�0�%� ֑#���h�<�Vh�I�(=FU��t�b�k�y�<�1���j�B}0p+�d���HB��x�<����G�\щe� �W����# �v�<����(JA2qK�3b���dh�u�<�u�M� %I��D�t���FCW�<YR������u�\���$�P�<�@,89�`;�@R�*2��DHUO�<�E'&	��0�%ғ)&E���G�<!� ��o�T�`�
%\�!���N�<	eAڑ
|ؑ�q/�1���I�<E/� ܔ��\Y'N�6`A�<�.�-pA0��#IT>�jH $��Q�<� :��V�ŗ-sf�0��X$�	��"O� �ˇ���`�3KŘ|@�"Ox�YEàT�Ԓ�c��?���I`"O�� �a�J�n ��mٞ)�����"O��ō�0 �|���K�9T�����"O��Yb���[~�4Q��:���v"O>p"U�Y�+ ��rG
�͉�"O
���ń�8��W�f̄�ha"O��9�n�o��Z�&�ik��q�"O��y�)�(�Z�z%�I3%c�� "O�LJ�o�3;��㋅ �pm��"O�Y+b��1���֪K�P��
�"O^8�)ˁC���a��F0Nr>0	"O�����$�ڲ7�ݹf"OrA�U�˽u��P� �X m��"OJ@ɂ#�Msz�8Q�^:E>�w"O��I�`ڑ@��2��U[)��j"OH�%P�nK�<Bf(H�	!�a�"�'�D]<G��N�0���@WGߑ*]!��՘2&JpG5~���wE P�!�Z#r��� "���`�X��=w�!�D1ݺ!b�^�"�Э�be�n�!��T�������"?�ۤd�6�!�$�++��	s"���`<ӴĘ@!�������E�k�@��&%H,} !�$��M���Dv��t#d��'�!�C;��	CR�/��X��� vS!�$Z>��ʗ�,%�m�F��3^ !��X`�� �f��W�̈w!�d_4"�\P6(��-��|9�%*$_!�$�FKܓ��T�z���%�C�!�$�����G�Z�(I�82�!򄜆3e�R�b��K16M��Dę!�+9Q 5����v,�t�P��5!�$-��%I KX�(��,;�!�*w�tpy��K�l4<�ؤl
�t!�\�12rQ91� `'�4# ��:\I!�V?�`�J&.�}z�U����f�!�D��C4�0Hш}Ѳ�����C�!�ĝ�W�$8 �!՜R��%�@�s�!�D�p���LQ3KM��&�!�X 5��OT_CJ8����+!��yQ���K3@1���X�XE!�T8�d�P�ɖ#P�S��
N!���sʀ'�̍#x�Jc[�0!�Y	kB�;7 �N$`�&a�n!�dF7!ń� Fa��_��X�ʱ��'����F�B�?P�A`D�;w�H��'MJ��H�k�F�0cU�?����'���$��g" �7K:���'��M���4����������y��l@t@*�K���xP�b��y�B�M���($��\���ӈ�y�ʹu�(uP�� ��\��"BX�y�| pX�T�â�-��ȏ)�yG�m,& �"L��{�R�3�B���yҊ�+v�\��C�bY�����y��_n��r7�Y�C�xM�5����y��D��0x�aKA�@!�b��y�߽�4�ih 91lEa�nO3�y2��wV�l�ժ����H1b┲�yBѵ>��I1�ڐgw2��P1�y2ٚ&��R��*e
[TB���yBƛ�
��T�W�'�� ŨҼ�y
� "D0P�\�+����a��1C�]@�"Olc� 
'�h��&�Z� E"O`��SjMg���J���c���!"Oz��$��P�J7�\<O�l�F"OX���O�VI��J���B�&�i�"Oj{T
�+N5 �6�\�Y��b"O�4���ڢd�(5*Eě�J��P�"O�աSB��XM.���1I{`�Z1"O@ف#ʈ#��P��އO��#�"O�ah䬗��Ѱ�$�z�J�"O�`�@�µu^�4�ҘA��X�C"O>T�
�N]�DDJ�6vyq"Op�c�n�*rO8<Xօ >�� "O
eC5��/z8: 1�e_�v$�4�`"O��@��Z�k����&䈱k&%PE"O��geT�$o�c�
�  �"O�퉅ύ{��aBH�n`
"O�L�ë�*��@���0^|k"O��)���A:t��L'�v���"O
����R$U���#�w��cs"O��)�%*�bĒ�2O�pu`C"O܅�'��P�r�� ێ�>hj`"OR�+`��LU@� �V�)���c"OpU���N�fi��⍄�<"ژ	�"O��V���tAg��.Cnip�"O�xŢܒl�����F� ��d��"O��̕ ��U�Af���ѓd"O�h��OMy��)%�O=d��L@�"O"���2�u���\?\}����"O���������i�M�Q`x�"O�	R��ԱS�*�+񭒂7H|�"O���fC	�
���"ǹD5�"O�C6%@�E��=���U�l�i$"O<�R�E�<1�bM� �I���ȷ"O�McX-�M�"yLl��"O�m��g�"g��;O����#"O��9c�&wD��at���"O��:�dƗD�s��G�)�[A"O�1T��$�-�U���
��`��"O~���M7=���+�#s�a"O^d��bş��آ!,H�K9�Q��"O�@"j\2zJL"�B�*,���"O� cB�]���򇪛""�f"OlT�O\/.��4g����"Ov���B�&
x^M�u� &}��mb�"O"�q%U��U���Ȳ�\��"O��pe¾�J�zSMߙ%�2Xk`"O���YR���� k� ��|c�"O��
��-|�`E�ׂPV��"O���C�ɧF��:aj�N�z9ٰ"O��&dL1*Q���ɗ�$@a
�"O6��Gf�@ 3�*$J�hk"O�I��j��g)�q�����7��S�"O
@���iƤP)��,d"OX����^5y�����(3zyʵ"O�`"��N�U��j�M�����P"O�0�&W��f��A��� ! "O��w*@^���j�t#,�"�"O��a���Gw�)k�Ð�C|���"O 49w�@�"�X4��a
�mn��h"O0Hq �	R�:��#/1��s!"O@"FN�
b�-�d�U�@G���"OX5��F��Ma�91!A,[:\�w"O�uX80�a�4��5�V&{�!�� r)�*�Xg�h˳K�����d"Or�K�а�&dHV ��t���x2"O���_	Z$�	a�ىZ��Z@"O������5���ӡ:t��(���]�<郦ѩ>Z�00��$b�2ã�b�<)7���_��܈Η�daˣg�U�<�H��0��1k�ɟ�x߶	3�m�j�<1/�*(6nQdO�z�zB�A�<a�mMeϦm�&IX�RPe�f�y�<y��G +� a!%ʱ[�l��F
j�<�(6%
�����0H�j���Eh�<��,Z^X�S�	��(8�4e@}�<�2b�7F�%!�Z��L5���{�<�h�� ��N�^6�0�BI`�<�`�J&b<0H!�G�~b��!�j�\�<i)�]U�3P�@�z0�	A�b�b�<�C�6ά!(��T	c!H�1G�u�<g �$Ijy���l�H1�"�u�<YE�R�X�f�%@9��x2�J�<���y0��13�2E�D��F�<��MD>c��P�u��$3�H`�A�<���1m�L5ȅ�p�Z$��Py�<�m��*�!�߄Ol�� ��s�<1V�^�mǌ��"�"���k@s�<��,�!��8!)�k��0�y�<y��6?|8�C���L��Q���j�<y�Aۑk J�z`��N�p�Xc�<!u��$4k�́q�ԋ9Qꍸ�`^�<�A�	D��Ѩ�He����]�<�&�Γw�0����Ɂ��q0�H�s�<1¨�=����3uo����E�<y����F�H�䒰]�rp�c�~�<1��\|������,�b|�3i�~�<�E��@��ĦкT����bPs�<���L!l��IGhT�Pမ��@�q�<)�]�b��p�8�$uQ��Y�<�R���'���ի	�g�"�ȗ"�S�<��*/,����-\�h���g�<���Lw���A��`\�hf�<1�oX�<ڶ8HD�r&0�#KV^�<��GU'�8B1��9:����*�\�<9"�M'�l��Ck�/i���K���V�<� ا1H�ٻ�%����]�a�$T��C��"�>D�gʔ�}%r��%4D�0#l�z��찰����B�H0D�QV��e �уv�������*D�`��,UB%���� ڶ4R1L'D�da��L��pH'As����#)D�,�֯f��HA��Ҕ1��*5K"D����f[�R��CaNҡXF���d!D�<�Va�#�tc�U>{�8�{'$>D���iO�ʘ�3%?���(�h(D��s���N��Ѓէ�����g&D��#�$�1�Mh4�ֺ+�ƥi�a9D���@�M1M�"XX��Աv��U؆A5D�,0����R����\���)%!D�,y`dZ�Iy^Qx��O�Q��#1�1D�h5�*_����S���@$D�0;DB�o<��iA��R�0#T-#D�D뚞�89��P1,D���@�"D���cV��\$�L`���g4D�|k��,m����iQ)&���s�2D�tC�ˁ�\�t��4m�ݳ��1D�|A��ʓN��� �?p��x��o"D�� Txْ%Es"ܜ��-��(�L8۲"O�R��߬ZȨ8!
S�ȩx�"O�}���@�lH����*���YB"O��O�
���hF��!�X�`q"Od�S�Å�W���u��>���V"O�����z�P=8��M�7
����"Oj�j2$5��5��R3��j "O�ؑ�
 �2t���癷� +0"O���G$GaV��J
�,ih"O>1�3H��A�B��v'N�4��=q"Ox,*qo�w'
=X�ֈ4�I�"O�0y�m_L^�!$%�|ux=Q�"O�y��T����65]�@�"O2i( ��3���� f.8y"O�M��K� �P� �|N9�"OnM�7D�"
� ���J�+Y|M�"O8�ˀA\=���c�O�(��Q�"O�Ha�E؀w�h����(�ƝY�"OZy)��VV�tkWI_!�D`�0"O\tS�iڨ�.�;��=�4H$"Oe��MX�*�S�e�,<B�"O��î�12���w�A�.��X��"O�<q	��g��Q�A%Y9�蝉�"O�U���!3�drU-��O����"O���w�1{��� �$�n5�$"O<�TAL�Rƨ�Ib�Yx��o&D��a��F���Y���;Z!�Y��2D�Jf+M3cB 0��˭ �R��"�0D���%C�9d����H������3D��䤛%}R<�6�P�ECޑ�V$2D�,�����[a�#�fQ�1dj�&:D��pC�|�y8G�� ^T���-8D��eW�0Ƹ$��
9]`��Щ5D�X�$a��(��1BG��+^�b��@�1D��Ȧf[�s�ĉ8N@�tF��D$D�d��C�80�(4�c31<�)c-D��H�K:���z�� (���-D�T�F�ݷU�$-�/W� 0	�M1D�$��E:q�Ȅ�!�6��ua"I.D�X; @�R�X���p�A
��)D�(�p��9�@c���H�u�'D�t�7e�)��9��k���Bɦ<Y����(��D(�e����%�%9w�Y��"O�� �"á[:�k"�T$3n�#V"O��w��Ǹd�a@7Uܘ�"Ot;�d��R$n��F���"O��*_=n�R�f"E�΅Bt"OHX�Ee��B��Ä��P�$$1G�'��'F�=�hI{b=�Ҁ�%�����'�ў"~4A �-¾mӳ�� �j2�Q��y�']1Pg�T���I|�^������y�"�t���/ABv8���ꓚ�y�ma�^����8���0c%���y���ٰ���+0qޘ�Q�@��y�IB���{b��?�F�����?a��*�@��h ����=nA:�j���xOۛ���R��p�t����߷��<���$˕(�������X���	�!��x�t�zc��2�n� ���!��ĀC����g�2������8�!�	�6-�� X�y�Q[u˟�T�!�DJ�U��)�7Bq �P�u��cx!�D��?.��C	�/2���y�(	d\!�D�� ���&��Q���!#I �!�� ڥJ��=���p��"%~�Є"O�rE+� 86 2�$Z4�"O ��n�ib��D͂5>��	D"OLD!+G�� ���/z�"�"OT#W�N��0�C��u���'�PU��O��sa
�_Iơ��⎔-]� [�'�ў"~2efB���M��+
^.�Ar�9��'yў�O��u1'F�d��s�E���q��'�(9����(BJu.!��1FN1D�@ K�WV�`VFS0V?���U//D�`M+�քP��^q*A�+D�8@�9�H�� M���q�*�O��CƜhP��o�t!Q'֕ A̈́ȓ=~���M6!�l��ʓ ���ȓQ���ط P^;��@f+�:$�I�ȓm>���4����Ԝ�P��oB|�ȓ7�2���֋/c�KՈ|W���ȓ~��أ3nN�7D���47¬���h
����f�am�X&)\|�ȓx��v-@����XsH������,h2���`
�T�H�x���4T���'�a~B�)!��i�j�2���Y���yBKB�^ib=����@��P �yR�L^�1�	0��\�aB��y�O�u����CI�2��[BD���y׌o�̉�A�~~�z����y�E�%6FD|`�b��O,A��� �hO��O�c>Q!)��&�92�HO�IBe�$D��2�.٬U��c��D�pY�WB!D��v�\�t��Dh�n��ˆI�{�<y��]��Lن�F����S�d@�<Qj
�R�����]i�i"�O`�<��IT2 64����;!H$1gMZ�<Q�صg������׾ffЈq�`y��'i��x3ϒ):2�)�+ګ
�T$����xr%�X(:�����bx����yD##by��C7�XR�$P��yB�
cd���,�
K�Lb&�M<�y�A�_��H�D�6m�x���yro`
�YCk�$_�Q-ŷ�y�#�R�T	3�H�#��l�cO��y�OW��X 7O 0űr���ȓ��퓵��1&L0�+Kh,���o¸��jʎ3:t!����b��//����-wʜPD@�Q�^I��y��ȑ�Nk�Z��0��#j#����*�x��@>�:���G�6�'������
1�vk�)�e
�/��C�I�R�b�HE���Le�S�� ]��C�	����6��,y��Pd�,��B�	�3���B�(v�����_�X+rB��Hh�$)�(�%RƄ�&,C�	�)�J����j��<�w"Y)37��$�O b�TC0H�	=����'JD�ӧ�/D�bf̓�&�\��Ҽx�p��,D�d�L�2�4hge�0�9#�o*D��b�ۛ<oR9IT��F���`�!(D�X[%�:xF�a��8^)=���9D�h��)��o!�EJbH ط�"D��)��ȍ_�$�Xv�˩*y~a���><O��$"�	<(B��5�V	r4��0�kW8u&B�I�ib�[��?ځq�i	A�B�I�P048f��m�xB�GG�4B䉭w�LC���P�l�c� B�)� �U��� ~�$k��-c��`xB"O�|Z��,t5ڤ��DB7�"���"O�C��d9��c�wVL�c�On `B�U-n&蘅b��8J�X���8D��2'X��z��t;V��G�8D�X�CPV�Rժ�4N�a��2D��H�� ��ҌC�}�҄�pI3D�P���C���1#�}t�0ڱ1D��PA���r��Jg$G���y�&$D����b��2h�����.0 r d�-4�`z �؇(R�iKö0�̄xɚٟ���lf�\�6,ڣ4�xAc��>i �ȓ|�a����{���$J�;wVꍇ��� ��/�`k剝;5�ڝK�"O��:4�̕9}ey���8ڬ�v"O@�K���
�P0a����n��@"O$%���A��n���\��y��G9�*D�2a�+bԭ�%� ��y¢մ=�XbD��u�P���G=�y�K��#���HEIW�6n��C�T$�y��ǋ6R����f��YXdآ��ߗ�y�M_�xw:lr�J	�AK6��e��y�Ύ�l�I iG:-Vv�H�bY��y�ː��=hB��zXBe�RB���y҈A���󤧘�w�})�k��y�.]�1Д�:�n؎e���"�$�y���7��pc�\$���y��X:;P�kF-@U ��rn���y"ޫ-�8���@��B��I� 	)�y���5WF���"$�3#6�#���yR�[�G���T��*��M���I�y�'Շ =zd���W�md��(�7�yb$�*%�Hi��Ê�h�G���y���-o*��D��#��]�����y2����M�*3^(�&k=�y�-M#+�����e.L���B;�y�^��}ీ�	*L�,)���y���&WW�d��hI�y�q� ��?�_�ZՊ�ɐ�h�~�J� �NA���'!p,�㈰?L���FE���q�'���I�I�#BvE3��F�C���z�'�0���Ǉm �T�d�S7����'u�T9�����	�mԸ5�bij�'҄5D�=K���-^�PI�'#�AҨ�&Z�|��Aj�/Fd�����$f�L%
�Ǌ����JL,s!��8�����	I�]�f�S�?��T��(��S��� !�*'n�J�<yB"O��'H�>eDܹ$ϝ��(�e"Oܱ��j78,�6���N��0"O��%�ɻ:iջc�ë �X�3"O�Dwß�-ӢE"S��{ru�e"O�Ij�l���cG��id�I�&"O�24*��^����o��>��T�W����x�S�O:HAb���!~R�}Y��M���
�'1�}�愕��L��3�07��yi�'�\�(��8EkJ��a��:�ƀ��'<�����M�KY�%�%V�/G�E��'~b�S�!M��*	 	f��'<�I�s�8!����[~%������O��O�">�5(-��:�痒I�<u������Ie�	o�O��:��mY���F%>���/ �!��þal��7!*6Xl�RK��u�!�d�TPQ�7�w��Q���C�!�� *�����?<"������K�䡺6"O�A��+��|``D���8 F"Oج�q-�(cx�����Nްm5Z�̕'�R�'�"��C��vVt���K�<������?a�����h���A��V�j|��b�O5|�4`�3D����H��.�12
�|fpH�&D���Ӕ)N�:�8(�����J'D���AgBrU�`��s����g-;D����-"$}���{[��Y�<D��ʇ��\8��Ξ-`���<��Wu8�#�,�P��]9#��!C�$��	��0�IEy�����W
���(T9~��`��*D�)$@�#Nᾬ�A�?n���&D���cE��ށ��a�#=���+&D���V��>�2�
�"'K�DT�8D�T*�fƆ1���a"� V ��"�;D�xrA�-]�!�J�BR���V	8D�p��B
��Z�)�#I�4ݶA�"�<����(H��#6`)$�.IH)�,�:C�I�E�n�S���DYi�{�6C���L�x0C��x4GK0}%^C�sl��0m��Q�L�4�TO0C�	�.���3���&�� �1.�BC�'{$��hS�V�2�Y��/;�HB䉢G��aA�]`���B�t�tB�I�J� ��L��DxTd٦3�B䉫C�ʵx)4�H��P��69vB�	�f�����7>�0`�!8�pB�I=
���6%�)9_��ժT9�&B�I6[��gH���c�Ҝ	��C�ɑhJj�F��˰����O�S��C䉬2^	pg-�%�<�
�ぅHB�	�.?����jV?|'�YI���WPC�	�<!^��ѨOc�8��G�RC�I�)�i��!^��;b��;PT�B�	��;��}_^]X�a��B�ɾ ��m�4/U�,�<M���4]9�B�	�L_��) +��6��0�ULE2C��C�	<,��\pM@�g��|#�+�;-"�C��##=@�+CO�o�r�*���g�C䉍7{��S �;jM|<)6��	�C�ɾO14<Ф�%�P��fT���C�	�8�.T�DA��I2p�3S`tC�I�6�j�'Y�f2�;�O�ަ�?�����Lt9T刌~�h��amg�%:R"OtycJ 3%����f�EW ��7"O�� ��*]����n�ri쀰`"O8eY�A�Vc~�k������"OxE2�$[t"�H����V��T�g"O�|DK�Q����$i���T�J4"O ��F�5"�Rsb�M(D����ӟ<�?1�O%��ƍ;�R8�Ĩ~b0�
�'��P�-�-#(��r��Ȳ((a��'��%0h@�t��%�?�nI�
�'!�]F�Ӄ3��h�#�^1j
�'���U�an]�bdK�E�r��	�'m�����7�T���A��Pn����'����F��^�u�@qHd��'���8���/{
]�-Jy�`�'�ԭ�C\-�9��픉��0P
�'�^q�3����j�U�u���':�!C�IY=b6$�$"h����'&��ە��cv��W�2Y>漑	�'�H��@�B2h�F�9�N�D~�x:	��� e����y���Ȧn�nEB0"O �i%&ϭh�ص����"O���#�<5�Qt�8  "��E"O6�{��-%���C5'ˤ(�0��"O�}�1A_�<�U@Or�&�SC"O���B�0��	�$D2�B�hr"O���� �>h�Q�i���N��"O~D�3)ݹj�NP��.�;=1FlB�"O�y�5�ũjf�AboL�	z��*T"O��q��S#V�(c�n��|wR(�d"O��3�"
l��R�ɓ6\dl��"O��!��70�y�լ�WE���u"O!��!�9h;b��+A�
�t(�"O�Prת	5|�X$ CL�> bh��"O��(���2|R8kg�D�!��a0b"O8��R���~��9ۡ���.��a�"O���b�)@p��/Y&K���ط"O��@�oD*�~x�hU-(���"O���c���mȢa�Sun�h�b"O��Z�#��1�:D;bd��q_���%"O�I%D«IyzIK!�{vnA�"Ot�nއW^��R�1Y���v"O������^żD��c�>�V�'���'���]2Nt@�D�v' 	����?�C�"<`%K-�$,�p�竟1.bC�ɲ������	e���6�ӢY�ZC�	�ph��Giʴ�X��6$W�<C�����KE<	�1ϫ[6(��'ܠ��`AO���@1�įZ����'�j���b�TE�@Jp�ܛL������?�yn���0�1F_�.t�@���y��I>Ofp%Zw��v�`AS�C�<�y� �.T�N�җ�[";ˮ�B�c�yB�'�m{�ϒ�~P��� �E�y�,(9ڨ<9��J�,.A�@@9�0?�Woʟ�P֫H<\���\�^;�Qj��Zyb�'�<$2d�/�Vd�QC@~��
��O\��񏍾hS��kؑ]x8�B��X>9�EA"E*��0a�)=���,D�P�`NK�Y"60
�סJ7�٠��0D���ƃS�j\.y�C�V�k1�=Q��/D��{��֏A7�X��ѿl�AR �+�O���n����M<;�ʙ��.!���d�O�B��q�3��X�.��0cF�_�FB��P����ۣ~d��[�bB��6Qd�S4�M+iJ���+��`!lB�	)�F��O���9[CY1:srB�	R��d�T�ڲ�*��hD \nTB�	��$�W���b�`S���4��C�	�8	�dI�Tk,@2�C�Z#&X��!Z*(�t*׫5	=j�gΘgB���ȓ6�rA��"@D ��5�+f:n����H@Z�¶u"q�u�Ǟq*��ȓi�2�uD�N���8!�L�@%"D�Tjƫފ�ֹG�T���m�lk�C�ɳ7���SA�E~�>�c�&��B�	�>�����
��x�Z���lB�����Ҳ+ֵzJ$� NR�7:B䉤Bd�|�CK˶:8�2�QO�&B�	�1XL���YQJ�s�C*&��B�<I�t�g)z�D̳���Fj�B�,.�j(@��+X&�ȃ�[	.�B�ɵde|��� I�e�J�Pd�Y�C-�B�	��z]+fU�w�z���T2p�RB�)� B��v�+F��
�#�D�w"O����`��B�@��=*h��p2"Ot������ �Lӄ��BN��Y0"O�y���4Â����@8}5���"O�=!��fH�A���H��ԡe"Oą1�Bޘa�՘��-	V��G"O�@ɐ��n����"�BH�C"O|���*Y�F�+Ĝ!U��Pp"OJ z�Eַ���Lˬ w���"O�M#D�_|��$���5�d
"OF��4d��_-X$Ч��$b �a�"O��yRNJ>)�xp�U]�$��c"O��jb���dM�(3�N.a�@�"O�L�0�^=N��� ��4O�@'"O�( w�
$̂�-�겜�*O E�w�YB\�F���z��|��'�t��/X*q6�&,_�w]Թ��'ڈ�`A;�.��uF��p��d��'�TukG.B�Zg���'N31D�L"�'���5hH�Rf�m��5v�!�'Y��	�,��eӕ�ۗ0��H�ȓ ���⯅����R2H�=�X���U��ir���0}����ÐZ�(h��TR�z`oa�����	�V��ȓs�r����>ZZ��v�]
�h@�ȓv�������2f�ԘF�
;�|�ȓ~S���V��REv� ���<�Ѝ�� ��8�hܒi�@���MH�bU���ȓpA��D�2F��#R�[,}���"]+��|���� i\�Y�|���� 	c�/�P�ģsA�_��ȓ.�(c�o|o�zA���r��b�<��Ĝ�9n�����r��+�`�\�<���kY��@q' A��ɩw��B�<d�� ]��t�Q'� �����Z~�<	��  
�j�M��h9FD���w��?���ԟ�t��n҂;���G	Q��l�F"O�����\I��(�iN:7�^9�#"O��Y��
?��  /�8l�.�`7"O.)�b <ZpA��&�H0h�"O�0��lQ=8���B�C;m����'��I៬�ffJ�2�g�
(��i�	
�E�L���J����t�.CcT�w�1j��'22�'ra|�/�R#�������+�r�˦�:�y�Q(*��۷��)y�E��y��ϻF�xc!MҬk@Jݢ��ř�y���+dh`&��w�X1;����y-4~Ht���u��9�����?I�'�~3h��e���s!!�M��q2�'���b�G�]�Y�0ɛ�ZPԕr��x��	%*{��%�dU��y�-ӗfh5��%W�M�ĳB��ȓ+:�P�Z�-�qk ���q��؅��ι�w�T��D�ध�J���ȓ�V�+�e����0 c�a�����<�0�*4q���\?sc
%�'[y�<!�ӌ+�,�K�'Ä��k�&Ory�'����@HX	�B�ƽS�����'Q��
�Ʌ}�%��[�ER؍#
�'_�l��M�b��7N
�Y]v��C"O4��WC��p�d����ԇQGp �a"On�C�@ߙp�L���OA�L �h�"O��X��U>� x����6�}(�"OjP#�-��P:�X��hF�Q%\ �"O� p��V���T,r��c�[/j�6��"O�D��V5d;fq(����B� ���"O����;_�U@ %�3V���c�"OL<ɒ凮�8�iD;g�H�V"O�4е�.U�,�RÇ�6s�Y��"O%Ћ�8R�0 ���%�a8�"O�@��mɻKl~�c��#&��A�b"Oh��F�&{I�]:�A^����"On��`D�4J��=B���}��!�"O���	�x�B�"`Ts�~5p�"OՓ���t��P�W�O�$�0�"OlI���ކ5�����L�D�V1�r"O�D�	?&҈�b"j�!�'v!�d
0���ŏU��4 �:�{����)b ��EŽX�^�P&��&y�!��Q�n�"%��#n���Òɗ	�!�D�����p$Ѵ!���Cl�!�DX(����f4��N��"�!��$ ��;���M����g\�!�DEg�] wՇ+�B]�F�w_!�DR �Nua61�~̪ ��!r[!��-Xo&�iƃ��_��x��4E�O¢=�����I^Ulhf�4^JR+R"O�	����=�R����Cn3J�0d"Otȃ�-J.`f���3VӼ5��"O�tk��ڮ,1��ACa�,o����1"OX8�1d[�,:h�xя&y6�#W"O�s�".>5J�B0�d���"O��#��<{��El��RɖT��"O�D����_txiq�9/�45(e"O�� �;�Ԥ��)�Lun��"OD��DU�x'�8�F3p�А"O��2�o�vE��i�|�|x�"O��@fa�#i,- ���ge�8�"O�Hi�dY?#]�1�,�*a*9FOJ<��M.(����*ن=�P�@j�<I-O����K�(�
r�C%q�	0c�&�!��K	o��Wx�������&�@��p950r͐>uX�iw�K7�T��K�l$���ѫ$��]�G�H�_e������	���P��-���F� ����ȓM3EA&���*.�I	��G�g��E{��O#`�j��*z(�ò��[���IO>����0=	c�B3 '<P�&�Ha<-��N�<�r(ڦ�p|�sn�
16��¶��L�<�4OR)�<	i"LK<y*�2��FC�<ifFƃ34:UZ��/�����j�<ѵl�S?���`[�j�$-h�Q`�<)��ۚ{�@8��GY 	���\�'�IP�<�����X�*�h�9��	� �65�ȓ0e���׫,]+����ƗE�����si�0��˒; Q�qq�@���ȓ+{TA� L+`���$�]h,`u�ȓ)�x�q �P��-a'/.Aly��750��$ʢu *���
 2n����ȓR�L�{���
�2Ԩ*n
���u�L�Zy{sI�9M��d�FުO����Gb((b�א*�ZD�D!�LȓP�� �t�ܹ&��g�z��ȓ~�jM�ADŢw%�iQc抮Q�N��ȓS�q�P��(\�Z���"2 �ȓ�����'?T���lR�Z�6m��t�v�ʲ��t�IQ� ٧0ߴUF��I�@y�Q��F*i�M���͸x���?��S�? �|�r��	3�Eh�@�Pfr��"OIB%���^ h1����F��H�G"O\H��M�^�9���K�@�=��"O0���.��F���0��O�l���h�"O8�P��)����C%lg��1�"O�I��{�<��R
�9^bģ�O0��'�<t���ar��vj�(���#�d5�OTp���əW0XUr
Ł8(�d8"O)k�e*q
�ma�+��-(��"O�;��ɘ!c�R&�ȿe�x� "O|�{@��0Rw��z����\����"O�@��?�xջe�*u�&�#�d=LO@�p���\�ӗ/G;R2�y`g�|��)��C�dA����"`�ٹ�c�4r���D9�O���u(,�	W�P�,6����B�M�B�"O8 �h�$�48�<R���C�/$Y��Bg˾!�t�F�I�B�ɔhB���`e��-���s����K�,B�	�hf�BC@��>>�$����^� B䉟g��t�*�:�z�����4v�ʓ�hOQ>M�fm0#ģ>#,��b�*D���2��.ݎuKP�Ĭs�Q�A�2D�t�� Z
H�Q���r7�A���/D�`ڴ^9c��h
�K^�I��B"D�(�hDN�Q�dڟ �R���i!D��"���:n�F��ů�lX�FI>D��S�EeV2�2�+G�0ii��<i�����O��d��Ko,��F��>���3b�I�<e�O���Ć%"�3�[�{�����9rq!���/{�m�SC���%�Vm��fG!�/s��(9qC�	z��EYm��q!�������H��G�"1�F�U!��ش8�1ǚ���f�.|�!�$���x���m��}�v�����'��'�?��)�r�
�	wN@�qGX�J��;��/�O�H��ÿ78���W�_������I}�O�P��AH[�uO��"�9 �Ir
�'+^|�5��m�D}S�!�!@��T2
�'Q.�{����Z�
�¾.�p	�'#��e�,x<�Y��M �0/�<��'LF��W�V�D�2y��_�����$�O#~J'�H�9�h�(e���'�
�����x����b��F	*���@T�W�nq+Ɗ)D�<X�E��
w�8"GCѿ\Nv|�s%D��J�!L�/�t8`��;f�4����=D� 
�]0 ɧ��hT2��0�<D�0A5�v��A���/�����,D�(�D� Y���Kͫ��5���)D� �"*�0Y챻����.%Cf�%D�Pc�^'qM����n����{��-D��# ����!�wI�*bu2A�&I0D�T"�@L�����r�X?�)��e-D��(Q �QP��.�i��MA�-D�|��o��R �M�B��$�,`I�I�<1�"�>���M L:�9���O>�<��d���b� / �f��G�F0aV�0�?�ӓf�`l�H_� �� �6�9��L��P��,H�%�:Ձ�MԭkaP1�ȓ;����g�=:؈���B�CrB�ȓ]ͺK�D�'E�i���
OZ���>$ `�t��N�Ly�uK�m�a�ȓr��<y����,��\E���m��BG�f<:e:�@Ù8�DT8�"Ox�`�O �:(�⳯G�"M�鸧"O� ~m5� �r��GB�;׈5�"O����7施�a��1E���6"O����͛&:qb蝮a�T(С"O��kɹ6$�����ּ;��h��"O���s)��=�<�g�x�z8Y"O�\�p����Qu'�S�"Mx�O��Ǐ�(.���;��6>&��?ړ�0|�#�ý>�2��ER-�Л�L�_�<�5!��="挘ĭ�X_�L� @�Q�<	!��7V?h�XPM��j�ܳ�� x�<�V��x�"��S���m*���t@w�<1��N����U��,L���k'��G�<�gO3"����s���By��E_�<	���"zμ:A S%բ,87o�u�<!E�MY��1�)#pܬc̋G�<�Ӫ �"���#��z���R (SY�<� ��)&�����8-[��TW�<����E7�9�ׯȭ,����@S�<��`�.N� D�#�3R��.�y�<�Q�Ț,@�K2�$'\��Ss�<��	MF�D��^$5Cc,�p�<	�
L�X�k7��yve�`E�l�<�"�d��u�a��F.�}2��i�<�pd!p��-�`�;���FM_a�<��ˈ�2F��(��:<�����]�<�3�L6_( ���=eT>�s-�U�<��g^�y�����K�i��dO�<1��X�h^Z(����/&��q�mPV�<1���c��г$X�����P�<9��100>�E'��#�ay��K�<i��̪i$d�bn�0�))d�~�<It��@�z,ze��.Wv��"��u�<�W�E�'^�X쒗��p��l�<��T�����3!~��S��L�<1����T��i^;�*%�D�<�gL M�%�օ�����d�[�<�n�妔Ô`��f�F��3��S�<aC�S��`�SL���qi�U�<�ABD�ԩrS���:����u�<92@�<�\�����r�d�p�<A�`ԭ?V���g+e�LQ$�g�<Q��'h<���U���A�\���M�<a���zZ��H�"�6e���R
�_�<��l�|�H���(��"����7
�w�<a�)C6�!h@k���I�Cq�<�������lS�u4�Ec��T�<i�
#:ʅ8�\�t�]1#mN�<aR��qQ\2$AB�3��sP%�P�<y���k��D(ĭ��7�<�@�^B�<!3�_2@����C�4�� +wfX@�<A&h��)��r!e�����ۇ$�z�<a�b.�$`����3�Q%�AN�<��k�=���jv!C`Gf���Q�<��b;D��Tq���!G�]��O�<�"�	a��pw��.����o�L�<QW�אn/%q��� Y��T	��Mb�<M8��(=d��� �fJa�<���E�U��A�ѿf�X����\t�<�6l�j�m��:D����m�<قe�	����W��^�Щ3a�m�<��G�:�	�ʖ�9�z���g�<I/!wi�t�tFL��	�\�<9�Dίo��c�ò��Q�DZ�<�C 
�Wk:%
6K\nb���S$�@�<� �հ�V2@�:E���H+\�I��"O���s��c���Ip�A�h�颂"OF{����o���h4ÚMJ�m	"OµA�k�O$~yq7X,��A"O�hR��u:xqh�2Cu
��C"OP��!Ϙ;�|��7�@�*�D$@�"O4�A��D�<����^�\�C�"O��aD��*�	��N����݊�*O�!���ջ[m�����1���'���賈щ`��� �g���k�'/����a��m��P�@�;#��J	�'`�qA#V
6��%ys��5� 9	�'5����G.��j��\%�q��'�l���N�3+M���I��,`0B�'t�]Ӂ�ƅ5�Aÿ>�4�s�"D�����1�
\;���@�I�7�!D�4�ݹ�R�0�H|x�K��!D�H*�Ґ%�h0�p(HB�^sd�>D�(*g��9�9C�@D�xz���¬"D�,�R�F�cS$�sS�B(���s�"D����R�(�1���'=tL9�j+T�����\"`��m	6�ޙl(�t�g"O|1*���2h=�V�;,�X "O�4{�-7=W�i8��� xl��"O�E�bhɂN#�ب��M�pY�"OLi���ؗy�8����5�^�""Ov�Ia�ӵ(��P�g'�7�>�kb"OL���Nٰ�.}��&�vlR"O�(�R'�/1�\�8�%� e�"Oac��>K�~�"�1�x�Z4"O |6A�|�܄�B�/��Ԉ�"O�\ pb�O�Ƀ����%�XQ�5"O$�b���;�F�*cA��ؗ"O��G�v���SR�_{��R"O���q46ʤY��&�zx��"O�%�����"�>a���Հ9֮Њ�"O�͠TE�FI)�bՌ(�L��"O: ��g��E(�[����9��D�B"OL�	���>
1z�A�e֋4���{ "O&Z�#Z�.ƌl �D��<Y��"OV�#�LQ�7���lˊi�r���"O�Y��"eB���;���S"O��j���kM���e�96�@q1�"O@�g��Yr�%+*�4M5���"O�%�D���o�I����b��"O�y�4�غZ��Th�o��SR"O���F ߀#�t����W;��Cg"O`1�@E�C��F�Md5�`"F"Ol��#O5U��D�"���<v2)�"Oՙ�-ٌq:��5�R2O����"O�e�����E�A�>)�"O��!�-�.�X\��랴v����E"O��Gd�t�j�W�zdMч"OV���dI�G�������|�@���"Oje�	ͶB��K���$"OVy�JE�;���q��?|���ځ"OuU�M"%�2��à�͂�Ps"O��"�Z�T�j���p�:"OHt�!��0 ����6U�l�ɲ"O�I���ѝt�}(�Be���:�"Oȡ�!�tܲEO��k�T��"Oшc%H=^��<9bm��{��@h�"O�]Jp���
��f�ě&�@��2"O�U��%���x@����+H�ZD�""O� D��&�S�Z̲m��`V�*@P��"O���J!QTr��o�'^2JRR"O��&��KW�/�a��"O�ݸ ��D�С����(�`|�"O�XQ����������Ii$�i�"Oڴ�gVR`$i����o���0"O2]� (�6U	��ె�VUr�0"O@�a'X��vq�&Oԑj7T)�2"O�e��KY�DfD%��A+��"O���O�~�fYq�MO).y���F"O6��!���Dڈ́�l��k��C�"O"eX2�Ӥ$����`ک-v"as�"O���SM��x���?p]�ԛ�"O�)`�O	Y�V�g��^>��"O̴F�ˈH褜v��
4A`�&"O|D)V�Z�=1��A7+�"N)��r�"O� ���n��l�6F'��h�<QŠ��P�+1�K���p��n�|�<���U^� � ڭp���D�d�<��N]�T�^(�IJ)O)�<�`f�a�<�1�&z0dq�Ќ�J���C�_�<qŁ��&4���-X�;�(���^�<�b *.���EŚcTd�j��W�<��m�h���D�±/;�D�k�O�<�!(����W�l|�5A�[�a8JB��&}nd��g�]]����х��c 2B�	��B�y���$A��2��C�"�2����^�j�Ɛ�W���+o�C�Ƀ9趱b"��0Q��vkA�S�C��eɲ �g	VD�tr4Ӫ6tC�I���X��S�&�N�k��BYdC�4[IX�brDԇbf��%h(�$C�	"cRB!��0I��8�,��
�B�I�#�b���0�"�FH׃8��B��!����ݠo��ȓ�9��B��8p��Æ9U�h����B䉐V2Yi^&(p4�%!دKTnB�	#�=KB��-8T$c1�W8�C䉞m��YY�
O�|�(P�v+V�Y�>C�I"*�\*1��%\�h[��m�C�I�d F���3�@�~(FU�*O���% "*�$��G� t�:q[�"O ���k%i��Y���c�T8s"O�U��@^��ʩ0�K�@~ֱ0�"Ozb��G���pHA�p<�5"O¨�⥓`�UZ�N*0����C"O��し�R`81c��&m�h�F"OP(:�P�
J(����*S.�"O��*�fDZ��18ċ�$�q9�"O��f�0���	�##e�"OhLWe��OF�-
�핮
 Q"O��v�+3`@�Єbڠ�;�"O؀�S&��?<�����Z tL�0"O���_O�Dِ[-g
�	pQ"O"��##�0{����/\>+a(���"ON=�VE�V4|�*�XB���"O�}b��X>x�#
�D]Li�"O�b!0���`$�Ɗ,?ָ�#"O��i��ܧM���y�C3�Y�"O `��#Nl��N^8*f�rD"Ot�� *wԺ�1�	:�y�G"O�K����F�������R��+"O�1�DK�?w��.M�!���ْ"O(�X$�ô�^�.Ya�lqܼ�!�� �ar$%�4*ic��H>Ot�$S�"OT�p�
R�@��,�g�M(���3"O��:�DH��^�B�,����"O�! ��c�t��M�<ެ��"O^䀒�Z 3�T�[��I�-���"O��'��+h�L 5c'V��9����g�����v���i�\�
���T�$9�O�P�a'F�>���`�]�b`��"O�!��, �sJҮ�.q*�O`�dB<?xABwcC&<���5՘xx!�ĉ����f^�IWx-��n�+V����ƭ��u����%��+v~t���:��j��%A$Xf���u������Vڪi���TE������|�Y��X��-R��T�����	�

��j�S�b%h!LU�s$$C�I&k0Ҁ���:�v�Q��T�\C���젲WZ&������7=���'��(ɗD�
Wk���0fӒ5�$��'�����؏7�*�Y	/�ޝ�'{VP����!a{jTR�ϊ.�D%8
�'�2=�P|�4p%A	*"����"D�X��$I,�$�1��<*���e�!D����Qv���w�Y����pr��>�,O&�I"����]��`����E�ʑ`���� b�C��*'t"�A+�&<N�j�,��oJ��&� F�D�&uJ� �F�&3'R�R��"�0=1H�8��6�HD�TE~�uU�_5��\FzR�'&�5�2d		�;��%��$����3�J�xM�D���+����Cx1���8�j�.QS��{�NQB��-̓��	x���L<��r��� V�H7X�-ƂA��\�'
�1)1FO,n:�9qf��rT��4�yB�/�O�qb�)�"*�}�l����m���'��O��w�P0�@90��(M�(���"O�|Ze�D�K���cɊ8cR��`��O(�"~Γ l�	t� ����"�� =��)��>���s�IyX�EȽ[��ȓ;Ǧ  'ED�&�x�IB��8�<��������_�����a�Z��@���	Y<�i�jV�x0>�*���h�y�ȓR{R]�E�b����[�dɇ�G���x�CYB�Y��-|D2e�ȓ!q���4E�W�J2QZ����_��ㄋ\IҐ��yN	�ȓk�Zlj�%P*������<V"���$��ţG�ɤ@� d�EHйE�t���k�b�p�o��(k��Sf��3P*��ȓ)qt8�ǁТ!t�m;���F*���hO?��d]�jϮ�1��ݗs���)5D�DP�.�.���sD������E2D��
K*x2FB��.�$zQ2,O��<��l�%>�l�(P�P�ĸP�`@f�<ɦiT,g�(��#�D:�e��k}�<!�+B�*p��H�LAFE���MX���	˟,�ɭ�t��������Б,�>1�6�L$��'�ў���D��N76�%
�F�!���#�"O
�x��D�Qx<��6d6��	Q�"O�m�4���z�BPPԂI�b��]@r"O�0i�EY���-��A�����#"O�� �#��a�X����C�*$�`"ODA� e�y�PЫv!�5)|��"Od|idP@���AE�&���
�U��r�O����<U�X��G���:�� �J�bG!�� X�S���bZ��:�Δ*"��E�s"O��ht�YN���wǋ/�ޅ�1��g���S'I�`��C��\����20i0B�7
�vDr��͊~�]+��y�"B�	:a��ȃR�p��)S��y� b�D{J|�0��-N� ��T��4W�z�c_��~2�'�X��#D�[����~4L��'1�0�t�ʘW�⸑��h��A��'o���yf��;���ML�	6�فט'<��$"��I;;s5K�L(Tzd}iAm���!��EV�`�"�`=>(G��!�D���+��C:)4�i�F�1Vq!��/X���qƃ-1`�� J�n�B�I9����ς�= d��� z�C䉫
mp
��N+b>�9�@-O�nC�	!<��x�%�����i�1l��b�8��	(;�j�He��7t�������JшB�I�q��s�J�2L6�����	�pB�	�+�����;F0j1���S��B�	ez�F���Xx,]�"�N<D��B�I�+f��5�P+Vb
�.��f�D��)��<٠��K�2́$��#��M�P�W�<	�'�Q<�a�ȑ'��T��V~ާ���R9%�Z,��ٵ�э�y�-�j�������(ގ��UN̴�ybH+d���e�r� UJD�߰>O�0@VE�5g�8�-ا[�@���!D���"+�2	x@�s�Q̔y �=D��Y�KѤ�\5��K��q��P0G�<D��k��åۦɉ�ğ��t(	 ��n���)�<��'����E"8�[iX�Fhd��럂kj���^�=-�q$ߗ jՐ�k��=��O��=��4��Ĵ&�����ϕ;���i��'O��(O��"G+Ð��F�V�>=�#=��YR��ʷʊ:E���ʱ���݅�2�xR�GI�fj�� )L<.��m����?�Wn2#Ota�r�צOׄC�^:�yR��-�� Agb�Wz�P�
 E�C��#��Ҥ�Y�W|��#�0K$"<IS-O�8����>���n/��m�L���"O��!�O8��B�J�,Y�"OJh3�
�h��dVn�o�,�c"O�$2��>�V�ڣ��g�~xk�"OL!���$L���ˍ?Q���[�0�e�	f�'nLD���>-�<��Ul�8�T�8�'̘��E�yy����y��`B�O��=E��N�a�(�烞�j��J���'-��S����4	�� (c#KN;h�q!+�
�yb�O6�"~�T���J�$���!�4A ���o�<�7`�0WŐ��p��:_6��;��h��<��!�.MK�ِx�2�{�ܝ��	�<�@�M�NI��"�hkc�\0��x�!�<.xL���K�H�L��b�+��O|E���I�|����6A�,D/��q�
�7`71O*�=�O���L�A���iRa��nֹ�5ˏ �!�ę�-�}�`[a/�\JE��q`!�d��W�F�"�$S]6�dD�ZU!�dF;z)������ ]�	��I2h�	hy�S� '�Е'Y@8"��nd [�f�
�'�d�I��sW٢�EP^�܂�'��u�W隃|	��Y��\Fk�U��')I����<_�XYD�O�T �*O�����a�4��wJ@�A�����J""Cay�剹Y\��C�(܈L%�	�eQ~AxB�)� ��Ba���,�f�r5�E*2�����"O�8oB9���� ��<|��R�
9D����h_�v&Y�����[N�4��a8D��+��_3M����,P�R*�M��5D�P!%�Rd�QG�/`��#�D2D��B��GvҠ#��,S�la�*D���Ğr�ld30�J�$��T�d*D�0Ӳ����-��z7ʝ`�,D�d#��3'����NуL}�y�GM*D�LX�ʉ4��m�6�M�C�Vг+$D��xw�D//�*���2\D<<j��6D�Dqa��%f�����G��2"0
��&D��Ň����k%��E9����"D���Ѥ̑@����R% ��فC(#D���	?lg��Ze���A�
5D�ܚ7��U3��  `��}.j���A D��#a��O*����8w,(ӡN?D��+/]�h�9h;8����� D����G@<�Sq�8>�}���+D���L��mn^�;���	�|)p�	'D�`��^�$�p
�!V�f_H�K�% D�Lr7aU�u�b����^Iv"��(=D�H��}L�J�Μ3X��p�%D��9i�}�Ӄ��-Y��R��!D�Pp��\$6�1[䢅 |p
x�$�)D��LZ�22��[%��UB$QG5D�`z `�.���3�g��[8�b�(D��Sa���n�h(�,�/\�>lC	&D�@��U�D����@�Z���I"D�$�@����rq�Ѣ%eNIz�
 T��B#�H�^tĈX bT�t��@Z�"O&(`��>X��w�|�lu A"O�=*��@�t  cӋ7�L�u"O� PC��Jt�pC���(g�ġ�"O~]�1% 0c
�Ӎ��h�Y*�"O� �s狴{�L����L_� c"O��C4a��?���*#L�0��xa"O���r�W�
�.��'+�"H#࠹�"O�Ds�l�1kD8X�J��z����@�X$˶�'�l�#
%��#��۞J�\|�
�'�~��"V�=�}(4��	��8�
�'
"��Zz+�d��̪7���'��=x��߳b�d�ƋW	zq�<�	�'��0�ꏙ %b&�>c��	�'���@ C�27F0�5�P1����'v����Ly���B�s�@}
�' �t�&M�=K:iò坖[�Ы�'�<���Ǉ�Hq�ʑ*]oNS�'�@�g�ћbw�䐱�� 'ZH��'� �����Le�!x�B�gϰ��'/��c!ƶC��� E ��V����']j�6�����!�m\BW���'�f�;��z�pu�䆃�?����'^I���X.e����%�K(��'���U.���t���L��p���
�'�h���6~Ҙ��$��0 Y+�'�Bx�L&�VP���չ��H�'�D:�jM�d�S"���4��'`�V�)Hϖ��q	/d��8�@�0D�X�e�P.�2����,s��`�D.�I9o`8P2�O��y:M׳J��!�a,�92�@T	C�ܧb�p9��
=p�	ѫ��}����8�x��c����>r���)�f�3d�H<qu����O P�)HPp+�	-\��P�V�'U�`�[�'�p=�gI�ir�d���f�̙c���������Άx]��A6o��'�x���π ��E/ș8��AU!&B�m
�I�,�B�BF��3�,Yh%H�u���'?G�I"k���1��^�m�1���%`����H�,}��m9�3���m�� �U�Κ"�@��'�VA��M�F���q�с+Z�ıC�.ؤ�|r��Z�4��!{��7��`���
Y�H�r��U icQ�-�O��*�#�$wv��b䆈�j|ho�.F6<YBw�H0,A`���I�"��	S$tp�$��D��jH ��Oڬ��L���W���!��}���'��$�)��2#�,c���5I�TA�h�:f1 �C(R�u��TJ��MY1#��(�beo���?���[���s��ˋ�{yh���$B����نU�����|��W��4�'Ǉ�U8)�dI(�y@��O�<X	�cE���S�N���DC#hB�5XDH�'�ꐡᨋ����#��D��K�NY���8I`�Ʌf@�0�bh�������M�p8��%'(��!��K��?���:.e �D!e��`c�&�HJ&�S�VEN 
։J65"t� $��ا+��$? ��l=�Yv�,n���c�H��c��`\r��!ڬ:md#|�%���D�Z����q�ZB��Ș�`�'lE�a��O���F5�2y'>7��x�4�ɽ+��5��ϗ�䂼���߸_ڼ�Ul��_�f�z��:xM,\̦�u��+풤���?�2� �||�}�!��(��|q�N$d�l�PFGߥ�T��X��U�x�p�;&ˢ,S�h��	X�Y$�����P1�pLϜm����A%Y�t`i��L������vH߬P�9GA4�X%��,�i����Q3�?ͻA�$���*"E�����Aa�4 ċ�:j�t
��[;N���C�"���j�"D������U�d�$8�˂�F7�{
܅E���k!��1�0S�H3�K�#O�����	�i�-�I�V�6�Tl�h���'+����>Y�P��ϛ!{yx��BGK8h��UKD�$��=�G�F(x����4|�`���6A���PE�= H�Q��Z4�jh��f��� �肠ŘgI���F6+m恑p�A	+J��<�7�B<-�v�	�h�2d�8;��Z�.=��)�c� �� {��sƨ�b��1�)2�H�01`�[�,Z1/>����_���#���[��pu���# ����U�3My嘍U�.�V3<�T��g?B�� l�
f��YCU�O�a�'�ڲ#���v.�4A�4��O܅|�S��ːm��e#�i�,:��u�'��1%���fN|�m��'�] U�ލ~��]�b��/$���X��7�^��I�ȇ-!
��ځ�[=S@���7��)�|�rr@����S�䟏]����ĊغW'h�r�$:���E*-H���+E"����q�#:Y�R��Q,p�"����9���XH`az����$^Y	3Q�CϺ����V�Er,
�"T�6��PԬ�^EzM*t��!*Lai�Q@ȴ��䖝X��[ �?@���*-v#�� 
8�?Y �B���2�B�Y�3?9�"ϝ[��H�Ζv�v��I]�g���JB#�h�0gl֢;���� fۯ/�,�`�n��p�r	�]<	m�ͪ
C�#�l��g[��0�L�h+*�:V_y���p��s�<��T� ق��5R	���9�b)�"��q�%�S�^�,��햑r+�P1n��?_�QK`�O9�x1yGBOw����4$���;�P��.��;�u"�%����U��Ove��,S-��q0�-�S8m�Ö�"9��J�D�2�Væ�)JV� ��]��oF2*�p� ��r�AR�Y�<�z@s�K7r�f���1��,��)��P�Rt��i�,(�6嘒���^�� (�H�7z�����R�/FX]��HT�F\�g�ˮ,�"��2�ՕY��8@5��s�B���Y0���À@IνO>ԃ@�AJȱw4�[���b#`��y�R���g��0�8���4�E��O�Zw,�i���%���:� ^{�\��'�*�`2(��7 ��u���fpX/�.��л�G�Ye|�F~"���xvt9d&:X`�B3Kޕr�v�y�@1*��1�ϒDX�aQgl�F��	��O�V�0q�%_v�x�YD+��2-��%��S�( F�T���3K��D��b4ғ��1J�!e��ɚ�d���@%��y�ʲ,E9/������0X�F!�� .�X���ȋ�jD������<A���>Hʘ��4��+�"�Pw����G��Q�2u��ŝ"��|��9A�	�	T�I��ʪB����7�h�
7Kݟ_Q��q�-�yBG�
�td�QKQ��x�@�B�4w`�����Ψ!��%	�"XxcF
�vd�aˌ�R��X���y��	�p��ӡ�J�����&���>��FY�1�!�D��X�́2<u�LU%ۘx�S�-�O�$��H2~���V��%�*p��ɛEpa�OЛ!Ӯ�ВĔ��Y��ǈr��AfE��_{�$�d��6�Ԉ �O��Y����OPصI����<_N���W�Gq�M��'����B��A�0��ʝ+��0S�)�.%���|:�bQ���Hҡ�H:���Ϭ2(D�'�p<��C�ؘϘ'Zʉ�0@���A5j�0.���ܩ		�Yx0ȟV�
�;�A����T��+ӱi���3aQ�n� �JE�*Jt����-gv�x�n�S��{r�я�6`��B�-�x�y�-�"��P�'J-8�*Q�"ۼ��QBɑ:|���-�`��mێ'��i݉���XTZ<��l�Ym8<ۆ$�c"THQq��m�v��P��t�`�D�*]7f����������Aʱ�E#V�.x4Qq	*}�P�i1�ONy��!��O�@��*�?m�p�� ���-֌+���G`�>y&H\l�ttt�?	�Q�#� b��A�F�FE���; [:�����4ݐ}!��3Q�8ݠ���+�j���#�T S��R/�����K�'g^ r�
Y�Ղ5OY�7���ֆ�R꼠ɵ�.\����N[-ibT4REJ�[���E�Y>3�͒�D R�~��p�=����A��!�&�pSmƪ��	�SN LOF��Fc�:�@��t#�s=�Q���3i#l(�#m��L=pKg���4�:Ӷ�G�?ՋS&���;Id<}:�4�M�֪�*C�8�Kѝg0�p��g�T�O�t��'[��y�+��c� ����{p�����D�E�8��o�	?D�/htŃ�+ͦWT��5��4^���/־{��dn�� ��7����^���
3�Ԕr7������=0o�/�ڠ�� ]���IHގ(�� MccLe3`N�o����0��z
�X9FF��ZL pCX#b�r�����Q��dx�oK 6�=6j�k|�#�̏A���P�C��`��'���@�#�#[��å�HK�pӆg�.T�!�P�L�6S�����jwF��b��U��p#�M@�)�>�xyf��14hM!����Gl��T���SB�חž��!�Q��T�.�q���X�!�U��꟒{IN�҂�9� � p�DZ^ �6�Y`�6��C�i�X3Q�� �h)�,\%4|XU`��7&� �;X��<k��WUb��t�Ҙ�lБT�z�ʆ�ٓ�M[��Z�D�
�[S� -K���7줱adآ'���ؑް�$�s��s�BL�FZ��`��֌?M��(�G
8p#��x�E��e�z���Dʍ�M7�ě��(�1,֮w��d�)�D�!L�^r�����  n���A�LĜ��oӦ	z�dLP#�-�d	�����y�#[�A�$a��$h� �aG�6]�mkЦB�:��l�� ��u�7�K5l	�Lp'��O�y�O������)��X�iP6��[��A=18`JP
�*%�*�p��I�U���c���Δ"�i�Q5��K =16Lz0��+'�&�p剎[�\�V��6��0G'K>��|�%K����Ζ~!8屰��n�\�iF���D��"�)ؐ�m֚("���ço؆�b��
G�t�ْ�.fb8p�&mI�a�ք8�-��*��¥j՜�
v?OLl3r$�)^����ǆ�e��@��d�	��V60��AS�X�0�(0p!�	�R�lm#s�ߛ2��{3)cӢ)Q�hD�E�E�f�J�!�$�VΙ%)�Z���Phξ +�
�k�E�2�E[y���*ML���'�\e���ǓT��W�f��񡱌T�k2hu��1mDd=#V�\��Zq�O��j��;<���p-B09�WJ�:�ԡ��jW�1N,�	$a��p<A�ƪY[�����Kpp2�c6w��LLb��  4.5��)�:H�}�\p7�� EbLBvÓ�	x�`�T	H�DKV
��Ⱀ��#��^bjpՁ#h#�UGx"�5i�MI婆d������E�R`æ��Wl�(�k�#--f ӡ��>м=�5P�R��5��B�3Ϊ\����Xd
�0��O,b0���J�;��I�w��)c��\�p�1��Vu@"qbw���"� �E)FW�~�hg�R%s��;"�
_�v��'tC*mB�m�\A\b�@.�E�o��)Z�W�$ "!�F`�qY��&��"�p<FeR |y���*�='�<PİbQ*�7Gg���GI��NV%��~~���> v�"���[u���=�q��叱 �9"�
Cm8���H�*�F�`���HF�13�����kr���hT�焔�7���1k�> �2�;��ƥ|NJ�a������;"lS���Ԅά9�^yYs �
Q	���NC)Q��Ē���Srh�9�*KX��g�p^�b��b�|����@8O0]��%Pv�r�׎����D5I�Y
��G�~�SΟ@2�Ҩ:zT1bԻ�8��O],8bň�O_��#Ŷi��5�-����@cS�d��p)�K��[xȪAk�?;&�9V��ם�r��i�@ˊ�|W������%�	���X��OH�!�s���Ӵ}T	��ԟ	�d0u���cCM�P}�݊3�\(5�1+�뎸3���9ՇX,:�ʅ2��0t��T�Q~�ђ\)2�kw�<l����OQ!90X���'�SM��󶈈19��scU�||M	���=n�qO��R®^7D7�<�Վ����!����;(���#��J3_�xtaЯ	aF���
Y871�����	��f�8.��S,k��QW�Q��l 4�N�W0콁0f�v�}D{�D�%���FT�~e0��v牾AGz�p#�� a
h�e/�mC��[�d�0��4b& �4\�P ��$�~����3 ��ҟ5�EA�%}�qJdN�RM��ab�M�I�SH���"\Z�x"����@� ]Ke�K� �����DsXT ��B�6<�����V���)��a�*C�-Ol1)!ʄ��D� Q�]!«HR#r��2:��%�FV$i뮽zD�	�U�T0��ސj�pY��کB��!�İ9��-��4��jX	`y���*��ߪ9�#�˯������(L�!�088���_�X8��*4�hO\�QAY=�`y
��S�K!\Pa(��ո�Mץ�2͂D���V	��؏>�hq
Y7�:�P��8��ރWWp�cJU=M1(0��NC�g��@%eWP�'uH����Ƅ%~�}h���yn\ԃ�M�S骝��l�9�E�g��>,�ִ"5�[_�ޡ�]&��I��q���b&���(�#S�2���:`HŜ&O��򨛖g��O����[�e�9�H�)�X�!R�I>%��II�'��-�'�Q��+֏G$V,ƐÕ叱7w�pUI2d�|\Z�B̹\W�<+��P�S��V�ƦS и��3�M�!��� S�*%�̍n�u��G��0@�ޫPq����mP�%Y���QDX�U��z��M�j�u)bY�H���@�דU5ȵ�e�zFP��M���S+�H���B�/��4ʂ�ݮ#�~b�dp�k��zJ�CR��'A��X���ˎKь�wdѽ�?i�/-�ܸč	"zI�=)��Rӟ� �0'Q�l�°�7�Wb�R�iʑ|E�f�L{QqO�D+'�<+���ͱU�|l�[�p#Ћ�*m�t@qCҜ^P�/��������::�)p�7d��S�k�hxa#�W
h{FoJ6��pJ���:�r(!�bFtm�GS���q`܅tF�9�%��7�� ��N����@	�'� ����ҐBd\8��+�_���XX�kU�ô)mN�`K \���(`��9Q�&X��f� �������Cj�+hD6�]�^��A2!�>➙��B��̝��^�V�4�3.Y�L%|-1��8X��ir�a
�;ꆕ�DbW�޹����Vа��t��"��=�Ӂ��Q��Pe-�=M��!�@�2>��Hh�WҶ��<A5Ȏ�S��(����/-��V0GU!_ ����@�]�pe9��A]�
(|t���TM��*$!��r7��瀆\�~�q��)k/�-�c�x�P��1��S�`�����V�R�n��fB�:{ �臫���`�)E� �8�F�B�259,cK�r����,)".;#��e����a�� 8�@��������Y2�~"@ΐ?YJYJO
�f�ʨ	D�J>q�\��yVd(k���=X�4�	�)�<=��F3Bf���e^�A%�؉2��' �(�R���Q^D��c�P�x	�u��Ҍ ��8���.>S9��P��|�^�#�<�#��I�NRl���՗&��Qc�R==�8�T Ą|�HiIB��4'�2��	M@D�n�Լ[b� &F0�"d��M�VdXse�$�
�'���Ѐ�
����y��J�tC^9��BH�_�Ds�ME�"z�<��f�`%��H�U��#����"IS�t+!mD<!|�0ʯOX�h�Ǔ7>�`wfQ�p.0+�fG�w�~8��$
zP�N��t0�����X�nLB!Xߜ=J�p6�+gAL���͉��ȱ��b��ZV�ԋ��O�����^���x�#T�9p��	 2O\��%jN�a4\����؛(�)���j����=z��q�B����.Ȑɣ��Te)p���'�V'���3L�|؟���)�9=o)��Ê��Ii��?�\������o2�x1����ཀྵ#�D;8g�6����}@K��S%FZ��:�L �2�r���&�O��c"C�(4i��p1 �.:~(�0�C�m��q�	���gÌG�.D��K]7��� � Y�8{"�($ϣ?���{��,�td�����q#��X�@9F|b/T���#TcUr%d�$�����d��,0Af,׬`|�3�mR�;�H{��`�f�Z��F�F�4��[w�Q�� � �$9kJ<Hi�%�����q��O�Us��J(���h��O>S��OZD����X#t���LJ
- �'�)_1(��6��)<�n���p?A�)U�0�Ȩ�ꚉY���jWdX-&�Va��W�J��5M� �j9�jBIk�0)�M�,]�F�Rv�YcRő7�� a�4W�0u��n5�OХ��ʢ^I
�q&-#VH��"+j����d�d�P� �ė%c<���]?\L �i4�s���3[��b�ڭB��R^���O�d1G�ٶi�f aH|J�0dv*�0�o&D,lp����F��6�����$脎kт��hOn}�QGIt��M"�I!S���Д>�TH:C����өh�ne(�
�?�D�Z��#B-�������k���1O�*g�<��I3
���YP@I>U�u�)��=!��>ftA��ГMVp��L�Ŭ��}���2���t;�"OVԠ�
B����CT��i��Z�'�$x*�.��G�L}j�
j?E��jW�����(Ւ�B 4�� �!��[V�ntj�$GK��0aB�ǂ
ɼ�O*Y��$I�,,��O���2":+6H��)U*�� V�'<�]�f�U�ĉ��`�0 S�P���"���C5
�H<����ʾ졇��
�`1ZP�J�'
 뒧^J�'[a�ݠ`�g@�h iC!H_
���1T�uV/תF�Ү4?� �ȓN�(���'�c��Rl���zu��c��i � ��Jܑ��垎e&�e�ȓ2*���e+E�O��i:�bC�����ȓx��C�x�H�ɂmǸU}�i�ȓ"`�L�U!��OHLA�	�4!Fi�ȓ �{���Eb$�@&#Rt
х�Ӏ\��	� <�l4�#�3b8�ćȓkB*u;��͵p<E����4=�fP�ȓ.���h��ݐr�E(��Ʋh	�5�����g��$F�r�Ɍ�C�� ��T
�qW0 ξ��$�ֶ�8��Npl���&�|��\t�N�^8<��6ШK�ǅ�`uh&�R�`��@�ȓ����'�n�{�l�)F3|�ȓ$U��B-E$,����K'9�����V����℈G4��[71�P��`�*��\�"�NY�#%!�8��C r+�h�'? ��MυUV�@��0�V����чA�&���*�T��nN���U�Y�܅D���C|�ȓY�\Hs�f��bh�x�J�6�U�ȓ1|HS��[h����Cz	�ȓh���iސA�j���#E�N?v�ȓ��,���VPR�킛�����B
T��!��U��]zCO(��	�ȓir�H�[� � �@2@)��g�zPk��U.`�	%���P&���:x��3s��\�����>>����Y�A#|ju٧HG�^H�ȅ�pQ��
�"1Ć�!2�� �����1G҈�ׄ�;���G烻�ȓ?�`�	�"0p��Ă6���ȓu���q�)�$#��\kC(\�C�T|��k*���q�I�c���5�ȓ~��� B�6���c�T���ȓ���c��)-|�P��_�ɇ�V���d��W�0T2S
[����g���Q!nځ3�M�F�\���+ظ�Ã� �P9�H��x%��_�-�D��ZY�u���xK̈́�}�	!�bK�*9��֑x����iFڈ�"#�씭�U`%;"O�œ  ��^-��H�3U�.1��"OVli�t:@�B���Vj�$"O�8j�U	V:� ��Ɯ�x���ƿl��	�	�g�? 61�Gbb�U���J?��P1bÑ3z�I)6�'�x�c�,	�[��0b��y� �K!�87ΐ�'�I�R>�R�OE�bv��6Q��C!�P`��튒���s�� �O�<)�N�$Ct���N�/��x� c�(p)t�� *��!�ۏXf,B�@t�	�'>q�n�k!Z�O���+D�2X4ܓ��	�Z�M����>��{3aL����'�eY���k'�kʚ\Q|�IA����|��PԲ𢂋-�3��܂w�Y�3��OҠ�n\1hV��n�=	t�ŉ�cɛWKĭk�-J��6�|J��� h�X��?�1fH�r( �x��� �O�M*ƊH�8�dE��I��g��L�a�_&f��$����K��uIvΖ<󩈓;�bq���`��x���O���@^'e�h�b�f̣[�K��'�h�[P,�:�9�&�T"���qh��T٩-J�h�Xi@Bˌ�Va�T�|ڶ���*U��?�����S����#ĥMyM~��ѣ�7)��XӋ�B]�'(��p��J�GW�0�W�ƌ0@ �K	4��d�ߤ��%���ݡ"KК*[�=�q��Y@N��)����Oޠ�dC���ͥO�����$W����rLN{C�	˴��:Jɀm"�/�+��,��ݳJኼ��L9��ӺC��ұ�:ūu˚��4s�䀅R�8-#Q
R?_�������UMP -O~=��Cj�SXX�}�pl̩i�B�֑K��5e]�δ�v�@�b�x=餁1�'M���4Q�``R�]"0�j@7�9�����~�@�W�1P(�iX �A�&��	� 䈍6�����,p^řG��B�G�F�m V�+����2�) Iv8�a�\�#j���O�X1A� ��2E�q�8� 
��.� y`�ɉ`��阣�<��!A# -�q�v�g)ڬʴK J�'`X�3����,�Ԙ�B�Q��9Vrj��bn�A�hDD�`\���V	(�ưZ�/F�@�;:x@�#���T�D�@0�$�#�<[��Q@�j�P�H���3>~H�3����%n�F� T#��M�c��F�ّ�(����T�Z�X�A@T!��l�l�XP�!eȤ�O�B�D�Ae��򉈿`�01��"RIljٚ�N�K8��;F�S*(]�T�ׯl��\��CH>c�>-�;H8��e��=[:�����Z��+�9~�YaG.��?Ct�0E��!�§ޔu�e��䁅[�s���֍N�&L)�kW+:��褀*OX��Ԍ$i|��� �H���ԥ�I�"�	&V�>������eG�&d��8A�+Ԟbx�sF�#�@!�QDͬPj�Ը�f�9Qk���O�<�s���J�ig��P��HkZy�_KD�*�����  Q�A��,�p�U�U�S:��K�P0�rK�_H^�2�# (���@�?�c��� �y����/�	��\+o�7��$2�X٧��`�z�{�-��GQ
�*{W�="��V�S��a#ĠP&r>�uS��d���ÀcN�k0�sW�5p�i�O	�=��V��v4"��b򆨓c�8i2�S�������=u=�a��[9']����n*r�w�[�Ѯ�CR�$����f�r3�AY1M�:!P�Hj�/� ~jh�D���7�NI�uʙ?Zh�<�W!��?q�iԕ]����%�ȡ�3?�5�H�~h����'f�]�@U�YGz�i
�lp�M
�a�gNչ%dV�x��vg�$c�E3֠U]Ml�1�Jl�Y:��NνBFdV�=�Xi�呧'� ���\k8� ru��C����G��0KV�ٳM�_��=h�(�=vZh2�$�>�z��E�Z�S�XE����4@Pعs�)Z��(u�O"���݂I*�����(C��(B�c�'�M9DN@�d��i-�� �z<yÊ�M3���j���4HD�y�Pq�Q��v`�,�v���N�T���Է�.M�'3>!r!&�.P�zX��O ��aZ .~aB҈0e���ߴ!0F\K����jO�uB���\�R�Y��6#NԒ��&k�ġ�/�#6�1z���y�=ڵ�R�Jsp�;���S�Lk@͛#��O@��]83�H�����-
Ǽ�zRŠ;�̥cs-E�l��ɚ L˫&�P4ʃ˜91�D��Fj��ʤ�*¼��Ģ���K���+C��HT/+I��ד1�
	Cg��G�ޱa!&�'@�X�c*9#���@�@ܘmbqd��8�ʁ���7
ș)���&B�T���\x�I�>dRq��_~>��k%��#=�f�6��a�v�F;�E��(Rn���9��ɾ~T��&N6b��m�ƈ���������\e�p(�k�����HV~	�Sn��ht�:��S����ʮCr�I ���"S��`��cT����t��D��bEj�'k8D�0�)F�Ya��v$0� F�
z@B䉤KD�e�a�}��H:6̚E��� �S6�9v@�4a��S�l�I@�%Sc�]P3�I�5ʒ��)ȸa{��A:~ڰ��DX� �@��d�%�Ji��l�3V�P�b�!��K�DQ!�U�o�6!K�kժ��?9�hE�|墈@��'R�"�C���k�'�����mXT�T�ӄ}��hU(Q�"H#��V��NAY�d��}A5b ?��hI>B�>�b?�B�b�9�������H�q��뿟ȹ�OΎ\�H�p�/^�\-I�h
k������Ʌ�X����dTb�~��-��X��M��H�O��1�c>c����h�WL��"P;e��iQ�(8�̙YE`$
��SF
PZ�� �cJۦ�"e�9a�� �؎^�p�Ap�O�d���;A&�0_���I�g��xG���n�"4�E24]X�:�ɒu����/ADV8{�e��`�� I7jA, �j�*\w��xAE��֝�L~�I�J���!��CJТ?���+Ib���KU8 #$�7�ŨcFA)n��Re���h�܍8e�y�bƻ)\����7=��5�m�"�� �� �^�F]�[��R�4&۠�0�2�� Q�'2���E��^%��Z�үM
E1��lR���P7S����E��(�% ^NeŎ�̟D��N[�	�ud�7R���Dz@��|j@����G%	��W�H"
��f��j`� ���~z��PR�ͬ~nJ���j$	�,����%�����hhЀk���QP�d�6P������	����@�'�`��D�p�>�iT��f���Z�c�VE(�I�R�C�9F��)��RL&�qW�RD�$�;}���޴�McgKR��Zi��A˷\�.a�Ǝ#$�h�O,e���Y��y��է�L��Ml�*�(�$�@�21�Q� �PyK�'E2��Q�Uk��)�!P�T�yD��
�妁��be�Xe-��,���闬R�X6� �k󨞌;��`�
���!q��7��V��3Vy�b?-1:F�z���0��/����ѣqg
��eŢ�\QR���D��5�'��	^TR4�.�$ �	4h {���5�����{����X��,�oz�ڕ� K73���5�8�T��g��
�&x�Q��_���3����̙��K�5<���e(�/[<x���ǅ�}\�UC�3�f��uÆ(}V��O�Ȱ��F�S��o˴im��S&X�`�xÊ߆�r��R  �C�����XѦ�㰣.^���6q��$kb��
3n����v�G�]$3ʞ�1e/�0:ɰ��&ؒ�hye�^3��7�~��s� �,���+F�3`p�uї덱!>��7��-�,ʢU=(ኃE��D%��$��m>*%���=V�4��
�"|I�AH1�� P1>7�ʟ$R�/��/�\�:����i��KҤ���M�8����S�ڀ�Ω�M���Mk���>rQ�����eSEE��s"~��ǐ�5��	��WR{",��LωaR�s���%p�0�4%���QL��uHp0��#?�"��� �� W_��Pь 	iϠ�Gb<+�r0 eE�����lڭr#�����FWY��H��A�oΠ�j����)�z,0uE�z�e)�N\,y���E�U�C�4�9�g_���F�}���N�+ĥ��q�x�R��>��+� 
�"S�A��l�)R�O��D�dc�e�3�"hЖ� Q�j���ʴ#R�	�i�:���<i����Vj��'fx�!��_86����P.��"�fV$��+��B1Pa�S'd|�1�K�	�#�3W�t�3�ߜs�Bj��&�+�i�;G8��	�n#VPQҡ�py��T�
\�'ۊ� B@5B,�`c�e��R����I�!fis�"�%[a�π/jٌ��O�88��_ \ѼQ1��LBh�s +�^���bТ�1?Ͷ��d���p<A�*��2'�[��<�% Q"�)��_j�"T3aHѱdT�-@�"�">��i�&Ib�
1�,�7�^�;'S<*�0m�bP��B�JӍH��{a�45��t���r�'�>�z�T$�h�g��mc� �R�bDE���,tV�� ���-z88�j�'�	~�Bw�j���㒭v��`A��uT���Ƭx?(�:pW��e���%���a䀒U��Ճ#IˡX#d8⎍�C:�U�^�;��8��� ���Q����|���Z.xp؅��DQN����ь<�X���Yд�a$�T8�ɀ�C%[q�xrC	�t��,C���k�^�3�hԴw1��p�̌����T;�HQCwc�u��$S�H�l�L�{�8O���7d��!WT�iq�x[7I��p>	��]�vr�2w홳T6�I8�h�		��u��)�:(sCZ ���� �/���{�c 2V0�Q (����Q�b��<8�)Z�&>�l����C$�p��#W��>�{�(�
c��)�1��.M�b��J�Ƅhv	�A^�ڴgŘp,��breT<4��u�*�,LxP�ǂܯ'UD�K��'�P����?�2J�e�<��Bv�e��gO;LQ��BƠ;GB���n��仢�Ǩ(V�0�I+�d੤	�<.�|���a�Cr��ʑ�g�A�;W�tK�C�0�AGS�lq� ��l�~\ȗ�ƿ�?A�펤?
�<�Od��.\'��L��]���hdb�v��`w��<��䣅�@+��1���u��c!��_�����w��xG������5��@<�c�I�r"Ƚ�g 	��,�� ��2=��wB
y��àbUE"��d[�t&�@�萊A��yi��:�9`���k��@��Za�*�3a`��n	�ƈ�	D��iA�O�� 1]?�O��8I�����	��r��M�U�T,� �t�'�d%��+�1�Ƙ;�nԽN"5�ʔ�y_�Ea&�֌����R��P�����a�~�Q�:9�>�.��C�F�Ww�����|BЁV-YY"�P(){�d%�\2So�)-r�H9���% bm��Q'4������Rq�E1,l��rU��$f��U" NZ4�@8�R戨S��ER�J�%�m[�OMR��L��Q�<9H�{ޅ��3�����i�D���	�)D��Q`SI����,�Υ:��G�	[ ]�8�S�(�0x�*Ⱥ&A��R�`tpO����!���.o~�q5j���-"Ќ��}�:����,i��E�gLA�&��d&_�5a���fO_�� �9��͇e�(�F٭l��m�7���&��@@���~�7HBE�HaP[t����b��!�>�DoT�w�d����QT"�pc2�je����N�nP�KV)YJ*�%W���V�S<ޮ��ǋ���U������W.>S��0K�iV$�0Bk4W�4]C���A�V��&��ä@�R�Eb��!��Mk��4�,xB�J���y"�&�X�5�&;�����Q'�jT��
�6X��E�̀8Xy
,'�@��\'8���1�Х�x|��4[�������xP�蓗�٢2�0��e�
�y]��7�˿z@�b�NB�X������}Z����$�"1�8���iK�6bF0A�(W��*P(2,p۴ ���Ғ�K\�ə� dԐ ,<�I4'�@��㞯g"���J҂]dD ��(@';3������2��F�~�X��S���T����)�?q�n9��P�^6��s���`�f�{KǓVp��E��ɫ9����a�_"!h(���:Z>�L��J@��tc���j/��a�^��@� �ƲP����b�36�E�'�r [��ۻj"��#�5�
�k�(�0zk&m;��)}+Fm`q�<��m�3e��X5�D�q�� ��L��Mc�,��"��1�@U^� �Z���̋�	1>����4������ �K�=�4���
Jb@,�����ē�I�<����tf�¦�B��Ӝ'&̙���e�bY(C%�.!1&�҂��;�|Yc�I�4V��*rc�".رҳ�7d�v}p�%��%9:�ˡ@���`[w��o"��ֈ�:��:@�̶t �� �j���ہ �-��'���� Y�9 ���bA�},%�$mԔ[n޸�Cb�9K,Xc�g��I�N]���
<,�����q:�TM�?��"Кjx������e
��F-����!�V���1�0�H�Ua�1�N�3s*�UQ��8s�\�>AU$�{٦�
4���L�POd��G"U��e����]�2)��V~Һ0JE���;B�P��+�"#m����� ga���\)��?his#�ңp�ph�%@�6�rԻ�A�6D 5�ʉ�r�`9h��҈Uf:�u���2.�49�Lփ�,�x5�[� u8�R��|�f�W<9pB�j��I�δ��`��hkf�ˣ�����aLʘ	ήĩƆ־=xL�B�*	Ʀ���J޼���4�����P�j[� B�M�P��'Բ��bF���y�<�,X��k�����O�<���#W�>9���]��	4�\ܦQ�Ãh4
�-;��p�>I�m��O�S�m�,\��af�5qk�P��� �ɘ�< d�5_�T�cb��o�ܔ�Xcو�h`,J9@�a��)Sl�(���ì�`!�E"��!�bE��џ��Α�?�Ԥٷ懍@raYv�b�p�#�M�xgd�`�`�a/8�(�NQ�>�����C
fQ1�"�	D�i�����d�6�	BP��*�+Gj)z1@�D�V�#tFHr��ЇڣF�$�U;Abh\a���
w�*DA�A�L�{�CLt�P� @��{�? d��Q*ȹ#j�k2���[��-QP�'��<����W6���pE��,�ɞ05�|U3�㚽J�Y�.��%��{#�W�b:����� � 
�ٟ���+i14��CE�{V�%�a��
�`#>q��7{�����K8G4d��a�R�|TIU;U�aPBGR�x1Z� n�C�T�sU�!~0�ۧ#��ֈ��ըO(E�ѡ�E���S�>=hi�W�O<!RhD����� ˓�S� �O'\��Á��x�>q�!��t��cD��9Q�h�x���y}�!'�;�p?��+q����	LjD�Ы��߲:���Lb�@Z���[vgS���C�A��$Մ��'i]>�y�g�(	�IZէ����ds��Eް?���σFT�)�$��E�\��A���ȉ��ZJ�|�� �6v%�I��J�9;�=�dk<Ÿ�y��+|ZeB"K[�P���k�4��O�x�iI�l�F�:K|�Q���ST� k�E�aޤ��FFv�7�J�e(��
���{�z����hO��PV���5���]�،���>)�C�.����ӮnhLQ���,�*�.C�(?�A6�ӪK'�@(��/P�6Ѕ�I�;���+K�/(f!�S�+ς�=fc�`�����[K���,iDB�^5pd�R듀O&Qȇ"O*�Q��ԿX�
�@%
�(wE�(q�'�H�lЍW���Rg�I?E��(�	FN�d�EF̔�t0;���O!�"pw����m�ax���Gޔ
��E���)"蒞{W ��O��Aa��G�
����&`�����'���f��.���b��G ��"厊�Y�Z�"
j<yw��OLr�8u/K�k�X�"p�l�'�<9�uÔ}�'j�y���	�6���ْk�n*���/����􀈅C�D��a��SiP܅�\!��Tj�7?��p�ĖE/ ��Uhz]V	Q 2%raק�$<�訇ȓT�p�ӭ**H��û%�D�ȓ""A�eC�%����`ƍ3dՆ�c0�8���3f4 `d�u��,��yVZD�,!�	P��
�d?:�ȓ+ �;�w�>Y��IN>O;���ȓnϮ�Y��SQ$9�W@W4Vgjx�ȓLT�a��V�{q�T 4h'�Ԅ�>��!kV\ ϰU��,����X�ȓuŎI����O�L�'�c�����h��b��
�:HKs��P���0��DJ�B�>wՌ��Ù!zBt���c�W��z� �GB�6�>��ȓ¸��'��h,A��6.ेȓhe���,ɰ)*�/X�1�jy�ȓmc~��;����~MN!��;�FXhVSx��T`��Q�\c5�ȓS�r�%-�Db���
�r��ȓU��]��,�Q���4�F�y�<i#a���� �&!t�o�<��
�hNXIiR*բM�ܕ��CTk�<� '	3*u��z��# Y��0��e�<a�
ȪU	t�X!e��Şp�!h��A���"e��M�'S�<0A�I��	�\�c�@�q��Y�d�1G����{��� �R�)ڧ?Ra q��W����ϕ<Q�|@�!��.3^O�?!���(k�ftڴ�Q�d;�y#��~��v�x�*Z>�+K=*���x��.9�2�Ӗ���'s�a�]X>ɸ2�V�j�% M,bE�1���)}$ Xň�k��4��I2,H��v��.YFT,��!��B�IO����!bP�e��	�C��`�pgmY�|���D�O�zB�ɼ<�F��5������f(�'}�B�-���ӄЪ2�hV��Y_C��4Fw@t�c�G�c���@� �7�C�I�>�np	�HU¦!���V��HC�	�=���0� /$c^T
R+��T�PC�I�}f���
]����0�XB�Idt�*�'�"b� 0�
/&>B�I�*��c�ȷf�xp�.G���"O����Պ;ҥÑE�6��Ab"O� ����O'���r�bMn�{t"O�hR�Nʹ$�\��/�y3���u"O�4���	�EЪ�1@��'3Of��""O^%� Ŋ+t�<�#��[�h�cb"OXe�G�j��G�H�$p�)��"O0����g,��G��<�S"ON5P�[�|��H��&�7)]�9��"OFŐC�H&^��aD��J�}ѕ"Ov�0��� bV��!1I�50"O���FO2n��̨� ��cNy��"OX5���dx���S@�7~����"O2���]]�88�&@Ԓ)i(E{ "O`	��O6v���.VE���* "OX���J��T�Ұi�F��{;����"O���7iY<{�����hO���"O���KI>����p���x����"O$��'a¥"��@u�*�E97"O* �%���0��y�A��M��=y�"O���E4jhz���'�vak�"O&�[�]$(^N�:c���*�� C"ON順�&ZA4�S�eS=O����"O�P��Ö>�u� d�)SS��ɢ"Ona���f��3e��SN��k�"O�l�=�
`:@e�I2�9��"O�`2pjّtG�A�A���	�"O��`.�z�TX:3 W�[��"O�� 
��i�,c�.��k�0zR"O�U��f�,�钓�о?v,T� "O*��d�<̮�i����Jd��u"O�A��s�<3"���p:*䡠"O���O����dύ0$t�B"O��a�T?.kB��%M}�(�"O�ȡ�`�4:b=�s�E4|@� �"O|1��h�5��\;���^��LP3"O���fۥuxB��i�;e�X��"O*�����MH͙�J{�
83�"O$0�'��
J=�&��O�V=(d"O�)p��YQ�^���ߟv���h�"O�D����j
�u)փ� �6��!"O�УG�ۜ�b�{	p�����"O���C	�A�{BKW(}콣E"O�8�a���L��l����8_b��"O0��E��6Lp	� 4a����"O����mP%t�>l�ר��A�N�.d!���9)����	��2�%���&�!�݁ 4L�母z�*%���^�!��;2��\J��Q�l�R��Y�!� �2���ROm]���JR��!�+L��4b��[�Qp��?�!�K\?�,�U/[�k^li�#�"X!�$X�K�\�AF>S[�m�S)+5+!�ſR}Z�Ô���01ԜE��h!!�d٨yy�rCKV-R�v Ѓìg�!�]�N��s"�8��� ��<;!��֌v	 �yC�����Jw��1\!� ! Dd��ĸE��;��ڪB?!��Zp !#�:Ɉ\ctl�&�!�d� J��Y���0�5FC�X�!�d�, y���C7D�p�e�@�!�ȥi�B��P��\I���5�R���G:,x���RN��	��� ���ȓH^(ȴ�B�f@��2ꇩo��Մ�onH�J���n���!J�(Hb���g=��bI	�LHy�%;��!��S�? |����R�����Y,�@"O��T�n�ZHu�?w�N��q"O��P��ǲ+_�H��m̆�.��D"O�t���̂/
���K 6g�Yb`"Or�P"L�[%P���RdRX��"Ov\
�	�����c�*w��+�"O� X'�)\m�&��9���"Oॺ�'�{�2A���='�AQ�"O���s�4�U�^�A�� [��yb�M^|lď_�<�A[���y"�O!9>hT��U#5�xS�i���yr��o=�=¤bZ�4�TYq����y"��jN~U�0H%)D.���B5�yrI����A$ět���;`���y�M�@�@m�#C�j-r]�Ë��y�N�^�$б%���hlE��MK��yB��5b���e��b	����W�yBB�$C�Vx�G��t{��7�y­�8F��k�,��z��'f@'�y���w4�y�U�	q���,��y�ɍ[�$���$A+y�L���ݜ�yR�Z(V�I[D��e�T�$�	�y�H�^�<��K�_���5�yBB���XZF +>���/��yBM�4'z�Q�/ӽ��`��̖��y2 �"G�̂��v;j���C���y�,I��<�W�Ri8T�+��yB B RNt82�3w��$�� 6�y�"(Z��s �ˤf�JZU��;�y2iQ�$[�*rl�ih�ӑ���y�#�	�NqH\,0JR���o.�yR�/H:���ץ�'f��ڸ�y)�4'��hc�3`
,(�@eN��y2�ˏ|�d�%��U�8\�G@^��y2��$y�t�����7U@8e����	�y�	g�����*�E��e��.�y�L�#0��(O?C1>܁t��y"h� n�
y81ㅫ/Z�|��c��yB,
!.��q���/��H�"��y�/�*Rve`D���8��]��G��yR���¬5�K%dB^I�g/�yR��@��l�_����p���y�b�hٰ���$�h�a=�y���'�J� �� ��p���_��yH�K^$����.ٸ��$�y�PP�ib2�@�шM�p��'{f��^8�64q���=@I�'|�� f( � ��eç�Î1*,��'����!�+�3'�[�0�<E{�'M�@�Q��Ɯ���eʃ5Ut`k�'= c�׍J�
2C�+^� a�' �4��@Y�l��0YwfW���i8�'�X�B�9l�!�f*r�� b�'�<��k��ێ�c$� �V��'�^aa'��}���6�D�
�'D�y ��N�9 &���z:�1
�'=F��'K�(��i�E�T&D�$(�'$���-M��*�Ӡ���P
�'�
�z@F�EYt�2t�n��'�p�G�3M�A��ʂ��ΰ3�'�	�#g�X	��@AW7ʉb
�'ߠmJe�:J����b¸��'Ղ!y�*�]�T�9Vc1Sf$u1�'�Q���ٸ2v4鐠I��D
���  X`BP/)�]P�JZ�"Xj�"O8�S@�.$Q�R�)5\8�0"O!� ���p��ʒ/6��Q��"O��cWl�"��8(�*D�]���B�"OP���Q+P#���o̠�����"O$]2Ϋ�X$(T�[��s"O�X
2�P����!����Yp ���"O�,�AB�?-}�,�����"OR��篗9�0)�Dj�� ��Q��"O2�B��y$d4�%�Ko�L`��"O\ȅ�U-5z5j���<Z���"O�i�fF�5p)8w��K2>��p"OF���.�Ѐ��Ԕ?%>J�"O��EJ�b{�c"�ޠ`��'"O4�#���M�$��)$+�"OJ�Ģ�(<)"xJ����i"��+�"O������=Y��٫�fW����"O��è�
n�T�&��5��B�"O��Xfĝ�n$�;a-
`\�p�r"OD19���ڠ#�!�(2_��t"Ov���)Q�|� "K�>}A�0p�"OL��0�Q6=R\1���9�����"O6�
�l�90���& _5e����6"O R�ϐ)[��BЈ�78���i�"O������YYBH:��T�\�6��V"O�qS� {x���ƈ�^�dR�"O.qb�Bj�� S���gm99v"O�X��i��Y�|�*�.<V��a�"OxZ�� �G���pq��t/�哐"OXԹ����Ps�D��o��}�G"Oܘ�S��&0��Q�v�Z��"O��N��ͮ@�cdF<'ef�P�"O�	A���1�҅�QD3��L�"O�i�gōLVf�*#�
)�zB�"O�A�6k^"M��h��A�����"O����'(��A�?�R�"O$��bˇ�k������#(f���"O�p��-6� @��ās覑�"O��3�k[(	e�����:�F��"OF�	T���o0,�Tl;
���z�"O���8��gkN�-�ld��"O��"RE��,�P�1��L��"Ojlr�>� 	��NV}x+2"O"��._8��K&[�ܕP��Ҕ�y�Ү9w���4kU �h��f�y�g�>i�9�엛��Q+bL[��yB����Y!�@���a���p5\C��Ό���eL�5rTL��	
/+dC�I5k1.@�ׁ�'����~���u /D�i��	%^*�Q���Y��0��7D��8�&�H��l���d�+�J)D�Ԡ��=rQ��X4�ǦDx6�g&D�Ċ$*C.,�ERvBǘ�ʨ DL"D�8��fƈN�Tx�pI�H��X��?D��:Ǉ\�^4@���
�(�PՎ=D��*�+���}�b�Á2(��*O�i3Ť��Q���С�2
�1P"OD��D)'�� �I� F���"O�)	����a8L�6	�
3f�yD"O0���K�h@%i��,�,��"O���!�6�
4�A�P(�ɥ"O���0��������"��"O�����Y��w��#u�DCa�5D��02e��QD8��8��}(��%D�� ������bG���w�l:��#�"O$���A�v�R!{���Q��pY�"OX�0�M�]�snT�`��ْ"O�����&u��� ��Q�����"O��;���K����L#(\2T��"O���I6R���X[�k�r�p�"O�*7��]�����lK O*�q�"Ohm#�$�j��+T�#�l�E"O^aj$%ֶ[r*�bE�J6I�V"O6erD ���yA7��)%:m�6"O�I���!�@�Y�r2m"O.���)�]�,�⤀U2IF�"O^��1   ��   
  �    �  �+  �7  �C  SO  �Z  5f  �p  �x  Y�  ��  �  ^�  ��  ��  =�  �  ֺ  G�  ��  ��  R�  ��  ,�  y�  ��  ��  ��  h � � �" - a8 �F R Z T` �f yi  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^r�Bэ]lr"����Υc���!� �u�e|���ȓ_�}�㧟���\a�R�i��p��>�
H�?Дk ��t�Tلȓ*��5�&5y�d q%G�=QG>ĄȓGq�E@ÀVV�p`!��[�H�h���s�`HqH�Y�T}���ńi��=	�G$D��@1ib���eG�6�,�r�o�0��I�&��p�W� =O�AH�� ,P����D֪���8"s���G
�oºap� *}�C�IYW@	Pd]b��10#_� ��C�)� R"0)R�o"\�"e���v�X��"O��� ��)" u�g��w01��D|���On"�q�Z"f����m�,v�M��'�n9Z�HVYڢШw��)�8���'EИ�Ei�
G��Q�L��Z���'}�ݹ��f�i�6�F(]枅�ݴ�PxBjTWNX�Q꒘L�L�yV���=9���P}r�'[:��ƌ&)�D��h�X�� �'#I&�;#*��iYd�&ъ��Mh�OaV�������W���hc�!
�'�0��L�Hz1G��o2&R,Od�=E���N�T|v�8��?q����bI,�y� �+v�.m֦dVA���8�O��󄏊�j���]�,�̭���M*ޡ�/sj�=z�A��2oB}s��>��}�ƓJ�L�@&O!5ʀ�3�μx���G"=OС�~�q��5+�L\k�,� 0�~�q�'�z�<�U�2PI��|�\��s�v?���)�'^���k#��_3���d�ђD'�����%�Y4hD]��E�g�@���>�4 3Ч��!��0�f�y�!6D�<B�	A+�XE� AUj��R��)D�Pе�	)���q�Ɇ�`L�IC�'D�����R��$�� �h���bB�$D���-���|�⃌�b�t��&D��[���� ��Y�5	��3ru��`$D�7�=%o\�B���I9 x�@�7D��
�.�ag�� 2��7n6�r �4D��$Q�>�0�*�y<0l��0D��I�G�yPz�1�� }�q��-D���m�����c��L2�9I%,D�3�
_�	&h�;B��G��w�0�?���&��iz���k�Jł�jU�V��ن�	
�R�'2�,��@.@�[d�P��:8�%c1�	쟬��	�b�끤C�g�T�4��a���'�,��~��$��`%kƄ9�P��&G�y�N
�3��e��2/���p@����'ba{�k��A�	�rUB&9�B��"O��2WfΠ+5h%)�%��-���IQ"O��jt���B��3� ''��#"ODIkֆѬ|7����od��AT~��'0��'$�-hT��$$����H��E{���G[��c2�\�h�$���!G��y�N��v�����g�	P�6yPP D��'��'B����c)��ib���aǩ�4izԯ7$����`Q��{%i�jR^����ï�yB �
c�H����
�3j��c�U��yBo��*تőVj_<tD�ʳfL��yrB	�������
w�n���
��<���$݂���r��	�� A�']�}|!�W�R��T��f�"c����_/��(�=�
�ZB 5iej�&y�B�'��MR
�'���Z��C�Kj�[g�a$��
�'J�q	�M4/�.���E=B,�
�'C���j�F:�e�+¨�M�	�'j������_<��J�g�P�`!	�'�*@H̓B銰y��ׄB&���'��8QAhF�mƤ��$*��m;���'Ɏ����^�,s($���k�"�8�'%��M�{��ikr��<�N��'گ�yr!T����K�1�������p=��}bFШW��H�p��&����"�%�yB*Շg�T(V��T�6[��A+�y2ǐ�=y
\����P��!'�M!�y
� ��"��5���ZV�27�����"O��WM�*t�C�G@?D���s"O��9��K�U)����"+4+�"OH)&Ƀ�&)�5H���w"��*�"O����H�k��&JT�Ce,q�"OJ�لJ�{W2�[$ʇa�̐��"Oj)J�-^;kh�Z��X�M
��"O��醌�:z�� �k�g�6�Ȕ"O:�9XX�5��cD���ŞA[!�ĕV@��V��fp0�J�B@!�4=R��^�-D�x����*��t�	�'E̼�W�'>��1ꧩ��h�0
�'�����0��y��O�m7V]2	�'��m�Ԩ�,����(c�	�'��Y@A�'M*(���E1��H�'����	ӈM�b�2Ϗ���:�'g�|
錷E����&�1]��Q
�'=�Mj�,٠Q���ek�%@� �Y	�'���!e����u#�K��4H
�'^ls�#]4Iz<�ŭ��1}(�		�'�H)��H�7W���U��$���s�'^h`��l I�XH�	C�D�B`��.�S��?qRd�D���[���>n�H�!c!e�<�R��$)T�k%/�6UHlp�o��<�	�.�@�/I�c�v<S㋉�#�L��	妍n�
�M��O��H��(kV�3օV-5�R	��"O<�)aJȨK,���م$��ɰ��d�O�ɐ�{���)�p.B	2vh�4!J5¥CB��y�ھ&S
�xU狍L�R�@E�-�y��[:�c,	=��	�����y���G�����6��	����y��Q.F�4)����0 �]Hs.ݖ�y� CR[���m�%�n�:d���y�GڷL��,8�e�1HQTAЃCT��yR�8E�q��D�ZAI�X;�yBݛ �`�"4L��<�[�d��yB I/�� @THMNxv���'�y�eV�� 3'U�I#���˕��y��V�acn�0gh�HmH�����0�yG^Cr�(�v��ʚ\YQ�̎�y��X)+��H>\"c�3*C�I�)rL�j�!�?Ԁz2��/>��B䉋bR@��k�?N�^y ��Y7,3�B�I�4��!���
UK:�;�/V��B�	Q��b2�Ѧx2䠋UfJ�}�B�I.y�f ��%���+OI� ��C�I�=�������<�� i�B�k��B�	�_�l�3�A�1�f� 4n��B䉛G��	�&֦����EQ:��C�<��l8�*5`ܤ��$ⁿ�C�	>p��\I�.��F�pQ�^8�C�	���a�ˉ�Zo&�0"iֆ?cBB�I�{ɾ����I�k\̩E�	oyB�	+n�2�)�bۣ��́���:#�RC䉎V�쉲aQ�"��h�Ti�`C�I�/;z�Sv���	Vڔ��.υ`8lC�	�0ΨA3�
Q�cn��+��
��@C�I$�4����DL���#`<C��5�"��2�S�b��)h�c��JC�Ɋ� b�I��2󰝩0��DC�	4+� |r��ԡi�ͩDj�-
�C�I��D�\�YC�V�h:�
0D��)Ǧ� ��ɘ0�ǌP؈D���(D�d�Q�ܘT<���C��G�ȍ*�B9D�� čY��*.�vI��`���!"O���z�~�P�F犑9�"OV�� "6�lMx"�t�:��6"Oѐp��)D���D��i���"O��k5
��l}�)�ƃ��*�N�b�'�2�'Q��'	r�'b�'��'�=����\�xA�p֪I׀98��'���'2�' R�'��'���'��C�27n1�2��'��L���'?b�'��'���'bb�'�b�'����cՌF�t��!i~$� ��':��'�b�'Y��'��'��'4���7CO�*@���\q�I��'���'SB�'%��'�B�'L��'�0 �n�/v����2�#w�R��&�'�b�'<�'
�'Y��'�B�' 0yס&�f�)ѩ�#=&�ʥ�'�r�'?��'$b�'B�'��'������מrEn=�-F�]},IѲ�'���'���'���'PB�'B��'���p� T}��(�Du!8��7�' ��'�b�'���'���'r�'G�U ��[v�y��+Q*�` ��'�B�'���'�2�'���'�"�'X��� ���$ܲ%�W)5�`DIb�'3r�')��'�b�'�B�'���'=n�[�BG�F�Rh���7� Xش�'7��'���'�"�'���'��'9�U�c��4����N �v���q�'�R�'��' ��'&�e`ӈ���Ov̊���+4B��B͌.n,z�� L�ly��'��)�3?���i"<)���2��uA!n�6V����1���¦�?��<Q�����(OhD���N�1�,�(��?95ǜ��M��Ox�Ӛ��I?�kE�WPjl�q�)CD&���%�	ߟ�'H�>EHG�ڽ.� s�+S/®���O�M��iVD���O��7=��١��ͷX���x7�F;�&����O\�dh��ק�Ow����i��D�N��5��BQ�� ���k}�D���k!.�=ͧ�?��$V�p����B��a;:���O�</O��O��nZvDFc��DF��sE��w�
k�� b`�Mx�
W������I�<��O`aP��
x�T$��Aءo�K����I�2��:��+�S+2��K��PQ�PW�I�e_YlbT`�D�Ly2U�P�)��<�&'�`�{Tb�ts�� �<װi��U�O��lZx��|J	8a��ɷ Ԥ-�d@HT��<���?q��>Ta�4��Dh>�q��$�
�ҁ�Gd4Y:T.C�n�8y�G�0���<�'�?����?����?�/!�T�HY�T�b`j�*Ɂ��$ަeS��L:+�����ӟ �S&�δ�	ܟ�T���r#֌(@�\����d�Ҧ͢�4,<���5�i���	]�576����7�\]s j�)#h����٫i�f�ѵ�B����N��ם$��?6t��1#|�t����+V9�"G��Y�	�� �����Ɂ\�=�'�67�`����E�](H���iL7qz|�FeλX���ۦ���Oy��'4����6E}�Bpnڃ&誝X�U�'��|i)Ԍ �}�������?as�N0D��Ij~R�O��X3>�^9 �T��T+���gHF��ß$����4����x��N��CT�%�Vj�W������p:�)�J�-�?���Wᛖ*36G��ş��	jy���z�8��6g��
D�4OִD��7-Pg}�ja�.�n�?�ce���̓�?���ν1@�e�uc��;$������#3�qH�D�O�)�K>Y*O���O~�D�O�a�-ʨ<Z�	 b���jP2qaĹ0&@�$�<�иi��<�&�'���'=�$�w�@`���[)G�>es"���kܸ;�'hB����Iɦ��޴*��O��$��l��I���y�
�`�fV��؆욫�|���O�i�7�?��M1��F�h�.uQ�Ƒ�r^�q����@�>���OL�$�OJ��i�<���i�zP��ޠD �Ē�hwk��e(�	Q�	�M�Bh�>1Ҷi��h��+o@�K��]����C�kӨ�$ӹ,6�r���I8t`��8Q�O�v�+&+ܭ������pj�������O����O����O��D�|*�_.ktvݡ�#�T �pa˕RF�fD2;���'r���'��6=��]��ؔe qs"��<]�@B
�䦑��4�y_����?%�I�B� Xo�<ɓID@x����-g�)3$#��<A$ޟYX�d������4�����:b�y�r�T�mG�d)#i��?��D�O|�d�O��qǛ�K*#q��'z�Ę MN~���!�3~��I�mJ�O��'v6Kݦ]����ؗ�Р��
´�kt�S$"���O$��7,�8�rDbs��h��zB���8)AB�R��m0�.X!Y���B3� ڟl�Iϟd�I�HE���'7&���`��E0$ə�����|k��'+�6-�1 �TʓQț��' ɧyWcJ�Y޼	�1a�V���t��y�g{���mZ��QS�S�}��6�]7y��|���h��`x�o\�R����bPa���.�D�<�'�?i���?a���?a�L�/hf�K�I�=l�<�k�����$Y�A��� ��ӟ��Sa2����`��n± ��p���>>�dX�h����_ަa��4��v����ON�t#�%l�YF/��L� T��7�~��������4l����;��O�˓qَ�htСz��ɒ��a(�ѻ���?i���?)��|�.OZ�lZ�F���I�R�̴ؠ�W*,��#<'�}�I)�M+J>���I��MƷi�L7-�)AD�<Z���u&��g鈁�����w� ��՟|0�0��O�X��'�4�t�� @�4�%/o�}8"�[����>O����Of���O���O���@�ì�!��eE�D�_��-q�,�'A.��5�Ol�D�Ԧ��HEyhӌ�$�<��jM��;/L9i,���@f)�Z7m�Tyb�ip�7���^��q�o���	ٟ�c��>=������Ð Μ=����R�,E���'�<%�@���T�'Y��'Ɣm��D�v���gF��PT�'`"S���۴R,����?�����E"�
͘S����2�ĺ{m�I�������9Iڴ@0�����O��rc͖���2�\�Ĭ!��!����L�}��'���&ԟ�R�|�A��GE\;AR�9��+'
��XRB�'���'��O���F�FM�I��Mc!AQ�r��(*'N�a<�WeC�^��9/O,�m����'��!�>ᶷi�p�'�E0..
)u��7w'P,ďgӚ�l��~a��m�p~B��-/i�p�i�x��X�"�D�@�|軆'̨9�$�<����?y���?����?�+����w��u��;��u��!�Iɦ�C���ߟ���ڟ��Sw��'�<6=�4�ҥ�ܒ�ǘ7g��8�$J��5�ٴ�y�]���?y�I2�^o��<!V�ވ+J��#�͕:["1b���<��Dұ#���$�����4�����a��I=�pz6G��,��O0��O��Hq��B�7""�'��;:6f��3j�������^v�O���'�`7m �q�N<WCM����I��S�!v���B��<��X�j�;�K�g*�Y-Op��\��?Qg!�Ox�؀(R0z7|�A�AK%|$�P�E��OV���O��D�O�}��@�&E��
Г-͐4D=rh$�c�9�����1��	�M�����Ӽ����,��	��nyC�P�<QӺi:87���i�F�������?Qa��e��)��G��X�����OP�`���°;���zN>�/O��?9��� d��A�M^�\~�5�a�M~�x�B1Č�O���O��?����F`�H@�E'�5��O�����¦���4G?���D�O��4��5�x���j٩^�pgM,h�)xӄ�)/�剟5��7�'���&�Д'�Q�󦞦}�����7h@f����'"�'ob�'�&�h�S�<i�4^��K��<�0��DE&b�X���.V��\���N�V�'��i>���O�m��M���i�N�³G!`��d��X��x�ի:=}��3O���t��Z��M���?y3]c�0�qč�s���3-�MtL��'@��'���'�"�'��O������`���#S�a7�őM�Bܳ��'�rGk�V��ɷ<i����w�-�Pm։]��i� �!�� ��i��6��t�@�IQ	_F6Mm����9o��ԥ� HW��2"ƛl����蒴EM��\񟸕'��i>��	ٟ���j�n=@FF����I�5x  5���+����'��7��_���i�O,�����)g*0����,�<�P�oU;:��O�5�'+�7-զmhش��O�К7GV�]L��e%C��l+����xQ�Q���6��4��<��b���Oإ*�f&	�xM"��R8$ޜ(9u��O����O��d�O�i�O�����<a�iM �����3j9i�Ǽ|����P��.���'xB�|�O|�I!�Ms�)�nXT(G(�(�,�t �����mӺ�H��|�Z�o�\`�(���Ouf�����=��ERtEK�4���'[�՟���ן(������g� Ke�R��Rj�5s������w �6��.K�N���'���ڱ���DȦ�1}K.a��#����Ģ+!���4r�6�g��ԧ���O����>)8�2O�i����~֤4b�ő7�h�?O�IXD�O!�?���0�D�<�O���A���:PLmАŭ~v6y��=ӗ:B�'���۲S��)2���<7P^�b��äu�O�'��7-ߦMaI<9a�5(L��j�dB���Z�<9���"
�)x�e[+Oh���4�?����Of�+C�	!-ؾ1@��HZ����'�O���O �d�O�}λ
�>MQB�_� �����(���1]���W�B�'�d7M-���O�L	�Q�h�"�~�C��W�N�FԦ�۴w㛦O��:���=O����8Z�.5��'��Ȣd��3J�)u��46��͡�$�D�<!��?���?I��?ف�_Y	dh��e���
���Dަ)#bC�����(&?��I7;7横���t�flQ��g$R`i�OH�o�.�M���',�O���OL��2$\@fP<k��ͦ 1ք�",Y��­a�R��Xӫ�;f;R��Y�zy2��iD��ʃ�< ZĂҪ �R�'�2�'��O���M�7�X�?Yt우Z��g�JH�T��S�T;�?Ɂ�i��'��k�>�`�i�"6M�9	`� �5�
}�P��9(X`���0��lZ�<���/L�)k3��� �(O������l�
'hP s� �>J,#��O���O��D�O����O��$�A���eh�ar���;
�>E�T.Q�6��g�O����OXQm�1|���O���5�D�<X⹀sD��x�V�!�OD^�1�v
�G���d�ަ�)�4d�vID�S���=O��d^�P�<���g�P��f�J"�aa0���?� �0�Ķ<�'�?���?Q����x|	���)���3�,	��?��o�������U�Uk��?���П��S�?�@gJĉR}��nA�}���Km����C~��'웖�f�X$>A�Ӆ{@ti�C�]C�Q9��T�(�Z��g$+�@��E<?!�']^��d����v�p��^";l�@�JL�]b�d���?����?���|)��ʓf���߁RI���.�ݨ���" �	�� ��?���?i����4��˓4��F��2~6���A�^�Vi��O�s�6��킅�����"u���̞�k����?�3� ��c)T^�hF��Z�T@��iy&��'�r�'�'b�'C�SY(����K�٘dóf�5�jeYݴ̘z�Ĭ�?9����Ʃ����O�.K>�� �Wχ�$Ɋe;��Wy�20m���M�1�iİ��|j�'�J�⏎�M+�'J����i�Q�VQ�6O�=v���'��
�o������|�_��۟�2���:��sJ] �����<��؟�m��˓w	�&���`2��'���/+p�Xi�6V��JT.�1t��O��'��6�ŦH<	1�ߝ9�4���%�C�i�4B�<��� Z���em��)c�+O���4�?�P�O������mVf�!�& �nr��Q�Or�D�O����O�}λ}�I� '�5 �i�"	�|�D���i�&ǃ�-W��'o�6-&�iޑ��IK+;�$)�!�5�T	�	���m��Mc°iӄ�	T�iv�D�O083�Έ�����!H���q�_��Ay��ޭGφ�O��?����?i���?��R���J�&^B�H�Q��L�A/OH�:Z���'�R�'���y���K���f�˩3{�|��ұ|���#X��AlӊU&�b>�B�ɝ7�Bނ�U�ji#B˦ =�ia�qy"�D,�����5��'��ɿuݮ IS��?�t$Yv�20L��IΟ���ݟ�i>ɕ'W�7�B�����
�dTq��k�2f�U ��Y�l���D�OP�O�ɲ<��iO�7-K�Q��[�dCVD`RFՃA�q�u}=���i��O@���
͘�겒���S��5fBU�Hl¸�dg�s�={U+_1�y��'%��'���'>��I�=��}!҂s}�;W�tD�$�Oj�$����QѪh>�	��McO>ٓ�]�P�$~2"�"�<:�'<`6������1C���m�<�99|-kU*J��2�h���Ƹ2s��'B�D�$Ю����D�O����O��ĒDI����/Ϧ ��-�fJ̻A.x�$�O��!�� 3$��'�rV>��(I�B�2�+c(wspA#?q�S��Sشr���0�4�:�)��`����C'ĕ��kR�ڸ�t�N;0P�\A�(�<A��*���� "��=�lt;�#k��)�������?����?���|:�&�nH�q.O��o��O<aa���	�)�ʽ^�>�W�֟��	3�M����4�4y�'"�7��t<I�d�!k�U޾�llZ�M;U�؂�MK�'4���&ҢL����� D��4!�G� 5�X��	�!a�d�<����?A��?!���?�-� 0����&�[�AB?f�ޔʖ��ǦU( �R�L��؟0$?��>�M�;4+�<P��
����DG���(A��i�\6̓{�i>����?ER�!�㦙�%����
��/�����4Dn�͓Y�A����O�ICN>�+O���O���IL�:�����S��ctB�O����O~���<öi�j�R��'�b�'�p���7����T�3���A�EV}��aӈ�o2�ē%���0���F�$T0�K�	�iΓ�?��M�h�8q�O�-����*�Y�B�����6r����N�\�P�M�2�����O�d�O6�2���Z"����OB=S��XE4(�e�4
�8��7!�Oԍlڔs�n����(r�4�?�*O:�4� �E���9�A6�d	�3OX�nڢ�MS��i�60R��il�D�O�ec�m�� D$/f� 겆ǅ8l��{t/6!F�O���|"��?I��?��xH�)RA�`�����D���#-O�l�=EU,��蟘�	q�s� �@�ɻ0�~DI��>��)4K7��$B˦��۴�y�����O9r��+)�\@��͌�!�t����1v������%Q�K��$V�O˓>��P3��:��t3Ԃ�:\�K���?1��?Y��|�)O��l����I�iL:�:�I�4������ڳK��	�Mێ��>id�io&7��O,���%7���0��[�!����ʴ�d6�v���	0q"�`��OF2��R���&m�p��&L#�x!u�ѡs����?Ol���O��$�O��d�O2�?i{�'��7Þ��U'U�b�x9٧E��x�I˟���4K�P��.Oj�oZJ�ɊS 
�q�#O���u;4�FNp�̓�����e@ܴ�?�di��M��' 2�3,�8��1/�|��K�U�i��� ͟��|�Q�������ӟ��&W��*�
s��/U�h�(�G�F����dy�s�4y����O ���Ol�i��rl���X�$��Rj�%�Vě`3O��$�y}��~�2yn0�M�t��d�Oi��K
/APV9y����rˀeI���@~�4x�o����䟪|��'C�O�|J��8=ռ�öe��h�Tm!S��O�$�Op���O1�Jʓ$��F��,o~�0��Ώ/0H2 A%+�3eD���W�@ڴ��'D2�B͛���O�h�� �u�}�A�[|�6��O�M�CKn�`�Iϟ@����Gj�t�3?Yl�Fty�I�ɪ��%��<i,O@���O��D�Ot���O��'cWF00+�7+�8P����v���0�iF���F�'S�'��tV>�	�M�;.�4����)Fh�r6(Y?>������i=�6�E�i>I�S�?Aʷ��u̓'�4顓C-I���A��dɔD��O�d���M�Ob��?I��� �C�i��o�p�p �4}'d ���?)���?	/O�nZ�Ex���	��t�	�	�B�z+��,����ᘠR����?��_��P�4m\�62O��F�p� E��hZ�[��D�p�l��?Q�E��g=R�BA�M~"�O�r�����RN� Kqʡ2�nͫp��a����"�'���'b�����]�7�0�a͘3
-pA�Ȱ�4^�6c*O �mZL�Ӽ���'ph|!u�˔y=�L[�L�<yG�iG�6͙Ϧ¶!��?��O4dK��)q�? ���
���h0���8�>����9�d�<q��sD��h2%��+�Z��	S��I��Mkc΀��$�O��?y��Z�H�>�+�a�ż�FH������}��4r������O��DG�F3��2�<@�65X%L��9����3���7�2�����'p�H%��'0L�B�Dˎ�QG��%qPS�'���'!��TY��4T�2���.��9R6���,�fNӇpd��)h�F���L}2D|��m�Ms��	�>̂�ɦ~����_~$�R�4�y��'�౳�d�?}3�S������%�� �|,8aΐ�F

Lr��}�D��Ɵ��I��D��ğ ���71����R��&&0D|����?��?I��i�>�:pS�4��4��4�z�Z��I+[O*�v�Eg�@Zs�xJx�0l�?ݻ���Q��?	C�M����ȡ��#�=3���Z��k�O�MYH>�)O��OJ��O*y0�-ů|�u1��������O��<9Q�i��P���'��'哅��ʑn^1'c�ePF���e܀�(��?�M���i���"�)���a���YPv)��l8Q��Ex�d�pܠ�5�������?}a�'ȩ$��+b!^�B�v0��DK���3V#I���	\�I�b>Ք'ٸ6-O� �0�REL��)F� dB��s��<�5�i5�OT��'a�6�{4ɹ4*¯	�*񥋶척m���Bf���͓�?�$g���V���W~"Af[:p��₣s�|	B�E��y�U�ȅ�IO�#4J�Xt���cAD�)Űe��4!�M�)O(��.�S�Mϻ���(��0B(~�"�LA�@��*��i�7��ʟ,ק�4�O��4ȉ� �v9OV�@��7�^1(PkD�%W���$=O�iP��?�r�#��<�(OJ�3Aa�%y���TJ�P>0�IG�'7�r����?� �d�2Ak��F�]��E�<�i�?)&R�H�4��Vm�OF�l�HZ����0s�XC4N�Z`�ϓ�?�1g�y�p�8��1��柾e��XĲ��ֶJ���``۹�>�0�ǉ=F����O�d�O8�$>�缋���;b���fnS�<h;5!�?�i��C��'�B�jӬ�OL�4���`��R ?�I)���O7$�V5O�l�*�M�u�i��m�C�i�����j���O�>-���VS6�h ���5�j�2�����0�'"����p��̟��	��X���V}�!	#�,�ԭ�F�E^fa�'$�6m3_Φ�	�D�O�����T�z�,�<!�B[�i��&�ס2H���T�'�ɦ�M+1�i��6̈́I��?��S�~�|!e��w���Yᥙ~#���t�F�QH��7���p��O��	N>�(Oz5C��Y���E� EU�O�v���A�Oz���O����O��<醷i�&����'\���$�B�U�Mz��4�NT��'ߚ6�;�����OJ6��Ӧ��wKɱmCH5�5LJ�nap݁f+�-hݜ�nb~��	���R��O ��?>3��0$�M�K����u�ɞP�"�'��'��'2�'u @zR"!/QT�G�=ԤQt���DR�@�d-�0I��IA��'O��k�̰��'�*Y��Oq�'�ܜG�#�L4A�]�d�:G)5B-G�'s>7���m��4g�T�"�4�yR�'� ��PFH�q��`	�/����"�lO�D����'M�i>��ߟ���%sE��!�hʳ\ؼ4�����ɠ�EПh�'P6��"
ц���O��$���t`tI��I�fIp,�¤FI��d�O��?��4\�� +�i�n�뵬@�5*�AY�aK�@��yȰ��eɦu�%�	�J7���?嫶�'�nh%��1G�[�5z�mCyR` P�ޟT�	�<��ӟ擦i�j��2�QybfeӼ]Q0�.F����2�	a�DD�':��(O��O���?�)O��l�i�PD����2��7)������y�ݴ(�� �ݴ���B,b���'���2B�̂W�2Ea�aJWc�!y��ly��'���'�2�'��]>�J��7%�j����I?D���-#�M#�i��$�O^�?�"����s*�8H!��o��y�� �}���a�,�'���?-�S%M+!o�<y�ok�Ny��Q�%��:�)��<�F��Ki��ޭ������Oz�d�U	�quG�:/���qF*�"��$�O��$�O�ʓ@��ɉ�s���'�b�߳h��"��5;^������x��'U�Ȼ>A�i��6��ן|�'��i�e܌9��qLP�X)�=`�OX�������� �;�IQ��?y ,�O
��Oioza�%�'�������O|���ON�$�O��}λ%z ��%M����b�c�pQ0��H˛�.�=Z\��'�B6-3���O���&A�5b執��E��M���HҦi��4R���ʇ�&p��6O����$?���')Ab,8r�J�vB�(�7*X��@aX��/�D�<���?���?��?Q���O�d�`��#Q(BM ������禩�3M�؟����p��h��'�p� V�
"FR�� !M�J����e�>���i�>7�s��G���M�Yږ�Ə��T�~���+c]��eɊ��]W�������O�ʓ"�|��Vl[9 Ы��l}����?����?���|:,O�m��̼�I
HJ�)���u;�5{En0B���=�M����1e�	�Mq�i2.6N!K��a���c���'�D��B��lӪ���$"��ȔC+�4._dy�Ou��̯#ȝ�A
]�j	�q@gg֠�y"�'�r�'#�'w��iZ����Pοk�N��%�@�\*��d�O�����-�oe>��	9�M;L>Q�,��sV�K�V/
���_�ʉ'�T6�٦������
q���	Ο�H6�5� �z�K�<X�l�&l��j�(���T+�?���'��<����?���?����f�0�b��Jb�2�`M�?����� Ŧ���%�柈�	矌�O��,aVo*ܸ8��H�7Ι8�O ��'��7ܦ�CL<ͧ���J�3g3�}K�p��
���X�t�B�̀�J� ixD��<���
��&�o�(�s"X..�n��U�z��tH$��9E��!���8B)�� V�K�R��,�4�7C���ԣV�`����/q���G�"~QRQ�3� ^<9D��aߦ���KЫ'I���aB�R����Yd�6���4<H$x
�3Ֆ�S��SI�p�Q/Ĥ.���#0���<z�?M�:�JS�0ȑ���˦9lR�s�-���(���"�D�;��%q��\���
)�lt��ك:��t���b�TP0�M@*I�ȍsN�����V����7�R�
����ǴV��bdJ�9,�C$��_� [2��:J��x؊}��'�'���'AH� Dg��U�F�F� �HHu.O,̘'+��'T�\��
�.�����Q`�8� ��e~�A͒%����O8��7�Ġ<Q0a�m}��O�9�xlrf*ܠk�ԕ�`k���$�Oz�$�Oʓ#��[C��D`��RF%G/M�\6�����+/:�7��O�Ovʓ%����~
4�؞V�M��,Z,�`��rBǦE���@�'�����/�)�O����� ���E�a����C�zxhD��x�W� ��d,§��tm��"�0Ff]�OL�ݩ���Mk*OVș�-�զ�{��@�d���T�'���{@F;+�8h�HG�� Bٴ�?a��=/�!/O��?Of�[ ��n�P|�D�ğ%)@�z׾i��̡t`q�j�D�O����!&��SAo���g�8�R�&�	zY�޴6�2��(O|���O����OD�ʠ�վm� ��.��v��l�����]�I�����&{�rT�M<ͧ�?��'�v��+$� ;�(� N{M��O^�)O��<��?i�!��x[���8'lX��Q�'�n�@�i�b*<��O���OR�ĩ<Q�
Ϻ��ק>Hd�	��JU�m?���'�(��yB�'�"�'}�-3�<�W��u���cb��T�|E����ē�?�������ҥ  ���g���[���C�ԑ3����O����O�˓F{��p>�$��Fį/0ꔐ�m�$}�Y��\�t��̟�$�p�'#�ӯO�<��\9N�r\R�ذ��P����ޟ4�IXyB#��K�\�%Hr�܄^��i[q��C��K���ON�D=�Ī<q�b�N�'"�`����(/��m 1��1o��5o���|��xy�ĮlX������kL�
9�Pt��W����i��'��I�*h"|��O���Z��S�Ks�2SQ \`H�4���"E�B�l������O��)�N~���+Fg�Dh�.�5�������Ms-O>,�����'����Z�Đ3'���!��-*?J���rӖ���$���1��ϟ����?��N<�'1���pO]��H�T��&yHE�[���4��Iy"�'�r�Ϙ'�2�'0�tr�Iƌl~<�`���^�7��O"�$�O0���˭<ͧ�?���~2�E�;r�!i�q�����<��c��A����ħ�?����~2�e�rD'\kOT�[�F*�M���.�T��)O@�$�Ox��%�ɟjZf�R��@��cLˊlq.�[]t	p�%�c~B�'�BS����;���	wb��<!�"+���ԏ�^yb�'�r�'j�O��$ߥ ��M��$B;7�UJҏYN��ہ(���	���IOy��'���{֟&\����Ud���]7c���AO^ݦ}���|�	Q��?I�΀��ءn��S0T����&:y(i����%LM��?	����$�On\2V�|"���]hѬ�[�d	!�g�{w�iLr���O� �bW ��'9��IܲtJ��L�;pz<X�������I^y��'����gZ>��'�tF�X`����\}^�3�	�1J0�c�d�ɕOπ�zI8�~R���.3Px��2,I��E��v}��'��@B�'|��'+��O%�i���q�؋>{���$-]��xq�>���q12He�t�S�'sZ�H�'O�9�yRsI;�dl*P���	��I��`�SOy�O�GB�y,ts	�Y?E)r��O6�C	8ܼi���S؟԰ E�i��3P ���9pԼ��M���?Q��"E�+O�)�O��$����P��3�LD���!"CN,�!���'�:�i�>�)�O��$������$S�d[��	:<�by�E�z�T�d��B�˓�?I��?��{"m<=���ڰ�;Yƕ�G�����$��u�"�3ő�x�I��ܔ'#��!u��A���YL��
:^�Bl{AV�@��џ�	]��?y$�N83��H%� �5i@)k�D�/y,� :��s~"�'��\���I�,�~��'OJrI)A��S6ꭈv� {tl�P�	���?���9](�'.L�A�!F%*�t3�(E�=�4 �>���?i.O���K�@'�'�?9#��h2)�(Ҍ	PuJ�ġ��'��O`�n���%������a������%O|�R!�f���ľ<��Fqt�-�����OX�)V�"�Ĝ��<<�ʱk0o�N��>�.O:ad�iݙ��� �p�q���sxNE*���>�������?)���?1�����V,��f�?U���A�˴9�*�B�W���'�Ȩ3�����RЊ��
=m[�5����"l'~6�Z8eXd���O��d�O�i�<�'�?yo
h�H�2�
��8��\
vjE	5�F��Y���)�y���O�� �� 4i� ��m�bG�C����i�r�']�E�4��i>m��ϟx�q�&%1bN_�y��iCdF������ �,:�\4'>���͟h��)���0&(؍a%N�c,�+sٜ%o�ןd0щ�myr�'[��'�qOxp�����G�͹ᣝ 1@�� �[����	�`���?����O^5�1i��|B�՘��ϭ�Ř���(6��ʓ�?����?��b�'֜����_7C|8i7N�;__0���V@�h�O��D�O���?9�`S���$��uK�hc���4{#ԩ������M��?����'���
��8u��4-z�9k� ֪޵�����9� �'�R�'��� е��{���'Ĝ�Y�"�,�~3��#O�� ���fӞ��0��ӟ�IP@ q�O�X��̊$'n~��,D68k�,�u�i��W���ɑ:�t�O����?1clõ��8�W��;d=�ԋҩ��'����8((����y��v|"dP�'~BŠ��8�V}b�]�8�I�$|4�I럴�	ҟd�WyZw���t�^�2�b�Ui��KR���Ox���-ʠi����N�Z�l�Fc=1�B����W�;"��M�-�b�'"�'���X��ݟhz7��	�s*
4JL�c'nF��M/� F����<E�t�'~P����ʠG��Ux�DЄPy�`�g sӖ�D�<�B����4����O��?P�y��iS�<��t�� �E
��y2�9�������O��	�q����oT+��t��E)���\9,O@���O���2�I7n�X�E�9�J���+��G[��I:�9��eZ[~�'��S�h���"�z��'N��RD�0��z�$�s�[y�'���'|�O��L�^����L�|<n�X��:E��$���7�	ȟ��ITyb�'��Q�$ԟ�����Q)6�*���/1!ݴ�
S�i���'�"���O�D9�̓�W���X""Ĭ���(X�s�r(Yg�ty��'m"P� �Ɍ>Հ��O�򈈿yT�"�	��d�@��
77��O����I�7=�xh�:���� ��dM!}�:�PҮ�� ����'|��ҟX����K�4�'O��O>4,Z6DI,-��+�V�-���4��՟x���o��b���M��)]w�h@����1�p��'�rl��5?b�'���'��R��݌T���(�^�2�f��Z���?&f�l>0�<�~*ALr�5{&,�f e	g���M�G��>�?���?���
/O���Oz�w�N�A��9�a�=@U�5��צ��"�\]��c�"|���n����нMs�k����1�ܑ��i%"�'��k�r��i>���������:�6JTn�e� Ή%XH6 ��A�Hg��'>�����+�X�"�9\���A��� t �qn�ޟ��gnsyB�'B�'�qO��W�!!;>����nhF��BY�4ұ٢����?�����d�Of2ơ�e���8�'�	q���h'MH��?���?����'��t#fM̭0���Ԃ�g
�Xk'N�}):!�OH��O���?Q�A���$�N�Fa�$s�jG�:Qy2�Y4�MC���?a���'m���n.�5R�4d7L0gÑ� 
��/Dd��ROG}"�'BV����^[�Oq�j@�x:��I]%|'jpp�A�?~��7m�OB�h�	�2�aS6.2�Y���j��c��`�F�'N�Iܟ0�$(HK�d�'t��O< �'����$dp'#!�ҽ�$#�	��y$�Z�1]�c��>+�`��L�	�N��`c�2b�lZbyb���Hf7��O���O��	l}Zw�6��0k�8(:��u��X;�Ձ�4�?��TM��Dx��iӁpC����*T�E>X�Vj؄K�O� }�X7�O����Op�)�k}�]�db��$��p36!�z������M[`NF�<1����d3�S���Jҡ
�U�l�n��r��)����M[���?���� %�#V�l�'j�O\���!C�lJ������*Wz�3�i0�]�\a�Fa��?����?����y@���d+ϖ'�T�;Ո M;�&�'�~��r˸>�,Od���<����6�lH�cEM-a�w
�~}����'fr�'L2X�ܙ�H�"�����O�l���f��+æ�)�O8ʓ�?+O:���O4���[p\{&��0W^z����A#�Uy�5O����O���O:�D�<�WΙ�V�I�v	GY'$�Z�K�f-�F^����VyR�'���'	����OP�	*�nl��)�(3��h�w�iP�'�'��	�z�p���$
�w�<dy��B/r׈}6oV�MO�l�ߟ�'��'~Rn��4��iV�H��$�C]�W��X�n���M+��?!,O���&��d���'��O="�sǓԱ8���L������>���?���/�r̓����O��)���[E��U����4�z7-�<!�A˛��'�R�'���>�;��y1�M�k}z��/X$4�JYm�ß��I�`u�Ih�O�'>�Ak�]<%D�"�|0!C��1��U�M;��?����_���'�Y�È��hb�ڗ��9U�h$*��x� � �1OV�O�?M��*��铣[v-ࠢ2a�Z�H�Bش�?���?���T)/�f�'���'w���uw��'�!FEݺ$z��@��,�M�����d��?I����������1ڧ�7I���jP%�=֌�޴�?����'��jyR�'\��֘�d<�]+��Q�P��J@�?��7-�O���<OP˓�?Y���?I-O(@� ���b�8T���
�ʠ T,@�,��Jy�'8��ʟT�	��ԣ5��)��u�G.يg��I���9K�j�I֟��IӟP�	͟`�'Ǣ���r>��e��
M0���A[�m�(cӶ��?1(O����O���޺"]��6Ph��B�o{0�&�74N��'��'XbR� +5I�����O��Rf搂�Lxc^?7�XU��k������Gy��':r�'�ڠ�'��M9$�Е�@�W��	����~I�Io�Ο���vybm�5�L��?q��PBK
lb�hE�83����f���S��	蟜�I��<��dg��&����EɮܙR�W/6�)�O�HĴ�m�Uy���~�6M�O����O���A}Zw���eʴ8��Jh��w	.8��4�?����`l͓�?�+ON�>�	�iߺ]�ll���Dt������h��1�kCͦ����<���?���O�˓S�Ԭ ��^�'�xXq
�B�`[U�i_��p�'"BX�����!
J����cq�A�/	�9)H� ��i���'?�T�����D�O��)�6E�1aۏ'��!��H	�Y/�6��O"ʓ?�
��S���'Z��'�6-�Ƙ�N��A*�݇k��U{a�u�����4%��'m�Iӟ��'lZc�8`@a�~|ã��n^��OH@8ד����͟,�	���'&
]��K#��Y ���GZ�	�⯒(!������Odʓ�?���?q�l�+�v`����?%;��z�+��`��?Y��?Y��?�,O�� ���|2��J�"�\���lVK�\;pl�y�'�BQ�|��˟L�I�@��ɖ<�4��0b�B�r�Q�E�7a���ˮO���O���<Y��L)�����@�	 �B�kC!��"��5���M+����O����O�5h�;Ov�'�Z=�e�U�z����th����4�?	����w�N��O���'���E�=ndPA�A��-�8=8�ol~h듌?����?�`M��<�(��?� #چ,0��[���#^$�A.j�f�+�l��i���'1b�O$�Ӻ�EKA}wB1���n�h�j�̦-�	�PQ�!h�%���}ꆩ��S�ĸ`, %i$�y����1Y���MC���?�����R�ԗ'eDu2�i�O��Ł���s�8��i~ӴuÀ?Ot���<���'֖��[��r!�d#��X� {ӄ���On��T	�m�'��	���8{FP�"�	�M��m���I:GZo�ʟ0�	柬��*i��'�?��?A��hȺ��"a�"Y���.��lQ�4�?���^Z��Ty��'��ԟ֘�ƈ��Q��:d������b�l6��O�8pg0O �D�O��$�OH�$�<q����2^f��dI�M��KwdI�u�����D�O�O��d�O���)��.ո�iթ3|<C�O��{��$�<���?������$��uϧъt�� S�Bռ���)�j��$���	B�	����'Z
��bM��"�Y:i�x<�E��h����'�2�'�T��35�ħ3�N�2��X<CDpI4i�f���i�r�|b�'�"�%&��xb!�m�D��$�WxՄ�¦	�	�ė'�"���7�	�O��)/ 
<���/��V��IZ�ǋ�i��(&�L��ן KR%h��'���'8�� �+�(-6*ɨ���Y�FXlZ^y�%5/ܾ7-�E���'��D�;?iuAX���M ��lpH�y���	��P*��f��'���O���q�DIj�"D!I�׃��	r��"ϨI�R6��O��D�O��J�s�j���.�'��p!�`L2y��i8"�iI6@C��$.�SП�@'G�ySR��Cfה1������M���
ٴ�?9�GE"7V�'Rb�'��A9H +���:0$Pa�� �&%�Ob)�$���O\���ON Q�Ξ,8v|\��J�;�r�;���ߦ���J�R�z�}��'�ɧ5�(Z�fx���d�ܻ^ac6.�����n��$�<���?�M~*爔$���j]�B�f��1�Q� ��M֐x2�'`"�|"�'a�$Ee+��$hʎ>�ѹ0o��@5ʟ'��I�����E��4p����Optd��0B�kf��w�xiM<9�����?1��#Ft9��/��M��E{��"u�����S�0������Dy�
G,YLh�ļ�G_�r/���'�3(bj&���l���%�������nJ�[9��#�F
l�����'R��nZ��(��]y�V$��x�����{�A\z;,�f������^p�����������d�S��ktF�t�Q!.X�����I�'���Q�r�0��O!�OM,�
�}{]Ƞ���F;u|�ٲ�~}B�'���A�'o]�b?}���Ù^lqC �x���v�'6>�P��'	��'eb�Oi��q�t��TwtTP0]7{֡��ʙCϪ7�@AS���2��:tLk�d^2%x���#Խ	��܋7�im��'72I�{���'K�����H~�8H�G�
Ix��i�{󤒉*~�$>����@��/�ę C�!�8�f�7L��4�?	wl���I!��)�OJ��"}
����)�HՂn�r�h�������v��O����OJ��O���֦J]l�8���;l���+�+J� �$�ƅ�<�.O���&��O��Șl���q4m�>� ��1�>$Sڔ!m��8,��ş<����I���+�A�[�a
�N��!8Eh�k�5�3��צ�������Iy�����	����	�,k���G�K�L�1��Ы<k���ER���Iٟ ��oyr��8����?�� Խ��#�l�NE�#�,B��$�i���'=�OF�m&�I���q
BMT L�^`äӲ�6-�O����O��D�'>���O��$�O���ѵ`�������*�h��CT&�����Yb�P�C�Jb��'0k��3cɚU�>������S::�'JB���>U��'��'|�tT�֝�G��%nJ�8dmˀ�J$:��6�O���^h.�r���	H�O��{g�Q��@�nN:P��LI.cU
7��O����O����a�I߶�sAl  _L|CC��4��h9�i�L-������!V��#Rй�F��<:/н��#�Mc���?���ܦ��Ӝx"�'FB�O�]�!���t�@�H�<{��@H'�ƎK1OP�d�O\����5x����!>�@�iD�V��]lΟ�
�A��ē�?a�����3VD[$V)CS���gnn�xDUi}�D�ܘ'��'�b�'��a�x��h!�斟d�>8�� %�RՂ7�'oB�'���'��'���'�S����C���+�D&]�8��WNԦ֘'��!�	�jo l���&��O�@�h��&B����~��=��'a�5�r��,�}�p��)��b�{�U�d�h)2ӎ F��]i�� :Jr��	�%=�  �R�X+�Q�t��,rl�q�iG�;�%�q��@�p�`�A[�$��U C$����
��1oJ�it�QT�9���(�G�T z��n�Q���c ��|k��S �&��V��.�
H�vaP�aL����m9�?ybb��Ha�bn��Bfq�u�G�?A��"����w���M��PiAU�ʧ��i�0���Ǌy��܋0.�'�	����D'R�oJ�0q���@ec�p
a��]��XB�QO��|� ��	(�MS���d��LKH����DL���Ҹ�0i޸�'��'��2��$a�Q�G.M�4k�-��S"��,�ƛ�$u���/]�^�p{2��3�M����?a�K]�9��蒷�?����?1�Ӽ�&��Q�t]��շ>�2��cT�\�z��oۅy�B�^��Ų��L>�减��L#�NG�_<��xc�_o�I���4���E� �}&�`Ǣ�#'&2aB"�ˠW~lÑ̄ʟ��':�����|J��dU�V\z����	��r���j	!�DJ*P�v5�E�X4�D�HG[�	��HO��Wy�+`Q�P`\c�} �OV��\J��^�M��a�	֟���D�\w	��'#�)�$A�&���`�/�<a�S�V�/���Hr��If
1���-	k���ժs�R8X�ʫ9W��C�o�*5�|�Q���l<�!��0�8��$Ș@MѴM�Bf�PG���os�%� �'�r�	U��f��0v ݴA.�,��Ko���mTr<:�eV<QrIh��_q �<�W��'B��p'�>���[� q�ϛ`�V,(#��,�����?s���?I����*���d��@�8�\p'�i�pp� 5xQ  ��d��+�p��D�Y: �-g��ದU�8�!rj!4�\��a攟I���℆���Q� !l�O8���<Q���{:�]��B�e�H�	��Bx���=�u�;MޑXd逺HZUI�cI<Y��i�.ID��?$��XNR�`�U�'l�	�J�Q�Ol���|�LD��?��q�xt1d�/��U�2MA�?�Kf�(;s�S�Td�Nv�*���'O� ���%�}t��
���9��ݧOH�����cW�9����tt$b�I�j	�O�F�cC�P)����"pp�J��+���OH�0ڧ�?amC[B�I(�E�:�P�Z6�u�<)q��	j	�B�Ɋ ")���t�D����̜Q?�,"�N�q ~Yz�]98���'��'�`��𧜗o��'�B��y((��<I��
2���	�� *BJ�K}���3{�\E��L>�F��+_vB1r�/��b�Rp?]RX����>���lָ�>�Oݴ/��ࡎ@�;�d�K�i�Οp�'p��"��|B��d�t��D���h���g��7$V!���7�$XI��^�ˤ��Pj�gh�	�HO��fy�,D
k?�uY���l[t]��:UҴfΆ����'�R�'6��]�����|zdԔA$L�e��4հy٦d�*?	��x��TH�����!D�4�)���3�V�iN��?����!_���yЎ�0k��*6�N	|��	 �M�q�i��R�\��D�q��j��/i��9�u�����V�<Q�ӄI�l�a3K���04�g�z��Hy�� +x��6��O�d>�T�[��1O�<9y�"�h���D�O
�K�L�O��$u>�:���%��Oz�f@ҜAͪ8:rB\ÎA���'0ޱb1E���f�\��T$�8,���h�Z�"��	�`���ݹ�4�?9U�
�D�7�=�T��������O4�"|����,p�ք��Ct��b�`�m<IB�ix���̀%M^b$� ï!S�P����6 �,m�ߟ���\��,�Yu��U�PQ��k&�R��vU�N�Y��'���z��c��g~
� �Ⱥ����VE釡�<D-����>������O����A�@"f����VOK���xAM�h���O|��6�i>��	�8��h�c9	�~L+�%�
Y�1Or�d;<O�q���o�"aP�OFG�mB�'׶"=���G�
!V��VO��%Y�p�NزL{�f�'�r�'�`��,\��'+r��yGjV>(�ڱ�q��%�H��-�1Ob��c���?�џ@��e�/'�X���nR>pV�V��y�V9�w1�3�$J��<��j�"2��	�T�7'�V���O����I����Y� �IT�\ԓ���� q[�'@zI����f��;�/O*SV����@;#����'�X#=i1��
�?Q.O�i�A�٩))�����6lؒ�:���:wH])���O���OL��x)����O��S@��b�S+�pQ;c$[�_���%!�:g�������|��#Řb��\�C��.@ֱX���>I{���I�I{@Pj������*��)'6V�x��O�to�/�Mc����$�O��E(�!v��@�c,l�R��;D���/^�i,�ȑ���K�b��cd6�����<�eĎ�6i���''o�7	K I�E�MVE�-a�ĞG���'��c��'��=����FGS�b<b� Co�w��ړ���9\�aD��3|n� `3H���?�5 =0�"����H�c��A[�O�K�e�"Q�j3����b6	�P�'\�!��o\�fKm�f�������F�%[�~�� ���?������ed�h�a���{�r��`�\~!�$�!�@�A �.��I�2Wp�m	a�J0�'��Ւe$����$�'���O���"�'fN�*V� ��JD
1I�l�Y!S�'<#��@[�W2 �Ic�F�/�������
;A�\m2�#,~h�ef_�N]�92t9��%1���h�n0~��H��Õ^�t�3���u��RZ� ����%2n�I4@�����1IdD"<���?5L-�U�S��-K�Ni�<I�ȶ�4ݑ3��dǞod�#���"��<�Wb�*}�����A�q���O$���������T��� ����7,¢0�!�G�G �:ԧO�yBt��뎲)�!�D�
E������!�V�
"�2�!�C�3���H�b��O���Z��֟�!�$��q:�H��/4�4��f�'}�!�$W-Mb}�A-d)sC晻:z!��@_X��R�Yn
LCr��uh!���V�8��,J�y_��͛�bC!�$M�z�"�����6��鸣KXY^!�dTUd���M�%FY@�6��8�!��L�pP��)63�p��R�@�q�!��ܲ~��(%h�"t������H�!�C),�!�#� �hn�ъ�fH?t-!���%m��HbG5D����<�!��:AŲ1�c��1�D��Q,��!�$;L<�C5i,%�ڝ�@�I!�D��$�1p*Z����P��B�!�L�N�2h�$_K8l��J��!��2d����&�B@,�xfk��!�YG�j@��J*���,T�$4!� 9r�n�XdHѲ?��1T�O�n|!�$�Z���%�:+�F�B��?}!�$1
��@ff[�r-��4�J�!��jE|-�Ԧ�$!r��d�M�j�!�DQ�:c���ђiH�pΈ��!�$�zp�4H� q��b��D!�$�,�A
r&�,4�j�a��16�!�DQ�7��4K�����{G�!�d��ju�D{sdQbξ�2f�v�~�<��&[�U4FDYuA%)ݘa��BNs�<�����԰��_�&�bss�l�<�N��XÇ��b�:Y�$Pf�<Y�H":���i�oK�>����`��`�<�Я�!��ᓪ�y�D��,�x�<��k������ @d)Gq�'4���%e�������@��e+�<A�QSa�T�)"�c�A�7%��;��L-U�Ld��S�? j��a@�^+$����V��@�Ĩ�)\���NZ|�-cA�/L��eH��$���t��wFx�h��E�|������)Z�n���'^p����Z:JLmh�N���H�	ϋ}��E��-m\�[ٴw���7+i�)2���1�T��'_��b�/�8��4`��܋ �y2�f^����K��� 	
kb}+R�(�0-b��8 �3�*ƗbU�ȃV �V�<���d�'6�8 �cD�y�PU�_/����IÎ��0s��ުP;,��`%P��$6�\M%�d#�_�)7b5���J�u�i�P�\��?qE��!@�x<ȓ�)G�$a# �P d@�ֱX	��1EF%0���#D�hȗ�	��9�كq�2' Ti���؍RD"O�1�D��r`�a%k�h\5K�� !L\�ik�,6rv�D�X�`x�	�����"�g�1���#G��s��$h�^�y�]�hɅ�ɋ|(*���G��CX9�(�T�f9���&����[�7D�5j��4��X)�ꝭl�4F�(	�T�xyE ��3�ru"�C'�Op���I"ri8��6Y�lĪ��J�aj�a7����
I�B��T��B���r�q����#�
U�Y)H<��T�9@���O9]��g�lq��\
H=���Iјey&ЁԷ
�L@ZU���缓&
��0cx��aEM�,}�����>)"@�'�����'����Ϙ'�N��E)�'f�d!�d懿Fո� ���Y\ �E�(&��jV�8��D!�&S� �b꟏&2���PP�кp\���OނH�^� �)�,�y�HB�@h(x��\�R�Odu����Z�65h��1��I�������kW�F*�?�Ц^0 ���L>i�#�%0�.%Ç�v@��S��N�'ʘ��ՌW�+��\I�[=v,��ӫO"\�oS�#m����H�<�
���#z6�9��_
d���Q�;8���d�I�?"��a���&�X��PGF)14�!�G &��qhd�+L��	1B�y�Z>�6�!�BN��$���
L�=H�I<��!�s2�|�<gƃ'�Ҹ;𩉄D�屰�P3�<y�'c��aeG���$��C�IG(F.�?��W( �/M)n�`Ա� S�:�N�:C�5�ayb�Q��2�Jq
�\��u2�)ƄXZ�yPg�.ۼ 8ALC���Q�u:8m��Qy"�Z�C��O�A�̳$'m��T��	G�!}a�f-�'�N%����~��_�\���r����DAӗF�ys��ڕN���'N�:O<)cc�4�O�h�B)&}ö؂����`l��韆ir`�3d�h��ֆ��',�)�lm!P� O���0�J	)�$̐��7�d��R�hء���^��d��UC�s���+���љ��$
T�*q!0��~���ԣp��wgO0,�JU��fǲ;�\JG�:,O蔨��ݮ%�*�8����,L)���<g���E��4
ڈi�uV���Bk9R(i!*����
o�	�h� ���S ��-ʔ�ՍeM��<Y���( ���c�,Ȑ��my�ʃ�v��"�~ӱBU6%-<h����yB�V#DO���D�ů���2g�>��. �#u&�
%"ڥReh"<�P��%N�|�S�M d��M�BTTy����R�@=c��-O�����ڰ(\�%�`+�MY�eY6b>c��{t�TAj��h��	 v�u��A���Nd�N	�&��qfH�-�$c������∔~L�Q³DZ�i��X�To�X$�h��	�l�q)�lǿH�p����;�� �" ��x�t/æpr��̞J?y���:��
4��{��`�Y8�D�w ��&}� �A�JO7�ģ�����0H��R%IK�_:��On�~�N0c�.I�
�Q���80Ղ�wJ4=��i3�E�A�`���.(����b*B�.j� �J�.��(ZV�ط3ӬUXdh(S�6��'_��d�� L�� ��h
�T*����^��,�r S
�y���фd��'&��POS�II8��Ë��e�.O��'l5���CO~Z� `K�=ip���F#h	:���5�O�MB�n@.H"=��.I*1:mbf��do5�,�3;l�����?1�w`����&�>S�8�"�EQ�U�"�z	�'^�|y��PL0�٤��4[v0aB�ɷW���p	��L��h3f$���["Lda����pn6h�X)@ ԅ��&m����ޗ$Y�H\�c��Y`Q���a�j��Ȍ5>
�$;"��%V�H"��ix��!��њ|��
	d0�1�C+�3���%��AQ�}��)$�0͗'�P� ����T�Ґ� ƍ>"��O>8� ϸH��p���|�:�Y��I~k�}r	�1D��zqO�D�hSB�9��R�HP8��Yv�])H��� �C�y�^�Qs,�?�4-�q-X������R
7$2���DÒZW�@����<E��'�<A�����	2���QR�z��Oe 7 ��v$��"t��H�԰0�1�S�Z�����0�ȅ�v�C�1J�I	 X�1K��M�*�>��%��Y ��*g�`j�F��Y���E`��v�9O��6��O �c����N�8�dRl8�S��1�O �g/؈@�(ŋ-H4.�
iِ��* ��$[�H�<��MCm��\ZLH�Q$�[��~S��h��28�6*O����W	9���$�ɒM��,k"�#:`ń�^e.�a@�X��RRDx�I�l����%�$\�:b����.�O�|P�Q $��䐔�+S��1����%!�)/^�<�'c˟
�0��j���fmځ>����$�8� Y� ̛1��Z�+T��g$��K@�q��@�QVȰ@�!<O������?"a�*�Ĉ=[�2�G�J�	��c�F���$�?�����ȉb��0�g$�k�a{�-0Z�]S��"�0�c,O,��ec�A3!)�H�2͛!/P���4GH5^Q꾟x��/�y¢��F���w�H��Š<!�KT�:�J��ңWh	N%�R��{�ԻRj����a	�"X�5̑�!" =-�
�CLɏ"��a�DdW<���f� �{D��*֡��vı��]�'g�p``��QK4�L*�pc�O*���`�D��B��:J�lՃg8O���A�:.�΍�Ĩ� E��
�M�j���s(B�me�A
T=�O��!" 8҉[FȀ�=IxMx�ЫZ��!C+��%�֦#���%*0@��DҾd46K�w���Q&|΅Ҧ��)+r���B(�\ �"ϲ`%Bex��j���Ƞ�
*p@K�*U�Cŀa�&I���bH�)"(C	�jeRA�<�S.�8�~5����(����o�O�ĳ�	�p�e{LI�;�n�+���d��i'K�uL��²#�uC���Dʹ6�Y�L�l�r�S3�^�'�6(��JESCLa�d�KN�x@j�O���`�ߕ<����P&�_\��f2O�}��a/mblRp�8r] M�^h��1��"&�<�!%� �Od�:�/��=�DGEѮv�V�P�LW�'��c�Q0��d�/a@d�8�'��}N�D��6pF�<�L�Z6� u8���ɹ%X�|���a��(���'.P��k��^$0as���D��J��*5V����5/�YXaP�:.ɧ��aQ���YQ��]���:kH�PEF�wVax��
4�ָZG��
rZd���$�+����eΉ�4/��ŉ�� AxTZ�|B���$Iht�y���N�6���oT�|1K�����D� r(��`�`G)VW��K��� s���?��_�N������q)�t�A"s�c�TPcA9�g~r(�Vq�=�#G�&F� 0���bmb��z�l`0/"39��z��4�|�䁊w{�dq$���t2�8u Ó\@�87GI�0>vH�Mʆ����up�A�Y�c���Ҡd�	)��ST=T ��;J>�?P(���'
��o�&~L�}���"m3@q����C�!�0+��ʢN���Ꭲz8��E�)�V1���^��DQW�;�	�Z��dס:��qq ��.&�XC�M�!Ne�"�V�t3��
*-�p(w@�wf�9��Iw�O�����H��<�Π	��@;]@�iٲIي��'H�I���ܺ�%O9`��������T�ڍK��rǟ*<��K4BU`�����T	R��^E�d�T��[z8#H�$�N�Մ-lO`떬�	}"D�r��o"-3��N�4�j��#*P�j�:��"J�C���XQ%`�#{�B���Q���.(+~l�4�<xm��D~�m�,�v@[�k[���i�&V�@��HV�_�?���I�H�]��AH�a"D����䃳F����ӈ�W�|�(�'�>�־l��X��W�}�N�q��I��(� q�`�d���O�8-1Tu��"Op�K7��6[A��@ � @� /`�	������B � )G�����S�[�����$�p�P]ۦ�GI�a"·v?�0q�K ��*��	ȍil`���O1#5a:���8�ݚ��'T��."�*�_�zV�����ؾ7 @���At���lM�A*���0ŕ7=-��A	h�X��I�.�FB�	�G��驀A2�@-s�dG
F�>�\���҂b��a�B(q	�o�U�iX���ɿ���̇�%h!�P����+d,�/���c�&1���a��F�]�"E^�u�VIP�������*5�Ġ�\:`6��u��#a�hT��{F��'�T%Z�KO	,��S�l��#L�|3�FD�!9�����'��,z��fKV=�H�@؜�؏�d�;``6��c��$�b�מ��!ׂ?�� {��5:�+v�<!3�Z��,����.�%px�,@`@��2)>��G�ݖ*�(���)4-���9��*���`)ϼ�Py�g�+A�37�Ԟz����i�^�6��,�3�H��	?� �I|ڏ{bҬj�����=2&�c��ːŰ?� Ԅ���;�9�.�s,�-A��@?qۊ���i�3Ka"�9Ê�2�p=a��6$����]�.	Ȅ��#Z:"?i�����ގe@P��1m�Xdk�-�vz�)c&g��{wZX����"�!�$�z�ҽ1�n��BP`�!2�L,5���	7�D���I�b���� iޙD�DlۘZ��%�d�_:Ul`ٷ���y�IW1C�8�Ҳ�����lM��X�۠��,�jh[�EH�H�%�ă�]�3�	�.��`F��c��;�E2e�B�ɒx�L�:W��>�z��f�V���C��H�Q" h�I!|�h$HӖ_bB�I�|����4'��h]a�T�\�B�	��2�x���;zT\�A��~�~B�	 LP����O�r�W��a"B�)� j$�G&�%\�cF�V�U(*-�`"OU�P�U5>�;��ְn5�C"O��z�L�)@Д���U)6����3"OD`1�N�:HQ��!@*��G"O�Aɒ�Ԛ9cIXp�֖X?d��"O�PȥKO�
s:%�c�����#�"OB؂1��3Q�0��bűTBYyc"O����ώT�!3C�<=�Q��"O
��7-׉\�����a�Z�mss"O���V	,�]�b��2S�t��"O\�R��S�urY2�R�dKJy1�"OЁb��xr
9���Y2~I*I�q"OH�!ui͡�!S�[�Y,d]�"O4 ��n� E�Q�4J�5:�1�"OVu�s���.<,�j(-��KR"OD9�&"��8O�I�r	P k|<ɸ�"O`��UHS2	�sG�1BJ��R"O��x@�G�`�6�"�KI�A�c"O�B�O>&�f%�fE�\U��"Ov�	 j�9	B �t�GR(]r�"O��)�lML�IGÃ�[���"O<\i"%��'�������3ق�x�"OT}���)LQ�
���|�0كd"O�������⬘�v��%6"O��`)�<`�X��'����2��S"O0�1Bh�3_cxu�D�<0���@�"O�0��IyHj(�F��]���R�"Of��f���-�6��4i��}dV42r"OF�p�H'8�}��J��
\����"O�5 �ǇfoZు�F1h�t+$"O��rr�U6,��%8��	�3�d��"OF� �Ց}��Qk��@�W͸�"O��b�]�4���Q�>c�ܒ1"O�y�&/֥,&qbǩ�H(hL�"O�Pr�ګz��p(�R	>���"O�$�ݗ!��T��&��Y��� �"O�%����!��:�γ4E��@�"O�ؚԭ\U�bdo�gW��h�"O���D^(~��<	 ��=4�<���"O��#s��Y
��P�+�D�2"O�aCT���,"��
q�2?)޹s�"O��bE�3,�����5x���"O�#��^�
�&�Se�W, ���"O���f��?sb��@�+`BQXq"OH��a�1 *��^�afR�<�`뒸<��h�U��+?"�:���Q�<q$�*�q3�BƽJ��j�VP�<qT��(J��W,�=~�L���N�<IaoB�Xj��K��9Ye��
��Q�<I��S�3�^D1��_7cL�q*w-^O�<aSiԑG����0�˺o6*����II�< 	j���@�蚋��I%�DD�<��Q$k�V�A��fk�	�ED~�<A6���#S�}�$E�J��K@�y�<@��.kh�e ��ӗK͸9��L�\�<Q�˥���iUG��A�dȵ�WD�<A�c�.9�T�X��M�D_��V}�<�1,� �کic)�[h6�����`�<�B�I5I�6����,����UF�<QD�Q�j&ك���������!��W�^Tt|��l[aGR)�7+C:,c!�$ɾ��x���U2f�8�iĆm�!�d�?��9�gN ?�=��mH'	D!��<���%N�1
�ktm��Y.!�� ��v��,~y^��w�]^�� �F"O�Tk4*��7N�	2ʊ-��u��"O,��F�I% j���_)e��h{"O���#DO���lz�E�L�X�3@"OPd��H)!�J8�e��%s��x� "O<��`K#JI��յ?v1��"Oz��wǖ(;=���4��wj�u:4"O��ْ�O�F�Tq5�_a��zs"O���ǁ�b�b���l[�K$��ː"OJB�/L@h�� l�!"O�£�ca�-�3 V�k���@!��J?VxV�)S���z ��fA;x�!��8uN2�X �G$\��q��g�!��7D�R��\�$�j6��)Y�!�d)|r^l3w�
�	�����ۣ�!�D��X#�^,�ɲ��%.!�D�;{�s���81�	P���!�d�0�Ƅ��)�>P�H3A�Z�n!��	=Q�@����3&��&��gb!�D�2�2Ā�B�u���!�VM!��(r�E;7m�
 ��(��_?~B!�d]> \�����t䀙��S-r!�
�\�2'},���d�ä!�¥R� ]���^�!�� Q�!�D� L~����(.=���p&IF0a�!��l���k��
�����!�$��}��h�&4B����0N�)�!�ڟ
�����A̾��h���x����)���:T�ڇs@���dM��Tp�s ?D��Y��\�(�h8�J�9`��{�l<D���)0ldxy
eA1�0�Fb7�O�ʓ[�mKS�1�P���]ആȓK���2���4q��G�lx<���<x��/v(]����0s��",����:�:���!��R�*9�ȓA��1V�F�>�*��FC�����[̌P�	(nJ�A�-�5���ȓy�2��@4@]���HF+kq�u�ȓ�-��JH<�5�と
B
X��$p�g*['5.�y
��;c�T��Wȴ�SRǽO���yA*�5{�<��Y� ��� ��̙���pH-��0�"�cdAz��A�L�? U ��ȓ,,�ՙ�NR�g������׸ =�Շ�CU��S��T8s��R�3���ȓ %��s��D�TDi��R1ibb�Eyr�'�ܼ��EƳ��%H�8�IC
��~���aS8	��	t�v	S��.N�9���nI03!�B�8�f���d*��IG�'
���oS,	i2%��! h0h�'�~�*զ�/ �1����	)Pȳ�'���P� [���t��o����'�J1'][ɀ��cǂjt�, ���.O��SI��:�����6Vش�r"O��##"�����
*��"O�t�FD�ވ����/jܵAc"OZ�L��&�b�!+F-
hT�g"OZ;��,p�\VD�# �h�g�o�<�����J���V3��l��l�E�<a'JJ�?��������3�JH�<� ��4�mZ6#V�yj��S�UC�<�pH�gͮxXA�1ܥKE��A�<i�	.m�\[AC˳����Qh�<�1�]����'G�?6H�����f�<� |�K�&E�7]:�̝,Q��th���Ħ�E��'"đ�Q��:(�1x"�yv� �'դt"�JK?P�P�M)K�ّ�'�����#��U�:�*�IW�Ow.���'=5Ӆ��o�đU)�}z�
�'7
�i��)_���lW�xI�8�'m����6HrqjW�*m'�\��'D�� 9B���&KF�T�qH�'��X#��(5�p�v��5�xZ�'{���p ����*ƥ	�I~��
�'7x5�$b7.�u�-0Zg�9!
�'[p��5O�'W]
I��	շ�2Y�'Q�dp�j�$K��Ib�L�("H�'�������F5�Ѷ-��oW:���'��rFE\�M������M[��	��'rF�T��\���� _�S�>���'X��pd�*K7B�X&�\:�Y
�'�&m����)�.�ʢ��� ��m�
�'x�,�&!,�ڰ���[lM�m	�'�� ���''2�]��ec>�L��'?�;3��*8b^h"`D�7(���[�'z�-kwؼ��7��/o*Y��'^������ ��m�c
�$崩��'۔rŉ��%��S%�ĵ�'#��I���)��آ��DS:8k�yR�)�6x�@K�&��Z��h���*K<�B�b0��'&b�zd���4x�B䉓s��ģ�ET�=:i�p"K�C�	�n�u��͈�8��!��h�C�	>�����Y80%Z�%�Qg^C�	=;���*��j�� ��mX�<��C�I;w&�iK!��7�X����,>C�	�:�V�1��Q)w��5�� SC�I-0�H9��IM��I�V�߶��B䉑>>�R�G*e��x`ϒ�dQ�B䉑w��X�qF*&��1��fJ'�C�	b��DH�׽q��<ig^2��C䉳)l耣�I�0f��RN�q�B�		Θ�����Tq 9!!ϗsp�B�n�z�CZ1*���ѱ$9�B�I<B-����[�Jg�*2Q%7rB��-ek���n$x�P
P'm0B�ɗY�"$:r�B8�9Q���??�C��-/ĸ�UcM�r�z�������C�	�&[x�¶�^(�0�NX�THxC��Q����d��N�@)ZH27�4D�Hq�h[*!�����4@\��aK&D�x�g��W�X�r���z�p'*0D�09ĉ�2V����Jl�n��Q�/D��)�F��I���	3�ji��9D�8CV�0'"��*��\��z8D��#C��0O�b��� -*tA��5D�؂᭐�Ε�e�ݼnXdQ��=��hO�����Ě��
�� ��E	�}��B��?!yb�B��� �T2�/�j�B�"F�hq�lR%��`��D�Si*C�I�\�t��dБ�̭�5�O�p���D ?�rŎ=j��HT�^���!gRZ�<ٴ-	� 4�ġ҃DY���OT�<E�E�2yhR�f�
��f�WN�<i����*;n5cmd5>��4 �H�<Ig���4��NЙ$���0��L�<�#��&��9h�j,T�^�oa�<A�A]�>|�DR�Oi:%aR[�<� �ԃ�V�r%�-8C�C+a�i��"O,#Sm��*2v��"��86��"O̘X�BҩO�h�/�'9����"O�b���FD�)z�N�s�T�It"O��B�V�FP���Ţ/�T��W"O���QD׾G1�aA#�U6���"OЀ����4�,����YcƠ"O.��R�Xb�؀ȃ F@�H�6"O��I�+X�V���2�	:^Rē�"Ob���A�=mu��y������Y�<Yi�z�TAD�N���X�CN�<)���P�r4xPN�&-6�51�@K�<�A�
P਩�#ڤ��'�XC�<�2�̱$"�1�#��
�Ђ�@C�<����L�tب�.��`���A�MM@�<)�Ղ]TE���AN��e[A�v�<�7�W<)��@�s�:[��Y�VZp�<�R�������� 3mc�,�@ Dn�<-����& \/ Ķ�X�MGj�<i�	Χ+�*t1iI(F���[�K@�<�`��.m��2�S��b JE%�{�<i֫O�(�S�i�r_�0c�Çu�<�Qe�&(S�����3a�Y0&��H�<,�B�:��v�H�kd��qf�^�<i� � �Y�e	�,(�I�S�<�̗�tE�iie ߫JgH,��nTQ�<0a���)�6���D`�@m
M�<IB.�
T\<��AK�$ ���PՉ�]�<i ���$B�]	Fȝ�MJ��h*EA�<yb�Wl�:��a�E ^��I�%/B�<Q��^�r��@������l)&�H{�<���\�8����]���AG�y�<�2C�4(�┦�J�����`�<���L/3�d�w,��\SbMS5�E]�<Q��>5,2�����}=*�R!�@b�<id)�/5%A���1wZ��so�]�<I���-�UXх�61����.	W�<	�Βh_��yc�N/[�:l�&c�S�<qv�h�HT��K�p�}r BH�<��XN��Л���V����F�<	"�.�8�� VQ�Ag	�C�<yj�!g������(V�RT�r�We�<�s�_�C����K	(f"F	�S�BM�<�"��3�D��'C1�A��H�<���m-�Y2�ɒ!s*���u*C�<��h�n��0�J5M+ �
ćKU�<Q�@F*fXfl��IŠ�Bt�U�<鐌Ȗ-W�YZ1$6���q�i�<	���6jv �K�3p�1���Nb�<y��I��դ�1Ғ���,�V�<�U�� gK`�H��W*}�udOU�<��'IZ��1 [�I1��ʠ�R�<��ݤKpl���Y���:eD�<Iu�
(eR�]@��Tn� %�"�y�<�sK��7���e,��B����t�<��N��_�Ҥ��V$d����am�l�<�ҡ��:�1ySN�H6�t��Al�<�@���ލ��L�&����F\�<���?���ȃD�/D�*�#o�p�<�fm�V�F�`���=.�A�DLk�<Qeă|�P�+Ʊ`��R_�<q�L[�\`e��i�:��}(�.[�<�ED�kӢ��׎P�r\qH#

]�<ٵ� !qV�A��R� Δ�c���C�<� �@� &�B���+;��m�w"O^=ᵢB �$�W� R���"C"O��*E�0Hv%'�^�Q!"O4��vƬ8.Bhv/�7v�J9�"O�tB�A��u���@o��_�vx �"O�����Ý3��m� �~�0��"O�YÖ�ԜO�xd�]p�&���"OP|�e��'kn�{�+Z 8�(ݓ"O����]�1̱KP � <�D!;�"O�`��a	���D��$D'8�(2"O��@���Y�4yK�G3L K"O�뇥���*�8���-e/��!�"O��8�i҄u�THgKZ6~��"O���KјZ���pc��*S��L��"O���тc0V�QS��qZ�"O���1	֧fgҝ!��X{K�m��"Ol�i�a�1p1Q��@�J�8zA"O���H'�h��1È7s4HU�"ORUchI�G�X�3���!0$���!"O������1{w�ဂ�ЮTP٦"OΰxW/�$��xxd�H#i*8�s"O~<����q������C��Y�"O ���Ü2���e�/���"Obu2!Y�{�F>*��ƂW�O!�Zq�`-�w��g:�%�!M�qa!�d�+H�uJ��ԅ$=�@	��?%�!����!B1�?,��Is3��&I�!��9*�����[M�Ƙ�cJ�~�!��/gFl�tl"q�N9���l�!���tc8���3��P�����&!�dҵuth�&��~��А�'z!����I�,��DC"oj��څjݓS�!��?�����&PM8m�ꗷl�!�	�	�n���+�n[Xy�`�INm!�䋺%��K3E)Wv�����[�!��C�6f�����%97�P+q�Z	P!�$�.t��m;f�O�\��� A�S4!��S��jW�8[�,"E°3&!�$Ъ7�<K�Ċ�]=`�1��
!!�I�KAJlz��[Ut�ؠ�B��!�d�68��p)�iԟ2&��2�gV�Y�!�D]��&��.1#�d+E� H !�Ҭv����OP�ʰ�׏u�!�L�&����EW;o/�L�d�j�!�$M� �JQ�eOA�d%���Q%X09�!�D�>���[3NԜk�a�5DS�$�!�$��L����T4Lbf�4%a!��;��@�G�2�, �̐6(!�=X�^�pua������!�d/�:(!�. ~�3aI�j�!�D]�A��X�T$�3�E5�!�$�9vݰԈ`G4Qf���
�!�W�;�,1�T�L��>�����o�!�$�#�|��gkWs��xs��[!򄘽3��!cA��Kw�Św.m!���#��Y3�Cк{ӌ�:��=�!��~fVY[�$�8	�����A�\�!�ė�z#t=�A	�:a�)h%��"R!��
ڶ�����o��LU�x6!򄉦-���$�H�~u�I�*T�3�!���@E,�"W�Yv0�Ș�x!�DQ�g�ukD-x����C�4g�!����Y��hC�u����(R!�dS4AU�D��2 ,1���dW!�� V)����:er�kA5���t"O�Y%�8��i��A�EJv!�7"O��RkP�@%��H��B�`F"OX([AHZ�x�Х�Î $f:��
�"O�� 5M��>d�1:͟+Y/R��"O��h'���(��E�rlR4*
\�"O�`�&�M��M���ǄM�� B"O�ٓ�P*
��0c��{Z���"O�,�O!l��1�6��1ڐ��T"O�-xQ��CO<\P��˸hb�	�"O�h
6(K;o��#����'|	�$"O���F�I�J��5�߬h�$b�"O6@A�E^��*\i�	�b"O�hrv!��U�p8y`*M)u��x2"O�+�#�ho��X�G��)Y|��"O(�f�������5��x�"O̃�ѕ/�&]���m:j]��"OfyCg�����EZ81�`"O�I,�X3r������b^RE!�d���X� Ň� =h�aĳ`�!�ė�	�H	S��޾�>Cvn�(V�!���ZLU�Uƴ�kM)sx!��ƖG�dYb�G9=��0ҋϞoS!��Bs^��HaH�09v�i��<*>!�Dl��t�$�B0-R��ÉضF�!�ʮV�ֽ����$|$m�0�ѕ0�!�$Ч'����E�4K[,8X���L�!�D�(D_D5;�R����%I:�!�č8�\�
�ӏ]< �J�䄻\�!�� 0�h6�C�`Sz ���{!�#rGh�؄F�ID`Eb�!�đ+-ôm����RA���f��!���c�n�z�/]�[,v�a��ti!�D��=����fn��BY�4�B�"O���ʁ^��Q�a�R{l)q�"O���M80w�l��`�=im�=1�"O�=H�E�Hd�9���$���"O��"�ꄑ@֑R��]Z�Ѹ"OX���;T[8�rC^�X�[a"O��z%���I�:$��BO�	qXl�p"OP�S�O��ô"vk�JU"Obdk҇�*1	�ě�h�
g{n�"O�#̄�L9�q�$�#S	��T"O6��2g�m<���9"�d`�"O:��u(�;LʸJ��n�L�&"O츇'�m���RE�ľ;����"O| XѢ�4,��	��_�!4� ��"O�1٦(28~
X@g8g'J尐"O4hʂ%V�zg$袲e�:Y��"O����2 � ��R'Ua��KW"O>�J���)��y��8e��y��"O�P�O�/Y�Ei�&]���	r�"OhwJ��Vd�a��S��B�"O@�E�*k�XU���O�����p"O4i�a$�M?���c\�F����S"O�sd]��A�'��%c�"O�,j�oM���� qy,YR��S�<��ۘ?ƀ��#���P4��Q�<9a�.fb ��`��%���(1�N�<IaF�"-[0ض���&5����L�<V�]����8y><L ���D�<a�+[�3�m3�C՞4*R8��<�G�	�tRNUӈ�,+nT����w�<���[32�\x��]���+�`Ju�<� z$q�H�{��r`�&1����W"O^5R�ݺ@�dlEl�իQ"OX(�'W���ɉ� ܄�����"O���V�.6�h�1׏C�|��yB%"O��0��,mH�T��o��4����"O����	��b{��: ��(���"O�ͨ4�ʗ=Uj����Kn-�|[�"O�AA@�]m����g�|D��"O���KA�H�
WџbvF����_�<ɔ�/9�Ɯ�çQ�Q��ј�-Db�<ap*�MVmh �T�]f e�nX�<��7S�dD�Ţ��*pce��R�<1�_7Pb�2��r���gI�H�<��A��ujY�`�Ñk�@H6��I�<��ő�z`���ŗ�Mk��#�"MI�<q -B�x:�!S�.Kj���G�<A2@�W_�ڥo�/j�h���<	kG+iϮB�S�zZH@��O~�<��HQ�3�M�&�,�p���}�<��˳[V��w�7{�,ͫ�k�x�<����/5��0Cm�40�-(��~�<A��F3|��tc���-mHT,�cV{�<aR)R�tx���ϨW0��,�x�<��ȍP���p�\�u�`e�lt�<-y�X���G��C�ܰ�G�Y��>C�	��@���=Ka��K��>H�&C�?v"©�u��P0��$\��B�IR8y���;'��[$�|W��?Y���?���d�Z�U���:��Z)N�I����y���1h��[�],(鐁2�#��y�ǉ{�X�1#F!k��1!�L��y��S����r��?s��q"D��7�y�I��;b�t��kӵe�x58d�ϥ�y��w�a��N�-X��}�!��y"�.�&��JY"P0Z���c@��Or��O	<����y�����V""q����'Bn�K��o2����g
�B��<#�'F0a�E�.� �"C�>u���';2@r*�6$�FQ���fNJ��'Q�L��Y.8�4!� ,�\��'R\J5O%M�QFV�`ak�' ��G�/.P)R��|�����Ol�d,擏g-�0N��,j� ч@.bMXB�I���T�0	?
ј	�3��50LB䉨4��i�
�fBB\�ċ��82�B�<Nr,�*�*զn*0|r3�^t8C�I�Rr�W�B��,��E�N	�"Ohl�R�÷��%`�C�h�ԐH`"O^ܢ$�&�d��B�k�Z=��"Oa���^G��%��.G��X��"O�A���K�M�Cf1O���3"OxŰ5I\���p%�5���D"O�HP� ,�^�h5$�jn��r�"O� ��#3W"m��a]�Q��Y�"O��0�L� �K4@�1��!D"OD��Bƞ�*;�8y&�� � �i�"Ov��k��{�@)"�ϳ�L��"O���RDt�Ƙ�V��� �赋@"O��X�d�|� �F�	49Aj3"O��yG��},2�� oO�O)Ɲ*c"O�u�r�̻D:x�R�ل$�U�"O���UF>i�h)���`�8"f"O����K:�Z�%d]�$L]P�"O<�P��@�G�.�'C������5"O� �-����{��݀#c�-!��%"O
tx+��q�idE<kЌ��"Oȅ1��وgZ�[���)c4��F"OԘ��\1����;�RM��"OPt���":|�����{�4�X"O�T�kQ)V��2U R�y�qH�"Oa[���R��X������q�"OH�B�戮7Dn��ƟS��UpQ"Op�CC�-�v����5%A�u�a"O\�A�iPv�!��nK<�â"O�R�D��Yb|� e��,T<�"O�8[�j�"�mX��C09?�i�"O�DRf��x��,j�hM1��#�"O2<���F& �����ǁ>p`��"O��)!��#C���ӄˣK�,� �"O���D@�df����c��Q����"O*xQ��	�cv!���V=Hǌ�"O��#���4����G��* 4�Z�"OHx��؇h��#sB�)�B��"OT-	F,O�m�E����|	�"O̩�G�� ��t"FGH� �	��"O����"5V�R� MM#��c"O-�b���pT\%n�7@B#�'�ў"~2�F��F�%M�k�l�T��5�y�N��8�q2iQ�j�:�:��@�y�i�	��{Gm�a����⇒3�y��ɰx�RP����Zr�ґ"�y�e������A�Q��J��y�Cсd���QE��PJ\M�������hOq��-��AV�b��uI�=�T])p�'ў"~zS/�+=p4,r�*�H����˔)�y2�"f�Q��c�%7�Z��kľ�y�b�`ۊ�� ��>d���d���y򤜌N�X�� ]K���@�"P�y'ITh��� C�B	�6G��y�!4b�!�N�,H:�m���y��$2���rG�*��D��	
��?q��4� #<QqL�
.6f
��:�"���L�<�	�
���5�Q��z��F�<�eh?e;�ȣgM?xZ`)�1�A�<���$e���{q�ܽ@VI���d�<ф��7|�a��Ĺ@�����`�<�%)�C��ո�-�5EQ.<zԂ�]�<�dD��A���ju�H�8m��ɠ��П���p�S�OVJ�(�a��Q ��0��ǥHD�G"O���K�^7f6�
��4�X�'��Cn�N*jY0*D�$��'��e(`�I
	r�4B��V�Q�	"�'�@ Kv�+"v6yh���~X��'\aX���4wvU��X)߶ "�r�)��bk����͡��IQp#���?����1-�lB���""iT욧��JTL��ȓ*�
T���N>P�pD�D�U��[C�!��$�#>�� �B?Z]���ȓ:�T�!l�!߾�1��;>/��ȓ_lTbgI�6�>%P�C�\TL�ȓFC�0,̪W��ɋKű5����,�`�-ɥ0�\<bU��J�FM��V����P�Ac�+i���6�PA���4�$D�БA/� �๑#΀#����#D���c�%n@�H��������!'D�`H`���r��*��^lۂ���� D��sӎ�
s�nɲ�)JW���ի?D�$@��� e�`!�q��t�!D�� �5�b�T�D���c ����E��'�ў"~�tJ¢\"�� �t� l��˙�y�`��$�(���3iŚaq�HW��y�I�9��<@ԂD�LU�%ʣܻ�y��O�4������Q/U>X�#L�yb�3N��#*T�S.с�Ë�yB���$'&�ZU)��N�|T�W)��y�����c`E�J1� (W�W��?����$�q9���
:!�t(Ѹ0"�=��U�v�� ��YilU�u�B�\�60��i��QѲ$��M5���ڍU˘��ȓ��ysŜ,;�^ɰ3�E�FH�ȓC����e��b����_����ȓ(���Ib�N&n�29agA��<l��i��l�We��73�;���,�j��I���?�'�Obl�è�5�>�"�g�9n��� "OL8���I
� &�2R�Ex�"O<��F� =m"�ڑ�ŞhӜ��"O$�ÖИ��W*�
c�.P�"OF6���p�Z1qԫ��|0�"O��2�͆^&��E*�2fU&퀥"O�d�r)R�="E���e�
��@�'�ў"~�$�G�I8�
g�;LJ�/[��y�aq��I+gi�+V�����yNK/px���B��`, �/�3�y�C)nPPu�`QhU���!�ya�`L\��.;_Q�AB��y�#L�
G�<��ԥt��� 1N�+�yr#\�rV]�ƚ&g\rUZ�?�y�2~-�q�pƞ�vٞ�����-�y�a�e1�؉4	�ks��*�iӝ�y"Z�#k$1h���5p��1��y!� '���z�ՙ*J���q���yb��/cZ`󁩑 ��`B����y2��N��z#���b!Kbc��yr��F��Z,�<1<�Á��'�y���!�����;P���sO��y�d�Y@��!e�� <Z�8��:�y2͞=*�0x`푖B� ;�!D8�yB��B8X$���@=�R�Qa%ʵ�y"`͔"��ar�^�`�f4��ˋ�y�N!4�!���6R#�9J�
�7�yB�_7)i`�@���=��x�g�-�y���#��AZ 
1:��8r��^+�y�=
:tT�w�G]n̫3N5�y���$��T�����<9p����y"l�?J�@t�§
Q8`����yB
�^P����-ۺ0�hA��*�yB���*⪼�([����c��y�	�25���_<^��Հ*�y�`��!��C1e��0ݙs���y�L��p�l���7�z1@�D��yb���
�4�B�H��%"W��y���W�����[�ԘyCC�&�y�%Թ+
ԑ��&��|4YV�ϑ�y)�88��x؁����P�D�X��y��=1u�5��	��-{Ucі�y���{��� _'�\�C*��AB��s�Ĩ�T�֫3��x�F��<L�C䉎Z��!�p���&��	×�.��C�ɇ(Ϯ�+���l�!"��7S�NC��:?b�bh�%
�ƨ�LQ�xZC�	9S�j�	��A9<��(T�5�C�	 I5
��'D8a���c&�]�>�C�)� ��ׂ͎ ��bl��J��@"O��F �!p��EK±jj�}��"O�`3`M�$/쎭�E*�(4�"��"O�|AGEs�:mِ���E >���"O"a����=/��A�%"��!�|+w"O���eHI�� u�� �X�rX8�"O�-"�N�6l,��B�;���"O�h��C��.��Ѓ")^
*�
#�"O*܊�L�!}o�$�wa�M���"O2|��Y�=�d�ypG��X_�46"O� �� ̓%8�<y���)u:~�ё"OR�F-��(вJ�Z0i3"Or��#� [FH���6�U	�"O��qPA�[-ڠh!B�]T���"O��`�,UqJJ|;�O��@F~	{�"Oބ3gBV n.̡�2hˮ��E G"O�����;=�J�)��l�$��"O0��A�,)pҰ�N�\��"O4�XCčq�.��vNO+`� a��"O��sk

n�ZQn��et�=B"Oh�Ԯ�k\�����m�$�"O�L�R �,.����K�a�|D�"O̭	��O�* |����Q?|�ޔ��"O�-�� @�3���� 4�� 0"O�Y�ӎ�\�:���gnhx�"O�<��m�����vM��[U��9�"OT|��.����˕
oH�"O6���
UR�	�B��>:�"O�I�kG�W�#�皸p�h0�w"O��;$F��K�r���-ᬐ��"O�|#�fïA$Ł񄟟(ƨum*D��;P$D�j$d���Dv��d)�m=D��"��Q'Ƃ��q�%}Ŷɺ��=D���K,pX��(ˏ�`DK�-=D�pZ���	P|l��ӢGg�N���*<D���Ǝ�l�|���GE6I�(���-D��H�aM5	�2 kq�D�/��$c��%D�4�$��>%�3î/%~h+2`'D�Pj5�B�c!ĸ�cD1XYq�K3D� @���_d}�&�8�0< X�y�E�*q���	�+N�a����y��A-O��uk�'��o]��J��֛�yR	���]��?h�옪P��y�D�{�p5�D���`�t� ��"�y�D����L�E@V����@a<�y�� �p49"mM�,h�	��y2-\t�Lڰ ]�E�2Lip$���y2��s>�ԋE	��m����$��8�yRS�'��Y�l��\2�"O���y���QyBT�Vo?VtHͱ�G���y�L�H)�Y�b�)YFtX"�	�%�y2���~���D�4\��@�J
*��B�%t(hJc�J�e"�� PF�C��"_8B ��Z�^�R����7.��C�	ay$��o� �\�g��R��C䉟H>Ȉ�ЮMe�!�U( �C�ɸt�уȔ�p�)j�;<��B�1ph@e�B�KE)��R4
�M�B�	���� -�#��apc��7fh�B��
Z�t�# D�6�T�z�k�vJ���9��|����0�J�Krh�����QAI��(d!�ӝ[����"�:8��!�c!��n�@��!-�="Ț� �+x�!�$@�sy�-0�
�j�� � `F?�!�� v ����3δ{F́8g�޶�"O|�������0	.EP$�aF"O�	��6c>���V�mz(��"O�A���L%e~��0U��j�fSR"ORqj$D�0ab*�"�n�9�F�r��'��I�x�j��4eȣFYr�el&O�ZB�I�R�����J741B�ת{��C�	�^������>?r��!��%��C�	+M(�� �� {R����&,7�C�I�aD�ˤK�TuQ�/ԴD��C䉓X炐��ɚ�'�Ik�h��B�	
]�Ρ[$��4uW�$a
Yg�^B�I�NԋE��'����#X�,PB�E���6���8u �E#E��B�	;f��5�7��7�n]{B��-S�B�	�]���B7ά
�L��ʄ�+zB�	���(��@�?A�HI�c-C &]
C�ɴA�"��s�\l���&ߊB�ɟT��3R��
c&h"�k�_�C�1Aph���I=d��T��;��C�ID}��r2͇�>T�uЕ��7Q=�C�I�k�Ԉfe��ޡ��'�*��C�	����q�:|�I7&Z��C�	�n�^\bAB��lEIP��s�����O,�"~zA��\�2	�%ΠOҒ<����4�y���]��K K�֑�b��
�y2�I/��9$?��x2�L�y��)�"YQu.μ�+я��y�@܆U�6�'L� ����y�&�
]ҌPNq6T�����y¢N/
Ü����.:��$�(�ymL�!P��#�E�f�°��j���ybo��h��"c!]� 9j  è�y��L�|^�W��3j���W��y�K�kƜV&˨
��G��y2+ϲ�^=��c�2���#l�/�y2���@�H:�ex�C^��y��˼[��:u�\�E������y��C���U�C�?`6 0����y�*��Lv��n��e�@<rf��ybhɥh&Pt���>Y
�������y�垸E�P����/��%A�h��y��E�01�`��~�r ���yr*�(�$��5��j�d�3O�&�yrH�j �@{'���m�!g͵�y�FH*7<�}���U�BL8a���y�"�.N� ���a�l�J��@&Ɖ�y"�Xy_�E���m@Z�Q��L��?!���v����W���F���qg%(�ȓy��Z��W�g�,!���*��(�ȓpPh-���)A1Q�6-�m�����r���A4w�02s�f��5�IQ�����Y��J�
u���-�%���ƈ��'.Ru3 럂�d]P�Ɛ5�y{	�'�a�%	E!�0�q㣂�k�"	�'А�3�-��$����G�b����'�*��գ '�������es�'�9c��&������ �'��8�S&ƵAl�y��K	�Y�bT(.Oʓ��S�'�y­^��8HHwM��"�f�����y��_���a c��O�ah����y�
��z�X��ܽ@m~!�3C�5��'rў�O{�[�@3?�F{�JӸ
+ �S�'lt�j�#-��2��A���� I�v#�/n�����'2��"Ov ��ˆ�ܰ�#E�&J�\�x6"O��g�M��-1���a��A F"OT��E$êr�"�y'-+S$Ȩ��"O��$ぁ9���Ҷ�׼gAP�� Y�H��П,'�"}J!��m^�Q��9�vh���3D�Hj  Z�wl�u2U�U0#�2�$2D� �$	�!=I&#�gO�"�X��2/D��2�@�`I��B�g��lވ#7�+D��B*�.A��8�ThN��P�2�)D�P��!�:lH���c_#c����T�'D��Eğ?8Mja*�눗lӢ�1c�"��V���S�D���0.-�������[�<B�I0,�b�*حC\��/TC�	7y�fPpc&G2^��s@\7 =NC�t��L�b��`i�t.ڎM�tC�ɔ�Fầ�;/l4A!طB��B�"krLY�.�-�´o��B�I�w>VՒ��ՙyk
���͟�1\t��?A���S�O�Dms1˃�n.~����!��)�	�'���p�gظR�d��RI�/��|R	�'�V�3C��X�:���D�)n��'#��R�"��Y�$R� ��\J�'�f4��Ĵp�J�*��#��H>9���?ц��?���H��H�ekS6�b�AmN��!�Ę2/��a�Ԏœr�(\��l�I�!���&@P�;�2��e��Z�!�,8a^%`JE<"�N\JƤ�`!�D\�S:N��vB��e����VD��a�!�D	�A��Yep0�
�Bq �ȓ_"@���\�
���TSҥ�ȓ`X�e%��g�l��&��C�b��)k�*4$�dadU!<^�l��X#�QX�!�t�:���Cx|A�ȓ gr�c���s�)k��Āo(Նȓ&2HR�?6@�xt��8CZ��ȓS�lp�IۼC� urNðp�p	��)�r��4c�#��� ��X�,i��ȓDp��6N�*x����+?eB����HSf�6���M�B8؅�HYXe+�Dɂe�4�C�m[+��Q��f	�%a""Q�P�8��V�S0�ȓs���)ь�b�j8 U�ɂ��ȓl�ڌ2c�!V>�X8��+Į1����Li�ǂc?P�Db_-/��<�ȓ�H��s��R��lS!(;͆��z~�=R��Ӆ��6}�P�ʔ	�y2��5�ډ���O!dɲ\�����y���o�X �JI�c����C?�yB��&E���F�����L1�y���
,�48�T�1���y�@ހV]�Y��T�t�r��aA�y�fP�av
�ϖp��ɓej��yRN��(q,T��ƍc@m	���y�N�J��d�@��)2��\�kت�y���5����J�'-��Y�-���yr,�,^,��&�Ƽ@Zy��B��yB�E*�,@� �����(:�k��yB燠��`7꓄}%xi��@��y��&64��ɴBX4u[h��5O���y�NJӼ ���Y�lrpɐ�!���yr���|�4ȓ�LP5:pP����y����L	.��f��Ipvt�rݏ�y�nP;I7*�0�j�>�P��FNU��y
� �l92�
&.e�@;��P�k[4���"O]��+[
M�Z����_G�5��"Op��F�.n,�t�Q�G ;�Kr"O��[�c7$���AB�B�	!�X��|��)x�乻��y����oChY\B�W��!�CYH@[&(�-�4B�ɶ`��yR \6����)ց8��B�I�$�~l�TEE�YK#֋P>�B䉔u*�P�eˮw$	2P�HTb�B�	�S2� ���+|���GǤ>j�B�	��Z%��F��Ymʔ���E)d��⟘��ß�G���!����a�zM8	�@���ybG	�>`U)'xfPEk�4�y2�G3p%���ƎE� 4<�� /�yb�4G����4�Z���RC0�y�j�m4�� C�%4�r��y���Fh\��'#�pd@���+��D�O.���բ �Nh�E��]r,k�l^��!�%u�2����%�*��F^~!��'8,L�;&&H�`%JH�f�!�KԖH+$�N�
�%ɡH$�Iy�'m���$�N�����E�C���'�����<m��찅-�9�̘
	�'�B��T�נV��uSd ��5�"��'���a���0>���6-��b6�\�n�`����J�<Q���\�(�����"�{�<As(;����
L�du�4%Q�<�ՆB�#��@t�c�&qJ$�L�<�� Gw_����×>Bȸ���Pa�<��#��Պ Nƺ|�r�F*O�Q*'
��B�H0�wa�L*���O:��d	*y�"y���g������9U�O0��$��E;� :aS� b�Q[���_l!�Dŵq1 T�fYz����ҭ�]V!��Ty��ÄǗ�S�ta�g�$J!�d��H]����h�<PLa�&���!�DV�64B����_!����#�>w�!�da.�r㇕]��#⛢A�!�dȚd):M�u�E(��B!��j~�O^�=���p��H�f���B7��:�"O��yu�@�u�ZlY�lΛV��"O<Q3�(@;C��Q B�K$Mw�Q��"OF,�!�h�2͌�R8F$�f"O�!KƂ΍_�,��L�wz&d��"O.j�@T�s�*��*Ը2dh�"O��V���,�Z���X8������O��Ɍ*x�<��p/@�w���rCb�"l!��s�xP[!L¿:f}�v�G�A�!�HW�l5��\.bY
rcD0�!�䝻0d��BL=n/�d�`B��!�!���0��`aO�f,,��%��_!�˖q��D�!�=�'ϖ�L��)�e� ���hǷH��@�-��pQ�ъ�'�V���2��-db����a�'�A[WN��~	�T2b��'�*�(�'&��õ��&a��h!�#�����'��� w�ȭ]o�عs�H�Ӛ��'^���:k,8���8�`���'������]5=����o�90�А
�'$!�cdӐ{���@�D�!IV�
�'ܨ)�gU�>(��!��(�L��
�'�j�YV�* ��%��C�3K��Й�']��pp��I5�E����0C�>X��'� �A�	؆X�`��ؑ3������ �a�'�F=k�F�� �[9����"O ��gԕC
H���^�i�X<�A"O�8%�V$}l,e��'>�dx�"O�s��	i�E!&��1"�~\
�"OM{��"I���E( �J�z�"OZ�x1���۶�z�a_�B��"O$hE��4F"�e8$����8x:�"O|U�5cZ!P����hߩr�����"O~�Pp�O1jz�Q��U���i��"O�
��A�zMB�z�F�� e"O2�0�CRi�d��P
��2��Y�"O�<�Ц�O��e�G�}�Ⱥ�"O��HZ
@5�0$��.H��zQ"O��P�K�Nn.t���sJ̈	"OF�E&bT�\���_7��r�"O�y�QA��!�n���]'-"��y�X���IX�S�O:���׈XSQ�X�$�9w�
��'� ���w�0z�Wh�x4{	�'�"9��C�G��#�ʕS�����'ߘĸ��ē|��u���ЎC2�A`�'S\���AԚ0�����<�t���'��9b6�;?���vD�W��:�'h��2�����&%�.Oܢ=E�J�=�2p�ů��D8����y����,�yY���
P����2�;�y/Ə�2u�æL�ܘs"Jԅ�y���>ފЫwi�z#����Z��y��n�L;L�a�D�h2kL��yC͋%+�}����Z��\�!lD��yn7�`8V��P+XYB� 1�yNP��R&R�I�$�@���yRi2��KU�FDjL�X�
��Py�ʽ/|Bx9�����S� �C�<�Umϛ.�䅺U�l�a�qI�D�<��4~���S��S�,  �L��y��vi��H�c���Ib��.5���ȓI��	�?a�Nx�p� ����s�Rl/M����#V'�N���?D��!��JN�U��Dӽ&��3f
*D���6 ZQ=ܹ�N�-YJu�d�&D���� 7UR"+틲}P>� ge!D�q�K 
y��A!g�!CPl���c>D�<�r+\�:��@�r.ǠX��`�=D�0��c�ޙ�O�aH � GD=D������A���B�aC�6���<D�(i���3��1��� $*� :�!>D���l�#b����5��n0��g(D��[!�^ ��U��<,.�	c (D����A�6A�� #¢
D� �$D�4H'��/��@4"�2[m:��#D��r�طa�����;,�H #6D���"�[�4<��;L�R�	 0D��x�����=bv������H D�D��~�Ƙ��āOQbd�U* D��;��F-t�:�*��M�R��%*D����Ў&��૴b��{8<�0D�#D���3ǎuQ鉰�"���l D��aB��7����ƱR1�Ś"�?D��%k2NNU�%	)6�ȽҀ�=D����(T}��F�g�b�BM;D�dP�*K��*���/Y�<2\��c@'D�d���@�Bn4�%N�b��p`��*D��5b	�Y�	@�K��k�r�y�A;D�P�e	��)��8�����B��� .D�� NL���6Z8,�I"�ՎH�<=��"O`�(c`�c�u���<a��Y�"Ol���K�\���"��8�[�"O�y��F�Hl�:�aô=X����"OL5�ԡ��v�d؁r랲�(AS�"O���'۩s�̰V�C
�8�2U"O2��
��Dl�]��+
 A�Z��"O�L��Ł4r�&9���|@��Z"O�Y��		�TȈb)@�AӜ��"O�y���O�Q$j���b�� Q�"ODLBreI"J,��¤32�P8'"O������6�*T��*Y/,� "O.���L�`�Ec"���+NzD۲"O��0L��/7�8���R����"Oap1a��qw8@#��Sm8�"O��!��;/�@����S�h���"ONt	󇇡%!F�A�M��VI�"O��BD̑?zV$ҢF�Nì���"O�=�e
L�H�Vi���K���"OZ��d��Kl���gdͫ%��Q �"O�:qKM�nI��cB,H�z�(d"ORipUj�D�����bK�:gVQA"O` �Մߗ0��)��'6[��	w"O
P9���h4(!㞗gV��!�
�歰&-��e<�gn�!�׎	͜��wf������3�!�[dk0�2�նmZc���1�!�$�Z��f��{aGQ���2#"O����6/�]�3�ɪR�,�R"O�I�#�+�p����Fn�pV"O��q��H�kp* ��X�B|ļ)4"OX�3m	X%����̽&|��ڷ"O�L�Q��`����d�ח*վ��"O��S�D�%�4U�)҆Q�*�+*O���2 ^=oӲ%��βcJj���'P� �ŽiC� ��o��2PP��'�B�3+C-Z�T�W�Ώ1"�:�'P���R�Й^ �MHB��A�I;�'���6Fh��+M>XfL2�'�h��HDi�`�QB�\0���
�'�Z V�2�ȡqh��w�N��	�'�=cVh�$0P�)]�wf��a�'��l���NuTVsE�^4C�Yq�'8������W��N� l��qc�'L z#��V����nW,��
�'�����L�[Y�yKŭƣi~�u�
�'y�hiVJ�Gܺ|�D+ؔax�
�'�I��Bm,c3jJ�Ov�x 	�'�@\+�PbJi8�_�>萉�'�=H1 ��A�ف%�	�0�.�8�'��$��%�^P�ųD�U�0T�	�'.��e\��vDs�ɲ�'�Ly�F��?�-�Ո��f�(T��'IB,�s�E8A��Z��T�kn�`��'��Y[3�<e1�9���l��Z�'��FḄFkPY[��#/�p4J�'m�U�4�0�ހ)P$^r��)�'�$�g��R��׈�c�8(Y
�'P�Yy��<|� ��& �b���'f�2�b�0Ȣ��7 FK����'�h��2b\
a�
Ы�ł�:�D���'.(�"�e�� !ƇJ�!�����'� �%���T��q��L,m�R,[�'�	�r�U*�u�w�Ǐ^�.� 
��� �M�� �&�<�ë]�Ҹ�R"O��b�m
><�dy0V��%G�(ȣ"OP|@�CS�d�`Љ�J�����T"O����ȵ[	��"@׻i���Sp"O���d·+<�h�D�
:�)�"O8� V,4ê���"'ܝ�"OJ8��+g��52�-��n�� )C"O� �E�L� aD���bʦW�����"OX�
�H�@��%aݚFٜ���"Oܔ��ǞY�4�w-ȫ(.X��6"O\p��W�=���x����Jw��0""O���u.��[��Uڶ@�"tD��AW"Oj� �E�����ю8�v���"O�A��������f�|��4��"OJX0ǇG�X�
M�S���Gs\�U"O��sc�4<�� !A���F"ON�	*âS�8�p��!g�\��p"O`��0��4p��� ŇYF�}�F"O܀�1N��A�h ठ4 \8ez�"O�]�����1���#jA�R#�46"O�I��"ZR�Ű�.ب"aä"O�+�k��f�T%l����� "O��R`&O�I�!��B�&I��"On��!�F8JMĵ
��Ư爨zV"O���o<p��.<*�E�"OX-B�Mv��L�bl�2q(0t��"O��Y�h�*FV�;�J[$��݀�"O���IO&u�,M� @݌s�H���"O���#��k
.5�e/ �
��"O`�AAW�'U����K���g"O���l���]}tZ �3�|�ȓH;�m��f����`jŬ=Rdq�ȓ(���1'i�fLX��$�+-�a�ȓzMZ� 4	� T��4��I'L�n���);B�YA��6y�
dcT�R+݄ȓ]>&@����a@
M�=�z��^j$���Z�_�V
�t
�X��!�IQ�
��viR�2�&#2q��I1����F�*�Y+�$���m�ȓo���s��@�H��92���x�N�cf��A6���.�8&a�ȓ�!�󆃹)�$�2Rk��>�� �ȓw �m�āBDt0�c��{��ȓg�Ht�#a)m�ʠ;5e��J��"O���N˼f�\8�cnn*�Y(�"O*�`�S�,�J$sf�Q��B�	,M�~8Ѧ3o�b@�,I֞B�ɛ�� ����0�� r��cblB�	=��P���%6�԰ō�"5�BB�I6K��!Z7䉬[:� 'π�B�2B�	'������Ƿ_�Q;pG_4%�B�I�=��psMڅ����&�.�rB�I0u?@$yU��	Ш�H�/�	W<C��;4-����k$�%	D�N��LC�ɕi��􂅔P��c�����C�	�Gr�y�7�	%'�,8D�J�c�!���:����b�D�/��p��l
�!�N
<��u��l%	xt���SgK!�B_� ���c_�Srv��S	�+4K!���Gk���æZ4g���0fذ1A!�Ė?�~��j�R뚩� F�U/!�H�E�r�K�B�6Ty&�χ'!�$@5}��PMχ+o��Y�kN!�����ѓ�I ��v��+X!�� $$34��I�uh`j��:�B!�"O0hx���Q.���B�G�'��9�"O��B%��'Ә��v�Ą�J���"O�(�&f�<sON 뒠O�{��YQ�"O�����.u�q��`W�U;��"Ot�2����O��goH�>�>�¦"Oh����4*.�<3�д"OԄz@��L����S0 �P03"O ���"�-��F�~�(p�"O:����Z�u*&��Oz�<Ȥ"O�y1G燿6hX��큩zǢ���"OdI����u����"Y$uML�"O��2�.F,0P��`�*�N��Jf*O(�5�\,h�ymFjQP��
�'dj�;�%X� 0�13OL�i\��
�'�b=s�jJ�Jb���fB+Z��� �'uXl[qiR j���jPğ?�Y�
�'�&�C�ɬM��E���167M�	�'׊]��E)�����)5���'n̕�#ڼY�P5��7,/�	�'�H�Ӷ�l�DT;2�� FU��'�V� e� Kexq���,	%��'���s��3G�*�cq���x�1�B �'4 ̉A�Y����zE�\
� ��':
���BF�w
�"�эY�HT�'�l ���H�I��,|����'�\��*�`��<����:�š�'|��4�ХPB�I�pc�^8��'���+���6<2����J7t-��I	�'"$��tB� G"l��hHg4
�'�b(�%9]	�C�íc�<)��'��Rv��2@&Θ��m��S��L�	�'��D�����%[��wd��E�0���'MdD{ĮG8I�.e�$/�����'����(�"�'�U(uL�ኜ�y���Ѯ�rN�j����͏���1�OPP��U!"mH%J2B��;Oz�H��t���	�qm�����+zi��A�U��E�$��E&4SS����Y0��y��B�hT洡�{亩�7f�1�y�a�Fm�=ӷ�<�Ґsv��3��'�az�N�$D,(,P�n:{>y��B�.�y�O(�J���W<�`Ƀ�>o� \��'0����_��F����2a�����~��Z
[��!J�oK�R�9瞕��Ey�l<��<0o�8���+qkR�Of�Jg�d��L�?�Ï�,����bE�8oL|�Va\�'7A��	+B�Z��ƌh���[�O�?nOң=�}���é\�B���,�i�� ���B�<yM��
.���7�7�<'j�A���0=��dL �qv$��>�|ai5&O}8���O�pɆGɢ$X��FHC��g��OB��q?��Oޱ���'%�TTT�ӾYr �0�Q;k@��Î�d��O��?y5�����K����Q�t��6D�Ԙ��_�{]�=# �^�f�W%Z6p�<E���'H0��KѮ`t4����@���y�O����ǽO%\	 W��$�&�QA�9��8�0?Ɂ�G0�&�I�� �E�9�_oX�8��]�|Z��� �޹�eW����u��>1��F́�o��}���DS@| ���N���J�� ��ԿU$͇�*Mf��G@�l��a���"��U�'#ў���2"M�X
�ђ�ĒGE<ѻ�T;���"�Oꩉ�(�I���2���"�x��x�$0�O� (`q��Ӹ���a¶k�t9#�"O�٣`"C�7
����n��)q�io�<扤����\��;mP�A��h�b�1"O�<+��? �@��G�X��a"O�,�DD�	o,�����9 �~$i�"O�Ī_%Lb �凖�u�L�*�Y�<�7K.u��x)*�
A�&Z'�R�<��ƒw�%�$	���w��Y�<!���,���;u H�D��t�eg�_�<ɃH�.!�A@���t��wS[�<ɃKP�E�2�ʆcԀmSUx�OL�<Uh�2�j�ID�fx:��''x��(���8#���(Vl�떡��L�ȓ'����F*��>��2 ��Qӌ��ȓ"�X���'�72邬R7N.Q�Z���4oҁ��py2/ƴ\hL���C)�N���[d"O�h$ֺ0J��h8��l�Q"OHi�e�v"�a�ԮA���0"O �r��q�D�(��\L{,e�IG�O�"�K䃔�D�@a`'`K16����"O�X��ׂ@����Mrx��"O�\�ׯ�5,yӆO�uЩ�"O)��$J�G�!�s!�$Y� "OH$�l xlT)B�n�p5�t`���ߊ��'	q��3��L:3hd�iel�/j1�1��"O� 	Ae
(,N$<���g89��Ol�Ċ7p����G+\�x�I A��O�!�D��R�D��� �;kD
�/θr�!�DΪ�R�8S�Td�-��ə:k!���b�H�Ip,�0 ��H�Ǝ[P0��hO>���ꅤrb\�H������9YF(D�|�S[3x ����ЬS0-"D�x�����Ȼ��K�m����C ?Y�O�b�"|��Z�fΤ)c\�{�f� ����'��|��Y0V��E���8�t=����f���O��@lحkH�:�"Ā,�j]��'f�J�GB�T��1��D'5p��xR�^�nEĵ!s��-���aV��!��=����<I��.����Fi8A1�Z0b�@M�ȓ^���Y�e�#y�,QqD��h}�E����?9��;�!���X=J8;�%s�<1��6~����
C��q�@�r����<����8|`���	
"N�`H���g�<I�o�06I���KB3 (����_~b�|2��
}ؠ�2��P�"��E :<�.C�I�]?�!��D'h�H(�$јL#=q �'ٖm�g�8�
���CX'B^R0����@
���1�' �td�E⋟5g�Ј�ζdf���ȓ0,ސ`Bf 7�B$zQޗ`a2���	d�@���  ��솈R0g��V�m��=�l��BL�7����Χ@w�-�'P��Dy��i�7t+f��OHn��Y'	.O!���
	cP)���X`���I�HZ�a�`H�Od��
�a�j,�b��e�0�X�ӯ����T�8W@,��`�n/Q�Q'����I)dV�с�A�?�r9�rB��B��cKJ�j6��Qh�ې���q�`B�0ɞձ#*˽We`�����6w�\b��E{J|b%�ƸL�D�b��.=~��Z��F�<���F����0�=^ޥڀB]B�<�gC!/`���m��6�B�@���TX���mܓ���D�_8)��M�6hF�s6%��d���sfc׫!m��0��9>�J����L ;�HE�zY��rG˙�l~��S�? (�S,54�!�ȍ�g=h銇�d���(Oz���ju�ΧH)2�I��#0ڭ���2�S�S	o�
��Q�S�;�Lk3��6LBC�I��
Z7k9���Y#�&kv��d�<aT(�	�@(R,NpN��E$�8�!��A�l�P�o)q6P��I��!�:y�쵨���L��"�I�5����F��nC�n�>캥� Ȱ�����y��)�o4 aw��)����f����X�ȓ�:٢�jY�~��u���3,���ȓVM٢b`3a�p�aa	[�.P�I���s�@���S Yb�QD�
(Q&��MzӪ��>f���{0!2e@�l��{��n�<�'s�e�G�A��]�'Lk��ΓbJ2t�0!��;�:Ԡ��ֽyF�?�ӓ6���([�U_x����54���G|��ܤ�1�32�.ԛ"տ&��C�ɇ.��l¦��@ ��"e� U�B䉅�
&�(�:t��Ɠ:3�C�	#= b�zB�7Z�Đ���KČC��a*�� ��R�L��"����AsVC�ɛ$l�QP���J�`T�S�|�*C䉽9J�,���=g�,]�BNC�IN�%{�,�Sj��X�b�E��C��*-��+�E�f�Q�w�ݲVhC�ɝ�d��``S�tjfLk�,�8�B�I>��%�2$l�'yI�@�ȓ5@�$L��d~�E` O����'�<XQ!@I�&(�Ȃ�LZl;
�'�z��BϚzmPpWfI�KX�Ȑ	�'�RL���ͅz��H9v.�_4�H�'���A�@W
u�n-zТɿqb�!�'^]ʕ,T;�| �N�9~�r���'���G钖R��1Ό�|�"Ո�'��X��m��O.�DKV./}~�j�'�`�ƣ�4?8i��%�c��5��'���E�U�Z���/@;V~�}Z�'uP�#4fZ�5�̽���*NPP��'�t�pbOF ��Tˤ�Q�=�(b�'!��d�A
=�쩢dg^Y�U 	�'}���I?�F��!B(���1�'�:��!�H7{�u�c�Ja��
�'V )낃��:�JiҔ�+E����
�'�<��UeU��b೴�ܼ�f��	�'<���	>8����{��*�'iֵbI�"�T��#�qK^��'̔:bA�8\ty�D�S�d����
�';*���u���t�Y�Y�N8s	�'��y�Ύvf�� 4F�H ���'
x��ɘ���ȓ�]� ��'@�Ȕ�i��-i&�F�i�ذ	�'��|: �V'�n1�.
T�|��'d`�!���p�b�#O��C7�t"�'��e���	3"�`bGE�mN82�'��ur��ވ,���X�`Mvq>���'l�y#,Ĉ%��C�P�j���3f0�\� �`2>�)��Wn AЀ+AsrhP1��_	k�1�ȓ�|-�a�[�
2�=i�ŕ a6�A��.$����
;:�$��!�:nd�ȓ+-@���SsƘp���	H��Ʌ�m^���7k�)x��Ƭ�A�̅�`��؁��;�h�3� c�zL�ȓE�� �@�)nq1�K�"RD8�ȓ��	���1�Ve��EZgf]��S�? >���ל�Ak��N=f�D"O �J�j�,�H � )�H&r%z�"O,�;c%JR)�0�7�� X�j��"O��$/�6���*�#��x�j�"O�	01��%Z#��f"R+,�"Y#0"O�<H�kңYF�u��� I�Cr"O~t�u�K-�
3�c�0�л�"Ob�G�1��	DGZ#v�01y2"O�P�(tռ�H��; F`��"O@Ҕ�X�p������`h��"O"5��͙"o碈1$�8V�QP#"OF͒4f��qk��SG�6-M�)�q"O�mS�̛C6)k�#��<4�0��'���X�n��1���M��6 S-C��(�5�ǘ<��B�I#�0�U(�y�8x
�� "!��O:p����~"�(!2.3�'!j����C�o�9���W�*��ȓ
8yqpJU�D��I���_�>� Ӗ�RmB�'G"��)'�3�҆�2D�c�V�#jA�NsC��D�V�&� �D�oZii�fY t�^�ʴ��q�N��u�b��'�P��&�c���g�K�������}����à��*�Q+���$�uw� /�	���
# p�JW���y"�l$)�5iW"&ZT���A�~2i	.H�%�"�ѷs� [��L7��"}*Q��(<1��j!'��R���*5�9D�5Ù�r;�� �8f��A�s2U>�9s'c�	��K�h6?�F%��s:
�	������j���$��U���z��y��G���u�[�x�4)ʗ�ɔ �>-�S!�N��G�\�=��dQ�L��>T��$����p=�N�|�$��D�i�5�FM�ɫ<��P���Q��"I�+�0��s�P�������4,�28£�LQ�G"GxZ�Ў��l�6<ʋ�I�-�8��g��y����d�x��	Ӻx��GL�(�~�
.�>��O�Pm�&���������(���O���d�C��}Z�R�钹x���h��^w�����%d�(��L���2k��\B�!A�� �����ӆ��' h��{���`N0zr⛳svV S� ą�M�p`̈DJ�e��HN��	��I	i���LD�ZU�ga��]�D�K�"N�Kw`	�F���K"��UE�q"�����o�O<ɱ%d� D�,4�d�ֱp�F�N'W��ڰ
��O_t��O����aT:��İ���ɼ��0$K[B�sp�J=��8�;=�)I�铒��!@���!o@dm��4��I_���IAbM�x℔~
2+s��"��P`w�P�S@����b��D�9'[�I �h�Z�I!��
ԩВ��i� A�l2a�w��`�p (hq�c$��(VL2����Ҧ��1E�����D1y���E���'�Ѡ��I���Ǉ�+�V�h��N��
"ϐ~tl��KDt��!�/_�F*�,�g֛-�@�xgϜ ��%r�B�O�Q��KSJh�k�ō�B>r�a�5�$��DW�#W���ĳ<�4g�X��hY�k�K�\��-!<A��[�P"��x f�N�&��Ѣ��^��A(�g���t�R("e�u�i�D��q ���a�C�l="�K����F������RP�L��.[|�@��"�K�E���ڡ��&o䮥��E�+��i��u�~����%-.=Z�b�b9�g薻Ld�Uڒ���f/�) ƃʀs���iL�|j�E3 �b��G�ꉨq�/K�Ģ�@5W>�$�
�T��D�A�>h%�Ҏ�ħYw6�Fꀤ���󡏆�(�8@�7ؑ{F�\��l��b�Z[�a���8e��	�!��-�=p���6��G<▹#��&y��R�	�t4f]�U��8uiDA�gL	)Д�
�c�7]R��s�&��~�������v7bY�EŘ�ul^��f�.#�8�q�+[�R,�NlV.�^�Ԑ���y�	�YHp]�J׶n��]��K�݌)Z0*�,}�"���A���e��F#�~��'IүM�TK�Ggt2�
W�|�4ݒ������MI4懢�z}R��C$>�rdx�]
i��)�W��g~���D)6��L.\q����|�k-���)"<4� Zo ��ZPk�.|=ƥZ2@�1e�հ�+�.�⇃+&	0$�0���r kS,z0�*t���E���dt�i1 �J,5/�rǉ��[V�j� ���j��i�HSh�Aq U;O����I>G���E��Gc�je	�1k���3dO)X~ܕ(�fA,Q��4�&�]�A���M<a�m@0L��<p��θC�>��i��)���k��uX�3d��0�@��B@��I��Kt��E��FҪ[Z�1pv��(E�-2ԩ�ZT�m1�@��,�|�2��ѡF�l���囗1On����[  ���C����&�<�Qq.ԃY5 �hŊ��O������H!��C�S��DM� �(��n_8:�8Ej�<N��˵  ��6�
0@O���e�E(#c��*��Oy,�Y�+Ņ
�
�XÉ�=PӲp)3G�r�Jl��
A�1���{�m�0u8�a�KE�?�H�	��RռPi�w#fU�b҈)�ȱ��ΓH��%�	��gKn��5�!%���5�_)�~L[�)1�!"�"�8Y6�тJ�7C�<!���ؠ"���c�,�qOMZ�I���噅��4�q�I$t�8k��Z�] Zh��2*y:'IH��1���
�Rb�Q:Kĭ���ޡ�he����,$'az���9#�0����n�D9�m���yH�\�ȡG���4�a��%�*��E� {g�lipm ��t�#��RM�]x%F	#Z1Cw'�k���jd�Z�m��k��ء-S%Hw
��!FW�0��6���>U�T�@��Ւ��f�4��#Z%O���>��Ug]�&��)u�Y|�
����>u�@e� ���Ԇ�"I�`!��n�;���v��Mj��4��z�6=��^�e���t�Z�J�n�.�c�Ɇ
��ᢳ'\�Z���A�5W�#>�`!�:X~���ʿE92�c$�K�,�{T�X�PU�l����?��8㓏��C��h�%��od�Ջ�n̲?�ay"@�t�d�@Ä�Xr����y2/ �<X$����['b��� ^�r�H��#��]y�)�%bǘ^�UhWM� T�a��$ҍ������P�У>I�i�6xL&՘ �H�L�uM U�P����F7Jd��5bS�1�0UZ��U
�xdC��[#*�
s
�$G�L�� ͇�5Hf��B�+4�&}$-u��H'��D�lU�C��	��X��G�� G�ڝK�
Dȗ�
�>yT�qi�"q��ٱ�:��T���E��dEA]hɦ���#'�X�f��d�bEY�cE�h���[�"L�[kvDq�זP4L�ֈ9&*�l$�+���c�,��sg���\�fF�1�|O�9q�a��ϔnc<	;! 
`�<������h����3��u[7��	ɶ ���-�[A�e0c	]�j ��Z ���(Oʘ���XF�i
�V"t˶e�� �N$��S��ڧ5d1b��۶zdU�T�;&ɤir�CW�rŨa��\�9�R�.���:�ZT3��oH,0�r��I�'e,��f�8�JtY���k@<,����l����)��*�T�����s=���u*Ψ}����>��0��*X����w��0)�Z���(q8���5JN(|��ȡe�#8�QfBr�ܨ���i���9/j�dx���0�$��3ˑ	Ld��r��#డic�S�;�
�#va�MTd)�k�k�n��"�ιa�р�b�|ـ�ֈ+��;F!�ORtƋ�M�	<s�ջ`�@`2*�ɖc/	�0�k'��?/hif�B�m=\�ꀎ>w����b;:��FCլ�*���MGpaH�+��FzL0C΋2�.L��e�xB�g��26�"=�!G��0|j2K��R MAĲ�|�# �Շj����U AT� �(��BI�f!�BZ9t�i���� ���*(sU�A����P�������u���9����]OpȦ�	Xֱ�#�9A��4�U��^T~� �	 1�N	���H0L&����1�
�TOj�<�4 �Y\j� c�H"4�V%��ɱN$�S��4�u�b���7�K�>�Tm�G�`@S�q��MAf��)&0L8KG��dAw����� �E��I��yk+܈(��!he� XE��d\7d�ҥ�ROYS�X�e�.�I����N�Ml����W0u�8�äiX*-(��� D�8�p1��8O����"O�Hx��#�r�.���IX�NY�5����o$��Q,͑�]�T�Xz(x��	�"����˳S
���Ny��(�W��Fx�DIƵp���Κz������Cq�Xq�E����6��#�6�xB�'̲<(��L7U��u���#E�g& U�ў�"���v���������u�ժ7�D��a�)�Y��D\
�I��M MJ��bߕ~M�	��u9� �	/�}�wĝ�a��m>��h�5@&�1A�c�=�n�`����\Tb_G;x�����Q�^"���4C!�-q��=�`�(�U�ō��F��.XJ�Y"�A:h�J��GjH��%���F�8Q�VH�7 �uE|2�N8�޵�Q�Ӹ�Y�F�=�����h��kt��1��td򡉳�O<�Э�&��ֲ�a��8�"b��e�,��3eO
�hP��홥N*�tk���h؞8��)�l�b=���ӃE��D�%��P�ꬓ3g�#Xv&	 ʍ�_����N�8tp�U�����L<�UHW${T�F�:3�0寯E���:��	�`4�S�?������$yP��'�h�B1�i�5 �j�[��,axj�Ц
"L�`UB얻Μ����m�T-�T��#�f�{��Y�|�,�,6@:\��ɞr��(�u≓<=,��Pj]�&|f`�uo֡ިK@��.���P&��}A>���˻
�Ԙ�^�Dc"t�'��M���)/��fg���#7�6H<2XYW��#,ۮ3q@]~��T�E]�I6�A8y��Ѓv)G*�J9a��4`! ��'�9{��0�![�T���yW�ml���oL�g��k%��\�����^�65�Bh� ,��12j�i���R` R�,��1�B��"�f���O�-
<%�bќ"*��b��j���
�H�e*�L�L���$�5$���mxB�@p��:�X�i�a�%@�Xٶg���de�3���lZ�@l{@�h�HW$<�B�9�ʤA�T�V�9���هX 1�ę�6�܊�p<1"�b�*�6w'��ЄΆ[��(X`��:1�x��ND�=x�D��i��+��[�cM5M�T���狕X�� H b;8�P'����'�!�!2�G� $��a1C$}B換BO-HCb�
7�[�B7@a���DP�4%r�P��l�b � �òZup 1��������1Z. ��GF�@�	ϓ%a,���񶃓�C:��2/J� k81��(�;i0,�ȑ�/����Ӳy���6�R�J$��boJ�!f&��(V1xO��ҥ�,7gLȣ(����?�Èְ"I��s�H9jX��m
��\}A2A9<&�ܹ�&ծ
ݦ|)�J!M�ó�I=cJ��p�˔�Lei���=%���%� Sf�
�FY+Na��I./�$Ȃ�0O��
�J�X��QfL1_����6��6ܸ�'T+f�4�5�٪m��s�
�u^��ц�^����jOi��3�� �s��"܀CÌ�:|n&�QF�A'Xr��x�b�t��c�dA�rk����a+���S�ƌrc��a H�U�.`00BD:>�t�H�� ���I��<	KV��~��� �7	����Y1&�~����mxI�P�?>��=K�+	�h��F`W5��ś��0#�l����nLD�!����÷ A���?�cU�(��ca��
<�4 �h�1����A	:�������i@�(��3�I�5�pP�ܾ4��ʒ��;U��i{R��03"dBWnPe �ቓ{@T�فa��w���� Ȩg�9(�@��o0���mK�2
t(l��i�F�,{Ӯ�ѐ��E��h��j>٪�*�Ʌ<�:)s7K\U�� 
.�M+�'��qd$]%�F����&a�v�+"�@F�}Q2)�rPQJ!�$a�����v�d������P���(M��A�.\O|y0����)C�X2"� 0ʍ�a,W�p�H�B$� &+� ���rYxG�@7-I�%0�Bⅵ24���Xc�����P�$�Ɛ����28u��dX�zAd�3��I��`�4*�(�69�������3��B��B s��X��*n��-�.N�c�:���7:����F�1��V��!9��4����r��ٕ?�6H"��.H`���!k�T?��Yv\5S�L
C0��A�2$���Z�"� 7>��t�+>L�2"X�v(�=3�;M:R�:A�U�!���<� �����*��BB*��p�����9O��ra�&�ج�/��>��ͫ"o^�.���
u�����	�+�txؓ���Du���E�"&����F�;(4���Z�8"=��aq��i�c ��@�-Y2
P��Yd��bn��Z`� �W׆	��匞@-�d@Vf� ��h��Y0[��1��ak��B`� Tx�Jq��!h��6AL�^V����J0!�(А�E�@6��~�Y8��9��E�N/p130��<Ј���,ܣYR����b�2 BV���f�x [��V;�$��e��Q��N�x<�P�'��,����
�;x�\��GË{���*��M{�4T.���O�v�J���F�B�ab��x��Cђ2Ъ�d"?$v���

0CM�)D-�T��"�z��L�P�1��'�H���ޝ@�4)�6U�Bժ�ĻiF��Q�@7�j@c�(T,9�Z�ۖ_�@�$!cǷP�P�cI�l��ـS��p��yBG�E��E
[����t��YH2�$D�qO((�3��T�8�yN�3�p�!0��\�Ru��΅�=�$P3�� �����T�m�N0���C�4�d� ��Z�LM�6�ă8�0tQc�>@�B��'ʥ葃ɶ{N�uQ���	6yI�]1 �Ų/�n\Q����<�p���<D+��I���1*q�ۜ;t�Ux&���7Ƅh9Y%�L�&�Νe����M�"[Hh��D�k{��9&!�j���	^V��4��1n2@YI���*5���@ԸKN�4�V�T5��YZ��ԟ��I�䕛�@@�§H�V���S����&��hs�@�Ј�p�BKj�	���B�S͒� ��O&����F�|`��*��-/���k`��.xvt�����6�n���_9� �◧�-zm��zc�G-/��{p��xv�u9��˗_���`(��=� !$��T�u�m�h�,8�(�<���í0� A��'�Xq�)�#,��z�g�d"�k��H�E����NK.Ct�uBF�=�@y� -��B�%c*
�1�IF���J�oڎ:|��c'�RP-0 @���hܓ�c�MU0{�x��3�]�*�ƬQ���p�J1��k��'Ò.N����m��eȆ%��ԏr1*�r$
>�"D&�١(�P�HGcR.O�ȋ�Mödˎ1��J]Rđ��DN0`p����<������ŝ*=@�Dc��nzV�C�
�	LQF���A�S���Ձ�u3*�b`�BQz��vc�\���C�� � �@�+k=�D����2t0,�z@��S�'��q��՜P.��h�+Эy��C��I�qCD�y5bȋ�
ъׯ�������R+��H�됭y��k a�t�i�R���d�H���}q	�*��*]�*�@�P�V �7�
!�� 
�e� HT<�0/K<[�h$�N7m��a���S�!����	���l�f��>�7e.J>�4��Ǜ6h�Ip�)�z��!�wl�lV]��C����鉄N��3&�iRMm��h.p�a�;f������ڶe�x��G!��]�A�<�юBq�;6���c�"���-�d�O��#p�ё^"X�p�B;bS��{R��*�F�[�nـ���D����!H,��	�CN����0�mQ=;<����]8� lZ�ľ!�W��|�+�hk� �kߟs�4�p���6�8��������1�'o
�E��O���t���������]�T����Le|lb`
��.z����	�?�Ʃ��в-��y֡õ�7MX�tǺr��0:�8���äVM���[�SŬ\���{B�J5p��$ ���)D�� p�����8�MZ�(6D����J��p:���c_���b�:�,G����j1�EQ �ʓ��)c7ҵ��&���T��@��li�NiC4=����oM��1���sD�A8�I%��5$P��/tzm�r�[��Iv�B:DT�ȓY��Qa˂ *�HY,U ��=�ȓ���������V!���G�6cq�ȓi��k�(T� �Dgm؝� ��?��1���ܺ#+@M��/Z|�Ұ�ȓ	V�ٺ����8��F�]>)�ȓGT������5)��1	�ͺ-^���ȓr��C���r6=�P��l�ҝ��Ov�hPaF=�̩ �씬rr0��[8�P�bc�2@�	����~p@م�E��H�q�P�A	lq�cސ
�)��G�*�"e�E1 ��/Ύ�R܄ȓ|hH@� s�R��t��81:a�ȓ�f	���� $���Ȉ��l�ȓv׆ђEIV5b��q`��vdx��� ��a��^ߒċ�e+κ��&��{��W2Xb�{��%y���ȓ 4�jX7v��xc��X�V00m��a�x�f�<o~��s)4����ȓj��|3� 	�{v�I�al�O$��ȓR��@�A3Ze���3���p&D�ȓl��W�X6��1A�͗%�0A�ȓE;^��f-D)���n�!W�\����V���x�d<���G�=��0�ȓB�t��!�ψN:�!;�%^w/�����"t�/�8zqJi�Ǆ_�DR�8��z��5Z%ʲ�ļ��Թ4Xʥ��S�? p�3�V�I؞0y$���t٠]��"O8��p���B8��C�'p����C"O� �	Z]�p-Bc��;���KP"O��� D� ��ig�/X\|)�"O� ��U�	�R���lQ+�� ��"O����	����4� KX7�v���"O&ݙ6�)�*`�@+�$J�H�Xa"Oz���J�M��P'���Y�8�zp"O����Q+�����\�r�t�@c"O`��cD�"gD��JQq�y��"O��`�*��[��5R�Hո}|���V"O�4JѠ�#59S�MS�V<�P"O��w�ִPw~( �F��=}�mR�"O�\���Ö2��!6��9h\l)��"O��a��N�N�\���'���jv"O�� '�Z]p%p��Z%,>\h["Ohe��K��d)�"%��6��:��'�@���M�k���4l�����",n����\�6��C�ɫS�r���͏;�b��'��h`��O`���]�ic��*�
'�':>�x�iN$P�N0a��#.��lHu���
Uz���ˌ6if*��!6<u��x�'g�E�6�3��I:X�0KD�	� �*ucJ�wr����i
<Y�@�O�w\�ԩ�@����`$c��B���H����Q:b���t!׮X��D
eb�OX�x�Oӄ_�r��)��m<0qa��ipج��(=����G��9��A�	�'(6���Xr�\�A�������O�ęcV�-ʑ�E#�ߪՉ���G�5F*�s���N;@���	�
�!�ĝ	c�b��R)�5����$�������.!")�b��Y/|9��݃	a��r2�1Oz(sQON=^�L���Dx��'�H�	!��E|�oڏd+�=�׉D/?.$��D7���2h�|�R 4�c�A�6��z2gݥ\L�	��y���QGO�+�ēY�6�s�.ޙU"ळ�K� �"����<2��1��J!vT�@i�B�Rap��l�)���ɢ�r\�P�:�Tp�L<U�d� ��أ��f/��sf^*}5^�3���KxJ��"{��S���T7��afo�>7����բA�&����'Θg���k+�H�$/��ם<`�8x1�%�1UO�98�J�'P��0R�CXbK���NdB���!c�(Xq%G0VK�㞴K�+]�;F�T�D_m�`�x��5gH�b���#}2+�::�GA�A�
U�n.woʀ�qň>B��9Q�AڜGG.%��M*]��s4X�G���>	���jt��7�~@#�h�a~ԠAA�Se����<?�q#.�����;l�AK�σ38���Rwr��f��lP�h��$?�-r'�.8Z�G��5��<�'���Y��?�$�@IO���?�y�o�&2րc���!g24��ʊy���0��M�W=`�3-����ϙ�'0��2�u!ť���5��.x$i �)ē\> ��NK�b����GSR�N0���j�`�l�y"e�i�����3�t�0���:	�!�I=0#�`%�"��LᱏR�1��b�S�d=�����,�Ac	<2$�`"Ui�O��#�#�<[�"u3� �rw$P@�C�P:R��嬓5V �Gg�<Y�/W�J�N1��C����ߴWZ�+���/Yt�Bp�N�?��m�W��<cH4�%/c��H7xST�+�D`Ӱ����qr��֯*{��A&�
�S Ҕ`�7LT��c�<Yc"F�(e	�Ύq@�E��O$Z40�M��G �+HV@� �9f�����D������x�sf���)���"AۨNZT6��.��e4S�8\�;*��A@'{�p�g�Z2imTԊp� sH��}��9�v&n�g~��0�u����K��$��u��\�L�>�K$,�y���x�
^�",�ي�R=Bϴ��')ʊ���H������!�%ѱ��Q�D��f�Ni�]`�"ړ�e�|�Bٌ�����W��A�5�5q�a�=찝�k�6b��1-Їb��وnZ��|;&P��c'�ιmd ��c�Y��`H�';`J0���,(�ԥ4Oټd%8�XS&���1�PD����eW�ȥ��Q���7�sȜ豁?F����3���p����M ��$�m���I��:>|���)��xf�|8�f,e��7V6Wkl���L�Gb&@��L�zXheS�&��|a�l �6���G�4Qf�VGf��t�̀f��l��ֶ\Xfy@4��N&�D�8.������,OliX&�"j�dQ��ߍp{�<;�C%�j-���V�d���P'J1g4��1"-W�o�~epV�^tq�'�n1:�M'�p�Q�B0RXs3Hߣk��Yr��$,qO� ��KNi��� ��D��3&H�~ ���
�>c$��&��yƚ���A;�$4�S��'� <�c�R�m ��'B��B�`)m8�z�G#*���.OB��pJ������ٓo����J���̹(K�`���6�W�ZPB�$���v�^=gVh�@�p��+�a��o���؃��ž ��53W��A���ñK��NRD�Kr��t/(1T/?������!��!7"��yg'�'�Dc��\�/��'�W �p?�5��^ʐhA�A�Z�B��E_f�w��!>��nU�orJ yA%W�xO�ty�A�_�X1���J��>UI�BZ�[�8e�5� �Q�á(�� !�5�%��\���`���`�8G�_|���m�Y�,I�׌w��I`q�ʿ:�le����� �A��e8��x���S4^[D���>OT��Q.�5�,m�5Eňy�i�W�T���d�0��6[QV����{Zƨ�a.ڥ*�k`�jY	�t)�6��x���]0X[D,�<N��`���\��1�u 7@���$��H�J���}�x���{�T	����+��nԷaJA�� Q&�<ȉRHߵMa~�� %���`�,���H�a#@�["��!ˁo�"Q�.U1mDʅA<�<��S�	�F�YS�^6O�\��?;���:,��6{���4�I*0�����6[K������}�p]��CޒJ���l[�@���c���yQ�`�$N�Z�yf�A�W��yG��WX���Ӭ��z���P
j,@���}����Oϣt4��vBջ;�݉c�|��<"wC��l!Z��1c\�9�`���c�6Y��1 �J@^i�p���O�hC�eZ$Թ$�Ֆ	7����#�0.����M��tJQ�Q�P��0��ڨ�>�i�H@�7%��7#��ʡ��T��PU�� [c�p�jtg�6�Ȥ�F�E(�]Y�'jl0��I��,5�!Z�
l:N=���Fl�F`Χ��8��ա\綤�4�Q�z�L�����;J��u�*M���=G*�Mp���n�j'%�%[��3���-�@�Y [H�3�Ӓp@���¨D���A�;c�01)W$ȏ-�F�iP�"_^�+�vL�԰"HE��4��GX&Q�R�� jM4l�Á���Mv�MJ�ND���0Y#�I�4d���hJ����	V���TE��C�A0y���c��b!b�YUdA�?����K����i�bW��$��?JP��$&N,23�]�U�K��p��s��*����05�}�3�T�O��P��בp��j���#8�j���B�gjt�Bl��|�����V)r2��'/�T)Чo��?�r�:�G�b``���~����-��3�t�ޞC�r�b�!�!;D7��b�N�����[*�т$�{o �@�I�>9�����`�*Ex��'fR�4: ��s���M�,!�Q����H����>�B��Dn�U�B�M�59��c�T�O� 	#I>��)���6�aԍ�,t�>�ZC/\�%x J��A���BwhC)1�F��U)���8�Q���.q�$�"�T��?���#6K�$����$J�L8a���	(�)B���y�DY�d��S�'&��qC�������w9�a@�n×KkX�	'xzt�C��U�(@�t&�y.Ё��ƾ�M˰ꝅ(�Ȉ��BO:��ȸ�A�N�nԣ"@����$��x�'�I� �G$a8�my��׉pZ8�V!�6r�b3oNVc�c��ˉY$2�E�*3��y�&ϻܲ���� `^��"��NUk�;p�J](*�5���e	�D_��	M:@N, �Ajk��-)��J'/$�!�hȆ9RYYA˟�5���q���v��p�'OP@bPÝ�=L��AOϖZ �k!D��7򣔜��@��A�JZLrP�"Ô��`o�G�ԍ ��ܭ ʀ`x�,��B</ Ѝ0�C��&΂xH����^ S�m\��ד`C0 qVL��dl{P�Hf�t���Nq0��7�ayR��5*��� �#c���*w�B�^qs��MLJ�ZJ�,q"��A������Ě�d���"ߴ1�� �ٟP+�]�f컵��Y�&0�P^6��E{r'W��~��u��$p��V��e-Վy}`��f��q�	�>���S���o��i��c��CQKK��?������APv)�<����'�x:��0p��DKBoI�"MN�`�#ɺ+�ȉ5'���K"dՉ5�r�,˱s��TSω�&DZ�03�� !P�1��������;&��A������?�w���ڔ3�l�zT�1����R���i����m���MG>i�Dy�K�W.�K���L�f��V�t٨u�*~�1H3��&m2�i#��'gd��*�6H�)�� �u�VY�FG),��d�퉊!���奇0��L��#FpOp���=YOn�qs���[=f�9�ǺY3�ك儆�4��|o���ēxԈB�g
7-r�  r��!9�`�f�Wq�'ݶ���@�0�ꈳqb؝_�R��W8.0,��)�4},�M
�!܋d�r�oZP:!��υ�H�:�k���.q?^dH �k�V��t�C9�n�,�$Ӻ\��pcԞ��&�x"��)?
�qRļ< ɱLs��,�P�lH�Sb�-Cx����,Q�B�9%�F�;&��*��ǙiR�
�l��R�h�IN-��'KRA������¹}ʎr�d����Is��v(�P�+��A79����شe��rªN�p����m/�z�R�it��t��&D�I F�"���ڜ%D����]]�r�H�쌰!ج�q"��U�ـU(F���-��&C���E�\�z�x�L�1#ޢ�IR���[~<9��!�
roR�6�].�!��� �9a�J@����+�0Y������=�4a�n�@�@�R���!q�^�NV��fo)�:U��Йh!�h1p��<�HE�e�N�l�Ї㉁ ��e�V8���{��7P�}�n����� S�x.�Tɲ�v��@JN8$��g�.��aɡ.��	�ꐃa`2�$�e(HK��.+l�U��AOK��]UЌ��炜8���@�D�e����9+s2ȁÉ\��B  � ��u��t�V��gl�e̝��^8A��� שŚ}��y����.&��`X�t��9�ǄV`L��AC�\���N@�C�f| %�D<(< �5`y��(��\��Ĭ��%$&PD3�K�Xː�1�Y����Dߤ$V��!5) �h���*6m�.(���xr��U�
􈆈)`Ӳ�B�Ȋ%L��%� l���b�-J,.���8d�W��}j8 `5
��gw�,3��')���됒f
ӳ'��Pڤ=c���@NX)�Ȓ�wT��J��
�[dD�z�61�+{�`!0A�=CK^=���S2q�'3^aʀ
�3������oqJ� �O�����%2������G)HH�V�9��uj�-++~���Yj�|�2v�Σj9�����)	.�m��O�,f\���JK�l��D��nR|-kpvdZ��ŧ*
 ksn�/5�����%�LHjp���3��Y�2��jxfL
Q��$ (
C�n\6(�L�RH
7(f�[FN�7�XTa �'�J��aH'���a��|��5[��ٙ}�H@�
�3�L�7�_2$����A�' �����Ηx���؛~�\:�
Ywp�<x�$
�Grr%h�l���0<��e�*&Y"�3k�9`�:�%l��4]�-���N�7je��ϓ!Sh���#�P����:�:A"BEF)�<�<)J��	w����|�&mCWE�z���3��m����q�N�˰�#�qPO^�n�`�l��&i��� :���RPm߯b�,�0 1��"9���r`-�o��db�i�5~��@����=S�M:V❧%��D���%];�Ā�ś'e$�y"R)H7{��l�C�8Y�I
Bݦ�5� :t�0D2xh iϱ�@�x��	#$���S� �L�؇���3�6	�TN�EyP�
�h�|KN�R��0K���x�'U�6�B����+1�8)��N
AsF�RH�y����E)���ĖvJ�(I�GJ�>#��I�"����~Z�"Q�lNjII��ː!s����Z%�H�)a��p�j��Å˚Ϧq ­E �8�I�8W��AA,�#�\�EyB��D�ް�4�3z�N\�s����y��ͫO6D%��HD<������A�̔���1~�Rp��i!�t��܄�$-� km��z� ̶|�>ظam�Mׄ�[�'�܈���n��i�A�]�Jd���.7�J���P�I��m`�D�.]3��*cʕWC��D�On��EcL�1�\�Y�d�H��i@��ʍ�N��	��n<\��#ͻp��O��Yw��ʽ:a����O��8P���7)�`m@t��a�����ϋ�p��I�b�ׇG4~@)vh��>�,x��6*�t](�C�d���қw��`�0MC�m�p��nE�Y[�ؠ��η� ����+�R�lڦ���#B��)cx��?�&\� ȧ�6�I���=b�1�V%�LAR�s3b��Wc���zy��@	%�,�c�[��3
�6}Fo�/ɨ���k�?Y_�4� oS�b�P��R�	Z�:铵eɱ�&Yjfo�.ͪ�ȕҽ]V�(��/R8j񖅚
z�m��F�*�B�a���kQ���'Mk¥�=�,S�1�D�X��
7� �#ݖ~���Aڒu�q
q:�]� ['� SM�:�p�㝖�%h̓3Eӆ]��#_�q;z!���ɉs:9�
Y0n! ��A�WR�o"*���o?炴x�S�o���f�>�v)���+9F��S'O�]���3#�FWX�!#�8w� ۥ�\;?�,cD��3T��C�ϱY��9�C㎰B^�@�/�Љ.)Kxu[AGϊE�h	+U@ȕg�^Y# �V5q�xTj2W�\������'�S���: $��J�؇�]d-��2 ����xґՎ���Y� %�$�@�Τ�D��'�ܟ`%��p�x�g�V}�7�P�j Qaۮ2x�!�@�����H�������UI��(�
V�hP��[.2z�!��^��jY��!�D
�!�OD�-��p�f%NgF�a��eH�@�`ј�J���F�?,θ8�	]�A5Nբ��ln>�R��1'�H�Ԭi����f��*��<3��]
@9P���Lޓif0��H
d^��Í�	B<���!��n�qO�����I5AZ  ��O�o�@0��O�	�Tkte�cE��RgVK���+/��K/wrP4Y%$��et�l�RBI�eN��w��VJ � ��M*,���ݫw�9*wn֬VR�P2M��F�v�B1g"q�h�B!E��$�ʨ;d�({�'Vl�μk�2g��Z��ƥ5�d�1E�r'�;�M�# �`Dj�V�W�N�h���f��B��F�7މ'(&aa��96t���!8��Y"Ӕ � @�#!� C0Х
�cK��Ĩ�;<"4Cݪ!;��q�⒗�@H��F�6_΄M�C�Ɲi� �as��\f�q�eL�=S`́��I�8�RMR�
L�BI1dM�aSTd�3�G�_0��H�T�E� J�ń�<jj�5ø>!fQ�. *�i3�Я�B8�R���#;6H+#���g@,R��(���@�HO��� �̨�M3#�Q�T11t�A���q���u��ՙTZ�I'�;�CD���Dҙi�,�PBLDK�������G�{��4�C}hA$� ����=1�őU��݈�D�d"|b�'��4	wl��t���#�׵ $^�iH��qŔ6-V�Qyb����L>1"�,"��Ւ���-�hR&�2!'V��K,M�,��ڒ�|�'�
�y�-O!`
@�i�H��>H؆�ЛV��
�@T��6���-'EJ���υ�8jX�qŨΩ���䈉7S��8@�͋;��zb
O;(��ib�W#J>���c���=9���<>`��G*oӎu8D+6���XF$�(=rn��F"O6�1h�xϦa
S�J�Y��Y���E�2�9�S�?ΐ��E�̥8�P1 �F�l��C�3~`jXcwf�1
���æ��
��C䉾8�f�+Ռn�Ԥ�GĀ8��C�I�&�$p���ܸ�����"�>V�^C��s���8P�μa�t�FG߽Xh�B�	'L,P�{ �6bPSvCɾ`FdB�ɰ,���e�N�q2#K���"O�su���(]"�g�mM@!p"O����k�  ��Х�� ?��3�"O�	��Y��i�pDDg�Xu��"O���.S&GS$i*A����
�r"O�x���<d�t�ը6���P�"O��㶧,� �c�΄%@b�#"O��)BNŴԖyHt�»,D,R7"OXsF�UAH�Ёɕ�/��h�e"O�� PI��J�� ���5��x�"O��`��կx%`��7F�
W$�97"OP��[,e� I����̠�"O>�`t,�%X*�Y�O3xҤ��"O�0�)�6�vtQ'lA�>���"OBй�a��p
t�	<g;�H "O6a`�ϧA�*L
��B�T�0�"OB����>}>H�bG� S��#�"O0yb��I1H)��:��F*'(��"O~����{{6��qi�!\La�3"O~�{�A��xk�x�Q�f$,(�:p
��G&�p )���ROb�'� 2��F�N;N�*���l޹��
G�l�딍���M3�!PC�����t�BUp���q������M��4I���M;#���"�:�)7��lY���<*���9s,ȍj����wJ��M�W�Q�=f��A�Oq��Iz��)n� e�E�ǜt���h��yB5�)6[u~6�W4�)�&� �ĉrW���]yJ�:(	�Kbܨwd�˓y� Xش���'�1�� T�AT��	����� q��I��Hp����(a�DBL3
8��5(�	q�\���N�$�0���\�Bꕺ}���S�C�T	8��0,?�)���J�
 �`3�m� #�X	�⃺�P��i1�)��Hp����>�b)B�A�)xs����.;~�'���O=�ă����+��U�V��a���ɠeM�Z�0QeOE�gx�I[Ԁ����'*�a��U�̩�4�����'!
��tnM'q���O�>Q3�V=~�r qc%V�8�-�q�1�h���
G�7W`�������e�J�JUZ�H({q�j�d�N]4����t��n��B�"|�*�*8 �
(��q`�	�OF��҄`-�6mU�4�<	���vU���	�3���Xt(-@w9 ��[�5�26��2��Ȏ���|㤆<�V����F�f-� ��[af}�Bձ�?i�H�"C�L�Fv�V�2F%���'^���WB`�`�_�f�lx��#H�ri�`Dvy�IR |VL�ç\7ꔎ˕K����CY! Zte�-O,A�Vb�e�lم��"|�d��O�J�q�VqLX�w ��<���>Fna���U~���_�\����N� �Qh���eo��õ�O<�U����[�f>�Zg�٣N�|� �ƣ)�a`���/u��	GR��H?gJ���c��x)�D E�o#��{����Z��@
t�D�𩍯�
m��(ѹ	�� b�O�;l�	"s�	�l߈w�&���^84�p�WO{z̑�O	!�d��ߔ�)��.ad>�S��[M�!�$�M����N��_(�l�bꞦ}�!�D�<��\8��U�d�PC�O��*�!�$B�)��CBC�5�����$R�3�!�$�vE~���˛"f�l)�2�DDt!�DU8NҀ����w��%�-�>Mf!�$2Fx���bbʽs�th`.ܤp!�$��O1���F!��o�,ph�Ƚ]l!�d�=w;�Aw�[�-���&lW�<M!���~AڄI�Vk��aA��[L!�D�-7&�1���7!YЈ{��G�_1!���?�p��w M:Gp�nٻ` !��4l�����i��%^В�n^�(!�D�'|Pt�!g+�Z�2�nF�T!�d��"�F� �Q>z.�W �904!�ߟt+�	;2E�.�Hl�E�J~!��ؙ8����`o��/��Hq�h�=a�!�Ē0U3���4�{u�*��� �!�ݖjS��[�9hN�ʕ�%<!��&[��$�C聚YV~��M��k�!�DAl�����jNN�j�
S�!�d�1X]���j��
��Y�)���!�0b��z��ܼDژ��S��r�!�D	�#�^p��!F+�F��vQ�P,!�)/�x)� ��%l�҇�H�!򄟢ZK�qӂ��6(z�Ȑ�^!���r��e�JC��)�&�1�!�2K��tQ� t���&q�!�D��H��X��g�b� ɓ�n]�!���ba����%�� �̽+!�d�h�^ir�A�)e���čU:N-!�d�[��#'�QR��`��7,!��+ܩ`��.���[���6!򤘭-Q���G�8�(=�(E E�!�$ĞfN�����rY��Ns\C�I�P�``�2��19B]����DC�� )�� �bEppV�M	GkC�I�s <�y���-1�n�ô!L`�B�Iv���ˤ%�:�w(ǛSv�B�1��-C��H��J�8�C�)� �	R�E�\BͺW�],!� ��"O�QaGD��� l ��S��zA@"O8xi�^z���ɏ��ĕ��"O,���@�'����&ʃlf�[�"Ol�[(�Q$8�֠M=^�	��"O ��+J�Z԰�
V�~U�|��"OH��Ɓj6����Z1�	�"O$�KR�-+޴B'o� ua$"O��u��=g@P�MG�8�L��"O ��� yD���3̃�Fl�h�"OT�" �):~��
�Y�Qd��b"O�$���81��a2NO�_�ȱu"O�8�E<w��ԛ���UD^)�2"O�9;s�ݸ"�6aJ�M�~Z6�Q�"O��ϰmz�T��M�:��jq"O@x��)R�t	 �̼e,i��"O��P�]08<hy�l
a0�x�"O�ejg���M��D2��ܭN�H�R"Ov-"SΆ�b��̘2?c"��B"O��S�˅���R+؇?z�h��"Oh�2��Ѡ.8�8�]�:B�0�"O�ժ��
�HH�iRh�,F��"O*����ʭ<�~@3��B�VT��3�"Of����,5dX�%&�6E:�"O\y��ǖ�1��%��d�2#3���"Oش���3dU�����X+Jm��"O��KH�,>�BA��[I�m"�"O�i��a)\*���#a����a"O<�K�k�u�5�sO�1^�8�"O�("	�?jZts��O"���"ON�c�d�/Wz�Huo͹t
|� "O����팲��$�ٯ��$	"OTT�`�H�R�D�ʁ��)��,�g"O�Aɔ ]7莐B�oRf���qp"O0�oS.s؄P���t6���"O�Q�E��9����ICYz�3v"O~��0��}thQ��J��0Z8�@�"OV��υ0wX<���G!h:j��"Orؒ`�	m*7�D*A���Q"Oƀq�׊:&���gd�]��P"O����ɀ�9(��e�Ĝ���z�"ON!j�D�[�0u��J9)�2�k�"O�Q@�ʔ"�=c�.�?X�np��"O�<XפA�8�����BC>F<��"O>�Kqڝ{z	�!N?���V"O2@;e���`^Ld�&��#y���7"O��9p��<,l*�O!YӞ�*"OF����9����W��0���"O�+cF�4VBb��-�b�l);"O�%�G(G�L�q�b��p"O�����$=�dm���
�`vD�0"O`����1.p�0�R'8����"Ot
t撀-DY��G#-��a#"O�h+ǬJ�Gy^��t��^ԂD"O���tO��� �+Yt�x�ٵ"O��C��X�^8a��]'xHp0�"O���jx�Q�IÄ
�r��"O�P'�Z�4�f��u�U���T��"O���J�O=�,��I *����S"OH�`�Ӳ( �!�� ,v�x�"O|�sd�H�XUѥ��'gj��@"O�I���ۧ�P�&�ʔq�X�"O�R�M\2�Rx����D:0Y��"Oz�8̔�b)J5����$��"O� p����9<��mCfM��|��D��"O�t��!a�- ҍ/m�d x�"O�A�`�2wv�Ѳg�]�#z�M{"O�Р�ƛ�S஝��Z�g^���"O����/Z�H��qOF9 iա�"Opa'용f�P#�Λ(X�^���"O�=x�o�4R�1�3K<z6M80"O4��3��
0��h�;Oc�M�G"O6��R@�h� R�܂+O��;�"On�2�ެc�6TӢe�K|U��"Oz�BӅy���D�HH��2"OpLz�)S�f���&��
���Y1"O�<i�H	���Aǉ�(|���r"O�Qg"ŋz�6�)���(Oh�P[�"O<\���#t�r-�ƧtY���"O�S�@݈&�|�����+S��`"OD�#\�m��@��^\4��Q-
!�ׂMh ����X�Q�F�^�!���h~ ���M�:k�y��G��!�� �l�F�P򮗀S�d��i��VI!�$A�9R���U��(>�ɻ`	Ŗ=!��\>Ɋ`��A�34
a���4g.!�]������-�i�x��m?;!�d��" ]�G��()����mC!�$Is%�{G�\�|������!�YM��(��� ���j�$^4�!��R.��Z7�ݬ�d#��ϕ\l!��Į4����̓Y�\]r��fo!򄕺�)C^�~��@ !��7s!�J��4�"�5.(y#�lU!�d�=0�X,��l��u�r"�F!�$E�]eb�	gծDJ���@ɶY�!���M6�ip�n�
2҄�@�"C�!�C�r@�����s���QHL�Y�!�8L4�9Y2L[�0y� ��G��3�!��D5��a�E�EwR���懊%!��A�b%��c���?R>�뇄�!��R]��u��!mC�M�e锱�!�'%0z�J"oJZ���r��U3�!��j�D�'?�v�p$_� �!�$�\@:�#���$���/,�!��>$I����4B��`���*�!�$�c�n�X��	W"*�#%�9{p!�d��y��2A��4^��z��N�To!�� Qs؝���)M�`u���,d�!�Dևu҄���>����@=E!�Ď)��
O��v��吰�R�3�!�؁S.�%���<����'�53�!��K>.����0`�$��� 3�!�<zb��"ڙ0{�(6�^�!���ŵ�{ �W`Ք�(UK��i!��I�|L�QB�%�(�2��d!�䋢8��\A���4�f̂��O�
O!�&^F���,qo��i�=Pg!�đ�b_�,�S�G:4Z��6���t�!��d�({PC]�$,��{r%K�
�!�D�1m*���H�f+��c�M�1w�!�D�:��@��aQ ��J �_�!�M	�R܁� �:���2�E��S|!��M�rm~5�EM��s��tŚ@o!�O�}yp	��vA�5��aF�zk!���,��s�&#`5@@U�Ŋ,O!���Y>�����vø���捽S9!��j��J�o�/�8p�1�7nC!�� By�b/ݍQ�֑)Њ��n�z�"O�Q��K�K���U�q����"O:�����b߮�J���5Fi~���"O�uȂ�ՁH�@)gD�	M����"O��m�ȩ�FY�/0>���"OzAP���E�l)���X�y�&q�C"O48���ͅ(?�xb��0"\�R"OQp oMV0
x���7Z|���"O`A��˄)d��@!�ˉ!���7"O|�z��M89�P�C�!n׸�ʠ"OP�sb��>ޢA�#��<Ȧ�
�"OJ-1��M����s��C��^��""O ��E!V�C����!S7jK:(��"O8����]�XuX��b��b�f�� "O�aq7�K oWJYJW��j�Lt��"Oиs���C*���bO �b_�9s�"O��7��Z��DaA�F=)���e"O�ۇ�EUքx"�̘�7/�D�!"O��0�)2J�1�k	�R�K�"O���J��0�4����S�Z�JP"O��*�l�a��&�4}zZe�6"O~Q���n�~�XgؿX Q��"O�9�'W�|D:�`P?Mrd�B"O@�[�j��E�!OZG6�Y�"O"9���9$�\�`�-�uĴ�S6"O@�p��|l�ږI]c�ԁx"O\xq���z�����0�$�I�"O�����V�
���i樁���۴"O쌹�g� 8�D���J	�^t0A)"O���   ��     �    �  �+  8  D  ;O  �Z  f  p  �x  e�  �  -�  ��  ��  $�  g�  ��  �  d�  ��  ��  c�  ��  .�  n�  ��  ��  ��  ��  5 � �# $+ 9 �G UQ �W �] Ad �d  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|`I!'G#\���%�T��'ItcbꀀK<�k��̥:O��'������Ǝ8�ݓ���"J�S�'y`=c �d���	%�BPiV��o�<)E�I�M��c�Q'��I���k�<Yb�`��s4��/~�����M�e�<Կ��رD�E�?�t�Жgd�<��j�aZ����Aّ'�F�r�b�<��"���e�ďfe��ѣ
�[�<Y �{�<Ԑ�[�0�Rѳ6aE|�<�ǆȕP�,x��H�o���ۀj|�<��\��!G	��lhP�qI}�<�cێ�,����ޣ��@�#��x��G�<��Fъ��u��Z�JQK�%v.1���� ׋� ^:�Bэ]lr"�&���I�-4��Bbʴ9[��g.A�$&��$@?�vĥn9zt�&D��v�����Z�<�5��@e�
I
p%j�a�L�'�Q?y[��Ph�d:�
�Z�bg/D�$2��q�HÄG��R����I�r�����䕘!��8r@�P�Fi�	� ��!��̲��u*4%#\l􁦪��,�du����	�j�����
���k�h�7EB���˃���.*����u$ML�BQ���C���C�I
|����d�2�y�e#Q�B�)� ~�ȠB�-Mx$5�2�	�-��a��"O5c�CO!	b�l� �, �6�q��L���Ovl9�֥��d)0䢧�L>"���'m�M��U!:��fG�+�V\
�'�0yVLʱe %[s	D�|�Je�
�'�|+��D�n��k��K�i]��Ėw�6�R��È4WP�W�n�a{�@���d�ONL  +N�Wu8�Sģk�L���"OH9SC��F���
cY �b�I��h�P!���2>ƹ�'K3c
��B"OFS%��-I�2L2��O�7�`�ARR��E{��ɚ�)�\��&�0f�p��f��7Y!�D�Y�`}*��P�Z��qlk��$��Iìb�Ĉ7N�6 ��2t�C�I-�̕K��>4��7�vf�1��'ǎ虂M��h�p��wȝ�"{*(Î��~�TЊ�$b�!U��9��	OnOf�( R�'�v�Y�	����Dоm<4��'f�#=E�D��A؄U+��τ$�6\��a �yRJ�;��"��ڝ�p���
S*�y��B�.b�SCB�3���݆�y�a"\�l@�S7d���'g�
�y��ص�i��	U3�M�t��%�y2d��ch��@����G7��F��y�-�%�<	��J�D�~|IƆ��yrA�
�0ճ���vL��5�y2I�{��$����q`����&�y�O�M���b�C�|�a�'͛�y2
  ;"d��`d�s̤�kFй�yr�ñ0�dXT"����@��yb�[�@�\M�D���m�@�%c�y��Z�U��ȁ꟬lҔB�
��eNh��<�O�dZ�.ڃy�:p��a�O�����'�>|�H�؋tHY.�N��7���6��M�aK����'Q2�'tN\��cĕ^���w�\%�x�
ۓT��	A?!S+�81h0�SC�ŕ`�v�aƯ�K�<��O;VTJ�hT*O
̙�6i�Dܓװ=�������h@�K�%K���X��C�<)A�ːa-H!� ���Ƭ#��C�<y�d�'Dx0����*Ms��x!@�<A��+eHR����<fW��%�;T#��C8�p�F�π;���[7G�=�M{7m<}��)�S�#���D#]��9:���Q�C�I�px���ē+g�5I�M���c�d%��Gz ��b��x�D
^;��x��:�xҠ�2q���PA�5$�)�b�5ApC�ɔm��Ȃg�T<.�x���Ȓ��C�	$'�I�%�	�36��%뉌q:�B�%o���e"Ү0��e@����sSn��4ʓ��J����H��I�fb����ȓR�`1��/=b�Yu��JJ�=ۓih�c��4#^)�@AL�/ؔ��0yN!q��EX� ��ƾ�0���y]�b8`�r� ��C:y�Ѕȓ�
�@�[�:鱓�Sd����8�fl�7�Ĭ[�DA�%��*<t��ȓT���*bdA�-�"��ҊZ*e/� �ȓ[���w�@S�&|����JM48��_N�Ц�T�;��I��V<RVT��Mە���<Dht��/͛�\�҆��@�<�4�ˍK�����o�!_����D�z����>���3e��tJB�5&Q��,`�<�rlU�!6�2WͥB����gZV�<�V0�u��
8;|*mѦ��z�<� ��4�Wp����#oT�%��"O�9��K��c�6}��ˆ� Q*� �"O����FT�VN���c+�8~N �p"O��X�j�6��l�g�49|��"O
���dY�9h�.¼

�R�"O��A�����@�T$�u^F$�P"O��Cc�V�x,�¾�f�B�"OX �D㈅:���D�M�4�.�@"O�IC���}�D��#^$��"O��+S�_�u�~i��C�ZX��4"OF:��,d^���c�Ⱥ|꘲�"OH�bq�^>l���m��p)�"O=��	�i8ȱ���N���G"On��FɊYʸ8��çU�H1��"O�ݩg��Twu�Dƌ����0B"O\0��΄<����7�Tz�"Oh��F�,`�]sp��3x_^���"O҄����J<:��D4A��1�"O��r!!� K�` )��I.q/V�p"O���Ы@��P��:�~�+�"O���DaG R� 	��@̹ R��"OH��؆U���!`�5	TM�Պ~����B�B�,�4`�C�>#�M a�y"�˰!�5	���p��R��˾�y�'��=��
<y��w�^�[;41��Mk�4��6���)5�h�I#aғy�0	#B0D�0��虈$5�����(-��a�-��P!��	X."w6�c�ΓK�J<��ӑP!򄖿IBb�1�Ε>��`q��MB�!��ҏG�aS�!��y�a	,N�!� ^?��P�`
	���b7�V�&#!��! "%�2D�N�`$s`�Rl!�Ĝ�C8���U�-��t�PY�!�ѡ=$Ɇ�V��<0��+��M!�������&U�(��vJ�~+!�d��Q.�@��CU�֔!�k��f!�$~"F���-�,m�Y��P�y�!�̋ X�5���6Tb�U��"��)�!��t��y��Q�w���u Q�!�MS݌�9�(de��a �m!��0-��=��'q��;�^8Uf!�d��n&YY� Iꦙ�P��!��'9Ȁk��E��sQo��'�!�DO�=��<���'Jr%�g.Ĺ�!�D�/]��=�&�F�E��8��l�:<�!�D�'0r��NJ%}��CrKK�[�!�D	j�HPP�g��z�H���
���!�0�ɰ�g�]��i`7��0 !�DH��:` �L/Q،4v(�8s�!��� �n	X�g�R��$�7���i	!��W�e ��5�"�2�Rg �[!���I$�A�n��r\F� !�߬S��Xy���1p�|�8Ѯ��p�!�
~�0����dKA+n!�$"aKf ��NĒD�Z��c�U+f[!��)z6���S�Y9����E &6D!�dO8F�(����D�
ܐ���D֗%!�!�fA+c��#�P�ѐ��!�!�$(���k"����\s�cл?�!�DH�X�:���%�^�� ��h�!�&G�չgLB�1��ɧ�M�i�!�LǆRN-�P�����o!�D�NPDt�w�h�E�pt!�?;��Q�n<"@pЋ�e
N}!�� ����Õ�:�:Qȑc��?V�L�"Of��w��. `�ơZ-.)z5�"OU��H��2��M�D1��r"O,����$m�!���n�=��"OD����&j�2�(B&R��R��'���'���'c2�'nB�'b�'���/�� �~�qJ���j�'&B�'<��'���'��'���'���bS퉸U\�{g$Q0�T��'�'���'��'[��'	2�'���'s�T�òa�����܎?5^%�S�'���'���'5B�'���'�B�'��5�A��4�� O�O�Hq҆�'��'���'��'���'��'}��+�5T��#V�&��zF�''"�'���',��'m��'"�'�^�h�b��~�`=PL<D�I�$�'���'g��'�r�'&��'�"�'�v����/�zD�$ ��r� �� �'���'+��'8��'�b�'��'��%&钭)���{� G��"���'���'~�'WR�'�R�'���'ߢy���

i�)�C>�X;��'���'c��'�"�'���'+�'	��Ye��*L�|p�3�W�_Є�'�"�'XB�'O��'�R�'"�'�����
�d�ˇ����pV�'�B�'C2�'��'���'��'�XL;B펚q]�x��U}��u���'��'���'}��'�2$u���d�O�x඄�=Vr�; K�9�Μ����GyR�'�)�3?�Q�i�y���G�&���NXW�M��g$���S��?��<��l�|�GD;u�Jъ�ӥM��p���?��*L��M��O���,��L?��F6N�2&F�.E`l(1��3��,�'��>��e)>+��c����A�������M�D��@̓��O�X7=�Ɂ�#I�H��IgRY{6�I��O�$}�<է�OДyñi�Y+>!�;�䁬� ��vGx!r6O���,�?�vg8��|J��b$Jݫ��B��$<��	�Fpع����#��������9�	�8,�joL9@@��7�A��5�?W���I�@͓��d�-2�ʰ���S0[�*��W���5������p@9Ej�c>��`�'k�I�I
�2���N��hvV42�/9�f��'o�Iş"~Γ2r��!���=b�\�s$O��Γ2b��
�
��dB˦��?�'ZU�l���8yb~���RBM��?���?Y�&��M��O�����3�8�b�\#d�!� O�K��Ol��|���?��?���V�R��5�(�^LH]#nИ`!G�<�üi	`D��(۴F���'[�����H���'/<� ��V����֠�j"��i3˱>���i�p7�����zL|��'�0��(~-��z�`+X&�!�H�6_GL8!w�ݶ�?�AG��|�T���u��9}"ǛeyrAA�Z�x<(�h\5?V��Q,F2�'���'�r��7%���M�B����)��T�i�%N�;��p8B�<�`�i�rW���I���������ٴ~���c�Z���Hp�?B�R"�㒤[�� ��ia��O�\"W��*�������5�_�HZ@~�yia&]8�Iş��	ߟ$��؟��P��]��A���0;� Ǉ:hlu�Cϗ"�?��i�V��9.{�ɾ�M����T1@P��#,ʪ\�dM��Z�h�^oZ���D���� �4��V���M3�'v���=��cHԘh�@=QK�f�B��U���􉦝|rS�������ٟ|�@��N-{��ֲ
t>�����u�Rd��zy�Eq�h�sm�O��d�O������`dƐ�W���*�n��q;O��VPy��'ݛ�hj�l%>��m+�E�D�нt޼�@m�!D1,P��e��[
l������n���\�Ojt�4l��C��5J�;<x��%�O*���O��D�O1�Pʓ
ě�Iȉ
�"`ˇؓ^2LlP���_��H��Y�4��4��';L�NF���Ru��L�/O�d苇_�V�$7�ѦuXbd��eΓ�?!D$��i���^<��L6hl�b;�l�vHɓD���<����?9���?���?I+�"�:��%G�\s��O$$)j�(F�5��l_ß����@�y��'�7=�|S�bO3ywp}�����y��������@�4�yV�b>Uj�&Oͦ�͓Ht9�S�E�50�H���Hlh�=U�q��A�Ojx�L>�*O���O�|y2�C�cZP�qd,ۿy��r��O����O���<IÿiF��;��'���'hΠ�Fa� y`�t��ȃ1?����'�'ID�z@�Ho�&%�L#p�����}����l��ej����=o8M���m_v|�'_�D'���@�!�'s�2R�� w��p��W9N<����'#��'m��'5�>�]��)R�-_�Th�ѻu�h��	�MC����?9�CP���|���y7�M�m�cj�ub�尀�
��y��a�̙l��M���M+�O�+C���Ԡ�?����cAx5=���P� �O˓�?A���?����?��E�H�gM �y�JH�ԋ�5K�h�3(O��o�bR��I������?E2����3K�L�G"�@p����+լ=��OL�l��-̲�4g��O����O������e�~i���O����3P  �[�
)�O%	D E�?�0j1���<i������E&	
�͐��?Y��?1��?ͧ����Ħ���jXڟԃ�F<d@���倭4w|����U��l�ܴ���?�\��h۴q��Foj� �R@��ұC�� �,xRD	N2f=B7�~����O�,���O->��'F�$�p�� `��@���J�N�c��_��H��2Oz���O(��O����Oړ��xk��ʈ$���G��'X_�L�0��'!�lq����O��d�⦕�7�myBbsӼ���<	c��,E��Aٕ �8!�p��%7G����<�ش��c��Y`f}���ğ�1*�;k�4Mbd�C�z<�@%��0a����'�8p$������'���'�Z�Kl͗V�ry�+�4J�:�	'�'�2\�"�4uvj�@��?������֭��Й�\�4�HB蜠	q��,@�O\�mzm�=���|���x0���g��Y��#�b�>��� �M�>�<I�a�\������$���}���$�<1��F[�&��Ҁ�# �D��e^��?9��?����?�';�5�%oE����T��ɒG��'hf ��'J�ac�ވOlt�'F 7��OD��?YQY�����7b��7z�"� �%Fн2��M�%�i,t��c�i��	-A~Z"�OX�D�@�fAǭj�@5��)��A�X�����O����O �d�O����|�%�3*T=s�P.Pq���'L�fK�7gR�'����D�'��6=� �y���
5� �kn,�Y�	Pئp�4C�����O���dT�[�?O(4q��Y�yU� 8 �%Wd8�ۑ2O�eu�� �?	E&:���<����?���C>Af�hk ��k�H�LQ�?	���?����$�ߦuɷ�ߟ���џpU+R�0F	p�o
�+�|���YG�Y@�I�Mնi��O,e��>�t��D��81�D12:O.�d�	[�¡�E,ˮ˓����O�,���u�T�{@(�)yU��R��C"��R���?���?9���h�����8W��T�%΃������ρv�r��
�!�&f�\y2�wӾ�$!�4�%�q���j�hС�j�'^t%d9O�<n��Mq�i���z��i��O�\;�%�*qA�"c�~�@�S�Uƶ��w��Iod�O�˓��O��3��Ѵe�r !��N5��``��d��4(��ј.O
�d'��3na�52Ӄʹv&� Ҳ�C=8����O�o
�M�7�x�O����O
j೔!D*  ���2����e�gzB�BT��dC�<m�
C�_y�� Y�萱���$�f�G��1c	"�'��'��+߷&��I>�M���1�b�H*o��q;�H%Ho�3����?���iwY��3��$�ڦ�a۴q�fAY�-e�E+� O��<P�� vX�p�i���O�P��ǰ�:����S��56�>|���Hv��L8���UIU�r�'t��'�B�'��'R��oB���"0ir��f0uu��&~�����'r$�O���O���m(�dҵJ[�5��%��W¦5RǆV@�8Qoڱ�D��ɼ�M3ֳiܪ7��p�7Mu�P���j㲬�ӹ��[F�p&8�@�	�,p��4�	�u`�'��i>����H��!0�t�H!	F�k�N��4�L^�����,km�5�'1J7]B;����O��D�B�I��;BD�D�Mn�����@����O�|�'��6M�Ц��ش"����톢7E�B����O01ȵM�u�*��@E(Ke�i>����
޺+��'���-z��B���N}de0C��.R�֔�	�8�	ڟ|�i>�6,ϟ(�'��7M�b<*�
�ͮS2�0�'B����':2�4���$�O��n�X�N�Zd�W)YX$P���9x���4P���\(p�f���R��-I�$�~ڣMȹg)tp�e&ʢ-���/Y�@�Isy��'��'�"�'b\>)4��3(����"�6ӱ�:�M; ����?q��?�''�j��OT6=�8���ֲw�X����(���䢎ҦUz�4<W��ϧ>�'����q�z�4�y���:y;ȹY'j��(Y��*vA�3�y"��t���	�b�'��)����&~���`�a�:*��1�I�pc�4n�>��)O���
6r�9�@�3#� ��ɘ�K�����O��m���M���x�dڸ�V)���A2U$��Pu���y��'�lB��Q�{�J�pP���ӊF���Qӟ� K�%N� a���-c��	���ٟL��ğ���˟�E��w&&�Dq�6��I�������')x6-�V6���O�0mH���]�W�Y��
�J�T@x��_�F扭�M�i@�6��=B&6-r� ��6p$�ڥ�OI�%�e�Ɉk�$�Bf�<&,���� a�	}yR�'w�'���'�2&�-7���8vaI�r���փ˰/'���M�����?!��?�H~b����=~��<�fݱ-Dh��ST�p��4�����O��>�i�ּC��H%Z|P�E+E~ú4)wK�s�URE��<��$W�cB���������++
X�S��LX��p%�Ϟp�����OB���Ot�4��˓4���P%q��B�i�2HI�O<:Lx�S0�J!R�h�,�O�I^F}�w�&HmZ��M�Ԏ/"�hQ��F�|�sᄐ>'�X�rݴ�y��'u�X��]�?y�V�����e2��,A10(���O>J�����e|����ϟ��IğD���%?e���G�Z��'�ޮs��d�QCڻI�A�3BJ͟�����M��oH7�?����?�I>�gW�5]´�Tk���c�I�F{����>���i�47����&Kw�\�	�,��l]d�v�1W�A�JZ�abT!"g~��Fos�0�Ify���u�ڟ^���O��Ă"}���6��0��M�H�=Z"���O���%Dy"T* ��d�O0����E�Shf�@�B�aĩ��H�M���Ɍk��Q걮C�<���M㑲�*����	�c�cB4m�p�0 d�K�
����]<92�3���
*�I�?͐gO�ǺS��'�剈T+�٘�X�\���D�\�Iܟ�I��
�`4+�b��	ğt���?	�]w�)a�
[/,'� e�'#��`�m?����?1I>9#��?<�Z��� ���DZVR��'�L%!'<Mh2���=D6��� B����&fЂ�J�Eo
���?)�3� ����@�V���A��V;J�1��i4�x�'3r�'���'l�'��S�Ь(���*0�$c�;"�h��شw�q��Y(�?���R����?i��?ͻ���%�Pr��4-Z�78@�b�i��6��ܦE��O�������߈DQ�6�$�#d��hH� ͥv�b�m�DAF�����U�Od��|j��0��<��n��14܉���3����?���?))O��ow_�\�	ɟ���;b��,i�&1#M�k�n/��0���>Y��i$�6�{�ɘ+x)q��ĪYh��"�����Ih��V�k���y ����&��O��!�b��G�cȊi�p��q	�(���?1��?���h���0i��H*Bk�?e/���8K�R�������Cyb�sӀ��9T\�)��� �B�3'��va��	��5�4gu�F�ѥU��8Op��Q��½C��)�$�*��_���k2���|ؖ�c�;�Ġ<����?9���?I���?aq���Xj��@�:L��A{��?��DFۦ!�3+Z��I�x$?牦g�R���4������i�/;��D��)Zش0Ή��O�,�����Tc�mخB�6HbR6!�3y�˓W��!�"�O8�1L>	*O�D@��By֍��̈́���n�O�d�O�D���<��i��Zw�'��H���Ώg樻s&8I�r�Ҧ�'�"�|�O���9�M���i��6��fRX:�$_�lcԈ)���|)�F�o�F�Iן@b�Ě�4���o)?���uak�ʍ0���9�"�
r��q�H?y���OT�$�O(�d�O^��6�5F(��Ӯ�!f�	��țB66��	؟<�I�MUh���^Ҧ5%������5{H�É�=U�f�������.x�h��8�M��'�b�ߖ��P���1=����
Pɚ�,�ϟ��|�\����������|�ꔼz��� D;��J ,Sퟔ��Zy�	bӂ��f��O���Ov�'n��}����(_uLT���Ҕ#P���'�T�3T��/tӪu$���?UЦ�G�T���S�z� �$Nmh���e
˥��<!��)���DU=�?)(Ol�p��;(����gԱw��Y���O(���O����O��M�p�8<zȽ<��ihV�"@�q@�ٺc�@�^-
��X��'N|6�O���|��S�`޴?�9��ƚU(�� Gۈh�ľi��7�^��7�c�|�I>|F�
�O���L��RH�x�^9�1@��v�ϓ����O*�d�O����O,�D�|b�� �V����^�UN@�!��6f��V�yz��'0����'J�6=���� U"q�&	S�\f!�a,���}#شD�����O��DA�/3��:O�<s1.B;���b��t$�I��0O2�s�Ȭ�?�G�0���<)��?Y�N�tv�|��JhV$��@b���?Y���?�����d�ۦM2T 	����I���5aؕYԸ��l�"u���`�(�N�$s�ɥ�Msǹi��O�x���"!�j���:�=�P8O���tҤ�aC����V���g�O:�[��BQ�w���JP�e���Rx����?A��?q���>� ����?��O�*)�^��U� l�%��Ɋ3�?��i���3�'3�������<��Ӽ3QnB4o���N� Fq`�.˴�y�z�~�m��M`];�M˝'~@�Ġ�S�hd��Pg�3!�*�q�(f �SU�|2R����p��ݟ��	̟�:�-�a���C�ǐ�N� ��H~y�-~���[�@�O���Oⓟ���]�$O��D�OG/v�̌�'�6�B�����ħ�B��VOm����[��с�Y�g�i#r�L"�0��'Ǿ�Vg@۟�2Ó|bW���aL�y	����!֖��X�#���(��̟<�I��gy�Be�JH���O��c�;Dΰ���9�ИI>O��n�Y��Y����MC&�i�"��Na��$kH"%�HZ9��h�'�i��d�O��7,�ꢙ���S<�56d�P�1kc-�č�����y�'���'T�'R�)^�{�>d�҈�
*�`���$���d�O ��O����� P|y��n���OƁ�҈+m�5�2�)k�^��զ|���' D7������2[�(o��<y��u�81�$��^���D��7�)q�PF�D۫����4�����O��$R�n��r��-S��� #�ޅsK�����O�˓j�6��R���'�"�O�w��
�p��b�	t��a.��yr�'`� ��vl�p�l����'��oB\��X��$/y����h�>m�����-ضcJQ�'��$Z��D�6�|r��$f,,��2��+5�Xu�$�J4��'��'��d[���46�L�e��}T�M�W������@h��?���K
���|��'��^���B������Jߙ٤i3��@�d��7�����)F(�Ҧ9ϓ�?)gďC���������^\��@��A�'3ȐbU+�#S��d�<)��?Q��?���?�*�4����J�"`���Y2���4LWۦ�����ğ$��ҟp��U��'1l6=�z���-�A)0�&*[(�TK@�ʦ!�4#�����OU�th��3��7O�xriW: �� �ُF��a{�'�ҡ��GǟLzW�|�R������#���52��k�?�Ţrf��H���x�	zy"KnӌP!V��<���ix������@K�@�r�OTَ"�>�i �6�
Q�I=��U��)�He�
�n�\�	�h��#�!b�T��My"�O��e��9#t���9h�Ĕ���� ?X���)-I��'���'���۟� U�Ҳr^� 0�b�b,���ϟ��ߴ�,�q+O��o�z�Ӽ�%Ł4OKfãG�[���ۦnD�<���q��n�,>Xj�l��<���]������� H� 6@�Eϗ[Ӽ={c$�/_�,�R�d+���<ъ�Č4*�x �@�*-6L��-��b\����M[a���?!��?���t��+�^����a<�C1�ۘ��^��sӂu��v��?A���pZ�'�0SXpU�޵9�P*��5g�'��0a��ӟ�I�|�[� {�� i���@��[�AQ���*[�@��ߟP��Ο�STyBOsӔ���M�O�e��*� h~ A���:s��:V<Ov�lZO��&j�	 �M;�i�6�AM��z%䁠x�=���3]��9�-y�T�	�.v_^ ���XB�ʓ�J�;`Z�;�]0E��H�AIE*�,���?A��?��?!���O'l���H�v���2E H��@�'�b�'`R6	)��O��n�X�	$t�f܊��E0v�P�ZF�D-�NMZO<i�i��7��}���Ӏ�I��dB�(F�-Lب��&1-[|q��A��+����R�'e�$�Iwy�^� �I��D����<�(]�_� 9���շJ<�2P��$~,b�Oqy��c� l/=���'���O�'LC <RLJV ��L��Qn�4�y2�'e�I�M�i\6�l�'D���2�N̺--���,�W2���A,"Cp(��"�D~�Oo����;	3�'��B��(J,<��t�n�r�l_�\�	ڟ��	�b>]�'��6����H8�l�=}2��v�͜|�ʥ;�ͤ<C�id�O*��'%�7�ܡj�ʑ�
���7�*g�$nZ䟘*�� Ӧ���?�V�/@�)�D~��߄S�%c�B1x�8�(pB���yrU�t��I,\C<�E�G�W�j�@�쀾�D
ݴ!�����?����O��6=�dJ��խи#������
�V�5��45��V����?���w7��lZ�<�@ȃ1d;���2aZ�r���K����<����;���=�䓹�<97� [��Q�p�X��Zp�CE�X*ܴ1�Ai���?Q�TS4Tr�(P�~��T��r��(�B��>q��i�7�����'܍����NȒ���H'Y��'A)��P�t�)S"D�I�?��Q�'�8$�Ij�@E:6P�[��x��I�CV���I��l��П<�IJ��yGa�J��|���0g�t�[�A�D��mӖt[���O�d轢'�4�iޡʁ��*�x1�աםy�H�!��|����4��V~��U!Ƭd��>�ܙ���L����@�wx�H�LQ�>�Fy"fMG3�䓿�$�O|��O\���O��1&�Lx��Ȇ
D<��*C>In˓3�f��=/�<�U�'6B�O�&���_��s���f�f��Z4`L�䄔��d�Ezٴ[��6$,�������Sj�̃� "pЄ���$8�	�2��<7���9I(�St�'pP$���'���!��/�,�a�擶z��QA��'�"�':����X�h0ܴ<�B�X��R2 �x"�3�p� ǻg�\������Hy�'��f*f�&���^� t)S�)>�c��Р+�7�:?ѳ΋?���i�/�䧈���	}���㐎��f� hT!�<���?���?����?���D� �i�����[< �Mk��X�eV�`��'}"{�𥢧��O���O@�O\8Q�#D?�p���@��,���&�Ӧ��O��l���Ms��m��u�۴�yR�''����� �@���S|�XJ A�&9+:��	
N_�')�i>���ПP��-2���.\�q��/��z�	@KىM.�ٶ�Ry""z��$@������O$������uL�&(Ѩ�.O)@���SC6O�d!?����M#��i
��z���M�ڸY0���b��\���ܻ_��xagl���G˶����&�ua^�6�1��R'g�T���jF�a�r�zD���O;5٣΅)��g���]𰈚nY�7�d���nC�u��Ɖ��c�n�� Ȉ35���;�U(s�y�p��G�$�P�+�83Z(�ɳ�Ӹs��Q�{����#dpӚ�s�Z`� :�/�{p�H���I7fDR��/�&0P��#J� �@����d��b�W�[(���`�F=rl� *�0D�5XF%G�4��dB�L�q�Y��	�1<���5�8ѤF������AA�":�� [�1���dB� W�����R�{H�i�!G=L�|H�J�i�� �` �}�$�7�����%�$�����+�%HDD�a4԰�a�l��"c��	ߟ��	Qy�KR2�擠kJ�x5�95X��B'��<-ꓻ?���?a)O���O�	�U?q���Y$Zw���p�#:S��h�&�>����?����T�{^�%>�r��H&]���u"�%-X@�)V�5�M��������3y�����䗳.�a�A[;��X�Ƿi���'M�I A�^$yJ|������Co.	R�"ϡ'��5X��9�P,%��'���b��i�?�h�-�<�z؉�^ J�\Y�FiӺ�}	U�ҺiE��'�?Q��Y��	>|�|]{@V�P���'n�>�6m�OJ���&u���S�$���V[�l����(�qa`*�/{30 m�R�z��4�?A��?��'*����e�5�r�����7���FT�|�7�!��˓�?	���<Y�p9�����͸[H�KS"4M�8QS�i$b�'k��Ϧj��O�I�O���8��D �m�(w<	`!��.�����A\1O��d�O@�Tw�H����ľm�Ȅ5*ן0v����Ol�挑h�i>������'%S	@%�c#��<A����L�2f�v�'+�<�y��'g��'�剝{�`�w��Q�8�!��]'Bhy�	,�ē�?�������dC~�b7��+7�pH�]�e�4ё�d�On�$�Oh�O�!�4��UQ�
L���i� A��&�{�\���	ğ $���'�䈬O�y���^+}��(e�O��� :�\���I�����yybh�M
�b<� ���V/A	z� �*���k����%�i�r�|�[�L0+;�ӥB�U�f�.F A��I5�6m�Op��<y�
���O���5�oH�G��JA!/�p���Bԭ�ē��D6z]>���d�Ny�X�T��
�J^ ͎�l�iyBh�WR7mM��'��+0?	�a�#ٸ�qM��i���Sɦ�'ҖU��O�SF�sӐC�Gs<�p�kĘ/����i��� ��g����O`�dោ�$��B��Yi�If�C$	Cԥ�ش|��!+Oz�d�O�����O�{�h5�`����[�ha�'�����INy���>H�i>E�I�`��
�Р��Dϻz�h��#+ 3��8P��7��'>m��˟|�f���cB��1ZM��F�/a��':p��[� �IПl�	k�Y@	��1��` �Y y����'\���A�ؼ����O��ķ<	�S�d��e��)�>�򠊒�gPQQ&����Of�d�O(�(��g��c�!wy҈��$�>]*i���M�I���?q����d�O��@i�?m�fIϵO��� G'�+&z<��g�>��O*�D-�	şBƷ0FBeӲd���E%`.���W�]:Sn��E]������'1�St�����H���<? ���&�Ƞ�LU�E��۟L��K��?�r�
>ְd%�|�N�3]8!r7�V%G�N��G{�j���<���Gh��+�����O~�)�&,�Y�6란'��Q	��>���>I��۾l9�"S�S�D��$f���2��+E
M�f�����O�X�@��O.�D�O���
�ӺK�$pZ�X7�]���Ajl�H}��'&�2�⍴����O�e��bX ��=��DAt�|ŉٴn0�;���?a*O*�ɪ<�'�?�ӭ6�ruX��~̬;�O�9"���4�	X�y���O@��"E�3Z��:��[\���xe\¦9�I֟l�	���ȗ����'y"�O�5�׌G�TZ ���o�2>�R��'�L̓I5�)Е���'��O�p!�g	�F��A���]+k3����ibReӤ �����	͟��=Q�ݾEjX��f��[:�<۱&^}bcV��� )�O��D�Ot��?��n?'���^)^��pd-8�2����<1���?�����'yB+��)H�� 6.��4���f���q�ж���O����<Y��7|�4K�O7�X��i��!�aƢh�����O���?��۟�Q�)�4]��7퀳��X��D�5�J���	�"y<�I����|y��'��A�V>��� /=Ѓd�$��5#Ǎ0����4�?��V�`��8�QF���T�R�$���Ɲ�4���'���֟�*! �h���']��O��h�R�E�/<>���*��l�&�	py�A��O�nC�uQ���S�{��⥅�"+����̱QG�����������?՗�u'b�����)O*�ڀ`2���$�<�6��K���'(�́ҩ�zR�2���%���n��`
8��Iǟ��	ޟ���Ly�Oq�mN�Ht$���C�E#.�b.�q��6T(���U���P�PH�]ӆi�3�B���!�:�M�����I"����|Z���?Y�'O,1 t(�"q�m��A�$�(�+-�ɍz�t�+K|����?	�'b��AC��d�t0���Gմ@�ڴ�?��G��$�O����O8���'@�KI��	��\352�Bqj�>G��dT�'Qb�'0�韸����Q'�!��M��(�&ގo��u�'��'Z��d�O�݃�ȓ�	N� �G��9f�C&e��`��4`�� �I�T�'�򣎤)�����.Z�ѳ��S�o����������F�'���'��O~��� l��Q��i��İA�>I�a;�㛽_"iЬO�D�O���?��lB���i�OlؐQKC2MC. 3gb� {��*��	����A��?�g/�R��'�8:L�[Q9q Ԕ4t�슑km���<�����.��$�O��	��K.9b�%�J=.�1��!\����>i�EP @g�h�S� ��8�F3��%#�T���KO����OD%���O(�d�O��D���Ӻ����)!--� �U�{��a��Z}��'P����<Ș��O��1�� �?Ve����ӽ ���S�4mĢ����?���?����4���dL5:��H9��	�a�0N�XNZ�n�E��8�n&�)§�?y!��e=��7�
)ST� �\$W����'�"�'{����[����h��k?��նfv�P���D��A+���F/1O!�n�d��П��IO?Y�V-(f�kr��.`E�զ��� '�8�'MB�'���� *l��ᰃ�8���i���(O�ɷU��<�k1?����?I.O�����a����Y�"��h�E�,#�<�4�<���?q����'RA_:T�L:#�ɏ�@4���	}v��*����O����<��,��\��O�(��!�R�o���Yg(��0r�MSش�?���?��'�ڽ�Ţ^��M�2/��6�����̓�A��4��b�}}b�'�rQ� �	8(�}�O��$ȧ|����3�L�e����U�Ce��'j�O2�$�<s	h	�x2ɰ4z�!S�T�Q�� P���M������O&4J�D�|���?��iin�PW�2e�L��թǷD����$�	��z2�Exnb��j{VL���/אI�h��$�i�'$r�E��'"r�'���]��=� 0\�NS3��賈:[�*@*EQ���	x�~%���-�)�S>K�SҺ�0!�֥�t~t(lZ�I��@�	����ϟ�S`y�O;BFгN@����e�(B����'J� 8["7�H��D����ݟHXf"��d���ԍY�N}�WȎ��M������owf��|���?�'��puC��WV0��#[�g�E�c3��8�J��I|ڞ�?��'2��Zd���)f��d�M)RfP��4�?��h�,���Ov�D�O@�0��H��~%�� �ܖQ;�H���>Q�G�WHq�'��'��Iß��D(}��`�f�5U�����ۨD�H��'���'��d�O$�U������W�8&~��&�
_J�}QƓ�D�	��Ԗ'�r �!W��E�8�>(�7�?C�	U�C:\����'�2�'��O����!&��(��iA�-���.��ͫ�m�jw��!�O��D�O`��?QK9��I�O�� �L�����tlۉ%��n�馭�Ip��?�TCA>�h�%������/�Y򰏏l�R;C�m��Į<q��0a��P)�����O2�i�	mN�I��\�V`	���]�SȬt�>y�0�(%�f�NI�S���I�P�J-��I�0 ��bc^�M�-OڡkSe�˦��	�(�I�?-b�O���(ݸxaR�T�4K�tzh	͛�'M�n���O��>%JG@�H��p�NGg����s��,�Kצ�����I�?��Of�$��pQi+m���#�;gF�ɱ�i�t��'abW��������0��:8by�FAɱ:�fh�иi2��'��#�������O��	����6��C��4z�W�Z7-�O�ʓF m�S���'��'ԍ��,B5�,�ThʵW�NDC��tӘ���>#��@�'��	ǟ��'�ZcF��o��bj&Y��	���Y�Ob����$�O.��O��t�N��!i�xơ*�)$.�9��B*c��I{y��'��	��t���`�&��9�nu��!
^�F����&.���(�Iǟ���؟l�'���d>�!#`&m�*Hk���	ǴY�tEn�ʓ�?�.O���O���И���4V3����x��}Aƃ.
�6-�O��$�O4��<�� <����R
91�R4��O�%o8� �M+�����O����O~ �s���sӖ���腖!?���#�t̙��iwb�'��i���r�����O���I#(7�$�X�y�P��`�3K���'���'�Y�y�\�X��r�e+C�(�"	�fƃ1�����&�Цa�'!��GCe����O �$ퟘ�ԧu�K�|_8Ms�2H��C��C�M���?at���<�K>Y���S�<��x1sB<pt2тN�M#/יIe��'�B�'l��Ƭ>�,O��F�v���w� 4����a���bJu�$���*�i� JP8j�p��DH8|�̲a�i?��'����Y��7��OT�$�O����O�O0o�l�Z$�q��@1��m���'�割}KR�)���?���o���#��H�C{�rf�1��R־i%�L޲1�������OV˓�?�1!ށC�		�f�&�[A��o��,���y��'���'RRX�K3�N����+w�u��o,���OL˓�?�/ON���OX��Ɓ-��EyAk�Asν�&
�-���=O����O���O|�ļ<A�b�8V��II0�0�6놜V�eJIo�S���Iiy�'���'VDQқ'7�� &ٱ>����@�2��k�>���?����Ĵ4@��O62;(�HyC�^:y�J�!��\e�7m�O�˓�?!��?�����<!O����*#�@�2@� � }S��}�L�d�Oʓe`�1cY?)�	�L���J��X#���;Պ��D%T:�H!�On��O���
E��&�d�?�K	)Tti�"Q$�<��Gy�`� �$页iV��'~�OŲ�ӺKF(0���7��(+����æE�����cc�s�x��tyb��"#�R݂��1Y��(��Q��v�9[^�7M�O*�d�O>��T{}�Y����χ�mF�|
S��oZB����6�M듪P�<����(������f���5�D�.Nr4�V�H��4I��4�?���?))�&u��InyB�'���
���!�@Ӯ� �	'9��&�'q�I�Fh��)���?��
�"�agD��G�-bw�p�i0�NʿSn����Oʓ�?�1-�P� *bܸ��	�`0���'<:u��O��$�O&���O�� �L!jc�DO�RѪ�jy弉#�f]�J5�IGyR�'��	ǟ��	ɟ�05�ڛx��t9��D�P�Y��#�%���	՟P�I��,�IӟT�'�ā�i>���.,5:��`拐�x�����Nh��˓�?	-O��d�O���� |�\�F�"E�;,^착Q�.���'#b�'a�X��0Sዧ����OD+���h�`ŀt )M )���Ҧ9��hy�'���'����'�J�`!HQ�T8�S%N�I�x�m�֟��IGy�jܕ%��꧊?����҃�U�R=�4��N�7]��b�BL:i9�	ԟ��I˟�ڒ�l�L��yݟH�QCׇ���FJ[/w�yP�i?�I"z5y�4�?���?)��Z�iݥ�0�H�3��VőN���I��d�d�D�OB �3;OV�O��>y��b Y?b �f#BiP�Tc�rHk2��̦��I��I�?���O�[�Ĳ�ʓ$1D]���
;�s�i�ze��'QrW������_��� �dY����de܃/�B`:�i(2�'�r�L?�듕���OX�)� 4M3�L	�X����D���sk"�"�i��'�2�,�yʟV�D�O��в c�Y!���s�Lɠ:���n���\�D�����<�������Ok�ڄ_X ����QHQ�և��op�^�Mkg��<����?����?1�����ΰ]�P���g���0�aj�z�"�ѕJh��?	J>���?��i�2i�hm��Q	u��zDd �ef�ϓ��D�O���O�˓#�dQ6���VCR.K�6�;����T���%���A����	�w���h1zKS`��s��5�aF.0N���'�2�'k�]��(f��ħ�,�9�(�1GC� ���C�q�؊P�if�|�'g��B7��>���?
�(�l
�#פ�:�!צ}���H�'��Q�E'�i�O����й����p�Yߐw<I<���?	%��<�K>	�Oa��3ggU�	
l1B�T���4��$ж
l���)�OR�I�@~�o��iQ�y��a����k�a��M{���?��`�<1J>�/���	|t��6ǀ/��s�)��?��7-W�1ӒlZ�t�	��D�S��'p��1�H}��AR��ۇH�.c"�7M�-����"��4Ed!'�P(H��\ �h�vj#hΛf�'���'��ek��9��O��$��4�q�N ��E��2s�DQ�8���@�ZI&��Iß0���:#��3f�
<M��҃�l���4�?��m�jV�O���8��ƜɃɓ)j�\�YŌ)=�$0aTS�trC�c��'�b�'3�O��cΐm���@EB]�T0��[DGQ�1��Od���O��Of���O�P)peJ65*I	��4./���#H�vd�<����?yK~�GB�Tn��ND�p3I��8���jR� �bȉ'|��'������	1!8�����3^��9wL�g�r��?���?q/OXp)�+�]�|���5јT=p$�FE��u!ڴ�?�K>���?�#X��'��I��"�3I��I�U �6�*1ش�?������W;j�t�$>}���?	�qi�)!� ��%��V|$�q��5�ē�?��k%ϓ��$���h���MKb����M+*Of�ch�������d����'���2���6��x�%�$k���O��$' _��d�O~�S�[�@�С�S�u��A�_�Qmڹ������I�<�jy�P>�I�N�Z��Q/��A��t"5�] �M�s�v�'���
�U�1r����6$
!�W�@ao�򟤖'.� �'��Z�<��h?�F"R,���ZVDďG�,q����1O&4:��{�ǟ���@j#�_5h�R���A*�܉���M��1v8vU��H��T�D�O��'�0�{C�O�3��h��j]:=�T9�Ox����*�D�O����O����O��1��iZ$�pd�)Mj���d�6�˓�?���?�L>����?Igc��w|X�����4d�ъ�_	?T,���/XJ~��'\��'P��'�+|�I�?�z0�G���7��!2q�Y�nP��W�8��M���<�ɇ=��xU�sӤ}H��>T���(G�3HQ�M�!Y�P������	Ny�����'�?A��ڳ4�`�b��Pke���7�P�*����'or�Ė�NA��80���#hL��e��,�`�#�p�4�d�O��d�O�-�r��O&���O��d�\ �f��2H��R� e�B�9C�O6���OXd�5F\�M�1O��%hB��)��Q [eN|��a[�:��?q'@�?	���?����*O�n�~��݀�ٿc���ҮO=����'q� ��$R�y��t΁� l�����s��(+�E��M3����!��f�'�R�'F��k3�ɉ P�P9��ǞX�E�vF��� h�4feV�Ex���O�Ձ���p�ΚT�f���"�����ٟ��ɜ.P^dH<���?Q�'�7��(g�\I��IC[�(5*�}�J��'o��'�bL\�+��pѷ�C�q4QI���& �6M�O���#Qf�����f�i�u�Tg� T��y�Si�@eB&�>a ��d��?i���?����?���
"��Ek���&%��I�uF��~����?���?������?���f�.�B�@F!X8$�7A�Sp8w\{�'-�����R�~y���F�ƸO��9����21������0q$�T��'D��Js�͘˰,�G��Z�J���{2L�-g!|x���Nc�$ �D��K�̈��C��/�T�i6)��t\��u�2��`� ,�p�	�ď:^�@q�ai�?�:1��/��@4xB��,(��[�*�D�ʩ����2�ک�uA,QF��0�#,+�n�#+��V�JbG�GU�3�͙�1�g��d*4�q&��?c�H�=y4��p� 4c+^�@1�+�?��[�Ē5D���l@[�ʧ��̿b�����OV�Q#F�3ճ>�OzrEѰ'�ѳ��1�k��B�L#O�n��ANRS�x`�O��1�'�X7�Z��O�!k*�z�ˎ�=�JM+�&{9:��$�OR��$H� ���Qn��^��5PAMT$rax�2����в�(�Ţ\�n+FtQa��M����?��8��@$�:�?	���?9�Ӽ�!��7 O��@� Ή;/� p��-$�H
"�3i�g�#SL����L>I�Ά'��)����Zr���3�,L�#���<+"b�z�\	�}&�Ȫӧ_}n����Z̈́|#������'��	���|ʌ�Dϑ/I���ě9YgF��@��)d!�� �乂a\�.:�RGع�, e�������?��'d� 	�l�]�>�JSŌ� Cn�!�D޸Qh��U�'B�'_�lq�Q����P�'Q����eˎ�:��I㬇�o���n�5mج䘀�	�����E�D ��҄(�8��ǘ"���qZ�	Vl�A��Q�4��
UlE��G/
x��'��+���1�fWܟL��[�'l�Oܔ��]�%�Y ���(a��}s@"OD�#e!M%3����*�/nB��xd��P}�[����g�
����O�4�A��YVNh`�H$b@j)8���O�䐇�v���O��(n"�ũ⪚=r��Yt/��Aը�	V�� 5M����Z��3O�1ڐ�Y/Q� * L�{/�5�5�!�ы��¨7�ɰ�A�2T�v�8��%�(O�Q���'��R�KPoZ�~bFʮ6$�f�7�	n���z����]u�첲*��sS�=˧"*�t��46X� ǀ�k�dq�G�5;0�d����ױ:����'�r^>Y��+ߟ,��D�s�� �2�ļ^�M*���֟P�	���h�fg_�a:���Ab��?�O��v�:��4�ЙS)r̛���{�*�'��4��Gֵg�"u�=�&���I���'|��j��)-hIă�;@�9�OT�(��'������Că��7��(�RF���@3',D��Jg�F=Y<$�{�ɜa�A�&e+O4Ez�ܬM�R=�d+�?�b���a*���?y��z`慻a�ɦ�?����?)�Ӽ6�� L9�h�Z�ٸ���Q,<��F�I�+��[�
0�c8�3�D��'�A��;V��	1�6P�ycd͇��䆓s�n9ˉ�L>9f-[�Gw�IV�P3�څsF���?��OX�������ə�Sd@O�?Ό��B���Z�HB�	�S�
�A��Ƭ,����al�
�&�����O:,�}���<xY@��5FF1#���#,``����O��D�O�y���?A���4�C�K�$ڗ�Ѩ35Q���~F���r�'aJ����V��i
��:�h�Y2�_���V&F��{Q�%}���U�L�����m���o�`�D�<a���'���KE�IQ�҈��� ��H��'�M���9W�x!��(�b�\�9�y�ƽ>�,Ol)0W#���Y�	ΟKR��2sr����m�tiyW�B�h�I�.�����՟�ϧRi���A�V�I�^w����
^<B#֜�6*^+8��d��H��1� �|���4��;$�&&���Yu��p<9P�T��T�۴*ݛ��'@ �J��:���1��Pq��T����u�S�O-�g��x��t韃2�"=��'��6M:kR�i��%]<�U$��2O��d�<��"JC˛F�'�B\>��g��˟$�G�^>O�ix�E�=͊{fi�d��f3���4☧�P����\Z����.:�z�� �:}2�Q*m�O�A)G���rǰ��j��v0��>��+�ş���i�Sa�('2�Bc�ߞI�4�!��.��c����@x�����c��~P��̄>!?L����p�'���y�ڔZu�!��0	�B���h~�z���O�����l�O��$�Op�4���B�_���k@�R���r�&�	e�J=
�`(��{@t�B3�W�Bs�񁣃Y�%�Vm�ybg�;����}&��b�D�jS�F;���9Č�r�r���Oh���C����Y�H��R�)��-ک~�VM(A��>)�Ɠ76X�u-͗KF���F:X�'h�#=q���?�,Or��g�Љ&�`��!�D`�H���
ZE�]�u��O��d�O���ɺ���?��Ov������"5v|�҅ �	���ui��(�0�'�X���>&1�,zT%]�I��Ԋ��A�'����[��Ԙ����z"�u���?�R�iې6��OX˓�?I��LM:Fҡ����6PS�Mޛ�y�c��H͐�o�W2�
q�"�'�������^%@�m����	1�t���H�&H
��E23��%�Iß���D��I�|�fNE�}���#��ͪ�D}��M�,�h9�%/T�G�2ȫvfE�Ti
(���$^'f��Y�c֑4&��!���nR��b*˥��y����� � �(��-�"4�	��M+�iq���jz2�ӑI�^٨ᓭ���I���?E�$�Rf`����̎�S�<uA�/�x�cmӼ�9�돗%�h�d�̨^(�y0q��O�˓��q����|b���?1�'`�ݣ��Vhv��0�5{����R%/"��R��?17�W�6��$�g	�E�@玨G�`��E��:n���$��&j���Ӆ�L0��	}������U���2T+�${�b IW���ӼAx����#�D�g�T�#h�<\�\�:�C�`����y���?��7b�4����!Q�M��.D���']�t��[��O?���#!F.O�XDz
� S��X��F�4�<�$����㟌���'z����؟�������i��S��@|�Jd��P�n���zu@^���H�TSvbV}�g����#-ݪ.xa�i�7�x�IK>q�/T����>�OER�c��ڹ8�e;j��	�0n��b۴�?�䮚,�?�}�'��F/o����k�7v�f�� ��pC��������#�M|����G�s�����HO�˧��4vLe�"dI9gL��"ƅ�fU!�䉨^ྍ8a �"5����%ϟzS!��	]ұ��E����w�KM!�đ|J�9G_�y"H��ʕ�^�!�V� �D�d&��s	x|��� D!�DM?X�h��Cƚ�$]1�Q/?<!�D�
k	���.YYf����dQ�~�<�䂆2Zg%J�	�*i����7mM�<q��_�p���S���khv�ҁk�c�<��d͗2~$�V�(���f�C�<Y�b�K�"�c$l���4���i�<�`��l��I������Y/�\�<�I3�^-x"H^n�Q�Y�<y�D��Sn�T�Q��>�ڠ��DR�<��.�%7v�,�v'��W�z2nv�<��hնpu ur�����i1iX�<����B�I��� ?�F��!ES�<yt�Z�	������s����Ӯ�Y�<	�햮8�Y�4N�&}X8 ��U�<IejÑ[�p�`t`_	IA�-���O�<��狱uԪ�9�,�J"���"p�<iP/��O<�B,�'v�TCefOn�<i�圹�~����$1J1���R�<��C��
��	��#d�@�H�,[P�<9c�u��Yq� {0�qGb�<���a��e٣j�[9����`�<i�_iz����{�9BC�O\�<Q������yN�iV��W�R^�<Q!�#jX�h5'�oS�T�c�Z�<I��?g���0$NV4;���`p�U�<�Bەq&(��5�-'����p��R�<Y�!L�=*}��MH.#qj�ا��O�<�j4��}�c��-n\��S+�H�<q�c�"p�~Ő��Wl� �$�`�<q�7/B�f%� \46h81�ST�<�n��J������ۡY��m��f��*r����ˁK�l*�1�?�P �?ZܛN?��ǃ0����(:oZ�����D�!�ه�<�sM�fu��/%t0|���ȃ8�4�iTcɁ�M��~>z�|j-;�OJyRH��?".��'^9>�K�b�0>��)Nw+��("��?/I䄣��#>��喼�>T�LV
 �;$�S��n�i��S5��OF1p0��)E�̃Ǩ.b^����ቔ_���!fl�3B�Uہ�I	<D���F���r�.�fe"	�a��-#vⅬ�gh�`��I1zc�ࡇ"��l��xG�|َ�3�<>���Ȱ���0Y��I>��7T(9Y��(����Bp��SL�:i��t�F4,�!�dU0s,���#��
'�`���+� YF$qC���;Z���]�C�9����'��(cQ��'�<91�K��^X���/�`	��kf�|#G��;���d�I(7[��h�d�%Ex�{��r��35	�b¦�֌��#�ށ#�QZ�'����Ir>t����It��؁��7[�T$kG��2n,���ue�t`�P�IM�VT�ba�N,��qz�.��������V������H ̙�e�M�A�1a��1>��,� ̄�?F\���#v]�0�7�� �ܸ���]�����ô�)>��#��:u5 �
E�k�OjA�����)=�aY`K�
s�*Y(lQ2x㢁�Tk���q����r��%�5"�|ZdC�:�X+`I�?��k�~&^A�$AɷnD��1+µ1���c�$����׌HW���1���wP����`�=c]����"E꺈V���).([��I�;c��
�ũ(�����u��U�7�_��\��'~1�SO�K2c 5E�l�:��ĉ-���a���zW�1�..�����b�,�P
Z�~��JƠ�2̊���l�2H%��D�$��(QĤ(��*Jnj�)��L�J`�X�@�k�l���F�B�Ne�*�5n� ��RǦ>Yw.Kp�,���uC��?�CFhl�5�C�s$J���xbc��joX�x���y
� ��� �H���HU[ߠC��Q�i!�	�d���) ����	S0��PJ�&���O��T�mD�9��Y���\��kE�L7�V��O�m8� ӂ����48���b~ȁ�gː,~R���bD��
��,a�"4V�R�'������3�$[�<>a&��mS�1)�I�}��h"��B��x}�2@$s�maVB#?	�.F�����"D�E�X�F!�Phb5Y,O� 1gG�I7aZ�,���~�6���h�a��f32p�UI�(s�R�I��)k2+�1�>�{yb�Ն�i�.L5T4Ta�m��x�LM$���j�I�c>c�D���Q�
���zW��D��2&%P�ON���O��xS��	��O�^�Uj��J�n�x���N�ʳ�T_�F��d�_.,"�oӉF>>�tY��T��È�!�``p�
g�	v�����Й��I,{ȁ&��y�)(1e��
��'lh�F+�-��iK��C��M��H���'1h�h4)6 T�H����'Y8���V��`�'d:i3�"�2I��U�N?���ɤ2I���֡f�L]ꃯ�*I�M(Gi��Yn�Ʌ~x�&�hRǤ<ybĒ3/���F̄O�P�!M�!N<O��4K�DK1�1OL�9@AC>r��S��	U��l�sĄ�C�4�!#�Ou��S1ݦy��)ʧ���h���E%�8j�����(؈b'a"��V��J���|���w���M2��h�}�n#�F`�&�p�9�W�(��+�Y��mh0 ́t���y@� �O�	�O�#2������h1%�����s �_�Q	"�F1"���C��D��<�~�C#2��8��'�>�ƳX�T�$M�S�������r�'�\,�֓~T� E�,~���*O�� Vn�+ ( ��CP�_-0�FS��� e~��p�
-&�����0ʓ4'\)�����E!B'f�V�%��ăR�LB���etb  ��<�s�p�1#;p���jt��<�$�[�″J/Q(�|"."�X�O��;�"���4bR�C�)��u~4x���<�3�	��y��  ��������$	�EV��x"/�-� Cf#�>!�`�+G�-+���	[�O!��a*`�)C�k�)�f&Q�O[�<2T�A'4J\��У��g���Qt�\��ԫ��'$U����8@��{6n�08Y���B�̻
� �ɓ1���V/�7:��T�`� U��=	�ʹ'�fm���%@�
2��@�'���
е3����ң�
 r�Oĕ�A��d�)X�"�}t��O,4�t�$I[�:��p4#�Y��DyFE@���`��⍓�[�'�u秘Ͽ�6�_�'��u��\�I�4�ga�<�U"RZP��p�F(K�Jt��h���"D�-�.�4��(O?�	5Rx,��f*gE>͘PFؽ���'N�}�5���;��h�B���-F�tƚ� �1JC�ɖa,y0q�،�yr)�t��m;΂'S��y�CZ�7�ݪ@�ߩ����a�+c���{׈ˍJ���%`��O�V�0��i�(S�d�)�r:&)�4��A���g�r��$�=2�"ٲ�k�I�Rl�F�=r˺���I&_n�͓-_ȕ�CfIޠE�a�G]�@O�$�֨鰯��BE���� 8�&ʳN]�=%�(6%�K��E飉Hb��p�m�0@ꡢ�=O��`�ny��
:^�D링X."e��r�e&��/1�Hp �X8n@rͪgH̙+0�	�0\����ǁ�w�p���)���I�u�;w���;VFL���J�E��YY�B��#��@���T�o"TPY�b�ux��A6�K�UP��ڲ�B�0#����U`K�4�%��mk,��cL�C2�[�Ђ�!�ָ��[��Uh��D��]���nA����:�V#S r`�'�Xq�
#ƛ�7�xp�*49��Fx"O� b�"6N�=�P�*�I��E�69	�h>}��I�d(H��0<���Y��ɻAD�GI�� H�b}@WI�$@�Ƞ��� ��q)�'4�H  ��X����H�(��O��+0�]*�4a�N\LK��ෘ�$kƢ��(��-!Eg �?v `�Cu��Ɇa�V| �Sh�Q1$� �E�5w�����H	g��KRl�� �-ɢft�mK�%W>Ob-����P�(��̖$�r�� \aN
�%ق&�����C1�w2���3������*S!%�q1�O��1���ib
����+-DpȄi�i}^�Ң��H����R�O�I��j�6uFA�p���B�8e�0U�<��
�9~�lc���j����1O(���m
�[�>q�`�A5D�K��K���$}ᨴ(��ǥ1 ���P��; �2��Z�2�~].���5#�M��<���S�3�Rx�'�lx8���� ﰄ��釵"��H@�'R8xHpJ*o�nxi�ʽf�zi{6M_***U��K?��i��'�p�p��D�K&�c�c�m����F(\��d��y����U&p�r��T��~��M��;*<!;�d ��c� ��S���]�< I��4�1�b�,3�\�� �͂�@h��E���ә'� �[*(��Ip�O�0��OD��¥��e� ��N������'�.�1�&ʾX�U�7��53��a�s��fu+�얊y�����!G��'�͡���#Ø��O��0�H�f������Q'I�P�i�Ob�i��Q�~�׀�YF�k�$&�t�>x���ՉN�dJ�J�0�` g�"��8�"|�'������	�aZ��C�ظ`W�H���$ �e��q2`��+��Oɧ� �XGo��{.�8�m�7��$B���u�,���'޼��SJ^��p��E�YLV���'�%$1�!�޴���l�o��'֤��Al���D@:~� 9�"H�m56�lݽ  ax�8W�m��!- k�$(�JJ�f� V�&�"�C��W�z�*7�|2C��S�j�j�y��dk@�?Z�h�ϏAx�ؐtB���d ��{fK�)Ҥ���6~�"|Jg�G�b�t��q"^�{��Ś��F�pNnt�<�w�G{���D�T�@�&)I��9�0�O�b����D�@*4�R���⌃K��+2��$�������b�Zi24uB�Mțe9���p띞(~a{�$W3^�nXW��	K=��(��S�v�RS�5�J���3N�;���%Y��3��q� [ro^�
`#��rM&-��0�DY*�y��F [���i6aQ�L�9B��μ,��`�"͐x"����K�-!1O����J�))a�t(�Z�8��MB���r����dF,��Eb$���.:J�4f�|�ѡV� k68��-
x8���A�<���߅lZ`��U�Q�tڨ��V�I�O��\ʢF�H���
,5��'>1�=r'V2@���x!�Խl�^Y���t؟���^� 
n9�`��14���`���nl'�1H�L=�IY
~�6Ɇ�	�P�	���hc�Q�4��"H�d"?��@�k5�eY����e-`("P�pU�q��}��`bL�n�|"OZ�#Љ�!�+D� �*�� �����Zd��℉D3#��I*e�P^H�|�r�3`�����RֈYr�i�<y�aO'��8qa��r7�E�����3��UPT��3WVNq*sI�-��h&>��=Qp挶`����h8Qo�1`�H؟ ���;)�쉩�1p4�s'Ǌ9��)� Ə�^S�PR�O7򬙅뉀A���-�Jy��Yd��	#�T#?�Ύ�,��q�wm� /�\9{�B� Oj�܈LK�7�U��KC��4�"O�5�w.C�f��Y�m�(a0|z�T�4yA��)�pdK�©bt��9��WS�O�f��t*��=�����WU�,�	���Ҙk�����.���. B�DV�S\���b���bIi�� p�t���X��ӽ 0�T��$Y1jqxC*�ObI�����"b�"^���`vGG�*�D���	b�!���-&�t��d��lml��j�l嚵"�gN�����$K;[��T�b#g�K�g~�Ib K�O�� �	]�H���bq�0[�ܑ���*Ʌ �-pO��#I*o��'	n�y�?	*Px9$�"��@���){��͖	U��B0fҕq��B�6u�qs�-�s%�� �ܠo�fiQC(G\r2SB_*`���B`&�4�ɜ�*M[��Y���9�G��;+U����ɼ?*pb!���͢tJUT��5lN����v��
'TdCq�'�|$X�HN�X�@j�5�s�'	�(!�@ٲpy("�_7.{���
�'(�����Q����ڬn/���	�'=x���┒e�
t�*�Y�:�3	�',���%�'Z�|�0O�'N|<#�'S6�%#��gmD�c�LT�?P��'�Xh�n���䞏]�d�z�'���
'�z���1�ZJw����'��\S �Z�g�2])��ԙ.`�Ԙ�'s����!j�t��À�aֈ��'p�0@(֍���'�-"H���'5�H�v�,�>�'���n����'�2%�Y�T�)v�Љq�'�$JR�¨;/Fd��iP%7%Bya�' ,���M�i��� jޅ+��'��Z�&<���t%X�Ф��'���+qH�*����g^�N�b\�
�'� �����%[S��!XkJ���'�l, Ci��>��܀W���R>�R�'�I�ぐ�1��*�C��E�}��'0JxwnD3"E 5H�5?T��9�'�d��Ί�l[��Ke'L2z��2	�'�L��� � 9Q􈞨4���	�'�&���$­&�Z�k���+��Yh�'Ә�V�ű�BP�BI�5)�tP1�'N�|Ij�j�tZw(�/,���B�'���D��[�f�{c�],P��\i��� ����[!djf	�g��<q"O�xj��b�h�#��}���au"Ob�� n?�B@�#ļ\��M �"O����cb��iDĀo�0�"O`���\�-�J���	@/'�p��U"O�U1R�ώAӪ�8�kX"?�t�D"OF��'i�6ƶ]cvJ�i|ؔ��"OjE@�ǔ� |�L��鞍x����"O
ur&��7)�<� �
Wf��1"O�91�6�@�c��@"FPL]ɠ"O�yd�T�gu6����0�;�"Op5�bG+#�� gM
D̴�4"O���FQ�B�P�G�;��*3"O�\
�.[�&Ȣ���I;/�*�R�"O��A@��(���;��|z�"O�EA� �6 � a�֪0a��S�"OFؑƦ*��$�2c$W��DA�"Of��NC�*���EO@�1�ԍ��"O �C�Cڍ`�v4H4��a�Z��T"O�jc���?� �1@��Y���"O���U��9��e� b�Kg
��0"O���F�*̌�ub�>+�z���"O̓�hK$G�<t�V�V�x�T�8"OV\�uޛ����e�[���(I�"Ov$*Ȝ@��¢L�*
� ��"O�d�&/�*����"9&����!"O�pxA��y�H}��!(t	�,jw"OD� �cR-[��H%`�	s����"O*�6��CD	�fDיa�H�s0"O�� -)F��M���
�g�09�f"ON���%��\�n��� D-S�d�aC"O�	H����$��i���M -�V�X�"O� "��!?ӜUA���!(�`-˳"Ol�G�L=-��:��0&F���"O*�J�k'�2�z3/D.4.bLy�"OF�0V�- �t)3Y-�>�;�"O������j��ƃ�*~�&���"O�U�2B�)$<�����y�S�"O�����Z��z�j2���Z����""OhQ8��K�|5N��O�RE��"O����(3~0�%
]�Z$.T!�"OJa�sሞӒ肖I�"�	�"O�8�Y����9�%�-���"O �ҶD�,�P8�E[�+, 1�"O�)���\�f��QC���E�1"O��2c�K�%<Q�2��#|�};�"O�ers	�& F�B�"؍G�. �"O∰�e�0cL�ɀ��(�"�8�"Or��W�St芰�1��\��%"O��9��C���qQDn�+[�J��f"O�A"C-C�o0�䓄mW&i�P�I�"O�|��̨~��Yz��a|llr�"O~�8Ra��K�&�;Ui]�`�đ"OڬY��<�֙�g��Wd�� "Ox����Wp|ℋ�!���S"O�l�AÔ�./��;Є��`�L�:g"O��{�I�-<S^�+e�ׁƬT��"On�a���u�P��(��J^���"OP����+m��X��4	���$"OF(�a�o������Y�	���"O4𡆏l��4hfJE�#���Z�"O���� ~�5+r�Ѓ'�@�X�"O��beH��Z�� ��/EK��bv"O23�NZv`���nQ8�)�"O� ��Q$)3~�ޭ:��O<k�Ē1"O�Pi�*ƻi!0�Pk.0ͳ"O<H�W�8�ĉZ[gɔPj"O�L���L|.�2e,X)��(�"O�+�.�V��\p�[!��Qj\�4G{��)6還��J=�,�S�i<H�!��K;S���j�&�4��BcA�k���x�����oޚ K~!�5�
�`bf�16�6D���a�<#�<4SnEi�0�귄5D�d�O�6����sI�y�,�YQ�4ⓐ���
 H�<q�x��G��Tٚ�"O��p�A0��3���M�n�a�"O�� �M:��)'����5H "O8}�$SI��}K���-�6�K""O�#��S�h��i���#tP�A7"OΑZ��ĥ&�����6k&��"O����H`<�s���fOv(��"O�\C1F�9m��i�שO�+^�E� "O���`
-�F%)E���(���"OT��c�̀4�h:�#� ��@�"O�aa  m( �*x�<eX "O:� �&��m���"hǫ	�V�6"O�x��瑯=��IVf��Y�%�"O�-��ER���w%[4i	�"O�u�A�8g5��d��}�S
JH<��u/�ȋBA��.��B\�'y����O�VL@��'~�H�@x�6+�'I�� u%Q<;�!S�M΅����O��=E��	X'FbUٓ��!�:��V��2�y2n%Z�8�	H�F"|Rf�[+�y�-��BM�>C�}31�/q��`H	�'�6��Pi��x�� �$b&hش�Px2�K�ri
ç��u��<�.���y�N7I���pU��>ۖ�*rM��yB�ͧg�셙�D�2!ȚY!ReU-�y��1eCԩχ2�ܡ��-ʟ�y� v�0�A�I��r,y�)�y�LU�he�X�shB�>��N߄�y"́7v����#Ѽז�gꄰ�yB�L�3T ��EGp��%�7�y↜�}�H��&f��a��޲�y�d��y:��ѡt����;T��X�ȓ+ƨpB�#@�:
r�hMR�b�^d�ȓO~N,�WlV�����n�^h6�ߴ�O>�?Y�K@9S�,�t
	T9�r
�A�<)a�˛<��*gJݚu�]�ƈJz�<i�ˍH�J����.>��A��t�<iD�ܱ0/^��H��%�r���kWr�<	w!�1��p�bڧM�\Q�" s�<����R\|à��/E�\X8V�q�<
\:L�b��egk%����#N�!��)q\%p���>}��!��7o�!����~H8cKХ��xb�ɍ<-!�d�/\xZ�4*��9��xA$�y!��*S�ޙy"�l�R2���!�բ'�L�+�t�v�R���h�!���s�zd�G�M�L[E�ֳ-�!�+6����T�J��:���f�!�Ćg�<�
��]@YJi�@H�3�!��[�ib���.ՑQ>��@�o�!��N�?��dQ�'۱dY ��>nm!򄄌Q䄡[��@���l���Yr!�Ժ���v��-��l����V�!�$ΕI�B��Wf�k����j��}�!�� ��CE�(v{j�z�h�'l����"O��)2CD�p�ˡ��wh~l�e"O~�1�B�~^�X�� /a�-A�"O*9�1��A���b,��0M�����jx�����%����$5��`�T3D�p�3�E!:����唬24���5D���j�RWb<�g��� ��i5D��Y��
z"D�!��,J}��@qO>D���晍 '�)�5!� JE�� ��?D�|�� ,+����#� pjmp�( D��:4ѣeJ
�!��+0�h��n8D�h���D5)t�tX��mMb-��:D����@�*{�&1+��ܵ5��tK��6D�����-p�����>-]����6D���@H2G>*���P��*��i�`C䉠Y���`'
 ̐y��M�u��B�IY6��z�Iq�j�rץ�W|B�	��f��c����5qN� }>B�I�>�+�x����"b B䉢$����
4� uJ��1��C�	�(}�)B�ӎO�>�7�ցh9�C�	*8N�u: mB>�.y�vO�/�C�	��D]ʢĚ2KgnP�R�ˡh��B�ɀE�Xo�4$ʓ��?IBbC�I�S,v��)+-�4#d+�	-!vB�ɇ>��y�����4����PB�� �@�X��	$� )▌N�C:B�ɟXFV0۠M]e?�5�PF�@C�	�}fD$SЀ�t���IL�Q�6C��-PZ�k5�۹v>�@�.̬A/�B�ɸlSb��RF/Kv�	�:N��B�	7��a��l�:U�AȜiM`7�-�S��M3�����>��I��N�Vc�lC�<��Y�3�d��Ɵb_X�����<Y��]3+ X41P�߰��t�ab��<��E=m��D�Q�z����t��q�'�a��LA�s�����NƷ~�"�@AZ��y2�V$s�v��#�y�~p@p&D��y⠟�"��u˔h\�H�����k��y��[�V��1��@BȲ	*���y�O�G<T�b ɖ:�20��B���yRN$U�4ZgH�?/IB:�'�y��EA� �,crY"����y�K��}�+ۀ,'J�R�y"��J5�Hi-E�x �1�Z8�yR�ƠO��9��fRDE��J�yb�����4��#tHO���ybLH�$47f̸�13���B�!�UF����6ۀi��͇�J�!�-)%��P�Cm���,D �!�D�3��]0 ���N��"'+�!���T��ģuCZ<	|�u�!C|!��/���逭ͽJ�ȲsK[,k!�<T�ACdF
i�@9��䀽T!�䟕��+sE�k���J����R!��F�3Y�L3��N�����%!�ē�=�<җ�څ{G��+W#��!�;'J��`0̂.M*�	�'c�u�!�d��tx�h7lڎZ'��j�!ߺM?!��۾v�P�$Y *o�����!�rf��A��S��(ׯM0c�!�������GH�ֈ0��ثFa!�d &V�"�c�늦V��	;C>�!�D �E��m����.��Q@WH��>t!�� �;�&�P�
0@i��p����"OZhR�힒){.iC ���`�*#�"Oj�B��� O��k4�Ɉ4
Tly�"O�P)�3ׂ(+��T%�ҬQ�"O@�t�U�@5bb�#���"Oq���Ίq�r��5�
��&"O�(r�B%a)���B�?O���{5"O6E�Wo����ʥ`�\��d#"O��FD�Ūb�H�@H�6"O8�[U�hD�Jb ����w"Oް O� ��!�eחH����"O(DY�gJ>9�-���I��Z$""Ohhi�����Bf#%t��"O�iZ�Şz����</a2�H�"OD�� �!oNȓ/P�$CT�A�"O�}B�җ|?j!�E�\3~�r"O�Q�#ԙ�h��A>|��$"ODq�J79�-���NR����"O�$�1���i�l]M��bE"O����)Q�d0i�l���\$�"OL��e�C�0�ʀf"m�Db"O��j2�/!di��a�aP��"O��@�Ɖ�T��8�Z�HZ,�1"O�ā��E[�x�ҕ�/ ���`�"O$�P��S�F�(t�Y
FxΙ��"OR�:R$׭=^�m���\D�جI&"O@���֌|Qh�c̊Ѽ���"O�dCG�,;���H���O���(�"O(1��.6���1C�*� ��p"O|����Q��SA�rM�$b"O���,^N,�� ǎnB��c"O��!q��
�(4PV�J��0\03"O�t��
"�C�% �n)4|��"Om���0��)X"�2��4"O]��	�.� �	�/��1CQ"O�X�.B�M��T�3b�0PZ"m@�"O��	�2��Ȃ��L�mZ���"O$X�S"A�w�H�F!Y�]A�	Z�"O��kѢ��}���y1|-�F"O89[��`���pF(�Z/��13"Oz�Z3���m�y+�G�k �)"O�����>�r�R\�=����"O|�	V�Ǘ�\��T���/���"O�੄�r:�=�u̒(�"�"O��J��'��u�E,���t�"Ot%���Ƅ09ހ��KB$)�
m�"O�`(AO�0G��Ԡ��U#�=��"O6a��#���A��k�8�P��#D��AAo�Y|��
���C���#��"D�H����rǰe�c�4	nr0@%D��"�ˀ`s�+Q���@�#!D��Rc�^�O�}S$Q����&J>D�8z#�1+Y�ljDh��}��O'D��(u��(I���bTlV�i�DP{�+D�PR��?=�@�C��	�K���vJ(D����$�}�n��Co�H��#D��zU��0֔�&�W-���3�#D��AL�	��Uԧ��%Ԉ����%D�P2SD���n��R;6�,�t#%D���%�\�'��4�R!�6TV	a�l#D���5k*RRH�S.���TL D�`��,�
��IRA�&��#�>D�@J���-X�Gʝ�"���+�C<D�$�sJ�3ఘ�m�](@�;D�� �h��.��p�I�W��"O>�c�j�I��k!K�ua
�y"OF��ā�~��d����Td-C�"O�Q $�N�Q�.�
CH�'"O"m�7�;	��y�M8'b�	�"O���X=w��y�r�����(�"O���]r�	�J,��"O����Ú+{R�a��nQ����"O��oD�]Drᱦc�"KX�Bv"OZ4 �a�D'�BC�B��y�"O��"���e�t;t��B����"O4�)���Mc��W���8�����"O��a��e6��!P'�B�A"O���W�Hጨ����9\ۮlZv"Ob�8#%s���Cb��f/�I�#"O��f�._]$���@C#6�x�"O�9k�kD2D�%k����c"O�a�O٫PI�АF@^<^�k#"O>!���\�f����������7"O�u1U �/Z�b�p�(I�)�>���"O��µ�H1d�	V��<քdq�"O���v�A�M*�k��.s����P"Op�R�F�2b��'��u�"�"O@<���R�e��ř�Ċ ,�e"ORH�ڃV��p+�M�;�q��"O*��� ��,k�,F�j���Y�"O���P��O���هa��]H"OF�J4h�k�8<�4��fj�\��"Oj�k3��rx�˱I,7$��'"O�aG���>l� c��"@4ލ��"O�����N7d(>��U��>!��d"O��ТA��rFR%9�	
 rb�Hf"OX$��cV�?��10�e�j���ʐ"O�����˭6A�a*A��e���U"OЂ�(
bȨ9���:���à"OB	����o�t�bܣV��I/�!���d"�1
5u��h�ĻS�!�./�X�aԯ���S� b	!��U&4��,�#ϖ1%T4B�_�O"!�d�5n�#6���z���nG'f!��&ER4}��!Ѐ��J �A�!�$�
*��x���.n�<��L��$�!򄈴 ��|r%DS�qef�z�iߑ%�!��2�z��b\�k��<ip!�$H*.���X�`P�a����2bA!�䂪6���A�@'^�����T!��(S���@�s�(sf�=:!�D��O=���I�sך��6�753!�_#��yA�mϝ|�(�k���w�!��C;S� ��2eXn���$
1m!��&'��ub�P5@R�|�T�H�ak!��24��㏽sO4��FAN�`!�EZ�Ԭy�'΀<?6��O�#U^!��H.S�3�.D�@������7[!�%4��"����ݱ��E�tx!�D1STĵ[�lܝl؞i�aL0R!�Cd���Y�-���H q@M	N!��3!3��I3�V�p��;¯B,S�!�D� �� ��Γ�I�¸�q.[>1�!�$�x�P�IM�97�[Qs�!�D��qj�u"�G�@���)rY!�$U S����ތ
G�X���2U!�D�?#�����5U60����(Qp!�U�&�[ve�~5x)dO�Iq!�� ���1qf6��C�#t5�"O��g��8X�A���ud~� a"O��`�n�1��I!$h��J�T}�$"OB�r�HFl<�P�1T�,��E"O:�C�n�p�8"��S刨�"OXQ���[�M�X�����^�|X� "OX���d� 4�$q�����4�jW"OH�+���"��h�e�"y�����"O
�AO�;��)��!W�(�P"O�(��GA0-��А��	F��xr"O���&b�8ش+0�֔w�X$"O�e��P":�]B�-$iȢlx�"O����T�w�<eb�l�{����S"O�	��jT�Ae�����/p?��D"OV�����*r���F�Q'
y��"O搱��,R����;B�L�0�"O�D����-|V�ȧ�P�d��i�"O��	���I�j%��&���"�hG"Ou�WbD�=���D�� ��!�"O�(�p��~�:]8�^\�|H"Ot|��d k��A����XJ�"O�``��ն[&>������q"O�P���M4\�	J�M#݄��"O0|[����~.���!δT���B "O�䘦��G�i �.ӄ�Ȗ$�y�IY�xF�,�'��rs��{���-�ykI��H 5쌏nQ����n[��yj��|��ͫsH��%T�X��G��y2�^�o�:C�فY�l����y��ؙrX���U"��kn@��yB�M�Zɬm0�3)|h�o���y�+��M?rE�h���� F�y�2<�Ti��0�l���^�yb�]$x2�#��јx�=	�z�<)3 ǲC�Y��D9D�z�4
�d�<���L7B}�7�I7j��T���^�<9�f��[����?=J�M[gHZ�<)�%)Xc 0��ʽA@XD��]�<і�ռBC̨���=.��\��$�V�<��Z�ipP���[��D�ɆEJ�<���~K���1�@|��(VQ�<I���� ����	l�0a@�M�<)V�R�����NH��Qʗ�t�<�p��$��ْ�G���Ge�<!��?�$E�!��
������\�<Y�D $dGm�SHA<Ū�H�R�<��
��fA������̰'�N�<a����%*�SPam˖�z��r�<ap�*t4@ʕJM�K4���oIq�<��	�J�.��D�I���u�v-p�<�VÂ�\rČ�p
B�IR���.w�<y��N��/�.%qxQ� ��s�<)�������8KX+`����{�<��M#+佁���&d�zكF�r�<au���"c�Q��ѦcpХ����n�<٧�@�m�������`,b�S�k�T�<S�ٰ�$=	�mY=�@�KO�<Aw'���`1� Ꮪ3�@�´�FK�<IdA_|��9w�LI
y*��WQ�<���Wz��6�Ĺ�5nV��*B�ɇ+���⎍�p�P�a2�θ<��C�	W��%��H� *.l�F�A*x�&B�	#�|�S"��`�h� b�/gFB�ɫ_j�(S)P' ���v��1^�B�)� ��$w���$/kW�<�"O$�D
ǐa��P��y8�Ѣ"O�0�f���3����	
��P�"O��R�'6�����n`�"On����O�Tp��+	�=�g"O���䝋���v�©U�H}��"O� ���W��г��1t��<�V"OX12pO@#k��I;��D&��l˕"O���b%����q�Ca�e��:�"O����wK�w�$4�:AY'"Or���ٹ@\Ⴁ䏬4���"O��	���	X]��B�CG�
��#"O�@B��X�t���R0�юa�(b"O����	g 8u�υcl8�"O.��!�%B����	28.U�"O���2d��lR��3�&c�H""O��{�X�$��T9�v��9��"O��!�I�:1bU F�O���"O08��(dHYP����2�ڴ� "O�e���}����U���.�L]z "O�-�R�ۤURu!���.j����"O*(��,�r���J��Ӷ�-�yrρ L�ⴺ����`��0RF$���yr���<�\�4'�-Gf:������y��a�������?;z ��\��y���	�,���E.0������Ȉ�yb��?j���4���
`4JT��y��=�00b��J3<p8 �Z"�yR�P�eä����;�.�1�&J��y�`�5o�H��f�ق�$�T�y�_'E�Q@W��K^�H	�ŏ'�y��'P(�R(C#�Qaj���y
�2skP$X��7ST�ퟬ�y2*��V'�:�D؇C������±�ybL)�2s
��m�"���DĮ�y���#\��;��ڻ_I�������y���#�0ɉ��b�Z����A��yr��&.>���N�Y�\@�o؃�y2I�6>��e��R<VQ�)��n�!�y�j�sI����#D|CL�yR&�:V���"E�T��qA���y� �(Q��!���ؘ�	P��yR�ŕ��p��@�����B�W�y����:v�;�Ң{�Ą��K	��y�B49_���d'ל⶘F��y��֠�E+�Ҡ�uJȪ�y���;u.�1��	~�*���>�y"ELwE����٨qA~�{B���y��V1LV��+�B>x����k��yr���P�q�Bǖ ��<����yҀ�jR�(�ƌ��x 'џ�y"J+KEz�)\?J%L�g���y�"�#C��H�a�E�����Ҳ�y��HQ�Pɉ�O�'��񃷁�:�yrIGIj���Y�T���A�T��yb#�:cW>�RA�"PrNM�q��y�� zPU�EaA�w���W�$�yb�NI%��!I=n�ְ:'�è�yB�*,�: Rˆ<����Y��yr��}�L:��^𸚦���yb��$�d@@"�!'�1a��/�y���@�R}����#�FS�c��y�E>Abd�{�(�;O؝0����y�^�
Qh�(�'��E��Y��y
� �Xp1�K�"����Ǡ*e�y�G"Ox��@OW2�z�Y�*�C���a�Q�`��I�5����C�# �a�#��U�B��St\�H�H�z ��ۨ<��C䉈P�0��ˀ���Zq�>@��B�I�u�R�̖@| ��f��y��B䉅|��Y�҇�;7PՓ���)�B䉷]��X�2����C*�㟌��I&�����CaҔ8�0���~ʓ[�z�0��EI���	5��)����<m �Ԅ�*�AKÇ�;+���F˵%1�|��+m�q�G�ߑv>�{c�0o8T|���pA�*�z�XsddC,fV<��ȓ� �������:S�f� ,�Э��d�i��NB�A�2�������ȓ~s��Y����c�84v���X�'�r�I^̓7 �+��=߲��t��.Ac(t��V�������	gt�[G)ǧ�m�ȓ~n������1l�T��aL&]�fȅ��`)�T�_�&��s��-C�u��O%>$
�J�SN���@\g�مȓ4�0��nӠ.S�AkDGҔ�$����b��(U�Q�î�7�h�'�a~�F߶M����b���6�	p!��y�OҀ2��	Q"՘J�3D�#�yB`D	4X,��DoPt�(��%���y�	R#P����퇇QB�x� �yB���"X�ҡ�A��	����yb%ا�j�9%f�	+ެ�c����hO����ؘ��-�� �~��KTFQ�W��	/�Ȅ�z3�H0l�x~"��	�4C�ɫ_���d���"�Z��v� %�C�
öl%X$hdX�Z�@C�I,t�(@��16��E6C�	�>���CN��hŸ�8T��U18C�j<`X���u�tZ��)"C�
�P����%|�d�p@��˓�?9	�D,bP	C��E�( (s��5N{�i��e�4T2���!W
T5
8~���,�ڍ3��C+d��Z1n�>X���0�~�#5hڏ��u�e��I0.l�ȓ#El��'� -���Wh�J��%�ȓT��y'l�&h,J�-́]����ȓt0&�AA1����ƓN�Dܖ'�a~Ҡ�@������J���Q�J�y"��2_��!���"r�YC��I9�y�CG�1T�t�%�P"k�X}{ࡑ8�yb��J3h��>gx��k�/���y���2|`�W熁cfd��!F��y�*jx,mԪ+i:X��f���yf�:@ab��%��_��æ1��9�OӃ	F�0�.ēKׇ8֡� "O�X�+ĕ<��h�� 7T�%"O4�`������(�l�ް�r"O4��w���������i�`"O � e��3���:��OR��T��"O>��1F,g����m�%�D-C�"O������'�,ݩ���Cِ�0Z����|���O̮4G�?�r��taǻk�B���'Q��P���5[y:��t�=�P���'�aS��߯K��TlH,B����'MV͹f(O�/��3q�M@����'�<ErrK��_`��ٹF�j-Z�'U�����]�U��	�_b^D��nT�<� ��@�"�:Ex���E9 ��qT�܄�I�*�p�z2�Kw8nu��U�I^B�;x PBUM`�@"�I��<C"B�ɧ"(���̛�lL|�Q '[�"HB�	(���[�%ޡ�F1{'`�4�B�	&~*F�s!#¢m� �h��G 1ԬB���VM!G@H8!ܛ�Oćx�B�&|Q2����(7����DXB�I�b�P��� ��uYg�n�|B�	�S&�8"U�
a	~X�($B�I%�@@��	�sX$R����4�C�	�["���aN��TЙ�"�6NR~B䉀[ ���V�c鮍Xנ �LΘC��61q0���O��q˄��>OjC�F��2��W$7Z��b]>,B�IK�����"�2:�H����El��C䉣�XAK�KQ�_���U큶Dn�B�	�,���1�M�T�Б�⟭j��B�	�W\�8(c�H1,��	�(J�>��B�
�ɇh�q�@��;L�`B�u��m��mڻ:WZ��v� 7�B��#T0�th�=1>�VB	<��B�I �0� n�֜r���"bC䉁�&	 �싪(���آ`I�pm"C�Ʉ_��uK4J�>_�ٓ�m��2��C�j�ȩ�"Y�Ua~0A
0ϸC�	�#R��V)B�`�j �L�C�C�I�or��0�����`�@�>C�	�+�a�)�|;.)�hE�]��C�I0Y�� 墆YE��x��R� C�6HN!���E=g��1�0 L �C�ɞ3s�9
��Đ�bi���QVB�I+7�(��L�f[.��R,��|B�	�4�v�"��{���
/DB�ɆI:��R�L4=���g�@
��C䉮.���P�n5}���p�_	m�B�:bլ|Jeա;���G��+IUB�?��e�o�D]�(�(`�B䉲#`Ҩ���r2��J7j"B�_~2�z��ں7[4+���@@C�	.M�=�"��t,�Azri�1��B�IIy�(��k�(@/����f
�J��'�E�OR�SH@
i�%}J�
�'2�d�A��]&�s�O��W�)��'�4�C��ɝ:3pQ���?w�X��'^�e�u��P��{"�յp7RLb�'\4�X��T�u����Fo��)@�'|���d�X�?/��ڷ�I^�d��'�<�����Hx�gAZ�\|N�H	�'��xi�LqN��ǩ	�,`��	�'���#�<l.���@�4@I)�'Z��Α.m���(��ֈ&����'8DH@��[���O�<0�F�)
�'�"�J@�t~��Gd{6\Y�'��0�#��kG��+�
 q�`��'}\ ��B�:*FƩY����pzĘ��'�*)�"U�(o�A�"Ă�fP�A�'�2R�-Z^�cB��:�+�'�	0f�''����'[�Ҝ��'M���f."(��J����6	�']��;%��E�^�ٖH�������'0��jGʘ\"|l�*	:[׎�	�'�n�C�A�n��TY�f����e��'M�T����0|���6�0������ $�y! �'>��q�l�t�\X#"OziR!D<Z�2��Vf�I����"Ofċw-�6����|+}�"O���ANB�B���m�	r��q"O��!��I� ��x�k��
�.��"O(�طE�R�X����M�7"O�y3��D4n��9��+�QJ�"Of��S�K�0B%
3`Y�iG|{�"Ol�2V;s�`�gM�8[�`�u"O"L��Mӊ9`Y�S�ܡ~~VtBD"O��{�ĭW��!1�ZB��s�"Oh���B�O��e���	"1��(D��%�L�c���ԏ |�@��!&%D�8��i�`3tU;TlQ�!�xKU�=D����E-M��P��*[U�|�! D��ȷ�гf��r�@��-t<U3��2D�$��o���S�D��a�q8�1D�\��cU%N�u�W�8,*�2D��<u�l����7�����p!�3�̰��A��i(� � Z�5!�M �������I �X��n*!��
B� J�O�s;��k�-Ļ7u!�D�\��y'�� !2 �v��*b!�ě!,ߎ�� &��[��1r�(.~!�D	�z8 ��ɉ(��jԫ�U^!򄆅~���J�*�V�����K:|!�d� \b��#u��:p-�`���� r!�d�AJ^�{3(���Ej��˒(!��̣{��"ˣ8����@`\V!���!Ne���/��ph��,���!�.�1�u�ݕ~}�P�a�@�!��9��ׇ�!V�(���(`!��R,8��q�P��?��"Iƻe�!��W T�|E��*�
\��UHBa�!�$J�m7dq&)�t��*S.��B!�̈Mz��j�d��G
"Y$�+5i!�P		Ŝͫu�B<��*���/Q!�DH�0L�ÀD�F�����T�/�!�Q�	WX\�c��}k
(�H��L��	ܟpD{��Į8Q�_�30.�C���y��S�V)�-x�9����y��eb�`�D�,�!�ș
�y�H�xR�iC�9D}*׀��y2��G��[���f@`s�y�A�����c�J�P�i"���yR�6[�b1ɣˌ/I`�@�Ь�yrô*�hɲ6�IC��W,��y"�A:mP1S�
b��E)�װ�hON��)RH����ż�~�ak݂M�!�䏈V��嘧�=4G�Hz�@L�@�!��]LȢG��_@>1��.T2s�!�DʗwML���'���A��և�!�dYnRmx�E@�y[ˆ�!X!��/)����jѣ*h>x�!�'z:!�D�;�^8���Phas3/({#!�29��ŉ��|ּ�ˍ�4!��T�2�yF)ҧhD"��ר�!�$�����@AD 48�N<O�!�=�f9
C,�� O2)j��*F�!�D
s�V8[��D<H�3�9X�!���M�XA#�LBF�+WO�x�!�� ��x�GΉV2*a�1O~�!�ĝ!cZ0��@�.͂�)G��9K!�D�]��Q�D�ZT�=KHUh!�� ��p��J�L��x��܅P�h��"O`�&��q�Q�7b���V"O��9U M�yg0d�de �N� ��R�p��J���5!
8b.y�#H�#�U� 7D��2!A�3���9&�/~��)cVI4D�"���>󦹉�&�+�T-c&�1D�`��f�0�Ġ ��(P�2�Q�0D���"g׿GϮq�5lԨ?j�D�o-D��Ҭ�
�p��6R�N����k-D���ݴՂ�#�/�Z����&D�����	[���D��aj8�c�$D��Kd�W$?;T=I�M˥y��Y��>D�(�f��8DD�� �> i���D�9D�H��q�8�1�Lx-#<D���gAX�����@ΕM��e<D�����Q �T(��螠w����	&D�4Bf��9�(qΛ�6�Ha�bD#D���C.�'P�������=p�4u:ea#D�8��-i�.���&ish,`ч"D�tK@L
 N�`�a�'s]d$�Qk!D��E�ƵY.��sj�.�>��!� D��C��ԋSG�-�d聘Pk($�+*D�Ȉ�)��v�+E#ަP�3!(D����A�
���j@/�7f��+�� D��2i�Mqv0�`'�ꂡ��H D������;�Ɯ3��Q�N="�*O⭳���-=M�H�c�]�"��͸^����{|:Y�)��Q�h���K�K��B�I�q��āG.�8.��D��8B�	�G�P�&�J�A1�r) B䉜6�P���gR'v\���ϡ}B���0?yʧc��Ђ�/\�C���#@�l�<�g흦1ඝ@Q��R��E�j�<�fd�]�*�c� ҭ!ò�� �d�<���}��i*�K�4+/�����x�<�7��KA�M�H�&t�b���Ox�<a�!E�w1�T�ag�J(P�Qt�<٥)C3iv�ŀfa
?K씁�*�k�I^y��'Jў4��\�02��Ce_(��(�J�<�G���W�*��ԯ��$��md�E�<�`�S;%1XeSr&D�R�]
iW�'Yax�`ѶE�r�G�&Y��镗�yR�ԈnE�2�c�3*H;���yBi�n �L�ǣ
�%�İ E$@��Py�&Q	q�ջ�" �OG��e�YM�<!ALu�]����Tb�hI!�s�<�Dm\�uxE ��O<~4�E%�l�<Q���Y���tᝊ`?j����AG�蟼��e�dB3mYO��9�Pa�Y��2D�\{��^���Zf���	�1D�H�^&wƮ�4���;�d���-D�`K�f^� �&�Y@�hl�d�я?D�[�4'D�I2��Ј����/<D��q�>fuT�iQGM�g��|jVN;D�<Qt$��LfA�g޾3�{7+ړ�0<Y��_<sTzH��-�]�3TU�<1� ���%<0���H'D�P�<��/\#
�2�� `B��m�c�<i e��l �k�_7S�j%�Vc�^�<�#��7h1�P&O���R�+AX�<q�d�U�rhF�-9Īìp�<�@bE|%�4C��Tsj���Ct�I�(��W�k1�[� �,i��)>OLE�F�<D��jG�і'�������=)�0y"C�/D�� TH`��}�>t�)�2�����"O<X���_&n�8|�QWI Ũ�"Oip�@J�vp�g�	,MP=hA�'��Z��'���
<i+��}���!���6��1�7d�-G����X^ơ	�Ƅ��z�R�H�U��'��)H7��l�P4���B�4�ȓ)~��v��K�"�N��T@���p`�$R"+�Qg��IR�A4��4����Ā��grv���>�Ψ���H7 (ր��Ñ�tm<L�	F����k�+)1�H�S.ޡ�
��ס3D�<��K͟ *��u�߱��y{eF=D��j�E�5&xY{��d)��;D�@� )_`cE֤M��7B4D���FU����	�H_
U��dy��,D��;-��Y���#�랞}����W�?D���ܲU����ħ�,e-��q�;D����]�_�tm
g@_�1�*�Bԩ4D� �,T<5��E���-`�T8Ea4D������\�qpv�	'�����0D�|r�F(r�DH���0F챸�-D�T8�NY-(`�F�.��Q�g.D�L�1,K
Y,���-�?@��H{�
:D�P���Ӷ&��L��F�e�
H�WE-D�x�vh?qP�4 �i�53���&&��0|B$n�� ��̑P���n �B�T�<��K`�q�cb�5�<ɛ�eOP�<����@��q�tɐ�1��� L�E�<a���g�uR�I=Q"��� D[�<1�o\&<,����8��L���b�<i�����r�噂 �Xh���f�<��FGk`�1�E�&N����k]z�<aƈ9�\P��G�I3!ٰ@Pz�<i��ȭ4�`U� ��%2U���i�~�<�	Qv���D*S(.�\m��
y�<�������h�AZ#~���3�t�<��/E0K�T�àIS��a`�Ct�<�0��B�`]1"�ŝ �������E�<	v��\�P׍E�Sw�� &#E�<�����C{���g�:R�b�@0�Cf�<Yg@B^\-��L�5ޞ�è@b�<�F��"}tB�Y�F^ '�$�cNNE�<����fE���W?0�����@A�<� �Y�m�����EX;<�9���^r�<�6�fLQ20�\�@��`�6�Ew�<i��A��ˆ�$�~\xCq�<�U�5D�R`�G�J�g�v<��p��0=�F�>O{ؘ���B�,��$�F@l�<����Bb�q�H\�`O�88a�g�<IfeMt�,h
�cXTD�`ENTI�<��D&�0U�u�Kyd�X0a�I�<�Rɍl�0@�A����@�A�<)s�ܹI�ʄ-Sv䤤���B�<)Ro@.\��h��Æ�+P6��Bӟ��	g�IA��~��'�|���]'?�6�:uH��yRFԖ}C���1�U�lz�%��D��y	ˮ
���tB��Z�6�!t' �y��.���a�蒿J�L4K��P,�y�g�X�U�!�M*-��������>����yrA����SC�L��m�1�y2�W:Pu~�Q�nT&��̺�N_��y���v%8L!5�#9D���j�6�y�1e妸�&K֍-T�E@e�I��yre��(w��e?�,�	��ƾ�y
� `���B\�^��d��#=m8]��"O�p�T��bª_�>��Be�'~r7O��q�e�3]�ԑҤc+ ը0c�"O��K��M�
}�'��N�j�"Ox�J�I
9P�D �
�I�xP�"OF��ed�6_%�%�����"O���h�X��l
W�Гw�>�bG"O�u�� �P����N
_��iq"O�
���#�$�rVɞ�3�h�P�"O�e�A�RJ�s��W:6�ִbO��B�W�]�2)��{�����-D�|
�&���F0�*���)D���H7X�(��3�#w�ŀQ�)D��Qqd�%��xi��E ��0��2D�0��%1��T(�Ar��s�,D��r��'@�ؕ�ͅ���)�M D���3g�c&�C���)p����?T��b$�  �33��F�I~�L3�G�@�	Hp�G�S�f�`C�;D���4(	<Π���!DG�ByHa:D���Tu?ĭ��. �8�ⱑ5�8D�BS�ݛ%�e)�õB$v��%�7D���Ϸ!��}iC)0��hA/ D���Ū��1��bW�L�0s�=D�����6X��T�ל,�R,p��O���G��'���#VK&'Wn�X��	�RP8�'���$I�&nєe��ɘ(;�q�'�,�
6�\ 
��@���~.�%�'i���n��W1��f�ۇpՖJ�':�����Ԯu�-	�E	%j�UQ�'��ţ����Ũ�6R�xp-O���P�㚈���٘��0ꁯ�+U�!��7ZȩbZ�F���U��!���* ���������)s�H	�!�1�hݲ�C��)ɴ�� ��!��F9��ĥ��Y��p� Ȱ�!��Y�,�D0#��ۊUi��E��.3?!�d��1", C�Ǐ��t�p���m-!�de��[� �)�P�#%{r!�ʰ}���j��Y�y�N�1�ڊMc!�Ȕ��b�&ȣ	�l�P��M (!�ĝ>6ŘriY�i�V���	ܞv!�@�f�(I�nV�G��J�g�"=!�d�B�R"�B��I�w�:�!�d�V�Q�@F4�Z	�uIѣw�!�d�(�X0��$\�8��+����"�!�Ę$��H��fæLP��C6Q�!���k0���Q�� 輵��e[��!��R'�,]p'JC�a��d��_�!�]1N��oL)+沔�p,K.�!�;h� �s` =k �K��;>n!�dA�V/Z�6)O6h@hJª�&�!��E��Rڧd�q`��̜;j!���T1���r��K�0�!�KK�.H� �C��H��*	"p!�$Z�a��X�aA��~�"iU\!�D�s��}3pd�j�|i�g�L!�D�D�|q��.�.��U�� `�!�$_��>d��*�lĨ���]��'��'�f�	��!x�,��$�=w�%0�'Ĩ�ᕇ	�%G�x�ndK�mFs�<�OXm��pySL_�{Lp���E�<ybN� ^� ����W�
t�D
�@�<��Y�Dg�]��O�/5 ة$'e�<� 8��� ��,��E������JR"O��m< ��bB�F�V�� �|R�'n�a�h�X�$�s����h���'�$�D� �pq��*�� ��ic�'���Yr�˃Z��R��w`!0
�'ֶ��4a^Ͼ`�ˊn����'��k�#R����Y"`�nК�'�N���¨�a������'�>��Q�K�*Q��{�/3�zUi�'T�i�!�Lp���kL����;�'@�.57�3�,@d�5BNl�<Y1�$���㳃A�X xӊS�<�qY�H,H���[^��VI�O�<�o�Ur��h�I=0{�!J�<���+�@�ҪQ�
p�S4ƞj�<q�C�*�-c�^�������c�<QfT�2��a����$�n��!�U]�<��j�x`�d��G#m
8�{֩�N�<1U��-6^�pQ)1�`��ŕJ�<A�B�;+.�A�K��0�B$�JC�<����,*nh	�R���;K��EJD�<� ��$9h���ҟ�ڨ)��z�<�d��\����jÀ Qa�M�<�4�ʾ���ڿ�n��2A�,B!�1rn�k@	K�B�&�D�!�
���A�J�$(�C���0!�]]�4�P�i�U�L�TIV
w�!�D�6T¢H��l�697�`�\ �!�Ď�{�����D�1Lq:���*!��U6̄k�{�.D�U#�$>!� 8{F�P�a�I��5��@�!	!�$Y�7pçjZ*'��I��<!���x�",�����)���z�!�Df������	�F�WG��d�!��m�,�����3fM��D�~�!�#CM�7�W�d��eb�"G�U.!�7�aB��[O�F�1��*!���2T���ݭ���4��"O� ��L�v�
e;�Na�Ƶs�"OX�1�����b9�¤�2k8���"O6���/H�8Ԋ�C#L?��(t"O����ݟlR�q�'���U���@"Opy�a�_P
$������*ON��L+N~zI�э�#��k�'���(6����h�*с^���H��'�x<�B/�nv@��7��%� ��'��m��X�Yܾ�yw�H�����'�Н�6��!5���S�����D%`�t�J�C[R�rWE[�~G�Ԇ�d��lF�]��HAhF5;���������0���X�d��
5)h�B�I) �{�KX�0٢@,� C�I$�I�%���!�\)���S9��B䉕��%�8�X��,� �B�I� �ʉPw�M�b��ʅeY��C��Kj����\������eV��B䉃#��h�����t;��%��B�IZM�b����r|6K8df�B�׶؀@b�
D>TjԤ��X3NB�	��fM٧C+� ��l �"�B䉥y�4\��GY&�ı��	�m�$B�ɰ,$`Z^X���e�=c.h���?D������M��Y���ƋD#Z�br,>D���v���0�Z�/��p�Z���7D�� �x�gAZkKN��4���bD8H�"O<AU�6J/Ƽ+Afˈ]vTc�"O(z���!Ph��2�D��6�x1��"O��X�F�9���a���=��t� "OҠ�`��QpY���X�<T��"O4����r�L(���ً�|ma"OJ�H`�M��b|Z�&P����A"O~�:���+p�`u�W2**��Q�"O��J	�q �g�@��p��"O�e�oE�>3���� Vcv�`�"O^Lq�G�o81H5 ˹USD\KW"O04#"�<C�Ԓ����^RȤ��"O��&�j,�� oL<-O�]��"Oh�p��c��$: �W=65�AҖ"OLq0��1L	��W�\�1Bv|Bp"O��i��M�m؂I\
Be "O�9;0D.���*�g �h$�d"O���@G��o���wƙ"��Z�"Oya�+S$qb���44-��"O��f�==�X�{b��.p�-I&"O~�jЃ��S|A���$(�NHp"O��3�./R�F��c�#%e����"Ov�)�.����h�"FL%�"O������	Y_���#���'IJG"O5#i��zݚ́�`@t9�"O`����Q
\�q)�B��;`"O�"`�13���:êY�28�" "Ozar`��{R P#���#{Ĉ!�"Oʝ�f�3NӀ�:7J�d(��"O`\!��@� �z���ɂ=:�P0�"O��[�+ۖt(�iҷ�9̬�˃"Ophf�ɏ]l�@�)d!<;"Ot�����W���;�c:�pt�"O�M �%M��� 2@>��c"OX�󈁒(�j�d%�(O$>ة'"O��� @'.<cץ۬Kr���A"Oz�ґ��(4���A��0y1"O����/�&:<	���Rz����"O��DJ����s�� Dx�H �"O�Ik��M^,$jWǁ4�(�"Ojqw�5'���*�E�'j �C"Ov��`�ZCN�x�	�x�R�"OԄ�)��v$Z5�A*[
mpX�"Od=kc�٨c�49B�KA�j1͊�"O�����B���up��'$�8�"O@9[v���Rd�ŋO�x2�"O�����l,�p8v�˛5 ��S"ON�b�ٕ)d�9��˟�#&�)`"O����'�e��Ia փ}�F!��"O��y��Ͻ8�,hс��8�D��"O��$֖:�� @qB��vIt"O4��Fʗ\���с�: ƹ:%"O����t�FEA��]\)"O`�z���#�n]8e�N���G"OV	��T)?���w���i��{�"O�} q�Q9y�.��4�^�gW��!�"O2�#&䟋�YA"�?w^��""O�!��M<�Ȅ�Ǣ��Yx�S�"O,��f� #��=RbB+J���"O���BZ�b��5�C��J�H��"Ot�y�/^�G�<PaG4��c6"O���C� |�|��A��3$�X$��"OZt�g.�a�)X�d����"O�#]i`�
{hh	�%"O� y;h��B�p-�↕~���"O |��� )�SFA!Aeza��"Ot!B�L$7��W�P��Bm1�"OFK��/D��+���8x��@�"O%˧%]u�OW%Z�漻#"O�a"��Ɏ'�L��mI���"O$��m\�tz��b�-�>�2�"O��`,H��L��+\�D�,��"O%:�%\�'L�Y�D*�zD@"O������&I�$C�{�N�A�"OZ�QhI�x|]�6܎��UЄ"O��rA�O	=�vY@Ѓ��"'�G"O 8 ���)	�i:逰Q�����"O��t��B3mȯ�q�"O�8�#�E�.�����T���`�"O8�{�Aܘ8]�!`H��a��i�"O�(`ɆS3�$覆I(/��r�"O�|+7h��2���e��[#4�#""OlE*T�o��Xg��C��R)�P�<)��� Ȥъs�N�y9^��2�I�<�dO�.��MhF�	;�f��%�M�<� m��(�zQXp���z�6NKL�<ѕ�L�`�� QD�[%Wcd��EP�<9pdöGx������x!` �#�M�<)�L���+U�#����`��t�< ��y��0��ǂ�`��eEq�<����X��M��,W�r>���( l�<	qK�Xx!%g�_�I�"�r�<�C 364���K}A�\Ӷe\m�<Q�OE��@��,d�
a�h�<�'��q��	2��,C��f�g�<�'��I>���JC%@���&�g�<�l�'@:��䓤')���Q�_Z�<�’��T���m� �)W�<I����c�ܘR��]@�U|�<i�A)\	+$�
H}��i�~�<�C*�7G�$���M9\�Ud�<�DJЏf����cn��̒�*O`�<�J�Vi
��' X�.��rv�WZ�<9��F�����Ӑi��Dr�m�<9`�	�f�fu��?� ���a�e�<�v��	JCp�:s'�.9SxD���Wb�<QS���u�[��@�{f���[]�<����o�ة�ǡ�kU@uA'��A�<i�.=6F�9q�M4>Q7\D�<Y�Ɉ]�|m����1K�����_h�<��� d���[�*��EZ@� T��[�<��I� 
�%z�蝩Qؠ�5+�X�<��R�a��:���%k��`�|�<����e@�HH���mhu�z�<��K�U�j(�3��23B���K�t�<�4��78o�z�*�y�Q`$��V�<���0ΤD�@*�7Z��7/�M�<��Ҧ$A���Y�4������d�<��+Q�d��y���B�z��x�GEI�<���F��dU�Æ��R����OB�<��

�c}�hp��	�/p�ƀ�A�<�R��$������H�Yף}�<A��m��Y�6G��n���C*�N�<�d�vH�����?}��� ��OK�<I�'�!Y���)Ԩ�9�RA5�|�<9"��'Ra҈Ɇ�O�|5�X{'@�m�<)D�(�z=Y�%ڳ.��8+u�`�<Y C�\۠U����0l��R�@�Z�<� ��*�*�4/��3M�"���v"O6�kR醩uP�e�ǅy���*V�	�S�Q��'k�*Hc�����>F�YB"OT��r��X%� �`�o|�`q"O��p�0?j�r�.����"O��Kb,�3A��Eb7m�4)d8�
#"O���X�]_��^�p��� N�y��x2�a��#�!]�r��rǕ��y2��1��ѲQIY?XĤ��Ш�y"i���,���:�NQ� ���y­  i� }ك Y�J���{ǀR,�yR�e�Xt���ĂL���e�
�0>YK>Yt�[�Aj��I lo�i9t�G|�<!D�ʳ;�YFhq��騐f�ux�d�'���B� �~���#���2Z40�'6�4�c*�*)�Bd��̀���)��<��	�fE��SDI	:i8%�����<���Ӓn~Э�R	�&9VL�
�c�.c7B�	L�"��� ����s��.D�C�	eLҕ�-!G����6�(0��1��{�I,D���L(I�J���i״�fC�I�_V������Դq'T�_�C�	�w��D(0�5|�	��	�.
B"?1�O�b?�dEC�y�N�h��J&N�s��b���'�'*����"$�� j��Q��YC�yb�)�S6)��ܫ2-�$L(�BC��-�d�3,(�@3��˧@��Q��=0䰸V�(�IQ����FI&vdXJ�E\�}D4�@�!#4����g@�u|0�C��T����fHE�<)��`��g�<6P�����ID�'�"=�'[
N���Ğr�UQD��(?��X�r�i��n�X�O��>����Jp���`	�_~E�DF�+�|������OL)�ѺG����TT�l�!�"O��r�I#~�Z��.Z: ��8{��Oj��D;}ғ>Y3�)x����4Nǽ-���B�. p8�l�S��|�A�;`o�y[R�3h�8�/7D�����Ίe%�|�G% �&xt8D�4ғ7���h������M;r� &/ͫM�z ��"O���DB8
jX]q���+=|*]&"O�i1�l8!��� Xu���d"O�A��נS�RB�	2Y��e��|�%%�Ӻ�N�lۃ�
pi�D�ѣ�K��]���%�O$��/$$� �J%,x� ��ب(��ąȓ��q�����@��T+.��1��IO�q3X��sd�t����Q��?猱�����+��Q�'��-���H U��i�*8��y��'
b�	6�څB�Р�dP4'@j�X
�'�e��TFle�1�� 
�,�
�'�<������)�'�  J|�'�@����'V�����  HT��'�P!���#��! �/�2�0��'�Ρ� �u1��a�ʟ���Ԋ�'��u ��K�J� ��%/�.�&�0�'E�X���ft��ٴ���|���'m^t ʖ�Gd������ �P���%�'B���Iw���{Q"�4	����Xh��BE#B7�2ͻS#.dw,ąȓS�P���΂�*|n��h֨YR2�&�P�7�����'IQ>ᙄ�Tu;����HH"N�2-PC�*D��BDjG�S.�E
�I�Nb�ikfe*D�0��f��(��2��"JԪk�E$D���@j��݅]6"ڄ"#��h��ꓣhO2�Gx�핞;��A�0K�%b����!�y�K�Q��*�D d1� ͦ�y
� R@�l�%
2q���]6zhN	�C"O|țq�T��¨2�S�d|$0"OjP
�
bԣ�h�4I)����%��� ���Y�p���ǀZ4�5dx�LA��&D��Q�k �r�@��xi�Y�b2OT�=�HN(H�P�3�H9�L�sk�v�<QvCz8Y�ǯ\�NT��%u�<�d+�:�ڸ��.�c����Gy����?�� N�y���o	 Ǻ�bCJ̓��=q�(E��!�6��(�J,z�KF�<A',��r
a�.�HaH���F�E�<96LÝEʖ��1���X�CLFt̓���?�<��'&~�Qԍ�?�Ԡ�dX�@����'�|�[��C�hP��C�\~�pi�{"�'#�i�����Y|����s��}����<��h���;Ră�d�[ǓY�<�k_
N�6�𶩞�`��I�Q�k ���h�rX@OT<7\�%R�CD"�(�B"O�ك#��,k������0�p	� �'�ў��g	8�$µ"�/{M���s�&D���1�J(�pdۂ��6l���f�7��w��� ��򔮟�":db`��?ĤC�	�K�ܭ�SE��AO�T��i�'+��Ily�|ʟ1O��Ss�U�j���g�+`���"O�\*��9Z��Љ"C�U{lm��i�8C��\5FU�e�T
)T�#t����|��V�p�O?�ɘx��i�W�V�t��-�WK�:�TC�	2z�Ri:F ~( ���= �^㟘G{J?E�f��<ypB9%F�)W�	PL4D�lۇ�6'����̮n�=(p+-�ߙ��=���K�w̐��|�P�Bv��JX��'���1O�IA��� J�D���ǳS�n� "O����@�Ex8��F���v1���'���ūoR)6mݼ���[B�ό,
!�O;O����""�!	�r.X�!��
o�9��݉D����CB%f�!�d���d�@�'U�E���[�g�����	V��'���F%�(v��B�	!]���Y�M�"AE�M�3��W;�C�ɉB��H�$䜷R�0,�@Ι�9�\O��6�)�uYx�2�N�,a�D�%��@�FB��8���C��` �P�t��H3bC�ɫ����g����@6�%�DC�	���@$�
?)`�8��n���s��7�B����dͫ ޕiDę�%���8�L��'�Q����I��H�X�O`-&%���ܯd��B�I ��3C��� ��7j'}��"=�,O��|��A#S�~@��(Ğ ��@����Y�<�)&u�(�q�@� \W�<!Ư	�AÌd[r�J�n/�M��X}b�)�'m�fd
&��!��T�*w�$�'7�}��M��r��H�F����y2h�%%PőQf_�x�mz��#�yҀ�&v������N���"Ѣ��y�'��H}�żdߚ��v�@m�%Ɋ�y��F�v7��'���9��#BS$�ybL�8���i$�ϣ5N�8��@���O��=�BJ#]�4��-QD}�e����y��R&9�lQ#��J�+8�}[u���y"�)�YqI��d	� [5)��&s�V-��f�|��U�� �B�p�9:�|��!O�ꄅI�ZS�M�@ ȝw�����%��4(��C'Q�x����.��Z�D�2>��̂4y���S�? �ЋV�ځEa(�[7 M�"��h2"O�E�q�S�����ÏȬ8����"O@� ��2��0���v,��"O����IP�|J���Z*E`X�"O�"�A�S@���:d><���"O&����˄A�jQ��!2�	id"O�T1�"X;؄Hb!%�/b-:m�C"OPd�W��	u� ��õB(��0�"O๚c��Q!^y�œ�N
���g"O��7
�'P���	.9c:}H�"O��X����{(�:s (j(Z���"O>,0���e��b�Pq��"Oq�R�_�$I&�2L]T�L �"O0��k.e*-�:�%"O�I4I��s�Z��e��  �\��"O.L�d��z�,	Y �1z���e"O�IC�B�9$2Ga[s����"O��P�ԗ@�nI�s� a����e"O���!�8����Q
p����y�(�_�d��k�=g@�h���U=�y�؞dlh�Z�vEZ-���,�y�G����2Qc@U:)ĈZ
�y�"U�*W�P��jP/�V����#�y�ˋ"~rrԐ�,�?�>쓦�Z)�y"n��$m��lS�~�4E`&�(�y��1t�nh�Is�nP�i]��y�Ϩ6�H)��B��j[Ps�ȥ�y�o�3�艗��)j���!k_�y�)ثr{�����Z��X�!S��y2�"7^F��1���A�����ڜ�y�%�x^����k�7B��d�u�Ƽ�yRˉ�Whz�r�E�1��)u�©�y�#�'�LT@d+�<�b�fgB�yrDR�P��-�l�=T�my���y҆=j�=h�Ä�)p�(��M��yL>�<8�m�!�ΡK5���y2AX���C)��˔��y"f9h���#��x~��i4"��y���0Q�H�E��1J Zܑ�֜�yZr��xC�ħW쎐��d�xA,Շ�Ts�l7�Ư5���#t%HWX �ȓYu��bU�#"U:�3�dD D�E��~{`�iE���x_^@�'�C,W����3Ʋ����N<�����)c�4��y�>}5nӥ>Rl:���,2d!�ȓju�՘��U��� J� �>�^чȓ:�:�y��P4�fX{� ��q�ȓ+�eze�E:C���*�K��E�ȓ?�6����M�|h�E��Q�<���KU�E�� �h,��M&Ԟh��_`�Xy�É5=�����%��ȓ\A� �P��z��	rg�<1-�Y��(����I'U���g`W7G t��=,$��R�@�|%.�it��,K�F}��
s� CBN�=A����%�-u���ȓS����Ҧ �.	3��ê9V��=��!Շ�~�2��	��(����^&�((����T�!��S� %�!�ʯ��˵83�8QpaҲ#�����Ol�xX�+q��@J��Zj�#tO����#R^���9�!xĀ�x@ W�,9(��hO1�و�@|M��	�s��UH�D7u��u��I'M�Ʊ+'�U���!��M����{���U;ܼaB��̖��`@6D�\k�ȥ80	�Ȁ�|F��R��<��"�eXE�K�"�ԡ Bi.ҧd���B�A�5�e����#��Ą�S�? ���FΈ="Kf5[Vϝ�b=Nu�@���o���䖳e����T%	.�'f�qO�x	v�/]��A�6��y�h��'Ѯœ�N^�(�@ ��X���H��ĉ:�3eLF=��e�A�BT�����Q�f��$�%V?����2�W�L0$�'�6�g���&�PB���+s��h�я��z�,0�%W?*@��R�V���ʂ%J|	F"O�\���;3g�"��4�6�	���z'F̸A��SG���I�p�ۨwd�u&�k�w���h�C�X	n%wJN$bbЍȶn��g�4Ѐ�{�����1�H-��'ױ~���T��--�S��U xsn�G�M}���rl��3�D1ڗ痰z��8yOm��g��@���;RD|I��5+k� ���pN>��?n�(b��عQBvQ bĘ>0�J��`
��$18E�$3�����:t��#�h�P�E�?)0J�!
Ll|iG�u�R	�E�
%�b�cs� ::�py䑟���FHD}`X�bȂ�cf�l�Z/g��Q�F*�6�fK�|^Z�y��_<Gr@��%�9g���"���0W��Â���>1�,�e� %���_&W��:��P�jV�0?��YU�@*3�f�q�ԭ��	S�TF���;��<i� X-������0���M�݀B��-}]�D@�bi��`0��Y�f�矬i�bj��U�n�jT	�&�%�L��6(��$����@4dnd�Q�o��a`@�hB-Ys��&�X�ə��!{P�;�H�!!c n�R�yP�ܳ,��k��՚6t�'����ıPdX�XPe[�ldSg�O�`�13��O:N+u����4SF�۲1�����~�I����3d�M�;L"]Kp�[�
� Kf��-u�*���1����2wU��3���x����ݗ<���(ոT�l��_+:����Cd��C�B�!��Q���gU�p	4�
�20.��42�T�C�+��h�w&f��iыr@�M9�w��&
�9]N�`3Gu�F1��n��������3zT�!�Ε��������\* 4>��1�J�V��,�C��
lG\��$,�,U��KJ�#96���+y������ s�X���ކ��'RʁZE��1"�"�^�%�&59��ϢpK��I��(g��Ahrn���J��[�=<�Zv�_�#�"99��O!vH��I�Z�m�t9K�I�P���Jve���FF%��녪82�I�H�d��@/��耂&�j<�IYU�C�3R0Q�HP�d_��iJ��Q�4cE�4��V�c��@QU���3S$a���>Q5GJ)|f�Y�捝	<��m��n�:sE�<���6.:����͗n��Q���Ne�b#��򩎾a���2C�S�~5hDT�uB��sV�L?$4�A��!L@mHW�<e���#c��z9@bD�pO��֭S�0%��@��>��Uag�� i�|�z��S3̼�*�uW|���6�ӕwRt�ƍ-Q��A�eDUj��H�4?)�-�p�$XC�ui��D�dm�3b؁˲iµ�[�Rg�YD�>٤��E����N_�����O�""RU� 䝝2
�镋��Kl��bB�	C��1�N�[������%/@q���'9̬� 	*B[�� m
AZQ#����bą�lRO6a�(K�ܮ��M!I)l�9�K�?5�nIB���*�vMѶ�R�R�C��i�L��%Y,,���;��{d���D�6jY���M�6�x��g��*�"�c���(��r�\6���,��B��61�H���vhN�i��4
Hw<  n�	�T��`��=�� Y�� ���l��HDy�	��JI� r4�'	�P���`ڃ�y'^V��h3�]i�@��&T�0�Ah�{
�F�O��.=
�|��%lA"!��U	�,͘1����Z�,	�b��]�.��q�ز p�إ,@�$.�$ʍ{�P(-l�(A���;ꄝ�f`����O��b����.��i0�0�l�*�l��`	�*����#���]�f-��*V�K���"*��<P��ɓ*|d�h$Gb=��K�@�]��ɣ<��Q�^j�Ū���8�d r!#o���m�2Y�)��g$�5;�h�GmF���V�"C�	�~P�r��t�6X��E9;@��@G�,B��P8��B'�Z��3�Q�y\�R��u�<DHR��;>I睾)����!��0|�cT\������.R��i�ć֟7���?Ƞ ��	���d�I�/�Ѧ]���3,A��c.:e�{�"�t�q%�Ԙ���>̺E��<Hm6)P�2��*z��՝cи|Rt
�%5�����G����8��P�N1D((	<g�D '��Gр�#U�'���[�� tX���ƆD,D ��X lOIY
�*#�h��ZT@�� ��H�T�Q*1���f�E�A
�`�,N�OV�J��ɮijB�z����mM�$kM�!R	�g�J.ǐxRiE� �@��$(���+6胥�X�	���0
��p.Y��	+�L&д�g��bu.]��2G:��;P/����Ù�^Z��. (*��'�xpy%�����c(�d*z�`���W�� �A�L��J� >H�`�_�t�"�����f�!��E��y��ӫ]�"��6D��^r�8O�Qk��G�G������0�j1���5'Y||h�/\!?�Z� s��/��YK�EGC��1�#(��3�|��k^6#P�lS��֐�����."#��{�	�&�|%��	I�I�,�b�|�'n�*�$[��j˥*�L�K��Z<t�|�g�Q�M��D�¯T�b����q�O�~
͋��
�,�H�S޴~1�ع����u�DБK�x�3��]9F,��[�w�'��}���H�v��*��E+��{���6mM�i[EB��;�\��&��<-.�!�3��U"��s��o�L���"�9��U+�8�^��)�=.)�=�c߷W'�����&�H��RhR�A���A�'=�yY�9*�6�Zt�[��+����"�X���/@�����8S:H!%`�7* �Ԭ�=�L���"P��)c"1H�������X�B5:e N�6.	�T�<��'N� �(���=Jl�񯂯`�XX�.�5f��Ė�6�zViĦM�� �#��?@z��aoC�f�D��=p.\��ֿz7��S�Ô(�й�C��)�f��ؼ�8�<A�/C�,�ĕ-2g�bh�m���r�K۪w��:�*`��yɦ
O�!���*��qh�
�8O��
bKڨp���"�F+c�Xpq�$HŚ�+v`��\�2���P�U+��"�Nd��!c�c�+I1)"�(+R��/ 2�B%r֩���D�.X��oۃ2ś֌�@;���eK���7m��t���C>��' 
F��h��W���g� ^$�P޴P�0P
�:8��X�D���8���� �0����OH�d���U�d[dv��q�K6yÐ-˷D� x�ሯ�I�$�ѾhS�O��J�W�p��ܫ�h�{n(T#�j�ZW�H��H��ᧇ�u�L�$�"J�f���)"�H`�� BD��&J�$���C"(O�S\�������,b��Q��'��\�˒�(UҴ�Gj�0�68�3d�� �T*��9y�451ӯ9C��H���'f����
Ӓ3�>$�D΋��P�z� �!f�Z6q�0Xi���|t�n:�p���:J�1eC[4(L0���3�X�:P�5D� ,s�'>��!�T/ �"Q;t+@�9��C�]=����h�~-06d� K ,h��3���h� F�)8F��c @��z���-�Of����:{�)�*N��P��F�-0V��� ��h��Mn�	4��2w3�a��U��."p�ΞCQ��ݖr�J!	Al�#���$�;�k��h ��ړ/FJ��T�qԐY�hNS��-�"��zcFEk��o��@Heڒ,G@��g�Դu܄u�F�ipr�p�dͯ>� �yc-��m9*h���tI����2��S+�;H`|Q�b Q82/�a���ɶ$��4账֗+�KÂ�˒xc"�
Loly��'#�i�l��hb#K�Nj!Ka.}2��sգ����>����2�>����J:R5f	�w`�Ml�I�Y &`�J]�vm��0��ؕ ��M�x �J��jw$�_خ<�4��!�ao�*^�6��ɦS��H�'�z1����$�@!�rI͡x�j�K��ף~��!�I��+������580j�G��q¾�����G��T�C@�!vT�
l�;=�
�X�I59��DA"{*���B�T���Ŀ��y����<��M�
�*ӎ�#s:ٻ��ޔU����_Vl�%P ύM�Te�L?8d��[����� �%Q�����&�p=���.�(�Ʌ
�
�.dJ��4.}��J@ʓY�� �OB�5*B@ےGޯ�&��J�
�&pb��.y��b���tq�@r6 �q�1@m�$��x�ˋ%~���m�lܜI�!	ධP��I߸��&͈�0��@��
'p���m�iׄ4����㴴@"�O�|>X�:�)U>�J4 `\;8�aybL��6yP�@P���s{���'�e,�9�ۏD�R(���1�Q��$5��P�m� �$�1/�f)�1	҃[G�Bb�Zf⌞Ql�8eE�)����0}b`
�$^��w�� F�T���j/ ��X1��>|�f=r�śE6,�q��R"DG�H�備8e��Ab4c��D�>�D��^+��[ϓ)�����>}b�;T\;`��!�B`ϓx��ػ�AW�G ʵ+6���-�0�w��<yl�{�"}yۥ.�v��3���3D�[D쟠B#���	T~���#�M�+TP�1P��d�"��m�n邥T��P1Y|~H�q�	6|��L��*�]}��8���L�'���.�VD�N��g�l}���a��r��'�)��˂�"�8�GљX!��!���RBX-3w	˽G?��{5�Oy��q�D��u���$�̼R>АT'��QG^9�I�>A0�'�@{�(��]�|=�N�ci0M�O��R�'�i��T��F_lE zeK�c���,�$n�Y�V�J�:�`�s���'Dh�%����/i��3�׺r2�H$晣9[L���iK(�լ\D=�t��#|0du�f��\�ҁ��1KW0���V�l@�E��	�FiKG�hԲ`�03 �m2v!J*��q�D�B%��I�2%���W�Vm���v&9qجSffN�+TlR��ʪlt�m�cg�:dg���%ףRd����Gڤ?|�=*Qb��v$΁wM�a�AϜ�9<��Ѡ�-O�C����၁��e�@[��	L��usTO֊Q2t��gIj��OX�A���8�MY&EmHa;��H��e[$O��1O2�$#�A�(�z1+ņ_� laƓ�T���	�|i�b��%�t ʀhS�\(h��k�(�bPp"	G�( R�,A:t}\��7�#�&�ڢb�3{��{�g�
{�,����r#4��@�ٱq� ؃��}��k�Bҝ3�=[��-�p��G���w(,����w�4�۲���{��#7B�U��IЩ%x\���Nb��D�M$�Sv�YD�i�u��h����=d�M)�a]�_�>��f��O(�{&a��G�q�J¬l���¼f�L���dϧc� {�	L���(��mN�t*�- ��<�F���Dt��FG#H��M�@	�*4ǋ�9D���4�	���Ғ A0Ct���äثH.�$���٠/
 Gxr#��[`� �N͸w�zh�d��1�~҇��ui��s�c�:�ՁeZ/5w�G�]�C5 P��!�^��b�����J�KZ�{� yR��Ǟs�
ma	�(&���>��m��gp���P���X���K4����HϠ~�:!���o�3�ۈM?������x�(	�� ����#J)������¼ ���&�,ժ�- 4$⧯Nu�D��Łf��4K�I�u�;���f@(J���5}e2�M�[8��;�AE a

h�w�'SZޔ����>gF(B� �7xQZuE�;]5���_T��e
/8G�@A\��x��E�+P�кd�~2���`���h��) X˳oH�Lh� �r��0��uN��>���dF��.�te���	\�t�/��Jc�$��������X	�4K��(�m�0T!3@C)e�l�s�'7,�=Aab>�:&iW4:�E��>d��L��e� �^��N�hD9�m^�MM�̸B�ΑI)�!�&�$��X�Cˢk��MZ�eвHT01�rmG���X3�9s]=��eR�*�V(�K�0�ԥ[E��KS8��mՁC�����;w[9�4Kі/�>q#a�E�� O�p����{�G	9\���:dE
�J�Faq��58|��ӕȜ,DZ�����2Q�1����z9>�Y0$I;6��S� ��	�Ԫ���C��[#˘�S �%�@H �0.�a�dh�=@�fP�4Q��g���VȊ����e�#�|�ƴa��-J�b x��P?5S��S�_/hY��� �2��t9���9C��uIF�)(��k��ؘB�\ r��C Yȅ��e�+��)rw�J�3@O���1
�$!�zA�!K+L�p��K_��q�V]���D�7���qJ�$&�da�qEK*A�\��+ݩ���A0J=�DR�!�?&mbE�$ 0�t���0��⑧W�1O�<���ХR��l� �2/�~ݳ�bH�PΤ�W(�T�q�RM<I"�p%aM�}��ܩ���)�z٣BH�S°���[�A�ҍ׽���`��AO �A�#T2F��P��#V7HŹ�+����l1Ĥ�"�#���(� W4k��"��9��x�2�
~Y�fʀ*�ȸ�@kH$-j��I��6n�
��"��
��p�����#q�-p��[�O	T�t�"B\��ł�'�a���XE� /(�yI��/w��KΟF��b���[b�h��K����sa�I�7E� �@W�Q��l�@��?`��1���$f�H����k1F)��8- �yu�Ɯ8��3#\*+�����Sxv̙�A�9Q2Ʃ��O�Y%gF:���(���F�X�^�(Vi�s(�S+�V�~��E�D�f��`g��<��U�>�dO-c�P����i�?  �#sČZ�-A?t�ĭJ!���~�a��+��k)\�P(�@�%yΘBѽ��eB7*���:Ի�N�69��k#.��]� ���ί�O��eO]�lq9�&j���a�[����F�k�<A�ʘ�gؐc BՌ#	b��'����F܂�japKT���sEl?��.����Z �͢�U6f4��'v� �%`�즹ڦ`L'g�Ĳ���g����t��9Rtq��FU�^BP8��Ċ0-2�3p�W�mj\��5$�boD� ���'M���eEW4d�4�IEg@�~�d��jO�\QxU[�OV���9O>a*�.��ʼ;�@�w�:��S�O�G�Td�P�L;r2�i'��j�����-ͶG.Y����v��
�D
?O��|S� RN�v�A'-�$O�r�QM�AL������%�Rǔ �L��LF����$�h��=
�H�*���`��CM��`��|4
��qFSq�<����f��\�Ћ�_(�l�$�Qs�m��9r6g�A�Z#}�����[������NF�ح���n�<���%
�0��ƍ8:S�
�_!�U�� �@�S��?Y�e�6r\zM�#!I��e���c�<��$(G���b�C�1�����T�<����
>PX�돹C`����z�<ɀcM 8�P�0vQ�5���Y��i�<�������d�5W�h���m�<Y�[�8�t!��ϓ�j��XAJ]�<q� ��uu��[1끰 ˞�2 �q�<��B�0>��aQl�/4��c��l�<A/́>�DБċȧ������n�<�������VA�
YĮ`p�L�f�<��������CdH�	ؒ�z�<�0�
Wp���#X�� ���C�<�mD����x����x�7J�z�<1���P4	�s���I�T�s��L�<a�LO9`�Q�ጇt��9��J�b�<!�Ӗ~r
�C�`��r��(BG%�b�<9$&\	Q^��p�kظ38R�@3��^�<y�i֢HZ�#�H��	�&ѳe	�w�<��(G+~| ��C�1qIz���Fo�<�F�^�V򀓴�����f�<A��H8�덿<JX�����J�<	j�R���r'�Hx(�qE��@�<�p�	i�"�Ѐ��a�\�j�b
B�<y�)L���)Cщ\�O��e�SK�~�<�GnٖV�N����}M�,
��a�<y���s�B��Hj�"����C_�<a���4#��}��U&0�$Q�6�V�<1��&h��t	��ԉS��x����[�<a�˜=�qF�ބ+�Nqb�Ci�<��H
���m���QE����B�<�C����"!9�K;Q�.��W�Yy�<��N�0g dq���� @t�<�ub�T� 5 ���)�9C"�p�<�5�!i>���u�K'R�
A{�$�p�<�V��� ���E)	��*怇o�<	�OKe`�F�B7
�x���a�<��-ʳ ܞ�r��;t봈r��3T���@��%W60�q���!�"y�f!#D�TX��<vV��vcM,l�Rq� D�l �j(��0��FF]6q�U�>D�l�4�_�(l�Db�N�M���A1�>D�1C�����*p�!j�e��a=D��R+ǦH��+�f�247Lɛ�L,D�d�C'DI���P��"Gw~��!D�ܲ��ŏS?uA��P@n� @�>D��uǞ�W�n�S�;II�h(D���O
R �J��R�f�\�׬-3}*�{��m�OX����]X���Qa�6*�
���>��	0���0�Y󣗫[��+���Q��'�jm[���>�NK�zp�d��Q��r�j�uH<���HUdLŨa�>�u����\���yf�"���C9|O� �#A�S26�I��(?nF � �'�$԰w��"O��1���}��BL�b/������4\�0�a���y�C�F`R,`HQ�Ka�%��3����OPd���h�J�OtZ(Tϝ\��0p�g����

�'yvY[uc����4�c�*![��y2'�P>�E`�+�=G�:�eʘ��Ϙ'��@��W�S=��C��&���{�3���;ҡi�|�Si�'7��D���Z���b��+P�Y:�H',l:9��펬7^�z�� �������G;�� ����G9��kY�4|�7��1Td8y!� ~r	�fO;�X�"��()��͂ ֥"V"O��
��Q4.�L!2�*��<(�@��E�+�M��Ԣ�±�s�L6mR��J�O�4��	oq�V�k�e� 5c�RE���z��`�1$I�	�4Y#�5�)�'p�n� �W�����<(�8�۔�����	����W��z�Ḧ��Ֆ9�����DJ�ت�k4�O5�~�7*Ĵe��
>G���I�h�i���'L�Z�ԑ:qY�)�t|k��"{ �LK$��:Z���S�j��bB�ҷ��Aۊ����+�	w�a���qƀT�d��Y���S�E�v$�!A�D	�����FX"H�t��X�~L��p�5!��9�kI ����m6w2"h*�-f!W�i�qOz����	�TQZI�va���ʐ�O�"�Vic%Y
b�L��)ͫT���O�W���H�̄�ڌ*U��|��LE0`.��؜w�h� ����up�D�'vh��J�u@>����~�#?U5l�CrIՍ���OP٘QC#Z;Z4�� [� ���+$��V�. ��D�M �m"P�ʼC@�Z�¡_6@V��i�س���Q�R��
�4�4CF/_�\��M�1k� �@�SK;vܢE�D(��+O(������X �O(�.��4�F5w+�h ��$��)�#Ϙ�qlD[��ȇ�b�[R�3;����AgF5t,��ֺ'��˓OY�x|\s��X�D���2��<�D`PiȽ2Ռ�v�z0@�� &'��|sf����M�.�c$<��������d	 ��DI޺k<�!���].$�q��ЎL��7�ǳG�X����1����|b���x1z�ݏ;7
1�E�̜lH&5�#iD�г�\!����`u�����ħ'��\3�M«uhj$���Vt���\H�T���A���!��צM�Kɞk�P�ص��:7���RǑ_��I"b��vJ=�!4!��Ale^k�Nu��/���	AO>�P��4�> ��/(*��+S�ըBo����E��	��$!���Q��u�&Y�*VrM����6���
-O�T�U��)#H���#*���D�/����pj8�ʬ���(����%u\��E��S]����Ö�rBqzr�>�L]��� ��[AC*ȸ�$�GMF.S�	Ӑ��a�H*EUtQ)FmHw�O�j5 ����q�Ab 	��g �Z�	�T�Y '��%�B��@P)V�~`�a��p�$i�d �2�wnr�	V��n���dKg�*�!e&c�XU+�'Y�(�%	k�gy�FWc�6TвN�y��Q��ciʬ�4nC�/�n��ghߧ3��fL[M�"d�B����q�H�@�@%D� /Ʊ�B�I�{	����� T�JP9��ܚ+�ث���)���W�̒UX%
��"jܫ�H%U4Pr3�F����&�|�Ly��e�4�`��!�xҡLl��Xq��<{���	�8bD�5Cף�ȉ��ƛ{��.F$��[�C2=�q�'�m�r��"�>�0����Cp�LV�ԋ]%��k��קW��8��1��W�V�� ��Q��ȟ���#
��h2ř!/JG�L�A�.8���Q�� �҄�����S�Y���4K�/HB�l@Q1�bEI��>c"�)�?f���`��qO��a��in�ɪ�7p�3��ʤP*�%����p��  �9 ڼlrEB�	�01G�^�?`�S"-��V&qOD���`���NB�%�Be�V�	I.���N��s�0H3∕$m^��T�U�G�R�qjT&bވ��ć��L�9�IĘQ�PMb�-�p=�@�2|h����BW�g"���#�h?Q��G���SqDX%(`�ؽ2�b�l�b)����胩�(���ڂ��� ��J��!��g�<����'��	��S%W���GN;-q>U"`��Q$i
�~���GR�����%�T�̨�.O�����4.�!E�G!K9�� ���z�����3�ΈK`�įp��;�m��&��1Cj��J�2�4{���@g$Հ6`X)s'���[/��
����-xW�τ�UP@�:Z�t��r�I�Q��{w��w�`7�U/P:PUl��k�>�������ʰ��0Vz %�֫:��O�yp_JZ��$�A�r`*�mء>�����·�!y�d�&`ږ5����I�l�2�'C�D�jLzFm�:����$N�-$s0`)�I�6���2�-k����2No"l��K��ᰤ�;k�LXCAڧ=_$��T�	
A�ˆŶ0�a�󅒿M��0D��k�FDK�!�$;R2��;m{��(A�m����.�=2x�'�!cp��I���eh�h4H�pa`�r�TF@.A��h��V����O�I��W�͏�l]�j�#���qQ�٭=������6��	"p��F�O����)ŤN��؊�"T��X����\=m�TD�I
-(/Bq�A�Ũ{-�����&J����B�Ԧ�N��"�>i�򐈃�2P�@�D���jf8q *�;@�S��ջF~钦S�'1�40E�Ĝ"{v�����t�|i�,�J�^ H���:Id� B�G�`�����ꅁVvn�ÔFO�r�xq�4V�@�@ꎍv��0���R�1�|�0���jo
��$�JS�'s�8ɳ-�-2�r��b�9ih��tG�=�P,��3\]�� �e����FE�l�zh���~ �HA��
�VfH�VM��0^U����f���*�ƅ�n�4h�g
`�n��%U-%���'~ �06��Y�@���ʣ(8$t"�gd�~��enխ$��Rョcy�}�˟G�m�D�'��S��7~��)�:J@�9���;7,�i�׫�F�q��D$���+d#����c�mG|b@�V�S���K2<�Vė� �pK��g$���oMj-"���U���J�y� y	e��7L=�v"6;���7l�rV8��cԲk%P�<�f��7?��Ӈl7Ya��r�R0`%�MB�OS�G�4L��&�9+d*=s�b��� �3$�ô]l�	�g*�m�R8A�6P��ڦ.	�݂�Q=tx�k��K���T�4�S��t� WΝ<7ȁ�0BߧJ�,A!� ���d�?DN� �����xҨ��nOx�ñ��˦�P��L9j�	�|<��2�fL,-�Y��4��XP� ����ʆ	����-iRh��Z#��8E�.5	 �^�#@44� b�,18@�S4ґ	��b$�#�����#;�J�D%�UZPD	���y��<��D�KQ>�eD�n����l>���C�#=P���4�q�&ƙ0>��E_;d_8�Ac�rfv�a)O�E��$ǏhK���E��M{w�O#R�s H��WP!��,qL����pX��Zb�0]��qt�s�<ac� jZy����� 8��6%� �V��O��<P�!Ɂr�2eCrk��jWE��� hW嘍H���a�Jh�v&K�HOx`�",ƌ �jI����>tsE�$.�xĀ�iW�U)��3f �!1f�M�V醄,�x�k�]�c �F�L<.�&ـ�z�\���lA9Ei�죢�R�|�ǨS�	��L��+�8���� ݼ�?� �K%k�2�ʳ�]���CH�:
��l�˂�:��5�A@�?;�(��@&�>�����bް5�yɡ��.Xg���h,�#�P�!\��F�>��O��Qe�6!���@���?�,QKIP��|3R�_�UR8q𰃋0����(��"���hUES9�S�	٦��$۶'2��7�
'i�]��lI�y[b3LO���7&�X���V�Kq0R"�W[��S��;TbE��g�#%��Y允�<�HܩS�w� 9r��~b�N�),����U~�c�	�t��ی�MJ`e��>\� �g��L/�ؔ��"VQ$�1"+�a@kq�>8z� j%eB�#��6��h�ɔf��rR�X�R�R�y��O�ġ�LՎBX�	���Y(���$T�h�f/QEj�82�ӑ6p�9[���Vh��X,���T�y�N	�,̦/M܁a��@�~0�h�$�p��d���]w���G���JF �ܟ�OJ�Jqa9����B�r�hD�����'�������(Z!>`'!�?SZ,��̦�3K)�r棍~�"y�E�ِU�D�2j�`<����J'Ye�zR�Q�-��v���)!T�3f���@Ł6�8��ccQ�'��\j޴G;�( ���q~|��$�IȐ�{ԃ�:�`�0�.��W�.ՉD�t�����l�� �0��qj�'T3Oh��J��=p
��	C
�avR�D�دFf�3� _�3��Y2&GձK`��R�V�ql��� ߣ)ĸ�#���B���)�GQ�a��Q��r=S�,L�p�쳖#�n�x$��b�d��+��m2�V��5�@�av@�}��c�o�t8Hc���g�d�4�(E�
��N {��Q���E�XC���7�@*�r!"��ڡ\V��I�,p� i��Q��z��e��;��y�D�K��V�Zoʤ�a
Yx�@
�G/\��E�Y�/��K3��9 � Db��Y���тn��6~�aB�c��B%N��5iY*��+��46�q�aF(U�X���nW!A08��[���a��F�> h�E��bJ p�!��~�	����Z�0
����MK�ON�xD��k��È P�®!��`3P'�n "��\�y(d8xw�*M��e��I�������8vSFAj�l��_;��3����u뢢�(0�kE?<���@�]7(#�p@B�c\����Aȟ
��U�b�I��Ml� �,đ��U���D�z�"*��k��ø!����	 ����`2��8@� �32�,/��2	��/�}a�M�t/��"�H�.�x���4;�<�bY+��<��дnEq�AJ[�[�Tb�� y��D�5��!��)A� ��|B@��hNU���Z�-Ȅ��HV�f���x4H�
%�	7�Ρ灇�p��R��{H�T�B�ȴT�� B&n2��Q��)��TK��"!g(�6cHJ�\�∉6S�� B�S�h9�0����*��q�I�^�ލ�C�	n12��	�H����g.U�iT\�	DH� ��Vǎ�2�h����ÿ!#�����h{��CS/�
l� �c�"O�^Ԁ����=0�b��m�|̓>z`Ea���l�b�3��&2UĘ�'��Ո
LIn��aGGέ,�n��M��y������K�up���2�Q�~U�h� U���Hq��bx��#��$�HhňK�����b�n�a�"&-ֹ��#��Qh��=r�"Rb�l�)AҌ^�g�v�C�!  &�6m�%��y �M	�ڑ�S�F��$�Ҍٰ`���$��C���� Ȇ`\�y��eh(Pq�<a�T`\4JQR����'���+��cZ�a��l!DYH�N�c�����(�f��4mR�=��������.���`p��1��}�����`�@S&L$L�� ��,��D�V"�7dq�6�^܁ �S�m�P� �M3B�h;��$ƿ)��)�jK�8��@�-V����	TX��q���a�n��g�a�5e�qa0�9�+�*}6�maPi�D��k�jS6in�"�'�r��)Tn�:e�0mG}r�F)P��I�C �д�I�����]f���4k�!u&��4��(E4v`����H��8'���OΒ�B$c�7Xl���d+��yW��Mі05�N<U��(t�!��'�*�tb\�u��9A*�]�'(TR)��6���xwN5	}�X��e0-\�3�؈t�L���*WT%��ž2����.��p�l̻M�H%W��~,��� ^���H��t�!�q!�3or�D$�ӷ9y�P0�%B��Uitɝ�F��������< q��F��D�	�R�iQ�Ȁ�P|1��1C���� 5�	*IҔ-H"Y|��"��U�4��ܴ�L���N�_,���VP����|�����tuhUi��n�b����Q�:�����-��`���G�&�<!�Oy,*�ъ{�a����
�&Ӹ����P�]��豤����1�Gh!%�E�M�ORDP2su�Ƃ0Y�����%��qGl)1�iO�X�JЫ�i�&k�P��E����h��B׽zr�����_NV2Q�0Z'*+p�ۧg,{'؁UǯMkp����!4z-��zcV�4�fp�P���pk1�O.=|ir��
��(���I��;%J]��X�sĄ�f�P=a���7Q��=Z�o<AF�MA�LD��mU���B�j�"Lߨ�R%NБ:��*��yT��hp�.x-�C!�,1}r�ş�"�J��V�9��rcgF�}\��XH<��d
&s�>�)6k�#Jdq����oK�LZ7�Cd�:<cDצ/>"t��
'r�"�Q�+C�"J`E�r���uIY���zT�������2s1����K�B.���Hٹ"< �<���Y�&(S�cY�
�"��&��-��7�}�p�N�d|+���
~x�3�Z'	n�D���!jj�hq��5�Eʰ�td)F�o�=�oT�d;e� &��fb�`�@�֥
�r<����z�@A{6C�lti���n�PM��'�[g� R���v�͈�zy8ɠ�Y�$�$�b�g[�O�Jy�W��2���{Z��%ۿ� z 0�/_�1P��'��#R�!�� ��Z�%��,]R�_�76`4hr/�)3S��'5er�p��8@�Z@�j	�,A~�0�,}"�[o� ��`�B$� ����A�8A�Rh��I�.Bx�H<⧗/hu����j�==!Z\���M%tb���H�-�2��C"MY�h��/iv����ʃ�?'T\ɴ��٣�q���
���U,Aw��$&���@7.��4q:�	��S�w2`@j�}¤]�� ʇ��5���[Ԣ�2x�ɋ6/L�jm9�?F%�뗁Y�m���D�V����sdb�1}�ś^w�&��5�-}��З�/�.]3A�*� 镌SM�'��y��O�	\�Y�V"J?@h!bkX����I�/���m3�d[2��E���R#��D	%ߘi�5�J���犉ɲ������\^�CSa�% �M�'ٟ��E�U�4��D�?+S��q�%!Z��n:�/R�>�2�������F� \�X��i��1����]l����+EM�g̓wh�t0�'�%�b8����
'�
�H�FNGr�jrOS?�e�%��<I�烷PGZ����[�r�����^�VtE�E� �8��eJG�.��zbcS\�&5@��7:q��X�(��e64����Ңàd�S�J��¤l�C�
�e� Rv�'����AM�gt�18���eӖ�IE؞4(��n��)�࠘�.� Q�a�˺2� ��!�Z����'0U�d�_�g���'��b���To8=�d��H��҂ J �l�;�� 5"Oι�Am�l5�0�揊-,��c��+��y�F���O
��bO	5|��f�	��`��"OT��F���q O
��%V"O�dk��Am��!i@ Ѝ\S
�yP"O��d�ԓv�p�/Ȼd�t�rC"O@Q�ɍ�
�6�y�G>s[���R"O�J��"6�Y��.MF����"OV��v�Na�e�5g�k�F��!"O��$���6�ҩ�E��;O��4`e"O`I3�
F5����m)Y��I�3"O6 )���J��B�l�rL�٠"O���䅀#���J%O��Yj0"Ol�5/�̨��0Ǒ"tŪ�"O��b�hд'��ۗG1Nf,U�u"O�򷢝*J��� V�E'DLb���"O1��쁺?�>}qn%a���"O&\���ۮe��Ŋ$��#
j�i�`"O^%âN�,F�B1e�ݦ	�%c!"O��J��B�ad%+@�C�|��"O��#�'F�)����%�H� #��@c"Oa��lQ�N]zb�ʄ[�\dK "O���� ��@&��Q�剫`�r�;�"O�1a$���1��35Ò�~�,�Y6"OB�P`��"X)����[�E��zq"O��c@�; ܖ�����l���"O���K
�cV^-��f�&+(�"O�E��g0v�Ve�f
V�&t���	�.�k�O�i�b��A���ҳ4ܳ@Ø���ЙQ"9#�a�� 6���Ȧ2#�O��ӂ��C"�	�$�/&	���:,834b�Цar�%��"@a��E<uK~�Ya���U6���.]V�[�ėڦU�G���^V��S�O�ij�l9>S]�ڞ�)�w���i*�G�#k��S>�@H�"=?��TkCf)���&I\ʦmY��G��y��0�&�G��e �TkL4���:a^��7KJ�E��C��d������z����OU����,�$H:���_3��9G5O��ʠj�$#m"����4��{���|���C�u�ʵX�#@=7<��.��?1�Y��|�����&���3����f�Φ}����}W�=�p��?�.�)�x%��g�}P|�;`U}x�@2~�|��<'�N�=�O�HH۶dY����v�(1R�TJ6��Q��B�Qc�0�ǧ	�f,���X�NDإ�wNUk��)���0q*��<s��\�h�B�: *R�K>��P0Rf i�.� Q���C�N��I�<��I��uG�7<�%�qZ))���򁍑o���y��v�6%�7^?�5:��O�������FiK�h�&"���z��oݛ&B��m���T��_��'Q�J|���L�"IB�UMT5n���ó�M�@	 ���B���x#���w�@����-F�J狄�Ni����J$m�J��rD�<�7bl>��!�*Y�x��$-
	Z��HD�1(���0<y��"��`3G֨UҸ��`bS�jVZ$�`��tss�&dԮ�@D�6�nx�֌���)��CR�k>�H�?O���w*ڂ(=&q����"~"4A��$���ɚU;ĩ���ȾB��X�j�j��]�0|� ^��#�߱G��e�Hò�r���8s�sԑ�`���!�pk�F+3�x�J3&B���!A7fX�IfM�4bW�#�3�	�����/�i�l��PH�<�`C�	�\p��$��<5SlLbE�2�"C�	^&6�:��O"i�:,�E�B�F�
C�I�2A��@�.5m?֜C�\�3ϠC�	w�%� H�+|���x�A�4M�(C�I�r^=��J��<�|�#� ��DC�	X��R>H|����Ռo�C�	�8�q;4�'I�ts��3Z��C��&.0�0U��;[f��SK��s��B��^��`ӁJ�T�*���P!M��B�	�f-�����],�����"��OƜB䉍g����AN��)�V�����L�pB�I���� �T;2�h����3�hB�I"8	������Y#N}!2K�%@B�	9�ء0w-և.�����
~�B��E���r�f��xm��&�� ��B�IqX�2V�� �4���q��C䉈T� �������f�`�՛��C�	�K�rԱ���7�Vu����7VC��4<!�I����X��5f%�%,�TC�*,����N�� ]�$a�.�bN>C�#�h��9`��<B!bE��C�]�����A�s)���%��I��B��?:^y*"@�!5bT ��^\��B��
f]�H���9Q~���Q�SC�	${n��%�L)Jѡ�a��l�C�I����SU�<i�*YZ�MΝ9s�B�	C�p��� ��pk��(~P�C�Im�n���"�i�0��p C�ɔ��l�D��HI� G�Jn��B�I�L�I�� Q��)@��*H�B�	[W\e��-��D@��Cc).�B�	�?�HX��P�'���aaJ�k��B�I�¦�j�-_���@];n�B�	� �d�4�U��B(�0�ضtbB�� o:��SG*L�.���iWG�^B��),�}h�C<ye���'C>B�I4�����CÀE��q��l�>D�B�="�:9�u-ڥQ��q�d�]'eD�C�zɂ�ۣ�ۣ-���U,�*-BXB䉜&ł S�&I:y��kwHPc�pB�	;`��l0*��H�\@D,<}�6B�	4+U��0c�? �Ȑ��*?5B�ɊQrV� ���(����/[6��B�	�P�8�:�7RzCKi�rC�ɨ?��D�H6/2�ܺ"�U�D��C��'.��!�j�'��B,$|��C��CM@0XꟖS���QvMN�V!hB�I� ���N�gu���v��Y�rB�b��ZtG��=]�yS�Զ+h�C�I�*��Uk &A9	�<�#å����C�	��Y��,��^��c��N7�C�ɭ
�Y� M�t�`�KK?=�B�*Y��A�Ø�Jx&I���ʑ��B��$"𤱩֎��y/�C@T=w��B��6tx�n�i�(qӕ�S88QlC�	�y�^@����Y$=�U/�z�.C�"��h��e���P�~�C�I�+�8���O<i�XI���/\�B�Ɏw`�ī K�(��,X��<�vB�	�+�tE[�N1������jB��&\���W�#h�@$+�$ݘoB�)� ؝�2�ɹ/e�*e!���|�a�"O�|���rf�DAt���j'"O�Y�խ�A��r��*�截"O���gL�6�
$af�1�M""O�Y�F>,&��׊A+E�G"O�8;��ڬ`�*$�`)m�"O����m��<�@N1�fL!g"O�l�G�L6[ǦHʥ,�5��-��"O�,�`�9�v�!�U?W��ع"O�DRRkL.J|Э�"�i<2�"O*)y�lׯ_�"m��]t0#B"O�C�ꊋ,�.�#�R�x���"O�Swf٦_;���"Ǟ ,A*�*�"O���AF�����u�(~Ύ���"O���V-8��-��V���2"O���
�N�����*׈^�B=+6"Ob�!O�$Ѯm� C_�i�7"OuC��:E���"YK�9�"O�@P�͐�)��ዠ#�N��XP"O��҈����h�+C��08�"O���B@�B�R�� EG�#/��h�"O�����?�0ю�� @�j�"O��2Uo�ĺ|@�׬  zG"O)p�U�]`��G��m��=��"O�i;PcŎ/s8�iWfX�E8D"O��:�j�P�x���EJ�+1�a�1"OƩ�t�_Hx�����d�d8�"O.`"a$Z<;�RXP�H� 0�)�"O�ثr�Ł''�A3s�X�/��E"O@��gX8�,]%ԕ��"O�I7���4�:!�V��}�p$��"O�@t��#f�6�b�A�%�*���"O�uy�k�'%$��ɖ�
�`�vS�"O���F�F"I�&yⴊ	 J �r�"O�]�E�ź-���r��PB�(y�"Op}�eě� J��"C�?1@T�r"O�������ا"_�M��肕"O��/�RZ�+�l�0ep�q�"OF2�bN�w�I�*�+)g<�"O�!v"�k���{�NE45@���"Op92���E�,¢�˴HI��"O���Fv��X��;G�p0"Ox�FHC�nL褨�"\����b"O&)��"�-L'hG�4z>u�1"O<b !S�{D� �Q
�1�mJ�"O����I��<��4h�II5p��s"O����+d��iŹ2 Z|Cb"Oxm 3N�3�����!*G�-�q"O&��&���/#�dRt�E1�Q��"O{qф*ix  tM�"vb�"O`�B n@&r/����S!S>���a"On0B0MF:�<�B�ҟbM�1"O��!�C�?��5�%���HE"O�:���R2�z�MћTNY�"O�]Y����,w
!�pL�i���r"OIB��?��1t��>����#"ORP�E�ŋ5��S�*Қ�%�!"O\M���6�=r����]��"O�L17(�G��$1'	��XM�p"O���IA�#�!��|�X��C"Od��bΎus�P3��E`�Rф"O"�y�Hw��ao�(�&p�2"O`�0��dȪd����l�Z))V"O�-i�A�����_�B#�"O� �l����;�8!w�:��A�"O\jf��D'z%qC�Hy�~�B"O0�p��HA�ތ�#�ƉL���"OdȢ�"w�����6J'4���"O��yR��}u��Y�-ΰ8<�"Oҡ20��
�4홒c� 8�B"O��f��Tw0�Y6cO�`�P��"O��a䄙+B��%1f$\�P�h�"O�5k�Π�Hz���9�z���"O�
FĿj�z����	t��ܰ�"O���D�{C0��1��	��� "O�� �@H.iWjMy�h�Bs"O�I�$/��8��Yҕ�l	xƎG��yr���	�p�P��_�Z�#�(؟�yR�!vhTz�CēQՐ\;���y�n�* p���L�R�KA��yb�.7,�b#g
@K��8���yb���	J�it+��p��'n��y2h�"#��kW�U/|l�+�솆�y�Lt:e�5�z#��;E�1�y��ɴ8�������k԰i$�"�y
����ũWK��c�%Q���y2%K&t����膶-�T)� a��y��գlq�%j� .����b;�y�
�f���p��
�����ǎ��y���h8��E�H�&.�gh#�y��p;�h#�N�$��11���y�O�#������	o�N�1Ό��yr� �߄�P��M�9�P���%ܮ�y��i��ѣ�2~�z���,��y"�9*Y��paj.�I�`���y�A**��a��ؕ��s�D��y�C�0u��;�e� #�}��Q��y#߃o�lH+$�!|�V�{t�΀�y�LL����C�J#af�bdeO4�y2j@�dbL�%��YFF`����3�y� �5*y�ӭK*TMX��qG.�yR�׷u7�ȳA��9�2]�`�M��y"hO:^�d�k�O8ľ��P
?�y��63�l9$!O74#X�YЩ�6�y�n��~�(0;�K���P!	��y�d��<�T�����#�a6�y2�	&�@�� �{.�˦�ט�y����D���J�|Q~�9'�P��y2�>a�I�Ћ�? �(�%�^#�yB��l�k�ɋҡ�G���y��֕vӾY�0��"����'$&�yR��2d a���S6; `G*���y���~e���O�X������yR)�5)sԃ��@�"��#N�4�yr$_�t�"��v��>E��t��yr̓rԼtb�h�n&�|�SO���y�m+*Bݘ�)c��u�c.J��y��{-�a+`�\��x�-��yBLO�X��Dy���b�)8����yl� tbE- q��	�����y⣆($��8w!Urmʝ�'Bʀ�y2c)T�~  ��)t���R����y��ى�@]���L5r������y"��Q��=��+�'�����K��yR���r
�T"���%PT�c��Ǌ�y�={����Bg£;`�R".]��y�O��Ri�A�V芐C �Q�T/�yB�y�P9 f� ��)SA�ζ�y
� �|��cY �& �N�:G:�I"O�]yp�E�EV�(g��[�,��"OHp��K>0�n�SEM��b�>�k�"O�U��*@���52��тc�<�S�"O
L
� H��N��l�
<?:e
A"O���a�
?W�6�R3ˌ�3�6��"O�xkؘE+��SFϑY���s�)D�@�g�    �P   �
  �  K  �!  �(  )1  l7  �=  D  GJ  �Q  ZX  �^  �d  9k  |q  �w  ~  ��   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl���2<O�1"�'"d�p&$�#f�<b�FX �~���$P�0�ȡS5�ʸ?8V�媜.�u� G�~�dM�r�Th o,�DS�F�"`���d�%�]pv���ZFZ-���[!k��ם�y����џ��.��:e����@������h�^!I�
R�?���kư�{��-K��6mB.D4B�'e2�'��c�c��Sw
B�y�=z`/Z#,��'���c�Dx��	��*G@^�?����0҅�Y�R{�1�0�C#H�Z�Ƈ�����ן0�	ݟ�)r F����N�OX�I�?����6j䬃��-������Tu��\ϓ5��@�`F���^yɤ�Țn���'��+�$���{� ]*��?3��  ���;QfZ�� k�N����O����O����O����Oʧ�y���h1��0��V M�6d��?��i� 7���ᩪO �l�+���xش�$1��� ��!`�	��#׀�Aa��q��R�����������Q���<;�� �$�>2)�`3���Q��]��#�THb�o�-�M�e�i����O��I�J�D>H]I��'1T���������t��-��#�5p��H"V�(�(�J>�j��ɦ%��4]��V�X�~�n���fι�Qs�Ow��3�ߌG/~|XV;�MC�i��6m�?�X��D�h��at��(S��|�B����pATN65�����b@.�*�� H�6A�D�oZ�Mۅ�i5$O�'r��qբS���Am�l�h�R�#�]�p������G�(�P��!�F�m��6d�r�9�IZ+������L?@�*�/&N�y�	_��?��InѪղi����\,r�P��P���RK�#.���<����?��O{BU��)�?}ɲ�±}����y+�<e�L����a�Ti�S�'�x)Ң�)s�܂�L{�� �,���鑧ľ`�b��#���0<�ħ�ٟ`��=��Dj���ɰa�k�,��eǜ�R���'R��)q�X�0��B4��d)�1=��u�.�O=lZ�m�4x� ��Q �j�ΆO*�5�޴��$�	_�tn�ʭ��H��DB�t����²M�R�;��T�[�	 ���Xr"�'H�1Ɇ�'Y����(���	�f�B��DA�%!�0��3��j-D�K�@%Z����	ѳ�h����@�"�\)���Dx|�q���J���OX�l�5��O��?���Z�
�|un��ņ"P�S��'>R�'i�I�.||Sa��h6|��k!  ��=��` ��Oy":��`#��)n�6���▤���g�'\�e��d��Q�`�`D$�ڠ��DZ�JU� �;D�d9����!�0č;.�baA��9D�L� ��c@F�'�,QXv�3D����6j�x���	3,���R�3D�,r� G��Pr1���O5�H�4D�tPD�D�%F=��j�QJ�<���o8�S���JI���&-V&u��`U�$D�<��L�:}�4ų�J�#�8����"D��sC�\�p�f��$�|hI��>D� @�76�q$OɒP���Į;D��PL�mE$��A�Gp6`S��:<Ohrt%�Ǧa���4XR���d�ѣH�S���B�h�I2Qʊ$�ID��<�R��H�Ϧ�B��
_,#�L��\z�e��q�	�'BP��0<	VܛUl遰�]'&�rh���+�����ȏ\P��B �-)�2<��ɜ?G����O�hm����Z�Uǚ�¡��9l�|�`H�FyR�'��OQ>�F��XV�\�fϙmԱx�I>��Z}r���MsקD|l�P�n�e ��g�_�x�v�|B�θ
iӵ������P�F�up)P S�9zf��X�y"K
;yGFQӔ���]{�bS��y�,��|e��������A��˽�yr�{���xc�]�wn��J#j��y" Ώz�樃�K�9p:�Ec��U��yH^�!����j��?�Rj ̠	��V�|R�N�F�4�'��'���NH�#�d92��Q0�B�N�� (�#�&�M[4�iU�S�޷ �S9��'��p�mB�#��'�X�0m�T=i��`��@�q�h�,����O����VM?�@)��C� \����)uFPI����M��X�@�3��Ob>�d�O^�$��N�H*�bA�{^����
/¨��dYt�m���K��L�����#B���'�7����1&���?і'\lU��`�n0i�V���b��{���t�����'+R�'�B@l�A��ɟ�̧ج�uK.��� �'?����+��k�4�ѱKضQ#�x@	�B�� Pw/�&V�
��FZ��Lh��e�C��S���1q v��ϓ@��{��
�7U�̡Tc^;9Jn��Ɂßh�	՟��?	���T*?p�H���!V��lr&��~ !���,�m���S�	9�5�'&�$_��'�R6m�Ob˓ �u8��ih�S�kc��a��G�h�NI���JmQd��<Q���?���7%����$�!f� ౑`֏�y
� ����nW;2�����2w�ʴ8��'�\��	[�v�-�H2�y�䊋i�&��O�-DH����Ə�0<&iN���8�4�?Y��k��\*�;_YR�����5Tn�H��?9��?Q��䧵�'�� b�ǝT�V\�1��5�D��#j�,ȧ#n�j&+ p40�Qd®�?�.O��aGզI�I؟`�O�|��%�'W0�#�N?-DI!�T��R1�'��C^8h��p��)6&��	K��(S� *����cV,k��-��܊ �S	9f�24�����52��EW~��R�o~<�O���ɒ$P�8����a\�=���O��;��'#�7�Un�O��)��N�.��� �e��6#��	�'�2A* ��Ԭ��/�J��TЏ�D_G�OB"zs��#
�Vϕ���m�2�in��'�R�A&z��	��'"�'�"5�v��!��	W�m꣡���p��۷=ǲ���aU=zTX�771�1OX\�# ��)������	�4s�E�-w���3e�\��@���(751�1O �4+^�$ʌ�*�R�0@�л��'%��%�~��'�ў�2���s���3ǉ=U��+�^�<)�>��E�׬7$(ɰ�!�Sy�� ��|����$I&x�Ո�区
��(x�L>?2��!C]��$�OJ�$�OѬ��?����$DC7p�&qi�	�<Af8ԡEƣ�����'���H0e��z���x� �0!#}�g*�MS�8���d+��bA�'T�8�t'�~"�a�!i�<.NZ6Ĉ;�?9��'6��PG��+6fB<�P�%Xr��ߓ��'|��)�G��$�f�A !ðUo�T�K>���i��'��-!��}�N���O�ĻCiҜS��p�0Eˑ�X�	�d�O�drS��$�O��$Rg���<Y�w戍ӣ�=j�.�b"��G�y�
ÓX4��T&�C�̡{뎌�?�GkJ4=����/�*�c�m[V��YdG�Otum7��d�y1 X��#˕V)�p�LO�{ �	ޟ��G��i�1i�d��㝖RԘ��͟0�'ў�S�?)a/l�6��� 7;�X�5)�蟨�'�658��>I��?��'�Ȥ{�X��������(���3(?��{��?���.1���c�8E�<����%���ST���c�8qэ��v���c5]D�ɝ%vf}�PG�(P�B���
͒W�Eq�G��s�������?i���5Ez:)ٳ�,��"��&?Y�g�8+�4.�F�'�>a��K��{u�x:GgۺXk���q�&���O����O�˓�?�Ο��r5`�i`�S��l�Py�V�	?�M��i��' �h1qA��[C�9s�š�X�#6�h�,�D�O>�dV�$Φ�ieB�Ov���OF�d��, s�
ɨ�Zg��]肥IJ�"�Z���u2�p˕S�j̺N<9�ϐ�UC`��-�q,�9/�Q�`�I�U}�1�XS�b��08ʧ*��ԪflLҼ�»�8��$�/ }L��!�T�M+��i�2+ S���Y�$��2m%V8P&��y��J�Ψ'ȑ�Iß��'�r��>�Ǔ �
Ms�DΨO>�u2��sy¢n�@nf�	|��^���'�!�J���H�2G�ԥr���/E������ߟ��	矸�ɣ�u��'��?���Cd�̼g��x��V�y>�}�1�L�.f��$4�����fW�'���!AA��(O��۴�	�#�LA�	<�封�>ob��H �B�8���֔!NpY�eA���(OJt9�ל`�\�u��!��Ƀ�K`�X�Gz��5B�l�C.�ڝ(4	]*.B��i�-�4��ɏنXR�|�/pӰ�D�<i��^�x����\�iS=�0�[��@&*ܛs�����	�0�����|�'�؅p���s�H���X#Y��]0#��
b+��1U��h��i�
�||iE�'ʓ~+�<H��[�P�f�$3⤀$h�)}eT�dK���\�-��z�DI���8�J	�u�	��M�*�P;��!��$B���R�ۮ-��&�@��	�y�Ց��̺N�2��B������Y��8a\���!��sئ���Ol⟈ID�$§�y%�4df�qi���R-ĭ!�d5�y"ꗷּYpd��9J���0�F��y��!�H��r.��5q&��\��ȓ9r�(��$(	p�+"��wQ̤�ȓ0B��b�R�+%ȸ"���2v�l4��4F�@2Sc^1=���R$�,4�B��ɛL�"<E��灦HQX����ɬaDp:wk�}�<y�I�-�T�@��>�*<U�}�<'���M72���+�����.�n�<	��(���y��&i�&��#��<f"K"Α3b-SY�D��![|�<A�=L�\�����~�ʌ1�-DOyi�'�p>I�`Ba��%���ҌȀ���]r�<� nX��Z�#Ǻ�H���9��$A4"OڥKR%S�t4�A W�ڍe�<�q"OR4z$Iv:���ٝy��U�"O�B��݄HbXQү;T�ـE�'j�${�'�8�A1!�-R2�q �.a,8��'TX���^!lg>y!�c�.��di�'@�@a`�8(��Q�3NT1:�$A2�'�6�A�ڳpX��`F�X*:���
�'  ��k{��A֯�q�TA9
�'|
�[v���:
�!�N�;l�:� ���� =	Q?��5�V7X��`0�lظe��� `k!D����U3'�s��ќ{����P*>D����@	U�,����pl�ȃ@"D�ܙ��Z�IFT�S0�L�b3(t�"D��U%�w�4�A���Y.�# �"D�L��(�:��aId�#!RQ��L�O�mS��)�`b ����:�H���G��K}����'�*�8t�:��Ӷ��>7��h�'{���Ϗ�#�\��vC��*s�\��'�$�Y7�8v�>ђF���<k�'���� 	�,q�����(8F�@�'����/��%՘����˥?�+.Oh��A�'R V*ÙqN���"���(�
�'��=s��*R|��$��r=LE�	�'%�i�� @�ڙ���9t���	�'&u��CD(-�
hz3LU�e���	�'�0ݣ$��'xsZ�m#.��M���'8�@�'G�rr.�/���BkJ�aۖ|z�'%¡��bƛeh<0�(S�Kǜ0x�'���B��F({9h��`� wņX�'R"s�*�(�V}A�G�)9�註�'�.�`�H�#4�I"�3|T��'Lغ�b�D�����q���k��DF�lIQ?5�(�Rx��Ë�+X��c�4D����I&�zux�l�.*%r���E.D�8[fG%�, B�z���Q�,D�(Q���VT�4A�Q��mrA�8D���عt �S&)�q^�Y��2D�d
��5���"ͰI�<���O�Ă��)�'P:�a�����hV��gOS&/��@�'`���H�� H�E��'Lh��'E"<� ����x�FD���l<k�'#RX���ւ��XZ���r�^Es�'�8�4%O#En<t���f<��k�'�p�����cq�"��Ԇ	���K,Or8���'_�=+g�CJ��l{��Ȁ{�f8�'Z���S�J�1� B��r��p��'�P����3��A�&�N �ܐ
�'vY2�bN�"T�ͺ�jA}���
�'c~��a"";(t��!]��Y�"s�t�#�5�c�O�/�,@��Ш:�v��ȓji�T95��WK��p�*_�����<�u0�*Q.�����ND�-�>��ȓ`-,,B�JVU�Qx�b��K�⹄ȓxpz��7/�&.LL(��@7����2�`݂�B��v=���/��S�L�E{"hӘ������g�B3#�ꥑG�		lʀ�"O^{��W�#-:ղ�ȐF�b�Z%"O��S�,ݰ>^�ݨ��!Cx�ē�"O�$HB��d���RG�h`��"O��sV#,4����PL�z��Y6"O�q����j~��Ɇ��ifUC3�'S�\Q������)��L"0u 0�c^!`�D��ȓ#���L9f�ֈ{�"�'SH-��S�? .��.�>Ax�N/A�쪆"O�Z��ڏyH�fT?j �W"O��A��5]��X����,b��[#"O��X���=�<8����lha٧_��	O1�ON���o�.J]�����|�0��"O����#�!G��)&�F7#�B�P�"O�E�AV
A�	'�˸pF�PR"OZ�C�O9gZݭ ���A�^=�y��>%��$`�&D/�Љ@�ɞ��>q�ha?	d�s�J0!'ß~j Xs�Sb�<�1�S%?�Bi���
B4�5�e�]�<ٕ�l��DZte^7��`�"&QX�<������`�׫@�c�`�Kl�R�<�A�7YA��cD	�.V2�˵.�Q�<Y5`ƾ{�`��
9 6q6�O�'���c�����}�J���&�y��p�����!�$g�
��&#�b������3I�!���_� 	
4�V���*a�<�!��� fU^̙P�$,y�9bAU�!�HI��\�f��
[r4��u� t�!��5#-4A�-��Krb�)��!!�"�̫�O?��%]�R�X̀ǄK3L�t`�*�v�<iSi�V���F@^�
�H����]�<��NKH�)�q(�'.��q�l�c�<��ɔ4t
A��eL�Y�$��d�<��h�}��QI'�Ra`3b�\�<I*Au���:e�J�G
I�B�YyBK��p>�3�)'�F�B�r��%X7'�W�<	���T�:B�Y*d'n��1�R�<1��F����c�=��̂%n�P�<A��,(��BR�֕V�zLk���J�<�0���GށC5&ҝx���:���Ix�d�p`������C��V�TK
7 �Bŀ��5D�T��?lsbɹ�j�U$���4D�lac��D�^�c�OKЭ+T5D�� �I_�:EKv�
3����J.D�$锊Z*��脥Y�\4�9�0D�@s�cD\%��Oݰ~)>)hb�-ړI/�D�䧏�� ��!�vUl�G��y�[�3X�e��
i� ى��6�yb'I"���1�)]SX �1	���y�	�<'�8��l�m;*-Pq��y2(��a��,k��J%dy\1�-�,�y"��%�����&�1`S"��?�� a����:k�j�h�4`խ[[u���d=D��i'���8H�}�G��M��8@�<D�`����K�V�*V�siYW�=D��S0c���Ġ6���G���gc>D�٣�ͺp� �`1FQ:0�r	�A�9D�Xv�ţ�p�KkS���Љ���<92��S8����m�:��f��", bhJ�+T�l�d�4R:���B��H��U6"O����>7p���b��xy�p"OL����;(�H]Z�ؿi�C�"ON��f�/i\�`f���Tc�,� �'�P�H�'�Td��&�6#�� e�C*ɲ(`�'�䜀w����L�fE\�1by�ȓK=x%���\&Zkx�ë���݇ȓ",ZdA�f\V��be��F�ȓ<4�L^�0!D����t�ȓ�.(s�U1I~���"��E?R�F{�DY���f|�A�Rz��JN �Z�0�"O�;�J��3O�h)��օ��0"O��%b��K��9C�X8�
�ID"O� N��H��o�� �3�v��"O��	&U&z��/ˠ=͆�"7"O�}�b%�
<� �Ҡ�-Q��j��'�|U;���~��4�Dȥo�<���DLHN�ȓ�rEB�
��8H�H��2,f}�ȓ4�@͉QH��k�.| ���23��a�ȓ:��d��
�~�]X��9F]0���9S"4�`(*8��)HP��9]�
ć�-���K�_I�f�Q6�ŵdu�ٗ'���`�'�t1j��8���v��ҩ�ȓ
�pc7�� A�bi�&�M*1ZH��J�X@��ȤV����j�]��1�ȓ *j@�wlD �*���iW0OT�i��P�"�-��{��`}R�gPx���v����BցN�ՙ$"]�|a���o%D���P̗150dY H!q鮄��"D� �J�=Z���(�y�rx�.D��P��؎B����Y�z�z!:��0D�|JGI�3�� )]Z"H�H�N3D� �uȔ����˙�?]����.��e/�''�ԝ(6!��{|�ҠSw����UQ�L;D��r`���^t��ȓ�8Y�!��7�@B�
�F�N��ȓY��(��@Ah�"���Ů��'���*� ��P�P�&NT*	a����Q" <�!��2"��Y0c	C�J��=�	�gM�#<E��䇘)c�� �Q�6$x�3�`��B"Ol!�0b �{>�׀\G	�@�D"O
U����Rha���D�f�`��q"Od����5��`Cf�	1M����"O�m��(_|��!�R #d��TQWO��F싱;�r@���۝�����OF�'��	��'�r̋@)FԦ�@B��?��S�]ƴ����1{��Zc�P f�P�Ƀr#�4��ퟄ�I�u�\�Q��ʈ[;���V˒E�'(������H�L��h��G[4X���E|@��$q�/�w{(����KB`��3Z�l����-b� u�"�f�'��I����|�s!�<�r��DC�0U�pR&�hyr�'��Rĩ����z�ƺe�JTq�a剬+�dH�W�D?1�Nc�ȗQ[f� �օ�x�����Wbh�թP�e�v�׭~�<��Z��t�R˒7b�V ℊK�< ��6����Gh�m�QC&ZOrP��W(�uhY�,�v��L V� B�	M�A��K_�'�\%蒡
w��B�I�g�\1`�1j��dx��1f� ȁ��{��~"b	� E�u�ͣ@Х
P����y�A
%���+W��8�U�"ߊ�y�B**��x��J�';{�-�����y�o[�@H�@yA��J��P���y�J$0��C���,J��� s�R��y"��ce� Ӯ�k=��P���?��)�M���q�G&U�n��({x>A@@;D�y1�8p�b�W*�30��+��-D�����=yV$y��e83�DaSD�5D�C�H�b�8S�Ϳ*�>-�n5D�9�ǀE�4����<��5��.|O2�2��>AB���0u;�g0d�~D����d�<aD�8&2��5i�>b,hأ c�<	�ǓjY6p��(;D~�`����J�<�r��ih8���J71����R�SC�<)T�LiH�qڅ`˴g��D:bH@�<ɔc\&�M�$O7YȊ�#� ��'{�i���~��F�E+2��6N]�1� |i@�h�<�5AמN �0uabZD��	�d�<!���u�F0+�V�_%	�Ea�<� p9����1�0� EA�*[@��
�"O�������B'g~�	�'��}ztiĠc�4��H��o�&��ƤX�'"�>�	 �@8����=
$P�fBB�	�u��{U��[���vi��rrB�I���d� �NL�l-�$��c��C�6_��t��@�H�F-��\��C��k��q8�g�2;p	 d�)1�C�I�r?`�H��}��Dj�.�+���1k��~�ɥz	�т�g�e�� ���yB�ݠ_ֽ��j�i�f�PI�	�y�O�I�@�HP�*+�ԩ�G)�y2Q&sS��㎝%q�*� �-�yb�O��<���j�ع��c˘��O�L�֋�Φy�Iǟ��'00�JI��'��	k���4���yӐd2���O��D�OJ��B��Oxc�擫s����O=HG>��%��v.>">I�(�F�Ow6�3����,��1�'G!aЈXQ��n� �I���Ox��i�iO+-a�lp�[�RN Ly�'������5G�9����PJ���k��I7 ��oيA=�i���=EN���?�����|�����YZ@7�ǆ4��9MZdџ0p���<`����2S�2,��K�BF�Ot	��x������O7�0�4��RI�U�G�ڼO�����O��K��\�O�s�̨!d�&v/:� "�H���U��$T��'��'p޽K�\YI| f�=Y`����0 1��ab�'e���S��y���$�F�)S�ìMI�p#'H�\d�%�M�ԫI��*�F3}rD�~��-T*~�V�;���^��U���K���:}�k֗��RM��h�	i�H�dn�Rɺ ��Ox��F�>ѥ�>q��RF�DS��!Sq�V��(l����E���@�<��RQ�D�\�OJ���e�
-N��]��b��䴟D�u-}*���B�]�	,9��x1"57�XE@ࣃ;#A��C��Hy2�����'$DD��,�MM"yt��;M��zV��?�4D��p25dP��|'?�;}����I�lD��� ��iC\�c8��d����?��m�r��@ӷ.�N�X$��\�<1Aɜ
{b�X�p�݀0�<�Z�K�����Iџ�'/��'A�	f�\c����$��.9��,q�;c6���4�?�-O@��F�4�'F���$�\�Y+,�2������PQP&��ē�?q��OH�MJ�5Q�A�G_n���B���ȓ-�x<�B�W1�0�A�b
�}�(�ȓ6#���A�M��})BM>Gz���ȓ^��[!H�K��9%�V0v"�M��c�Ddq���6r���_+?3����SF D�e�K	�����H&>lpt�ȓh����B���J�VE��B-lf���X(����r�|\#�+ا-�1��L����h�n(�)ǝ�|�1�ȓ%Դ!�⎔/"��֍I�/�|Fx2"4�S���~E�4'�3rGpDp&+إ�y"�W{���d��m�����9��'�v5�2��]�)C@��]�=�7�U�'���:a�G�x�[��.o���a��&f�EŻ���/�%��!!�kȨL���4[��#���
�Z���/&<�)�@ޢ	�����o]9b��#Cќx�]z�K	<5���0A� F�`��R�'�l8�0�З2,QjشF�܌J�C�+k��}��`Hx9��hT�'_"��zmLT��E2�T>��O*8X�������xZ�\Qi��J<�v�!.�,8��	���c�Uxx�$J"� �<��i9QH]*@. ��KQ�F7X�'8`��b��ot�(��"�>�$��F�	�b�b)��{|T��IzX�����	^��;��.X��!,%OޅFy��4V�����R�!!L��|Ia��O��ą:$�Q&OZ�X	�x��#Q��G�j�0(�r��]6��(j���y��+g6.�Z��J_D��G�yB.�  ���9D$�
SV-1!惝�y�ȃ�z9�	T��:0ژk0�%�yb�D;)i��yAT�"��t0��	��y�K��>~x�(d������x�쁫�y
� �(iw��B�b���A.Gn�l`�"O�p�dS���U�U/ĵnsN�c�"O(0x��ׯc1�p"���p�Lx'"O�1Eγ!)��Q�L�.�j-��"Oz���O/ZR٤��+:��)�"O�}��EK�1�����A�W�bp�S"Or�)��1�9�/
	S��`�*O���G�	�徐��D�dnd�'1�Q!7��.W�Ь�11S�%��'��3�lŊs�J��b��(�h��'B��bdX%~� 'Ă�:�!�'`(��C�y�"튕&�8�Ł�'y��� ��l¼R����~�;
�'W��: JJ�4	���*4�tJ�'�0Tx�ڢaZ�� �dQ*�Hp��'���Q�T�{�2�3�j��'@���A�3LnX Y�뇉d����'y��Q�F:n����DL�o�B�'���ņ���-�c������'��X ao�ʵ�Á]�ft���'�$IC��ݗ[���§o�]�� 
�'cj��S�K`q2�\;(�B�'OX);R�̂U� )2���>QO���
�'�lu�}JM����S�1
�'|�yoś���q��Lk��	�'�����'��?�!cA�]�?��A�	�'\���"c[�̪І�4?v ܹ�'W��q�%N-
>�xs�5��a�'2y���:�P��h�0`ʰ��'�-*3h/;��i�s�7u�6��'�\��v/�!`���AU�5~�y�'�.0c�ĺT��rMG,�����'�&�'a���ڡ[��^�%��y�-U.o���E�)f���Ĕ�yb�Y�89��.�� I0d�ҽ�y�h�>y���ÃV^A� ү�y���n��`*BA��za�`	M�y�@T9eAjM!����x�ઋ1�yRO&"W��R��˭4PS��'�yb�߳ckа�V��,~<t��U���y���E���8� �q��ze&�!�y�mI.�ޡ{��h����I[�ye�\L�d`K����5�yrl�" ����*ՁQ�:0���V�y��B=9xd@�mE�G��-��A��yI0na2���F	*p�vB	�yB��2'M��!&�V1Q�ʩh�����y��LN����'ʙ+`ڍ�R'U9�yb�S�{�RP�3����z�ZB�M�y�B�2[��Ht�������aH��y���4O"�%��׋8��I8a��y��r*t��ǫ2�,��ԅ�y�aI�O�8H�.ɶ"��]��W!�yrF]"g��Ź�j��F�*@�آ�y�H֔s���3ɛ+1����O��y���O[��X�jI��@�qN��y���F����/�Z���H� �yr%��V�Bi1�]��lp�A��<�y¦A�^�z�pdi�/�D:����y��)Gzvʰj��[D�� �,�y����ԸAJ	[Q��������y��RPޥ��7S��L�`�L<�y뀖xܠ-��j�35�b)���\��y��`^�@���(}.婴aT��y
� ޝ �`��;������M�vES"O�!�Qƹ)�X�k���{
(P0�"O�h��hD:N���H���2gY\���"O؁���?\h|y'�)XL�%�*OJ�Z�I�q��J���i%�	�'VF�y2h� ȵCW��Y��'[�Ɉ�C#o!L1Ў-{m�8�'$�	�L�J�����vx�8�	�'�z�z D'�}u+V"͐Ĳ�'HB�EI�<q�%9Ta�,��2�'&����l��,i�`
�n��'q�eA��*�asej��T)hu��'�t$"#��6dj�B݌w����'G����54ۧ�@	{sh���'7^:�ƍ	��<	f훉L�pc�',���HJ�v��8�e�H}�̄b�'DD�Qd�(R��5c�+�,�#�'��IѰi�:|�Ɛ���3u�M��'
^t;�Z�5H��d�_;Z��{�'��̰#EĂq�Np�$D@*U�!!�'x��j��}G�3D��{��A�'	�,��E�d�`S���*E���'|X|�0Y<�+��>rƢ�i�'v�  �ljy4dU�p�b��'��xu�[2V���@�?oZ�'4d@2�c����P���'c`�
�'��1!��6�
�`�RI��Dq
�'uj-�5j� ;5��c h׵H�b h
�'�vx��m��c��|�wcO<^�Z
�'":��o��.q�u����;4��'v*��%�	I>�%���3��u��'����`ӟInj��L;W����'��p�!��t�<A��Ʈ8���'�1Q�%��T��C-e����'��ice�(^����/�7bn��	�'%� 9R"6D���@f�J� ���'P�P�3/ˬ
�2��R1>���'�8(ɤ�''��c��Y:4�����'uxX��<j�0�Aܓ2i�t*�'�J��S��2Xi��
�L�&A2ı�'��KW�Ʌ9��YF� ��i�',�}a�/+b�F�AQ��C�l̡�'�P;��E"&���AK�4+����'� �B���DE�1aa�H21Ne8�'���)b��' ��݋0���' N)��'68����"�B��
�%SĹ �'���OĴ~|��A�'L�:�'���w(P�t���j��G'(�z�'ԨKD$�֤1b ��0t��'AP�aң�=fX��W�7	�����'	�u�p�
�Hj�� ?$� �'��ҫ�kj�9�K>s�D�@
�'�x%Kq�15�� ��eZl2
�'����ea=�l���
�'݊�S��V!dPv�B�ִ}>u��+^�9��*�g��\�2�ѻ]�L��ȓ6�vP"'%ڙPs�Hю;D-��'yʽ('
 S�<pc4U}���ȓx|(h�5] ��wl2I<��ȓ  �c��v����O�B�2l�ȓE��,m�$@B�ª	JBm��8D�0B��Ӈ,�P�1�,�f�)v()D��"ǫA�!t�٨�MżKW���%D�@���)����+d���RJ#D�� �ؙ��E����塆&l��P�u"O�������$(�!��[n !�a"ODE�+2kf�� �V�m~�I�0"O ��n�T;�u��¾Co��s"OT�k�F y��� �F�J[J��"O�+P��
������i.h@�q"O��ac�:~JtP#�Is'2��"O��0jD�H�8�@�o�� #F9��"OH`�"�:"50s��.D(\�"O�)[b�:160k��U�-�� E"O�a��D��Yӕ(
����D"O����Ӥ�Ј���R�~T�5"O����$o��m�Q/ћl�&�jc"Ol9�î��H��C�#G��82�"O"h)�����*oU�O5(�T"O��E��4(B��@��C%֕��"O>8{���<tXP��Q-�`"O,MZ��1�lMB�L�T&��o�<��$S�
fr��W��y���8m�<I���/����#	,#������R�<ID���*�8���"̪2�>9��De�<�գH*L��i��w��m 0�x�<i�N�^�sk_4�`h0R��^�<�aA�� _�QQ�ɧT�<틡ǉu�<y�͚�l�DI�צ<5�}��_p�<��V��XZ$�g�~��F�LC�<a�)K�d+��_�9N���@!�e�<I6�8S�2Т�	T�S�6)p��Y�<iMN�&>j����,�@��fF�a�<��B�a^�EsP+H3tA��;,Qe�<���;Y���k �m��TC��[�<A��.��dHB(8{Ȅ��I�o�<A���WH�h�ɢ_�xi!���m�<q��
vTe��N~R�T��j�<��C�e�A7e��^F�@%�M�<�qn�V�zP�7�
�;�*s�B�I�<��@U���- c��``i��_�<�&�/͖m�FJ�ɺ�6]�<)��ݩmݮ��$�61D�\Y1ZV�<Q��S)f�X%&#۴7�F<��fDj�<��h��h����b��G�b49v�i�<a�U�:�(�ɅAW/`��ŉ�a�<�&I���d;�Q �0�"LI�<�ĕ9v�\P:�B�f�<�G�F�<q��Q!�Z ����j�0�q!NB�<�&Ct�����eO���	�|�<�ᕤWňq�X?�R�E�^y�<wm����sH˷%V5�vf�I�<a��Ps� ]���IK��w�
M�<a0c�C�P%����V9脀 J�<I���l�N�ao� Zs 5��N�<���R`=�1�t�_�f����r�M�<��	C�n�VE�.��7l���_B�<��kO&I���c  K[��S�d�<	��ڣЬ��2@R��,��V �^�<���@#�f� ��+���:�[�<!���'H���A���|�D("&#�T�<!��]�0R$0	����;"�Uz��Q�<鳧կN�>� ���:���&d�I�<9�H��L�������f�`D��'D�<��=K+ ���[��y�;T���ӤU(Wk�P����]S��?D��@�����k �`��Ah	d�x,�h���	���nx�|Z@�32|�Y�.V�VR4j֩5D�� � �AO��DT�SoF7łS"O~@�w
���	��W�p�Y�T"O�,�𯆛]F�}�f �^gX�Y"Ov�Su��dhց�-͵Z��R%"O�]*�A$��L�LQ(>�ΐ9 "O8\�4�-���hӂ��d&�rD"O>�s�)04�sA��4j�D"OF�iF��Nh20�E��#Iz%ʤ"O���!��4�|	ZC �˒�B�"OH��'�^dJ("�կU8Vr�"O�LI�� alF=�g�-;�p��"OH�A�c&-(ue�f����"O�в"^��p$��U!�"O����ˌ�E��e�T�?��Y%"O����قPD�0G�I6{��]��"O� bC��	CDH�+���p���"Ozi	�:8j�aq��0?4�c#"O���6�V�
ܢԤ+M*l��"O��0�˞. �����x�X��c"O��1da�&�f�sS`�� V�*�"Ol��5B�d�"Y��G#q
���"O�x�T'=`� �{�Q�
O�`hP"O� bF-rH�$Hٴ|K�=��"O�y��
��B �X�&���R"O�`�S������ؔ��	? �e�E"ONǇ͎pa�j��(o_|��"OR[�D�(�>�"�A�UD�X@"O��*'j\;]��E�<����"O�}�W�SXn2�+��J�~�t��"O�4�n�F�]2�+��(t\�"Odi�
 E���"�!Z��b�"O���P�_���B�ML(F$�:A"OX8���hԮ([F.T�^`&�RT"O|`�'�2R��BCֺNX���"O��D�ںX R}ӷC�yW�Y�c"O�Ⴐb�[3�q��/J��k"Op�7�*��XIb+֠�>�R"Oځ0��u�����k��%/�d� "O~�(��
l�1T�@�Ay���"O0a��Z'u:�	a�>Kw|�I6"Oz��BáwΝ��]�R4l�"O(��gڃ?!���7�< �P�Q$"O ���!u(PD��)�b"1"O���׈6�,a�H��J*	��"O�	�F6�Qɧo��\�H"Ot	"`��#����n̈́�`�3"O��rM�y�y��j���9F"OZ`��J6^H�#I�͈M��"Oh05��L�E��-޴?[@\z�"OzM�K,E�& �0o��k�6p�C"O�A�Qj��%��!Ju��=q��0YR"Oj%b��Q	� ��e�!O���"O�`-W���lR�|�f��C!��Y�	���#�OՓ���'�[ +u!��I.5[f|�`�S�������"bl!��My-��O��Z��QQ*C�>l!�N,
��a[���'l-;�]F8!�DCl��Y&(W�ʉ#��#Nd&��ȓb����&,]�)8dI����(\��1�$@�f	U��bӣ��>��Ѕ�4�� 	�c�M*���&42���S���y�L�b�j��N[,�lх�#A�5:��*��鈷�!*F4�ȓhRtM�5錫4屮����@_���S�? ��;��Y��}B#Ҥ"�ui5"O@R��J�s��D��I�/�b"O����`Y��  I.A v���"O�:�����Pb�'̳t���d"O�`E�/�� !G	`|���a"O*��P�F9�v�""F�-=c�P�%"O��Z��5!d�����~��"O��`��%��#1
�<t`��"O �۵�����G�� (0"O �B"�ٶ>߶Q��\�Vޘ��"O(�����*a!�J[{�m �"Oj��&&K r'Լ�s#Ǟ>	�W�f�<a�*~���p����¡�dO{�<)B���8��}ʘ�tB��0[B�<ɳ��Quh�qW$ل]p��Gn
[�<)�)�%${T�u'�:Y$Ѓ��T�<��(��FtA��L0{$V��$�HV�<)dD�*W0�����t�����(�T�<�0��L��:��2I~�]�W�	R�<cJ�pQ�b�GT�x�ʀom�<	�ٟ
��-(F��w��6��R�<q�K��,6��IF�hj�J�P�<��BQ�4� $Y����W�R��ōj�<��.B� �!8%@Z�R:�m���De�<Y1	ȧ*�h��
z�4��<I�! ";�(��e���p�`�x�<Y���N\��K�蘋nSݑS�C@�<�����1��$�A�W�/����$�F^�<�u�M4.�li��ǰ0�k�W�<�)v��f^�/�.y��_~��(��{�u�E��lT�{� L�v]��M0������=�8�r���E����f�<):2@���l-2��K;T�v�����M؋,�����
��=��"O�͂%X\�p��@�4$���"O�q��� ����'���`��"Od!��F�+B^�`%M�L
ٰ�'���@	M�9s��k6H)�8�p�șD��B�YZ͐���c �����0��">�%cR�Yr��a����k �=�W�(�4�;�.��yRb���؆b(l�d�%I:6�U�2�ȦZ�(m�\�"~n�-X:�I8V�M:Nu��h��� CtRC�Ɂ���M��]�Tz֢
P�B�(��V=P��	Ǔi.V��G�/Ll�1f���j��	�qd}2S��W�R<CC`˵'`�4#�-z'
t�bm�t��]���(�dOФGt^��s��	=<v"<9��׮m�2)0����	��I~��.��\��A�(J�N���NL�<I5$E�i�4lC�BI�6b���(���R��R@�$���8d+֘+�	G��'�r h�n�-~Ɉ���F��z\�	�'�r|�Pk�s:���fFWv�ѥ!׷I5��2�+ڪ(��cpm�:�F}�!�9+�]HtnL=Sb&8£��=��=�cB�$�4��#+S�3ִ�c#د��J��[AD(�G[�|������F=X�	�.��e�A,
��Y�>q�8�r�hd r�0*����6+�mq�a<��E�ҏ`"xC�^Ƹ����]� jj�s+P�	4>�a�:Z��d��F�y7�D�3�'�~RiX$gMVzv�	�D<�q/��y�HO/[�M���>-@)d��5	�U�ɴ+^.��
԰�(Y�]w�Q�Y�a��8@Rm� ��DcH�b#4lO����`	#�l���Ӫa㖏�	^��Tj�'�-[%��مh .yx��$..�&���N�(3�	8 �Y�}�Oi�cO�T8�A� ��Y#�� �0��K$_#@ۀ�_�"�1��A.�y(�����rQmɱ
�H��}Ҩd �WU�����d:`Ћ��O�d�Þ���p�E�L#b�$��Q"O���˂o)�}��d�5g����Y�> ���5e�8�L�F}
� �$pG �?.�a+���qo6�Q!�'�DK��D�����H����O�d� �#�DDI���Qj�6c:�|��"܇^�m�/�Y%�l1��
��|&?��$`��k9X�L� ���)D��0���G}�! �hS�UR�ṟ<��)@�@E�N<E�Su$�Z�p_�y���x�<)�R,-�R8� &ʔxq��A��X�D\�iq�Y��o8�pyԋЉd4+��ҍ��-�.�O�t��ۃ���_#/$9WɌ�M�b�� 4�$���'oF�՛ՋK(r>��r�9�8x1��	��d�v�ZN��!
َW-!��;���"��ҧS2�!sȈ�K�!�W���Ii��O�S{2d�g(I>%!�Ğ(��u��G�.urqc�܍m�!򤗹d����ھcj\iRa읚Q�!�ʓiu(D�7nU7~i�4:����!�$A$.#\��ǝ>[����^�!�D	�<�D�{��.@"�u(́h[!��(I����`�d��5Iկ�3!�DF�b�=���m�\��� �D!�$����<�b`�n���p
�9!�Ċi�*��JK	�ycqM�R�!�	�!�Tq���+�*��d��,!�ϟ�mDZC��~�:�����t�!���&ˆ!UA��Xl#t�	��!���������s���,	.!��K��╅�5OfB��a�F[!�$G!L�x�1U�Q{Sĝ0cɁ=�!�d��_A���V/�
��MB��88~!��8�x]������ �T�+{!�$
&<]T��>Mb��2�*ߋCb!�BFc`��^�aCz츐꛰}c!�D��4��q��EK�+�����*\)w�!��	�4�:Wm��T�"��6@�(�!�dע�t���M�_x�x���j�!�$E�n��,0�KYm�6	�ȑX�!�dm�ޭ��nU�l�t���+J�!� }�`ݨ��ߺ,3��@'��2u�!�D֎>@DX�hֳ3%^��,>m�!�]�&���Y��� ���,Ǔ{�!��=��@]4h�$8p�F)5�!��|n ��cE�����a�^��P�ȓ(�ΩPw�H�7�V��5��&#A���ȓC�(%BP���" "|T��J�-���V�s��+wgޗ:|�=��f<�#挎(GVI���K�\�q��2��X��8K��AD�&4g�Ȅ�:)\�Rs��fo|p����%/T�ȓx�@����84�p	$�/����l!p����Y�p�"�N�\����ȓ}�Jq��eN�YX�-�wI�4uC  �ȓQ�&!�u�Zx��UΔ�
KT5��K&�Qt.F/eS��B�M�9I�I��^mn�xw��<=4&A��4q�e�ȓW�X�B�;6)~��AH�2��0�ȓ\m�Uc���9�pr�̇p��i�ȓe?���T�Ҋy�6<�#��2C��Մ�r��H�\�)oXLR�U�LG������u����I�]��M��!/��ȓb�����Hs쒔"E�@�%D�dZ���0j�x����	`N���/$D� �mD�x�`����P�-�`���D D�B�'̽�����D$��if�!D���ݓ]�i�����g.<��.D�� ^E��"-"�j��$� �"O
p*�)>w��r��rP-�"O��Pc���:#�T+��%٦�F��٩1&@��pAX�i"<O.,��/��d�e��+ �氱�"O):���8\��q
��=D��53"O��z�+��D�	��,B�"O>�[N�����(ǒ����"OX�SfB;X���uE-mGL� E"O���"MK�L?r)00n:G�0�"O��p�ڃZLh�凙�ez���"OB\	C(I:b�X8�f�'bx�9@�"O�-Jv��2���뒃ؼV��1��"O���ŵ`�F(�bмhh] 4"O��k�h͘�؂�S xO�l��"OV����%^�(�Pm�M����"OX�"(Ԗ>���C��2$մ�	a*OX|
�AD%Y
S��Q�f&V��'�V���H�6��@���X��I�'$�����(M5�tR�G��$M4!h�'��Y�jɌa(i���?
�V��'�dXLB/��`� �ؽ���;�'&���@U9x����^M80k�'9���樔a	
vJ��x�n5�
�'�耢�&�;����UNZc$X�	�'{�D2�zyYO��+�`�	�'��l�h�!�D@(7ɲ� ���'�4Q��O�6�.�!N�˲ 8�',�ܣr�����3��J6A��R�'��DO��rIH��Mu��E��'�й��4�x�{Q�X#����'�|����_/z��ɲ��	�P��'z���b]<��i�ӒH�(��'3j�Z'��T��d��KR;#~QQ�'�TY���Q ��efM
/.����'V2D8�K��<��(�d/ݗ!�~L3�'�aC�)m��{�늀q�`���'ޤ`1�K�4���V�׸_t0�H�'�$�I�K	)Bb��V[�"1��c�' &Ya4WkuP����<��
�'nT��щ�YF2�q�H�9�p��
�'�]�uʛ+c����Γ��D\�
�'�&�23	��w[
a�@B�f�P��
�'����m���Q�+W�dȉ	�'lVe��F�80H�ɧM�x�")K
�'Ў���C�7�.!F�ЉB�J�S
�'��D��ߦ�Z��Y*4���
�'�B���D;�%p5��4����	�'�Q9��M�:e�5"%�]�`��x
�'¢	�c*�0Ox��c�i�p�X	�'-�����e�'M��	w<��'�H��"bܼpÚ�R� R�	����'���D��2s8Y��j�}F�80�'�b��)bબa�݂^���
�'w%�ph9*�T��K�XÀ}Y�'O��ET2)e�)�+@8&����'/j@��	HT�� �㋘t�����'�p�T�Ϸ3H���`�\7vdA	�'�\��ᜆmB���P�u|4$
�'���&N�>��!���U�ql�y��'�d����@�Q�	�d���'��P���=�>�״�3a���y���n�z��!b��j�T�����y�*�J�\�3CI^�s� HAՉ���y��V�q�|h�ƀ�q��H��hM��y
� �P#�f۩Yqֱ10�؄�d)�"OHL3p��K�Hk���zz�,�"O�ɓ��Kj�r}�v/�,n�<�D"O8����+o���W.D�MVT�`"OjE���R'j��:nM�
dD� c"OTҤ)�	�̅B�&�5cڥY"O`��&���:��rfМXj �H$"OH�pD�$Kv�gK'[ 8aF"OT8���DS9���_uE��q "Oh0�� �b��WDT�N%B�("Ot�蟛+/ܨBƃ��a��"O��B�l޴��D�w��1K��0�w"O�hG��M�pCg���1"O��;���To����I��Phv"OZdH�,^���Q��ɰ�Q"Oba�vF�Nz>,HG@�3�.�y�"OF5���Y�?��q!ϋS*�A"O~9��+�V\E�>#n��0"O.e���4�����e�+��س�"Ǫ�we;�NA1���.��(d"O��HCDTW���Ԏ	*��Q�"O��*fDǐI����҉D�MjA"Oh���i	�n�sQ����J"O�`$��<-:�hx�,�����V"O�!b�\/�,,Ac̍ ���"O6P�A�/4����$_R]�2"O6dr���x�`8�7�ĝn�:I�6"Oĉ#�ł)�1���F
aں�@�"O�)���H�L)QC���F8�"O<����4s�< �q�Ť���"O�$�G�.�Z(�ȋ/7x��"O�����B� Qp�j�0'�,�"OPU{��Ӷt@$��H�%\{�"O*e��ʯS��=l�9B�"OT��Q&�5>�	���E�om����"O��F�ڻh���@�ܨ	[V�#�"O�:�'�		����uG�q/N�a"O�(җ�Sl���� ;�M"ON�R�k��0�~�8����h��"O��S�J)�l�JWC'a�\�8"O��o�.>���*��H�%��xI�"OR墦�)7׆�0� ѥ3�$t�"O����´5�PQcuA�K�i�"O�ѕh[Qkb�ץv����"OJ�酦��Op5K$��.:h�bt"OJ�@�/�?p����6ʘ6$��[�"O�IX?L��<IDo�Y��{dO�Z�<�tC���B�͉j%�f)Z�<�Ư�@���+֕X�~E���GU�<��.q(�)'CG`�,I��U�<�����/7�Hv�(N��=�'��R�<a����P���ص���bPW��v�<��/Z9�*,�v�������1��x�<���>���PEy�F�y�<�f�Syd���9�z�y��t�<�㊜�}��ġ���ze��Q�m�<Q���\s��J0�B�H{�p1!JYl�<�E-ʞT�b�S�V/�& �	H}�<���#"�0�Bb흊�T��@d�<�lB�c�vH �A�(��X��'f�<@�V�#I����Ѕn�ZT���a���=iv�ë0��8�M��pI	�j�Z�<�"�	Q�j�ѥB�-B۰q8�	OS�<ف�͗B�ҡ���Ѩd�e��\I�<� ��򮜊��1�0����"Ov]q%C���`��ʉ|��� �"O~�$$�h����p`F����""O.���晳�l�����tQg"O�dڕ�A�+��̫�C��:�CA"O��I1/��G� �z�)�"x�6(��"OJl�r�E	On��$腃 ����5"O ��k8;�ub%GW08�F�:5"O^1�����Ўt���$颬�"O ��1�� g�R��eD�65��ɖ"O�)a�R����³dP� ���t"O���E,�Nl#�Z1 "O0�g���t��_i��9��p�<1����h|a��Y0�����n�<���F`�恙���;	��us���B�<yah� 	s�J#�/6��]�f�CE�<��&�{I�Q�U�K��Mk�"�V�<��T�r�Ԩe\A�����KP�<�c��k�nJ�`�ڌ �N�<�p�B�"�dt"քǝ`zeX5�SH�<i�vj�چ�CB�(�A���i�<a�A��*|�}(�
%�h�C��f�<Yw�֧0�r5"�,G~ �B�~�<ن��3����"�r�3m�y�<b�J��a�Qb]�KRh��.l�<����+M�"HR ޯ�,���	c�<�e��0���S���PD`�2ծ�\�<!�@ԍ�RlS���tX�Q�+n�<��C��bդ�
��������m�<�R?uX<A�Po��4�I����k�<ن/��]L�H�`�.\k�%��V_�<ɇd����� ,[�"��$�Z�<A���1\��B'.��t����A�n�<1�Kيo���0�cAY�B��Og�<��dN�kh�;jP�R���&.�{�<�Sg�zZr����B���w�Fv�<���4i�3�K��'�e���Q\�<q�J��y���hA��(�XR��[�<�0Ď9Gd�;�C]����S��|�<q��2"�`��i�Q j��ԩPO�<�E�G9 ��@c�Gi���¥�O�<����30ZD�GX���@b��OR�<�5��^���1'�P��F�Q�"��ȓz*��¨�&]b� bn_�{|�a�ȓG�Լ���8��� ����)���I�y��ۼN���)����x��u��29����m�+�2TYWk�)K$�ȓu��u�
Y�8T04m�06�ȓw�y�c_��i�¡��.X�!��tQB0�7��w�>x�	+l6�!��B����d+"�B)�@O%4�����L�ۖ��;t6�
U�ȓD����w�ы7�z`�%��4b�`�ȓXJ�r%*EW%�-���*�]��H+�L� ��&-CBY ��W(#ц��LăG�Oo���1ЇZ"Vu��ȓR��������4G�S���\��ȓ0'N�r��� �(ٔ' �H���.P��`1�N�n6�=#� M*J�n����q Bk�	�
��ЀR�l�L�ȓ4�݋�_"5q�T�B�H�FL�� ����C�n��90D�]��ȓS�N� ÿ�r-���"a�M{�"O�s%`Q/hLӐխY���"O� ��BS&�Q����#?@Q�5"Ob ���?b��G�@5[����"O�Ӥ(�S����O Q���&"O��u�@�rW�@��Dܷ~%@���"O�5�\�,�T�����1�]�F"O��jWc��$DH6C�*u��"OR��!Q�	&�	�N�"a+A"O��@��Z�C��!��N&N�9�"O�*��P�N� f�؜K~NAKP"O �D��\���PՕwl�]+E"O��K��	R.��`oR^&)��"O���!.R�O�E�Հ{�����"Od�A�h� E�`
!n�	4$���"Oʠ������"S��*a�`V"OvE���@�{;J9vV�"��X�"O�)H�H���X�K��H���;�"O8�q�E�Ur<��I�,d��k�"O^�@۶y�.A��o�3|�> �"O�YT��.2������9�����"O�e����X��(�à�S�D�C�"Ovpr���)�*
oP3�LE��"Oj��r�[Z���T.�G�j��s"O<E��^F���
G�M+gnV-��"Od�)�HWr� +�OI4f��j3"O�c.�q�4ib0��[��7�1D���c/��[(�Xi�Ι�CVB�c1D��z&I
�5���2�*Iu�UB�K-D�4�fz)A���
b ��M�5�!�DV�b�n�"�(?@�Ѕ��,�J�!��Z w��a�@��&��ezqJ'6!�Q����7 �p嘕ʑ�a�!�DV�S\9j݁n�\���If�!�$R�^S�TS�E�%htmY��ܽI)!�dǂ��@A���Q�B�:�F�+6�!��=ӰK�@� l�6%ɺ6�!�d�*�|(Q�$�����WY��!��ٙ@��p'(�9���P�匕n!��V!�]��ْ(�4	jd-V�!����!�*шx�E#$E<�!�dM�d�
�b3��rP��JҤq�!�	x��۰j*<E����Ȍ;p�!��4 �N�;�l׮e��q��� x�!��ٓ�T�(&㛆(*���	>!�A�aS��U����)�G^^Q!��h�D����JB��
5���^b!�d��#�R��$�H�7aP-	�R!A$!��^�n���4�Jf�1:���<'�!�$�=�v�Ic�'Vlt�*��~!��2+F�=���k�-�4��Wu!�$��)�=3rJ]t?d��L�-�!��4c��`B��q@*h��S5vX!��6_Y�������1��/uA!�Rhv%(�oC:o R��u!���f�&3�͓�s⚙8E$�x�!��ȃs��X;@�Y�/͘���_�	�!�䗏1ڌ	d/L
O���8�f��G�!�$I ښ5K�H��Z,��'L��!�ą �$��d�
~d�m�����!�$_%X�)C�B-Ny��ϔ�{�!�d��U�p�ݡL^�5�VNCl�!��A�&�,�dAJ	M1XYZW&X0�!�ВOXp�zEc�M L�IucM<Qb!�DB=c.�T��H Xn�Q񦡟;0e!�D>l��H d�>9b��4�E�1I!�� ̔۠�E+@^��@1i�R��Ht"O�%a�b�%[}�W��wv) "O q ��թ`�� �U�'T^d�h�"O�]if�W�N��4b�8vz��v"O�hH�� 
���'�K�m_�=Y�"O��vnӝgZO
y�5f��,!�䚀g>͓V�]�#=�y׎F�Z !�$1g��i�66x��h��!�$��s'�}	!�R�D� %"�9<!�D�<Q�\Y��M��^��c�D�i�!�$�9��8�2fƀgQ���`��!�9	`~ՉE�ҌmI��%�ǯx�!�D<x�$-����j-YP�ڂ�!�DƟ}wԉ�ƥ�� ��uJ��-�!�DPcGrq���R%#���W�O�!�䘃b)bĨr@�{�fH�$M;M�!�F5�Lآ��"C�F�qv��jL!��^1Db<�[0�ĺ@u��Q��HI!�d&M-��`A׳$�t���H�%�!�5 ;���̚��:�6'�K�!�Dڧ~���1��l)�֌��Is!��]�����M�p��f+�	 X!�D��0�R7�[�d��!�sD�7|;!�D��7��xC�m~6���� <�!�Ę�|S~	���y`ɩ�ʇ�!���Bąp�e��p�&J%�!�D�b� u #צua<�����+l!�� M���E�L�W��-�S� z
�'<�t��`Q/\������ E�HB�'�F�#��P�!��]��옰D��P�
�'7���V�G*V�)�䗱HP���'�� ��VbƍA7랏��	�	�'����ϛ�4�ъޣU]���'��˓`��B��"���E�^3�yR�K>2��*F[E���d��
�y�d��M2��C�%:�5q���y��|�*�3����ʙ�����y���:��E ��<Vt��H��y2�Uk�i7�D�ȬXFަ�y¨����F.��}x��w`ō�y��W�9�Uz�%2oˬDpVѮ�yB�5u�Y�ʘ�c-i���y�ֻK��t�fA�C1���d�R��y���$b��"9^��X4W��y�nB�G`��E,h����y"�5���F�ܝ$Ց�D��yBo �1ըܹ�)��+ !�5��O�"~Z0�E�!�4���mMH��1:D�E[�<	rH$T��0�sPfb��SET�<�F�>S#��P��j�֝�"*�S�<��(\�h3�]����=�̭`��Q�<icK�>̠�p����)�Rh(DJ�b�<�@D�3�@\�g?=bB��t�<�C޿r���E bx�ЫdQY�<�VF�� em�Qc��pf9���S�<���\0/�j���8C��xy��JN�<��I7�؉	���6:x�Q1�B�<�q-O�M�`A� &Wq��l!� i�<Y���.���BȄN��99�)b�<I/I  �Fm꓂·?���#QaQB�<1���Kg�a{2c�v.����@�<��.��4����Ĥp���%O�~�<13-^cjD��8O��lFS�<!C��&��8p�*��;7��I�<� p�¦	'O0��iBh1(J�C�"O�""üi ��`���`͘�RA"O� D��N����@�ŴX]����"O�q��<5�Q�&Ÿ'B��sB"O�=��Ț=e���I	 TL�{�"OE��Ϡ;���8d@A�qM0��"Ov��H6�`�Do\�I�6Չ`"O����L"S�z����Y�I��(� "O��J�i�'��d.B�6�nt�5"O���&���&��� �#�J��$3D�`0c���T�	�M˶2^n��� /D�a�*�E�M� ʰ8�&��
,D���F5+:���C���a<i��&D��pB^1J�x�q��/P��=���(D�$P�)S#��P�1N�:/��˰�#D����N�|��h�  	wE���E"D�{���-V|@/�Mx(���?D��adDҴ
�^c��S���T`=D�����	)I����]�j4�M�j-D�Ա���7bt���F��[�xcċ)D��b�,��0���UJ.@vԊ'3D��	!A��W��p��n̨F� �rfa0D��x@��x�ܴ�� &�����e)D��@Eȕ�9n^����ï� �p�<D��:%�6Q���7���lO���`?D�h�T��.>#�� L��*	�����)D��V*�	�2�۴S�"��0lZP�<�&�u��(������a& g
!�$U�N�`��k�6E���`��t�!���s����M�i���dԢ�!��X߾}��N+��8�ƅ�v�!�6c�l���D�%�v=i�eZ�S�!�DΊSU2��A�>pۚMk�EP��!��h<��X��q�V$��^&t!��'�ZP�X/'OB!E�];Ig!��
}p^�*Ɨ#	gx���ر?X!��[�F��0�A�^�EV��P��W0!�Ǵh���q��P�HQE^�yE!�	�4�Hr��eSP�qw� E@!�D�����c�Q%H9��Ή�H>!�D�#����j�9h�	�6	!��Ŗ+�@!��N�";U*8��iN!�dǹD�H0����:L*�K���!��Vt]ɴg��*P�5a��!�$��&��Q�nX� �L�ʂ�ѝf�!�D�Pv0��� V�R�.������w�!��G,���Y0JV�S`�x�T.�,Fk!�D-mHL<:�C��u<0�ڗOÞ8!�$K�t��-�� 	@*:�a��N"�!���8w@>�������y0�ԛ^K!�^��}���ܓbx���C�a�!�FY��ɘ���*)`�pGW�b!�D�0p��ʴWE�%�t�^�YO!�������Ǒ$D8� i$�E=IH!�$CW� �po�8ҝ���	*]\!��i1������HhŲ�pt"O���nO'#���`��B�F�c"O�l2$DP��/̥W�0	30"O�EYr�ҏ~mR�1r+��Mu�`��"O�*�M,p������-a����"O��;�(׎2�C��I�?����"O�(:��:R��i@�U�0����@"OPu�b,̬��@��*{.1��"O\�� �s*�S��
�8	"O� 4�!��ފ^�D(�%̜��h%h�"OJ��$���q��,�Մ� �B$r%"O$�j�)T#m�t�8'M�f�@Q"O���v��3=��9A�Z�x�D�"O]	�c��	�����o�*�Z�"ON� g�
�8 +�$�q��Q
"OViRAI@^,�p�4-�ya�"ONt ���> �|�V�[�)8�"O�]��@�"LP*0�aCW�I���Q�"O$A�����d��A�)�t�["O����a�_��}��+m�T�ᑆ�O��e�\��Mc�O?��<F��	"�1A��)�P�j���k���FL2�h�U)݋��¡r���>Q���@�(p�8���͖y~D�`�iM���e��l����$��H8�ʋPvpH8��R~�s��(���9\����L�%[ՒI�wӒ�;��'�"jz�V��-�禵r�.}!��z�"D,7��$��ȶ����͟d��	�9�ȥ�Ô�q��S�.µ05�<��iU�7M?��ܺc�K���W,[-���w��)v�', �ˡ��?	b�'���'���]���l�	1h��%E�c��(C���d.��[czz��v���J��%D�����a�Q�`�'�샖�M�"�=��9&�!1v�#h�t��,[�h���`"�JV�U�X\	�#�)�Z�+�'�9c2̒
gY�(P��/I���H$��O<�x���O~qn>���<��'���D�
5�mz� �	#l�j���!��Ģx�lu�A��@� ���8SmL�1޴(!�v�|��O�t^������|�^<S�Շr^�1��b٫Rw@4z��Esx�4��+r�4��H�Gv�;�n�!X�����$�b
	�.#h�ڍ����$x%��$� N3DY��J4�_�=�}(��!���H���B��=�ڴ���
C�$�HEy�n�'��%�H�	�WP��B�
 ������� U��=�񌁱�M{�����Ŧ��?ydџD@��/Ŕ�5 C�-/@�ٙv"O�a�bv6�ӧ��/M&~0)��O��oګ�M.O��aºޛ��'�BW?iP-A"*�x�r�F}A:���-���%���?��u�����hS�<��1�� �] �L"Ժ��D�K�L����ᮞ�|>�I9�.��Q�d)sHƀ\�n,��FMT�H�)]�3�vDѧ�դ,���{��A� 52P�T�-��kqnԧ`�
D��O�dAg�':7������1	у�9k�����(�5<��ـ���?a����'�(9j���t��-�T
څo�k
�4�v�'����|4�@�*^E'$�)f#� �~��΍`��6�O<��|�0`Ή�?9��Mkq��O 83�����g�6p���th��"l�1`,|h��B�Ó'����'��Yc�}
���"�^�Xp��-5��̐ߴg�P8ǣ�*+P-�����*�n�c'/	wo���RF����Ba����-i�"|���UY#׽iR:8���:m���M����~�s�<]b���xـ@���H�v9I�OH��"���'����ŗ!G�@ݐ���\Iv�K��$V���4�?��i�"��^I���Mqd%Pj�͠�)Կa^��I���d�aiB�������	˟��_w�r�i (�#"D�%܌u�o�9IBf���d_""6��2k4߶���Jo *�i���N��|�˄/������"=bqP�GA$Ap6m�):f�C��" ���A�p�ăʌH�nt�G�Q7���Q�~����a�1S\1�(�e��.0���		�MC� �~�'�[��[���/A޼����u_\a2Dc���x��#�Uң����<"�.G�M�4-���|�^>Y�>�i7 >  ��PDxªM�c�= �%G'($
U8�C�0>!U�ҹ,ײY!Ӫ@<p+���a�3;�MR�gT�U�Ќ�T��QN�y0�'x���	Π
�b0���7B�h���-�s�
�%�:�#�A�k��re	�GP�\ҥc4J���y"/XW�V�i�"O a��7���U�b���;� J�P��d �4���i�g��W�A�`�5	�1���>J|g��{0 �7�
|�!��V�@��9+�-GtE�fg�(z��HD�����tHN4�V��;��8)�	-I�1OT `�k�fg�@0��݉1�A�&�'nN�z3�M���A�:[� B�� ��!A�.��`6�
 P8�A� �0=�S�Ј|��I`る�>80��C{�'FZxj��Ƒq9��:���5w��]0ଔ�rr�=Z��ۻc X`��kّ���IcL���y��¹N��!�?���{sM�]h,��B%��{º��e��WtИ�ûJ�(����w~�K7★(���ŋɰ22�A�'�4Q��J�A#"�i�_�M�t�E�]$T�Y�.[�Rp��2@����B�㢥j�y2�&*�l� bT���3rA�0>��叱k��a�fO�aƎB�Z!<�CEb׉אi����8���B?P,f���ɏ>�tKS��:2����@"#<I���_�4�3����*N~�a�N��$�^�_0��#b%Iu̓[8��c���)_�=��vI�<H�`�ߏk��D�'��Wd���L<&1���s����O�5Qv�c���'t���Ƭ����'��+���2c��S$Q
TBۋy�����lWߟ|2�I� ������-/��F���,�8��J�:&����Oם:����!�*,OLQyae��{�d�ѣ>ti1 �3^Q�6M!eU���k1��<�he9��x��	~���l�̌� K��Oda+5�c���W�9YX`���@BEH^!����6���������>�|��ʑq��!����=�=�UkVA��� 	��n��/O?�I��!Cp)ɒp0���U�zGJ�k�}�ߓ���I�P�0DP��L�~�*�� ^S�I$:ʅ��?�
���!���N�e$(8K�㙒X~��Q���.��<q���e1�5{�OV���q$A�*x��oX >��� 4ثO<� t�:㌒+Lj����>s5�!1!�	2S�t�8焂K�O�8p��"��Ds������y򠑭��b�b>�Dˁ�,��G
�_;N����'D���'�Н]ͶPr��\�d<���-��'G��1�𙟸�������rE��6+N`j�4D��KE��`in�P�� �8'.P8�钽P\X<A���XW�Ҟf��t:�B��&t���I�{T*=(I<��J��M�5J�&C���IBY�<9�F�|�x�� �bI��a�X�<a��P�U��	��(, ����P�<��8i�$)���ѻfh�dB�	�	K��С��6�*��d�VB�	��&@2��=|�	�2��f^<B䉯��i��H
R���'ғ,���D��@�t�q*Gb�.q��f!�"O����R�&Ɠ�Es��3�"O�xx����oژi#��X9G~$� "Oz�E�#<��}·�r�]B$"O`x� �0/u�y �$Օ:@"�8�"O����:{����bQ,�*���"O�!����#@(�AŁ�Vg�YKg"O��f�Y/M���A.��hM`��"O��P�1+��=�D�Kۜ�(�"O���ȘV�1���o��	�"O ����ϙs�V�c'�ԕ"�*h�%���
GN�k��|�\�^K��ӄԨ���q��(�O����Od<�qK�?nh:��#o��"OLM����7�Z��U��{�N����9�!F���=~C�Ũ�S�f���ƕ��0=��^�^�#cJG�<Qw�ο@��肤�/���c��<��DK������,S��^�9�h�A�gߒZ�n�H�dސ^�~��K�01�?防W��"�x��@.�����)6?Qq,����=$���~���yu����R�q
�?E������__~r�����	 8���Ӳ$�y�b�@1݅=C�ɐQ��q���|I4! �#R�-Y�A�c���D"�O��H�[w<z����
!�`t�W�'�F��
��e8���'l���(�u�\�;�j�X����'�=l���S���Ӈ�3 �蒌y�1$��҄oہ���:�B�H�.L&��ROIe<x�0"O�Q� ]5,�N�?r3N�t����S������1�g~�"Fa�4��ˇ$r��P�@C��y	�O����#N�WS�H��x(˄˥s�nm��'�i�`
��O�@S2`�`�#x��:2�!LO d����;^F=�U0Oxy�6��,	�b�"�.�<U�\B"O�}�U�==��� �@�16D��A�5>T�B��ٕX]?�k���0Z�ۆ�"�"R��?D���S�P���\ 1��>tx�<��^8M��`n-?9�-����F��ڽ��f�;N��s���W�zdۑ�܉k`a~bjťy�tā�L��!��p�F|�GOF<äЁ��4�<�{��0c����}k3+�� k@l��?D�0FB�=3�!E� $��a��>�	  ��!u�?�"8 +�ZP��(�v��0"Oxl�#'�YQz���:��|��Ƥ>z1O�\[�3?�QkЦW�z���F g�=q���K�<� F�L�� ѵ@7&���Y��p��(
P��|3&_*p���KB�d=X�J�	"LO�C���$��-���acX)J�f��� �&B�I�R�V�)���w�>E�mF:���?�Bڎp���<�}���1@x9�g�J�� RN>D�K�Z&ad����3 ��4�����@��c��p�'�g~Rᙍ�H3f�# **8a��yRb�_�L�	c�4&�ᡇ�v-��5���0?1���t^B	���@�zۀ�k��~��H1� G�i�������fΛm�0����C60=���S�? n@s�B��k48���^�sX�*�"O��G��
�X�cT���5�
�q�"OP�j�?�V=����=r��"O��Pk\�2� �YD�[*_NU�B�q����'\��ꂅ1�3�R#>�@�W��i��"PǞ-�!��*FD�D
3P��M3��S���"��K�4�[P�'� �2!�/WŠ4��^�A	�Z��a)+>�>t�'��`�+ �i��iu#
J9<�I�'��0�$+דm"��d�^�2tЊL<9S�U�@m(���iU�O�0QB-ʅ������VL(h�'vr��3 ��u���B�-
',�L���'V>��JPĹ0���xS[��# �V�pJ� �.G��x��W0��0�'i��c~��`F@�Y��$���!}��z�2m�U�G��>{��u�P"��I�y�����$<
�"�*�5H\1n,rl#GF�m��ȓ��(+3f��y;��I�oѻn7��%�XS�ޠs�~<K�#2�$E�YPs_�b�jeف���`Ԓ��ȓ7:
`�CC�x������^��ą�0���Y�H��=�L8�Ǘ/�d��ȓF3�8
��g���J#ْX���ȓ���઀�f�@�Ā��W�Ƙ�ȓ?+�<Q2,ܡMv�M�5�� |>��ȓ=�&q 򨉺݀%㣋޻�4ɇȓbπ1���]ސ�҃�H�Pćȓ	� ��M�4w���k'�9B^��ȓ>��L�e��fB�6`dq�5�ȓ�(�:UAֲ.���2�<V��ȓi�Q����~�p����r� �ȓ5%��� �Q�4[& �2�J���>����Ci��VM���AO_���X�ȓQ}.D��G�c\�2#��Bx���ȓX/��/5C�$���UO�dh�ģ&D�����Ɔ6W�<�dB��$��2�)D��т�_)d��7�6)el{��&D�����)&��٢B)<,8"U�%D���"�X,)�((���-)���#�"D���#k���1;�@H�x�l1�f D�L)��.}��j�E
&l$UHԫ=D�Ce!#.Z�#���ɑ�I:D���GK�f� ��S�]�4l��	�,D�(��i��[e$a��o`��`�5,+D�TA�J_R���"�\�6����b)D��*V��i�d`I��Y���D�܆�yR]� ~�ӀK�Q�^D�F���y2����8���^�Q�ڕ�B��y�5'F4�(��=����D�
�yb��%(��Q*P�/�>�qCL��y2-�3�Z�����'�B��%�_��yrj�9Q��0G*ϼÄ�j�㏋�y��
f�Ҩbp�ջsHL򃏘��y�(�(y+րp�e-*�h�
� �y"E 8�Tb�ռo��m�
�
�yrAJ�+vX����a-
1�E��y��#�����d�Wd��ť�y��*(�8:6C
9E�h�$��y���\-���ԈX�'����@W��yR��� N�����\����z/ �yB��B��<��cJ'M@��q�
��y���Y�����>U��t��;�ybj��N��q���ĔG�"x(`& ��yb��0��pk�A8>H�y���&�y��-H� 9Q�n�C�q eC��y�=A�������j�X� ��ybD �mJd�H��Y�W���a@D*�y
� ���Ѥʀ
�q3E�	{�{�"O^��N�?vGt�Sa'4}D\�W"ObUyV�@�RKv��Vȑ�
$�)2"OLr�'�9��̋���z���0&"Od��O�jf�BO�+lJ�"O�Qbd�������.b�2%"OΨ�WNO>*'�,T�9v�����"O��3��D8� ��$.	q0�B�"Ol��ǀ43�e�4c0H �"O��B�^2d�U��\�f�~�X4"O8�
�G��Z���T�U�T`8q"O�`�Ѫ�V����e+B�{eйY�"O� ��d��)Ĝ��3醍W+�5�U"O�P� �[�xI�d�˧,*��ذ"O�1(�d�B T�x#�Q�R!�YF"OK���Wy ܣg�)336(Ҧ"Ou�bi��:�D�M.���"O\�t&�X{�� ��5+^��Q"O��	B, J���,g,8�'"O*�`�eG�J��}�d�,�d�C�"O��s�iR#,`X�ZF�Is����'"O�來�TOB��
I�Ѭ��g!�],v���������̍Q�!�@1>qM��I�[����FjO�q0!�M?;���{�O<q�T�	��!�M�X H��ԉ�0f�ƀ!6��*�!��ݚv�@�p���%�zAaԦ��<�!�dĄ�����Jw-�� ��éx!���2�:et��&H�ԡD��1�!��X2��o^)L�,hH��2!�J� �x�Z�5Ѐ)iG�1'!�DB�}�H�� Ƈ4�pU{͛
!�D�ch�k� Y�S��{0�/�!�Ā�	g$���g�.��-��Q#!�$)=R,aP�-̀P������!���1���r���l�HiQ���!�$��R��%y�ʍ,-���*Gk�>$�!�dA;�2�QS���l9У�M�z�!�d�	��Q�c�8݈�P'�Q��!򄐌6���'eT5'2t��혜^�!�$Z�/��9�G��ZsReӑm֑F0!�B��\���蚦)Z�d��ŕ&3!�d��%���)a !��U��Ŏ2J!�d�A�<YK��-�f�fG��T�!�	 ^�0#B[��9"5$�/|X!�䙊B�f1��j��]}%�fA�I!�F. �@0cT v�у�A�[/!��N�r�A b�i�8��l݆-!�d�(xu�׮Ov���-X�!�J�?��]*��\�r�gT!Ux!�$Բ|���`�=w�<,(�e�*�!���Tꆍ�TC��n��� e=\!򤘿G�ŋ��_�VK�x� o��O!�_6���ꄊ��U:���c.F�
�!򄏫"1�B!�/r�<=��,��4X!� H�P��Ah�pn���K�&nW!�D�@ 怪�wXhZFT]k!��	K��1Qwaȫp�� B�67N!���Msp�S6U�����*~�!�ĉ�H_��`c��%�N%�R��=4�!���Tl�y`�B�}�.a��}!��#�@�����x��lh���B`!��S:QWba�����McU�=hK!�"`��[��7X�HA�W��'>!�� ܭ1��Z#AV@@
�9C$��g"O.x��̓/;A�
�HA>y,,p�"O���� jI���ӜV]��"O�D��cS'8d4����ݻ53��D"O(!�O�7-�C�C'y+\�ْ"O*��
XM��M���X8p�#�"O�}�%�FLiv �w�;���"OV%�B��	QA+#���{&mP"Ov ��ִp p�M6'�会7"O��sff�jP�����1c��"O����P�>w����-��Jh�!�"OF���֦+߬��7��1 9ry8�"OZ���I�t�.Ua�,ʵs�4��0"O����䛍G0\����/@.F�#�"O�Ɋ��X.Tb�}��e�X�x� F"OX��Ċ�t|n�Q��%)ϮY7�'Oў ��h��eF�CQ�N;\Lv�h�J4D���K��<�H!B�R��DI[G	1D��*0 +{Ԇ�{�%Oi��y�@*D�<Qk;(�<��%�5����B/-��p<y iKv4M���K!y�80�&\W�<YF�=��pA�	�c>X@�V��H�<�q��j��C٣����+[`�<Y�������!֣O���G/u�<�U�R���+	�qC��¤�Rw�<A�Ί+
�$%��̄�8qZ��t�<��[�����zn>�+��u�<��F!%�Ҍ�w�M�D`����y�<97c�$�2�ja�;Ev��CI�|�<�b�G�rM �� b.�ⵘe��z�<Q��1^>V����Z�VC`�8�Ɣ]�<a�k�U��y�>=D�S��	B�'7ў�'Wʖ���%8��ˡ
�<o|���ȓC�>�S��X.4l񄅻T~Э��;���y�I�<��ā�.iŅ�Ic�%5�(�%G�-{��3�I�(3��E��R�1��޸�l��b�I�L>���ȓ0V��ړNH�e�����W0>	��-�0��ΎQjK�lZ�/	(��'������" Q�x{�͂��\��L����LQ� ��m���5:�X��ȓ�&m�nSQ:N���AB�i���ȓa@ب ���}�V�1�U5.��A��($0�C��ͤ_�Da���d$���j�r�82��|�4tp&ӣb����8"Ds���u�)�(������&��8A+�.q�b���͚N�lM�ȓi|�y��^���"`і:"��ȓ����KJ'_j��p����5���u�������'tЄ�M����$�ڸ	�^1-��5@�g�1����q�����M��W/�)o�q��z��"E�T.]��G�(�
�ȓq*�eH͏7xD�s�� ^Q��ȓ[�8Mi"�3){��SV�;C<���+�����8tr�	�clO˂#�[��hO1��Q��o4pur��ŤN��� �"OT�A���l6*���h�,��a"O6M3�kޢ]�*� 1G��X\�"O$�p�(k�"�¤�8���!p"OB�T�ح�క�+�P�	R"O�(�#n�1;�T��Jݛ>�6���"Ob�i"m�8��s�E�p"O��#S7\� �L!�6I)�"O� 8Y�6�Űh�֌r�%W)4�¶"O�e�"U&������^1;�$��"O�0"�,���x��M� b�P�S$"O&yBU'�/eP�8�˛�M}<5s�"Oti�̐	vs�\�d��/�x��"O�%s�Z?u�&�qedˁ5��Q�"O�b�^�MÏ�X���"Oz�t�LG�@e ��]�(+��2@"O*QK�h�_���;� Ӽ)&�q"OR���7 �]�ab�1dh\�"O@� N��.����M�,8�"On��B�37\���#�<{����"O��
Um]�j���!�����Br"O�h�l���6K�T;�!��"On�K��^ 9��� 4��/���0"OzW��5!3j�	���1#\�3"O&͚ �P=$�%i�mL�Hڭy�"O��0D��- ����	��ȁ"OFĹ���rK�LP@K��f�u "O��xPK�+X�F�T�C10�5�"O ԫ�>lԩA�̎Kv	
�"O��ȁٓ&�j0�b��
#; =��"O�}��%�)���)��O� x�@�"O��%�W�D����$��(�	���'o����� �Q�|8�A�!��U(�B�I$O�B	�B�z���HwFɢlJ�B�ɸd<i �f��C���jQM�1�B�	�D��m�,�p�{�%��?TlB�	�UT���Fe	%+��A��[&�6B�I�RSh�{ׁ�5P���S兜�6Q:B�	1V���gЕ2x"�!Y�j��B�	<)m��%I�6vp<�3d�+Z4�B�ɬ?�j�KC� �ib�15nC�	>Ұh�e#/5�t���>4~LC�	h�NňF�>���K��+�DC�	7L���f H�Kc�HȄ-�;pC�	�	�|�*�6E�|@�a�p�B�1]|h)w�B�*��!
�5BʰB�ɪYg� �7�pm����S����`��<����fur�E�?\ub��ȓ1z�}�Vl
=	# ��!L8h&�-�ȓ`��-�C��	%��L�t�M)5�Q�ȓd ����Y�b�j
02�Y�ȓf��Չ3n��fB����	��e�0��ȓz����)H.* ΍!S�W�i�����رj�#��>���Q5CT�ȓh1"	h�I�b' �&�ڳ%N�U�ȓfn�p!�H�r���(Wb �cL����D{��Œ!�]iD2/-�-����He	BN���Q'�ij���ȓXiN���T/z�ltS�φ�R�~��ȓE~x �K�B<x�� �W>n͸����|�Gׁ9M��j��C�`Lh�ȓO��ŲGL�*p�r�J�b Q�	������'�Ę>$��RB��G`P��� �"�@�%%@ܜ�p�H�~����ȓ58Ƹ��\�1�ƭr�&�Q���&�P�i�ibH�:��G/��I�ȓ���k�(��I�~ȡv��T���ȓB����P2�>����f_�͇ȓZ��J2#N3T4p���ͩ6�D�ȓ��h0�̛2]R*�c[�k�Є��d4�`-�0 {~i�� .1]��$cr����H=c)b��D.�m0܇�S�? *��.�Y�	��`'\�Z���"O���B�:h
,k���@D��"O*��`�\(#��j&o��@��"O&�:c��2qb5� @6�t�"OH�  L���D*GÞ/N$�5��"O
50��ʑt ���, �M��� "O�={��ZCb�Dr�,��H�̕P"O Ii��"a����Y�nDyW"OV<! ��R��樌	�&��"O��c�̀ �4T����0W����"O����`�5 � !lH�)�JQyG�8D� ��3iE���$��[:E9��5D���G��3u}��Pw��3>X.Ma5D�Hc��A�8/��q
֊Xg��4D��[�KM#I4\II�ԫ`#�e�EH0D�`���L:��0#���+G`	:�-D�l�1o޺6s����Ϙ�&�||���)D��A�&�9|�{��C&';DXpR�<D���$�"����R��<d&2T"9D��U�UđbǊ\V�U��$7D� ;s�>V���q��m�g�5D����Ҕs7�x���X+|-���3D��RE��AB�Dsa�	3H�,�W�=D�P�$���ty"���F(N��� D6D��B-�:%��P��ŽkrҴʧ7D�p郇�$@6P�5�4����+7D����j��ִ��ر^��9ӠH"D�``�"��-�r�y�$��H��-�-D�dB�/�3�6�kH*df���C>D�X���5B�p$�!F�~���=D����eɐH�]�B��Rv��<D�Գ�@�e**q bb����Q�b:D�$ ���@���+����y�Z�Z �"D�09"kԢFC�T�wg�'�\�꣮5D��a+�&x�4������[0���M4D�4ca�P�L��,c񁅚S�K2�6D���S-�'�N�����"o��\:Bn!D�$���[v��P6J%{UҰ�S�=D�
��X�E0�sD�]�`�ڶ&D��"e�J�ME�Z�-֏o�b�p��"D���f̌Z��Q�s���T�@��!D��/	?�0Q@s�\<UD�$?D��A	U<��ds�-�aVB���n*D�(��c���t�7��;]6�³c5D�����P ?��E 3��8�hI�K D���D�&R�<�f��?Y)B�[��>D�8�1i�-s�(Q�wǫyw���?D�L�"�շ~|e{���,�
�H��<D��h��0T�x�G A( ��t@�'9D�,���g�V(�f�C�W�>4iC�!D�$��/��hPR���Tn,�`I2D��*��G�-����kug:D�l3�G�O���Q�[�0Z�8�%4D�d0�b��w�9�*Ү��V#3D�l{Ԯ� E5�BC�L�4�S�I%D��1��L=��xRw�۱y�N-[��-D���$%,_�j��G{9TTr �6D���(^�;�Ƞ��ڨo�2�@�c6D��c�_�O��s)�3&���F,3D���dҭJ/PQj51Tu�
4�$D��+�̖M� !�A��'��8�.$D�X�i�<����"G^�:j�\��#0D�8x���^�h�ia*iܤ<��!D�"ҏדo&��! ܕ	�b��wf+D�� h�5�Вjqd���ζP"B*�"Ov,q��@�{�Q�d���>,y� "O��#R��Hl��FJ'$�A�"O�Y8�+Sprxhٳ��V�%V"O��{b�V^�
و�g�Ic8�"O����9Ii�A�FT�%xx���"O�|�̗�#�n}�҅M3)eD@" "Ob�Q�D�4W�0x���]^^���"Of9M2��A��/�n�V6n?D� ��GD�I��B�O$�u�� =D�Ш�W8S����̓'3`��':D�8#E`��d�k�'�W�AQ��+D�P���ߎa/P�S��;�@���6D�t[�̔��Y�F��"Uܱ0��8D������TZ���D�?3��u�q�:D��hC���D���F�K�;�Tc��>D��زDzB�#��G,rN�A��<D����(q�H[�BF�����ń:D���/C�}?��0�B�pD,E.4D�sQ�*V�x}p��߲<m�ab"4D��Z&��$Qmx���/V���%�3D�@)�M�8��=�B�%:�vX���6D�0��)��N$���.�3^�`��b4D����.}�d1@�%�"�k��1D�Tѥ`�:?0�Fj>X�V��3D�<�h\���\k�
A9vk`A��A/D�B!I�a������s	�.L!�dV��"�!'�\afH ;!��C$=f- ��۩ D�6g�}�!��9J�`s� �6R'\Ȣ0÷m�!��;f���`l�\PŪޔ"�!�$�	l*�q�,� "�H��e	J�K�!����� �)*-^�iI�!�Ĕ�5*$���zh�ѓJ��!�C�L(Ӭ-/J��r���H !���hb���w�
�p�����i�!�æI���+5h �2��s�����!�$�4Z�l�)�i�� <#!�T�l`ZB��g2΁��@�!�D]8G�3i�:M~��"��3q�!�+	b���C?eV9��OJ�!�䍑T�kA��a"�����E�!�$��(k�PY."���.9�!����ꕁVh:t�b�֣�8B�!�$A� �h���3#�ģ�%� Vl!�E&/�H�&̤0�<��$�V�RO!�d�7w8��$hJ�A��YB�զ2!򄟋(���!f�IY���p�O62�!�$4RG����G��j�xv�٧[M!���Z�nICF�S Xr�b�5:�!�Ĉ�7c�Jv-ܘ����R!��n�X���:�p�v͡o!��]�T�T�P&K�I��D�o!�$[y͂�����c�V�Kq��R�!���[?����,�~�v
�k�5&�!�d	=B���bƊz�n�#���H�!�DU�LmT��"iU1B�^�)��ͷ) !��$?�ޡӓJFh��G»V�!�DK��]8��э	n�Jc��7!�ձ[Mz}ڷC�(V�h�7�7D!�$πCZ����Q�>R�]Iv�##2!�dQU2 P0j	</A����
"!�9k=�e
A�]�-H�R�.��Y !�DN�,�`Ycmޠ|�M*�#�1T!�� v����?X��+ʘ-v�$"O��ڐ���U�.��#+��:����"O|�
����~���&)�1#�~`�4"Ov-��#��
�*��D��½#�"OҬ�E-
#K�� �T�-�~
�"Ol�ӧ�m@"Q�a$������"O�]@���$��J��T(�D�Z#"O@����T8:h���Н�.�a"OT��WF�6M|���b�$����"O|%���[��0����ݮB�:��q"OP񩖇'c&��G��5t�@9b"OD�!u���)e4��O�PIyw"O$�3��!w�z���*�V䩠"OR�0�Ɲ�tU�=Ф#�dA	5"O\��}Kd�BQ�	:�<��"O�4��D�O\�Õ��.���C"O��cIV�����`B�p�Ҭ� "OT�&��gnT�@̑?�b�"O��Z�@0�F��RV"�bT�<1���#d���n��]�yCǙg�<a�`�r��@�t��s3�M1���e�<����f=x�J'!��-Li#�M�<a��V�p�X�qC"�G�\DIb��E�<)�a��
�p� AL0�XW�<Q��C0 0 �A�u��QeE�S�<A��A�S���`@�ϋ�r��N�<1�M7-�>�y�&C�~gHaj�h�d�<Yl�0=D �W��8�L�@�΋a�<Q'B�i��=�2�+<�r%N�f�<�&��>@mR�#�&]��i� �h�<�a""���EE!<�u�"B�k�<� ��Z8qf�ğJ~,��!�b�<Q����b������@C&�[�<Y���s,.)�#�_�<`̥A��q�<U�I�O{|YR�C'g��U�n�<�%�7�\�B�!¤y�����)Gh�<��fO�W��!���)h
��7��e�<��
3=��s͉�F�ၧ��L�<��o�8
1h�p Ļs[�0S��P�<��d�?Y�|�P������L�<�fCQ��3��9)����f�D�<��kA%T+��c�lۏFr ���~�<�` ;|�iȀ+ր���R�|�<����e9����GQ�:(�pb��u�<��40 ���*X�Q��X�䭇u�<ѥ�� 0H�1�T�6��|a�o�<����n��Qц�UWr@	�˜m�<!���X��
��|0��HR�<� M{)��|	@��ao)#�~B�I�1:�@�N�5���e#A%&�bB�I�?��X@��@�_��C�ɧ|��I���onX�ZE�BE�C䉌2G2 �wNH�,T��N��&4`C�	,G�uk�"c04��BIP�6ÄB��/ R�փr��U�fL?j~\B�	���C։@�d$��Js�,	�"B�I��&4ۂe=Qx���AQ�T��C�	S�4p0V狔]j��)PNLM�C�Is�B|0�(Q,"3�̑Sk d���?��?����$$@F�ϬR�M�D(�
�y��.�j�'A�O3䨨n�6�yrm�U�②�d�/�B��v!��y�6 h�yj5%��R�+&����y2�N"X�f��E)�\��Z�0�y
� ԝ��&��@��f�˳i�8���"O`yaDE�^�p��7�^�j=�t�A�ILyR���X)��g��$�PbC�Ke!��O0o' Y8U�I� � �*g�ǀ~T!�dS	���Њ�<!�8Q��GC!��	�[ލ��ϖ�h�����,'!��#���¬N�\ϲp1'KX�!�dX+dA�xb��Q�y�d��jP�r!��Ӗ8.Xy�ri^�*�"���FAQџ$������|�B6�T�{P����D:pM�P�<i�C� ��I��M���Ź���J�<i# ��W��Dr���B���S3�G�<IP�I�4�:���ƃ�4����ĨJo�<	RF�2�6@+��D�0�;Ьu�<�SJ�6t�����c0�	��@�m�<B�+ .p���ܢI�2��b��l�<���R8���Is�US4jEs��'T��
Ս΍kf���1A8s#`٫U2D��+U�}R.ðj���8k�J0D�|�e��4�j��^�q��Q��/D�p���u�ƨ�p	��YC�]��/D����-j����4�וhx)�4�,D��q�[U4$:��Ŷh�4*D�6��B��k���V�X�b��NL�<a�DRCR�ڲ��9u�x�9 ��D�<�Rg�<�:x9��R�����VE��<94C�x��
'Hҽ+�D���V^��%k1D����h����G�#iI�=�D%D��yg�Q9\�.(@��ً��-)�A"D��� �@)�J ؿ
���*Q�!D� :���{X@��A%���A�	-D�h�j�q�����D��l�8�)D��rV���~����kK�hsׄ�<�+O����#��)�A��&��c$.��q�!�ĉ�FA��㳧��#�0��G�#�!�dѾ>�FaʳxhXl�#��wt!�ڿOzRd�!�(� TsD��
b!�D�>\4a�����A�f�ZsU!�D�o¼�K �C��!�~H!�r{F�!����h�d�ʸk!������rr�ʑԐЄ.l_!�d�[�I� �L�Ftb�ퟋ,�!��Dm@��! ,	�*"Ԡ����W�!��X�ıb�R"	���p/F�E�!�4c`�(�jӬ	��xQ�ěOg!�d��a&�!ye���^b���.�.D�!�D\���[�I�|��bpm�)|D!�䐿f�@�0��)��(�k�|�!�� S�z(���WkUd24EܒQ!���r���(+7�r��Tj�$C!���	A���ED�<��3t�)!�$ľA�\�A��R nJ5Q�Iў,��I,9lK�.�0u�0�TJ�3�B��e��p`0zībkK�,���'�S�OR�e���+phf�R�[�	>4�+#"O�2���*fm�I�G,lPJ�"Ov����{����P B�]`��"O�P�������J0"�&��"O�,��fX	Fl�h��"9�L4k�"O���ʓy��V��-����d�|�)�G�"Q1��"e���Af)@6���?�S�O���S�Ɔ�|���:�c�
)�F��1"O��pa����`���Eu����q"OB]�PC�*L�u��)\#��Q�"O� �!�(=��(S�^��<M9�"O"	��Ɏ�Vk�d�C�Y�)OL�X$�|��'���>����0HI$��d%��{ c�<	w���p��y��H0z��M�c
�4��|��|��D��
´;��+�H�b�m�<2�!��5��d�(�����pOF�s�!�ϱei�D�c�Aw{`4�$�"!�d��� gM�Ye��"��L
�!�$E�������� D��!���'�|����3WW"I�U,�8���Ȳ�4�vC�	*Q#*�˃̒����z��U:���d�C7�"~��bC�����'����k9�܄ȓET�ຄ�,^$��B��Tk�E�ȓw��C
ٿuo0e���%�Vd�ȓ1�0��e�U �Ar*̞W����ȓv�2��W`C�ΜMQ�l��l7:��?����~b�%[9(��j��
�`�`���YB���hO�'
8�9�DA�.q�HU��'o�6�[wl����<E��'�0i
�(��?��=[0B�\�b10�'�Xܳѥ|��GH4M�>���'�yxЯ��n�"�����?�4P��'sDt�Q�ݘ8���C�31�t��
�'�l�@��ؙ@e���@	��W��1���hO?!Cg��b���4`}��5�h�<	c˂�Mhek�ծ=((�BT!�⟐F{��ɚ;;���2
F�M!lUcD��)FB�I�'^fܒ�%E�c����C� t$B�	�?/���m��P;�]�Sn����C� S&��\ %K���C řS�^B��dM�$�Y��a�jX�˚���;?y&%�rh=33��K6t��ey�<y&I
<��qӁo��e���&�Q��`E{��)�h(i9u�P�n���jX�4�|C��-$)E�R�)���� .�.x�C�I=!��q��/͗ Z�M��C�7��x�a�<$��Y�GB���C�I�E���w'�*ފ�CIڔrӲ����O��ɮ;���y7*
����B���0�zC�Ɇp (��Yn8�@�V��.,�T��/�S�O��Ic#I�tډrCL����v"OL����Ӓa��u�4��+H�:�;�"O0�Pr�M2d�,�R�� 8DV*e"O���q��)F=�HDn�$��W�'���"G��$��J?T��w!�?qbHC��<	��z`n�T��`��-�#�nC�&�*���ؐk�h|�Q��1˞��Oj��{�'�v x�@�YI��Aqc�g+�'�f�؄��7Y�dq�	��� ��',5��D��4aES{.�L��'2�0�ԂXH�AP\�o� y�'���+�g#$�\ P�,P`��8��OP� f@D��Y'��r��"OL�:�e�]&V�Q��&x���#�')ў"~����)
0d��L4Z�đ��P��y��H�>��£OB-Pm��9t���y�)+G���c��	<I&��/I��y�A4�z���K�lp@���K֕�yBd�F�ڒ�!e�����%�y
��Nm,���X3gG&!q&B7�y�hC�<~�c��\��BA��y�A�|��ԤV�\� :���yBd@�Xc�|(�B�Lx� q�ė��y��?>X,�`K�G���U�Z(�y�h��
hIрǭG�"\p�I[��y
� h�c�"�.��)���c�J�{%�	\�'8�hCF��v��:��
�`�+V�'�ў"~"��W'7��k��O�y*ѳÜ��y��>.�	��_ o�
�R�H��y��=C��z��e��X���y��ٟV�^l����[ P�1
��y�cܐyҔ `���L4$��)_ �y"i�'.��(�"U�w�|!!M���O,��?a���T�UB�P�������$P����yR-�V}H%Q�ʊV�|�nS(�yb�
�7��iy�D��N�\17`�<�yBHݲ4��5��,G��5	4�Q�yRUd(P9RӤP�:;@�s&��y���?.T�i��o�<1�M��g �y���38�]��#4y��t0�����O���.§4�d����L�s:��d�א8%聇ȓ���� b��MU����&��v�z��*�.�D�Y,��f.��[�TD�ȓi�A@$å��8ۅ5"��1�ȓJ� i1�@@�~S�bƯ'^�����@�ۍ7j�D&^"�6��ȓK%��q��T(Rٺ�@,�,�F{2�'W?��/�3¨H���:@s֙x�N4D� �Ao�5!���4R�Sg��2f�,D���D,��A�������A�%D��j���8Ch��z�$0D�� 2'�h�TԢ�,R�1%���7�8D����δ;g��� #���8U.8D�,��	J�~�z��O��v� �<D�X��ȬTDZjpKLI�J4���:D�p:��Q�]0�PA�--$��ah9D� @�nÅu�bXɞ�3�ꝑ�<D�@��E]�IX�0��m��bd��b	:T�02fF��4��cQ*u��`�W"O0X Џ��"J�:C�
��-C�"OP|ۀ担q�N����J�n��Tc "O~-+�^��p RT�U�]u*�d"O���j��|j0��/8y���"O��À�M�E���FN���F�y�"O:5�W�g~�5���ϙZ��YA�"O��0��5�~��2Iމ;�%��"O�8�` ȡ^^��g�"���2"O��J�gV�oh�:UȂ|�@��"O�C����M�ȍ�1�S�K��l+�"ODi�D�0�"��䝩5�x���"O����>l��*��C�Dn��hF"O`���F"^�A���3GLL���"O&��j�V���[����d�0@"O���%&9^�F䡤oM�[�d��"O�<�hu*,m*g�A�4��"Ob����F1	}�H��Q�&���k"O^��C�����H)f��E�x��F"O��c��#�LxP�NRV����f"ON�@3ژ1�H�$�;z��r"O�%b��3D�M�#/�N�����"O~�)�+8(Ҩ#�.��'���6��Y�ȳ��i��}�����nPS�+�D�O^��� "Y]D��ކ4��3d"l'!�Ĝ�JT��|����#�
e!�	V�T�3�N {^X���aW�%�!�$�0?/hC���z8|� ��
4�!��лz�|�Q�똨%&��z�V�1W!�;c�nd �Fk�8�"\;�!�$%�Ԥ�v�4A��ҁNC������Iz��� ^�J��E#p5f��$��2ȂuYW"O� ���;��a���W,���	g"O0�+�5-�B����MB�X%�"O�z�
S6�hL`�Iʜ�Di"�"O���f26z��5N�%TD��"O
��F��5f��r�,_Op�"O�Y q��+X�5,���	H%	E�m��Q�H�S��I�{a~@� ܋K��� �ϝY@�C䉋A8���СZdJ`�4�K�1/�C�I A������3��١'ʕ�(C�ɹScT(����!p�!ܕX�FB�	��H	��ϙ/�ڹH! �6tB䉺b��2'd��<h�xP��;:$:B�	�L$re��G9�,l�c��	v��C�#Q_����L2Yn4؁@iԉ�jC�I�_�F̱�J�����w(Q"�dC�	�k�&H��FS�	[ȉ��,	��4C�I�Gz҉���Wy����"!(�C�� Ӗ��W�V.|�k��Z�Y1�B�I*����`D� f�6K�%c��B�&3�J��2�ۓ-��@�ǓNFB��o�ٛ!�	9L���d�+Q�C�	����G"A� ���ƍ�Da�C�I/���!"-ҋ[��*��L�Q��C�("*�����	��8à�
�uaxC�I!<Š�R���b�\��cE��pC�IVT�(���hGv��򤈡z�t��>��|���
�jw�u`��]lGƙ e��8�!�� y��y
Q�Z Q8��wc�8H!�dџW��Y���%wN��RGiM+!�Dч�Hy�$���K2.�)�I��!�U/0�3��_�z��Xy��R�!��ؠ|��Ĉ��;�l��%��<�!�dEP�!�E�$A��vH0�џ�IO�O�B4!��Q�N����A�D��'�Ĥd
�Q���Q�:	�
���{�J����`K�+��u�!�d�&<�&���d\>V��ѤjαXD!�J������\�EE~Ux@i�N!��ؘ�����M�f��E�ah
��!�D����f��%7i�Y�ӆ��'aa|�
9¶�ӄ��`B���y"��(̜� A"�����2�ۗ�y�Dޛ"�0�Kd��b�D�B�Y��yn�8�����j��T��\�y�����#�9ic�k�cF��yr��$e�-iv�(u&za,��y®��\��5!�2jʪ���g���'aў�Ov�
� �1-Ju*��ڤG����'�d]�
^��J��S2"A��	�'��ӷ'�
�a`�#t}��'n��Q�M4$H�����	�z���'��=PP��(p��3�k�#�<��'R�l��L?~씋&
ӡd�V��	�'e"ećX@���EW)Y�X�A���?����������K�� 0V
ŀ�K��һ B��m��$�*F�7i@�f�.�C�ɨ+�0l�sD���	H�Ş�k�C�IT� E����8Rj��OپC�3	Y����C��	�̀	dٮC�	{E�m1 "�̨�d�W�B�	�3�ni��� ~�t��A	����E{�O��d��TT�(A��f*��B^	_3�)�'*
&�
���-h�@��Y�\��LX	��� >h�4E�"6���ffI�II"Ox���bE�E����Dȴl��њ"O޴�ƣ�(4�zfe�(��=�"O�I9�Ja�b�"A.��.���"ODW�h|H���Xj�����P�I���OC�� ��aqD�%@_)K����,O �D1��p�'� �c=&�(e���ݴI�$��'�n䢥��WHTh�"l��Cs|L!�'	ɘ3��uVH��ʞ�?���3
�'�nѐ��C+|���e��>hZ� 
�'��ӧ��� -���5�K�2>�h��'(Y�h�jؠ& (�̂��D*�`�I��B;� ���R����'�ў"~r��Ϳ4�v����(Cff$x��yRH�j"��Y�`K:wz<P�Î�?���S5X�|��͓~}fe�Q�Y�^�B���a�8ѸrG�) zN(�D-�J��ȓ&z̅ I��S���(w�U<z1L���F0��Pq��F���S��R7Zj^��Io�IVy���G�(&�p��+[��E2�n�(��C�ɸ9��UK@�ΏU��Y�a��e�B�ɖ
W��dd���	aFA]�wp�B�g�(�rC�ɒA�H�h�ۏ ǸB��5JN��¤�V  m����^#�B�Iie�)*��Nh�TiiA�A4��B�I(#�����!M��y��ԏh�|ʓ��$��)w����MA38$e*a�"�R��A%D� ��S�(���1�dةF" D��kp�Z-_�T̛v#�"�h��ad?�Il����	 Pp��#i�2Eֆ��adV�LvB�I�fH<�g㍊)����a��#�dB�I�M�����K^d�Ԏ��38B�Iuʘ�zv�0*�L�/�:C�I3_zpuHs��wmn�ɉ23�B�ɝGw��rE-�fi���H
��B�	�K�IH3Ɛ��P=.")����?	����S�O ���rAX��Jq�RaNd��'��*@��#�R0/�=X�&�P�'zv@� �R���'E%A�*m �'��	GI��V��9�3���8���)�t�������'�59��x����䓺0>�5��	
��\)s��V��v�<�`G3F𱒇� {����b��y���hO�'��,!̟F@n\��VD�ȓb]�qG(F.8�az�J���LɆȓ��d�3*D�����e�)Br<�ȓ,�Z���)�*�
q����1:�2��?Y���?	��IL�c�
Ա���� �sp�,(V!��4	�!�e�߹&�j�al�  Q!��(W�[ԉ�(z&a`5���Iğ��IS�)ʧl[���%Z$&{p�Q� �N����c�� �S�NUjM���X5:D�ȓʖ)k2Ϙ�EP$iQI��y��1�ȓ8��"�G6�j����(�G{B�O��1��i;I���Ë�f�ՂM>y���?�t���?�b�ձ��Os��H��<J�Ju���Z�B�H
�'�0:4�
>z�mX���.>�^I�'Nv$2�I��ܽ��� "=e>�I�'����8\�Z8�J�9#&��'<�ɣW���kN��# ��>'�zY@�'�&���́	�dç�ėLR�9�'Q�aÐ�@�C����W+�t���S�<dExb�'���xp`ۀm���#Aٚ�y��G�}�(i�6,o��\�@���y
� �0+��L�s�� Q�^�~�|�c"O8Mj�'�i����C�09��i��"OR%��m��T�f�h�m�"V<:02"O�tу�'���C�TY��T�'�'�O^��!?�);���ᢘ?{@f�E��P�<1f��6N���J�	�:Zl3���h�<a�$ό�@�!L�cDݺ��{�<i��X�lRX��	��z�e�\�<Ѱ�{�0ZB�f���u
FX�<�QÕ�=��PL�|�9p��V�<a@�K0�ҴB��Jz�(]` �V���hO�R^&�a5�$�Q�cLn��x�ȓH.���J��U�F8�-�Zo���	_~B됪W�J�R3`ʴY�h(�t�^��yrf� h��[��Y�"��GE��y�'ՠjƔ�Q䜛W�� a�)�y�[�M��9��P\"�fٵ�y2�ΫN��@2��[M6�kl߅�yRn��3U�T�'S�E�ȹ@5%C5�y�N�5gs CI�P�h��DGۆ�yrd�2ڢ�(�ʜBt�X�êT�y�Hٍyr���@ϻ?�Q�")��yB�лz��Q��F�<�t	{�$���y2IK#M�A�#M!6��U�a�X5�yҬ�df�#�
)3��	X��y�Ƃ�v:���ֳ1�$�Q��*�yҢѨR����������B��.�yBL��z�2�A���a��oE��y��L�!>9Ġ�*>�Q����y��έ%��S�I9N�QF虑�y⢅)Gtz9��#�4�ڴ���yR�؀EX���%ɕ@r�����y�!ߓU�ܠ���t���aumM��y��)P��Cr��>���t�P��y��[w�D��46�&�s����䓒hOq�n5��0��)�F�i`���p"O�)��"��\q�n��r��"O��j�b��QrT�Ĉ�"O��1��E��Z踄J�?��p�"O��(��\8"�Ĕ�E�PN���B�"O���a�R�`  	f���_ƶ�QU"O$eB0�F�q��oS�f����&���O
��&�Q]~G�FS�D�F�Z��	 	9#��Q���5aC9A����K���Q*		N���b��o^9�Ɠg3�"Q��6om�c�oT�KҮ0�'���v�K����Β�<5J���'\�ppU# X(�Aē�/�ȹC(O�$/�O,��M�
�z�j�G&EL5�5"OZ�r&�O�����:5t�"O�(9��_5�
]k��?Q�=z�"O��� ܕ0���񁯄4D��iy�"OJ���h�
^$��R��U�:�(��'R�|��اdע �� �4��9sdF>D���&V� ��ȡ�G<<	����I!D��� �_�p�p��--�n�H��,D�l0�
3R�`�ǫ�s�`��4�,D�X!'��7;��A��=U���H�*D���'�ْ�ĵ2Q�Z�	,%��(D�p�!j�$�NE	ŮĴj�V�{u"�<�I>���O��k��i ����ƙ40�tB""O��Z���U��\r#��z���1"O@����L��
Ɓ�AR�3"O�`��C�&!n�� �;H����"O� D�`��W*ty�$��&]��ku"O�4iVhJ�*�z�#��̑VV6��"O�\``E��U8D�B:!Gd��a�'��|"�)q�ƿQY�]����6�x�B�5D�����i�z���D .e�f��$�1D����  �Uӳ�\��N�K��/��B�����c�n�SS���.�}+VD1�C��	f� �@/θ!wzy��Mr�tC�I�A���� �.ٞ���+L;H�~B��xON�x�n�[ll���G,:B�%BĺI���Ww7ZD��K��+А�	H<�'$�k�P�h�b���|k����<AQ����g����#��� �q�`��J֦㟔�	>!sU�'qd����~{�~-���5D����@�� �۔k�`���!D��
���Uy���]�\�2�C��;D� �����]�$X��nێ5޼ᨦ�8D�8:#�X����*""M~ VPS��O���8�O~Xg��O_�	#R��*o&����'!��$.�Р��˹C� ���aéL���r��`b1�+:AL�͏�_ɬԅȓ5�@��h�8���i��z���m��c�9�Lиb�\F��E�ȓf��Tҵkɐ����ǗU�Ṙ�Yq�\Q&���
A�,y�$`�'�a~�n��`M�H�NLي%HS4�y2A�M�89Q��w��52���
���hOq���x�6�
i��	8�����"O �0ǃ�����P̏ ^f��A�"O6��cË29��"�=6=5j!"O2	;���>d'�KP��o?�MZ�"O�<����\�HФ
� Cx�3"O��)�G	$M�V�P$�ۮ%�n�(�"O$� ᄆ-x����f��X���q"O����c�#��41�U�]P$"O�e�� (-��8cJ�1U��c"O�i!b���}�w� w�,�"O ��a�4��	�#(R!Mn��w"O@� �� �Bݨ@�ӌ9 �(�"OZ��d�8=��J�>a"0PB�"Ot�hN
`D x$�_$%��d��"On��r��!4���dH�e�1;�"O6� teπT� ��Ħ��D��"O�̙¢�:����H�'Ά�{�"O�:�@U�+Ɣ��N�&g��1	D"OX`���4+Cv�k0�_��΅�w"O�tk�N�>e�*�Fѽ��c�_� ��g�S�O.-��	�z��Ր@�+���'����:"�ڹP�ˠym2�C�'�,,ɲ&Q�����A3�,("OJ��Qn�6L�P-�ƯӚ$L�)��"O��� V-%v�Ń%�I�FMd��"ON-�S��R#Z�(wMĂC�(�;�"O�=���(���ap,�v��FV�xG{��酴^��H���G���B��~T!��A%-u�y .���0y@`�S!�d�?BZP�) B:z��$��[�!�N!p�؅�� ÄZR�W��1N�!��>mܪD�%N��$Y�)@W�!�݊J��E��)�;o�:�'+֕k�!���K��E�ʹ
�XسhY?c�!��HZ{�Y �p��uS�4u�!�$-/�u�aϙ8���IW���S!�D��*ފ8p ���ꨲri��%�!�� �c�Αg��t�Eg�8%
]0e"O��Y��7ZT3G��2��Z "O
!�*Әg���Ae�U� � �"O�,�"J�iX�	@ �N�B�b�ʰ"O��0d�#F��l�s���fc ��$"O�D�AE؀F�81#Q�\pd�0"O(��"�X��tR"��r��	�""O�5��E	=�ޡ�� ��y�6,"OhQK�%����G�*��A"O(<0���Д�T�I�N�p�{�"O��{�瓥%� Ba�F���"O�H2�ȊdP #�.�=)^�D	�"O�2b`
YL��! ؒW�"Or w�Фw��I�P�Z�l���"O����ѕ?�|�ޒ"�u��"O�a �"A+Qתm�UHT�
�P`yA"Ob{ǚ�-�f�RF M�.� V"O��@��4b�Rb��}�$��"O�0�Zi͆�r�A�=��G"O��4�l����L~q
�"O�qB��f@�:%�=#X*d��"O���pc��2B��Ʌ�V3#U���Q"O� 
�gO#� ��ᐚR8�U�"Ol�Itg�e���J��/l�U�"O�ei�Âg�<�5莝����"O��9׀�`�,��጖�pw�(��"O�,��l�6IY�I{Em��|�c�"O�X�h[�M����l_� ��A�"O�!��9R�\|�6ҹc�j�z&"O�Y;���CrE��
�"�B"O�$�f�5g� 9xK<jp�)p�"O��*&k��a��U@qj�o~�-�p"OĀB%O�.FP����!z�%x�"OP�XP
�O��QE�\֞�S4"O� Iw��:*}pXk�N�+a:H�@"O*)9���Y����`�Q�l��C�"OTM�R�
����v(U0n�x�h
�'������*�LLq�6Nq�
�'?�E��Q�l� `�*Cz8(!�'C�A�
�!	���0�W�@�fi2
�'o\�+GBU#R1 ���`�	�'*`��EʣLf���GF�t��'a.@�똚�R�B��T79��Uz�'���	�/�*%�%��$578`�'�R�
��9 � ��C1R1�' \y�G��0C���*�T�Y	�'�d���%�Cp��Z�F�+´l��'3<����D)W����V6X��qx�'Vt���b�$2|S�#ҞI.�h�'�pᠴ�ʌ���[whG�P�e��'clh��`	�I�q��?W�z���'�Ԭ�&怫t�@0�ը�?z����'�
�a�S&�5�HO�k�\���' ���7H��uޤ �,�h�(���'����.�Fȱ:�� *h�=��',xA;�ϥ}�j���SR&	�yIS,�HrQ@j�};�k
<�yr�Ċ�d�+h��f��HX��ȅ�y�a�6�2�j����h���tGܼ�yF�N�J��W��]�� ��NZ��y"e��A��툱c���i%�Ü�y29�ر��`^Wx�sSeٛ�y�N�h�f���AI&#����R�S?�yX�;�s��L
���
r�*�y
� �h)c�W�"
�y��Pn$�e�!"OpĢ�B�nc� Wcm ��&"O捩F$K�`��P�mO�0R,�Z�"O�!���V�V�:u��_��x�"O��	�&g8Hx�3.�	e|2� "O���c�<��1�l�-n�F"OVB�a 0&���1Vl�r���"O�/��[��s���df����!D�Ԁ�M.7W0�qbD��oj� �=D���G�.SXY�1A�O�����!=D�p���>_�(��u���w։���/D��K L��2)��-P�D,D��0u`_(#^a�a�KV���rr'D�ܻf�N�`R�QC@�ǒA��y�&D�r'ew֥[�ؑIp�sB�$D� �IYjoJi�����V�@�g>D�l����v�$dQ��B��
�7D���Ҏ��g��ٹ�L�*�@��ŋ D�(�@j�8�1��B)hTF���<D��H�d��d mJ���-#̥B�:D�D[�F,M�L��N^���	�:D��J�W?H.*���o�SY�6�4D� �t�	 mq1C\�)u�4D��c!ξa͆Dy�@ 0�A9Ѡ'D��c�o�x�2���
Q��$�g�:D��p��]l��j֫S"r �H�6D�p����F�X�	c��O[*��4�2D�,Pa���<`�g.�0��|��%D�(��tFΌ�꘬b�T��-D�h�%�ۺV�ɐ�B�Ls�|��	.D�H�n�-|��+%�Q�'f��2P')D��
pȀB���ۓK
 *�����%D�0� ��5yl���e	�8B�a�!D�Ț0+��XP��
v/�(a6~\s�N>D�$Y�O�*Z*��bt$1M�����<D�4�\�#*!⒩���z�"M D� S��t�:���/aO,���3D��u��<�{�,�5
�m�C1D�HY�'�, ���+�̍�.C,�.;D��	G�b�r�bŊ]�
�@�7D�Ġ���L��=�0`ɔ�YZ�!D�@�U��>A>%��-_� =��<D�P�f$P:Z&Jȹv��Z(�Pd�<D� �b�<4�I� �	����g�/D�|���d{HA9��0��0"�I1T��If��yn����ˇ�k7!�4"OhEBs�6F��㇊�-Mh���"O�0i�#�9+/İJ���	Y9*X��"O"��-~��ڢ�߳Z4��w"O�!8W�E!�zq����7�x�%"O�YG#�1wh�2S��1� �"O����
2"������"!Ҁ"O<< qKZ�JT"wV;E�Đc�"O0LhO*6H��2���;\d[�"O�� l�4T��b�CBSG���"O$=��d�YgX�cĉN����yb�>M����sfD��<Yچc� �y��k��}C�A�y�80ƧC��y�ܓg��sՌ�-��0�բ��yr+	���LS�rh�%���y�F�Kl~���膗k
$���ᚶ�yr+T�3��웄�NZ.�Ce!ߍ�y��1!`D0�� \�6��TrQh���y��7f(8�k�� �X��f�]!�y
� 4u��%D�^�$���IY7���"OhYrh�%M�&9��̎���"O"q)Îԁpl3Qf$��k6"Op����/b�0|���&"� 1"O�d`�f��o�*�H6Mܫ9� ""O�9�"b�-z�Ġ-Ʊopv09"Op��.�;a�<����54T�y��"On�s��
}�N�a�ٟG�e0�"O�T�D�،OV`BQ&Øb=����"O�H6�ѣ�M�7eL3}04"O�\9��62kg�Cev�[q"Ob�&#&:��!e�<Z{^��S"O��`�i� �6Ku��k��B#"OfD��E3!$��d!ւa�.t�S"O*K.��;L\`@�C߆�y"O��3caF�gqR<xP@�r����q"OMxT�5_,�M)`	о{�"1�g"O�5� �"N.d`�F�W昐;�"O4�@��~���s�%��9"O��HE�-`!���	k�>�3�'�Pl�p$��:���ч<u�l{�'$�жcR�\ AKW�dI�	�'u�İa���V�H�p�j�}f�*	�'��4KlXazu�ǅj٠|��'䲌`𥗥  �뤈��dq���
�'�ʰ�4��+	 r��dH�c�@@	�'d��sf�| ������_6����'�	��`ۆF�`@��Q%�z���'�Y��b�-,��@fE�4#Α��'ښ	��Ā$����G�&�y��'|��QjH Kz�ɷdB)S�e��'�>��V*HA�������0�=j�'Ҳ"���.(zK7@������'V6ra���豙����U
L��'tv+���}�HE���R�	q����'%�2E@ѧeW�tF�{[^aP	�'�u0���7�U��O�8s��t��'��a���g��avi7q���'�p����4@���z`*	�'�=W% �5��2ix(��!D�: b8p�i��!���a;D���Ƌ_����bI$���)9D�0�C�ߍ#�ڬIe G6d>��[e8D���R�.���G��D�5���5D���NxI�#�,!
�@aa@?D� s��R8T��@�RE(qi�i�C?D��8Q*A"#YhaI��";uxhɷ�)D��Y7���8b�Q3�m�\@>���&D�tKU�!")H�pB���4�g�"D��sv�M�1����5�@�`�٨��5D�ȓvĜ���b��K�l̾)C��2D��s�I�{
^ �,��Z=V�ra�/D��B M�j�zl!��@��hP�2D�������4�F�O��h��*2�O<}�O��S����K���gj��~��̋A�2D�|�5lF�K%���?g F�2D����G�d�8�'቙H� E��O>D�T��'�+u�aX��=@�(Z�#>D��	'kN�e�� �&E�j�d?D�l�Ƣ&\�
���G�Q�XX*��9D�p�̏�/�$Hjbf"k\��M7D�pҕM�.��@#b#���j�0��*D���Bg׷sfN`�p�P�te.��T�(D���Vh�1g���mK�a|ހ�si%D�� `��#Źd�� 	���rM$S�3O����]�Ԍ�ĂW�#�蹱#dS�n>!�$�2�ji����;$�ݳDҡ�v����X�r���efF��@�o,��hO���+���ڂe�m�a8���y�x">��I@�<SܙB@�%����n 1!�ǘRG��r��۽Q�����)!�dЎ
dȜ�whU:Ǻ)����F��O����5b�B���w�ΰ�f�2��7�O��#�)O1�*�R�����}�"O�X
cj��o4���eȯV��	��'��D�t�>Q�4��z����I�tn��*��DRn��yrI�o��q�+�@^�鲤)L	�0=y���W:5fHhAgKٶj�bĬԮ�(Oi�� ڹ�voW���p��hV�vn�%��E{��T!�
B�$z�߄���KU��y�`�!��Ѻ%��ީ9����'?az����T�؉�W!6�^���'J��p>i�>q1B�5��Pj\��i RƎßLΓ�~r�'b?��O�N4+�
�>��f%Yۦq;��ɧ#ĢZ�#��!U�	%��W��{��n�<��!CI�$�����&dS�ٕX!��Ey��)�OvXrf�ɞvW4���E��9��Q2U�@��	p�p1�W��;r���y���Ysh�	�a~2	�G�t1��p�a������>���<��d�Hx��Q.��YGXix��	D}��'�icfg�N�[�,�R�1�'A¸# ��6�p,Yf�J!H���'��M3�ǵ5�d���H�@-v�.ON�=Ys�Ę�.�@w�7��]�QmR73��	a���;��DC��	���/��q�%�7�r�L+5�O�`崽��)!����(6D��y��;=�HHS�+ {b���#�uӈ��m̓e�Q?!���ȍ"L|�ad̚Ίɑ`O>D�(2S&7� sSO?dXEԥ<D�ܸT皣J�fM��K�4%8�$:D�h��Ȇ�n�P�[��	n���o7D�pRb`�Tl��@#�C؅Af5D�,�pFۿ-Z���hHH̚%C5�1D���a�
�/�R �¢�(4d=��;D��pb�W�%���|rdX4�%D�h8��$��
��Q��H�T�#D� Y �"3,�i)�`�' �@g�5�O�II�F��T!r֪}	1��+?"�B��HM&E��Z�[,@�F��0��B��)�L�K"K�*�@� 蕭-E���$�/U���<ad*J!h,�"q(�{��}�؞D!�Q�`jqJ�G�e��I� ƀq'!�P�/R� ��i	*�d��c�!�D��7�VL����a�B��S�HD���D��,T#Ԧm`G�H�\�����!10!����B��E26.���P����9+!�#0�@ԲLG\8��C�ߗp!�$׳xsT��Ś� u\h��b��P!�$��x����C�)6���8���)�OpHP�{�����&�Qwo�1IGh�!BL�:ǒC�Ʉ2X�ar�B�&V<���g�mfC�Iڟ���G�F6er�AE�Z(��
��2D���1�]�/�
[d�C�X��;f`%D��ȡlB+'@�5b��η��d"��"D�4��ߋT%�T�G?V�N�6͟jy��)�'I?���!ʗ�8��T�����K�jчȓ'�
pH7�� ,��@���Z~��� D1A2�]�%<z`#���BD��'2��z�S�π ��[��a��䭟7M�R�"�i���o8�Djs�Ϧsf��Y�'6h1�2�(}�)�ӫU`P�A 2^p���һߖC�	%m.t�f�\��z�#�Q5#%���&������?8|���Av���(lO�Lyb�'oX�%K����!Y0����	�'4Xt	�B������2fp{�'L"�I�`l8��,B>UX�bO&�y2/�W�B�*��F�Ѭ��1c���=��y�X?x�`L��BK&I���!��N��y�L�{
C�	J�"�qAk܌���;��&�'a���0�ǉv���`��Q�;�L�ȓQ���!��6h�L؄�Ѽw��<Fz�g2O^���'�#[��8ũ̻b �%J�በD��Ix����Hȕ@g��P��A9E�p��"O P�G�B�enp`��^0X�QA��'f1O�PL��6�Xc��W$V�bհR"O���Q�D�a�����F����W��;��)�'M��2�C���([�"�M�rl�ēR�J�P���
� a��Y�"�8��>I�`+�OH�wj��p���C�ɋB0H��"Ov�eH���R�P��V����xb�'B�0rA�I�{g�"&48��x{�'�h$�7�
��>U�� �(��p)�'�LEӕ���8LXǈL�I"ы}��)񩇘N����kFƄ�ZAMA�2�!�d�;w��5`#"��`�0E���["=�!�$�O���Eɐ�̚Ē�K�ay��'[qO8��4��%W�A��툐A��ȥ"O��a�FгA�9�r�P-N^��"O��� �ϟ2�����q�.���"O�����,� ���3>B�0:���3�(O�c>�j�&�
�� ��%X8H�����$?�S�S�k�u�s�W@� ��b�tB�	n���bR0Ն�q�C�;�^��d�<a��+W4Aq�JE"(��+�W|!�E:6)r�҇a�'o�PH�-�/o!�c ��x���;��S�?$o��XF�d�K:SR�ܘm��4 P���D/�S�Of�!@֏�y��0�S	�2#�TT	�'�hI1*�7k��p�+p�h�'G`�A�#�3Z1�8��%?����B�)��<�hT9�, "t���Z��&F����'�a}�J4x�4ȗ(��~8
YzBJ�y�� &~�XƦ�eGɹt� :��?A�'����G�Q�m1&�_a��
��'�>E0�iq]��c'#�2;[�����5���2��3�޾4$p
	�T�(Їȓt�<Q�G%O��!1@� �d�dH�ȓ4O,|&��6q�z̐��&*M�)��x�.���.�� 2̤���l�D�������9��m�2J�ݚl��{���*'��L���bko�D�ȓA莌H�郭iR6H*w�g���ȓn��4[�L��,.�`Z���[R���ȓC��@[��ˣU�|˕�A
xt���'4���AC�h�8DB��d��B��a�r'�8lET�qҭ�i��Y��
L�)�B�Y=!A���[T���W���؁Ŏ�D�ũ�FA�u���ȓ]�*�䚔Jæ$z���c�V]�ȓ}c��G���Ň�7)���"O�U�G�(I��!�\x����ʡ�y���*$�����)�g,Ξ�y
� ^l���TPґ�jL�+L���@"O��� D�<:N�TKR��j,ne)�"Oz����5�̨��T�(�T��"O���`�Qܰ�Yu��n�ف&"O2ܺ�O���
V��?R+x3f"Oh�k5σ�:H�|���˖u�v�9G"O�-�f#��5������K��� �"O��ң�k��2�"�f��EJ�"O����G�\�&�BV�N��j�@�"O�a� % ���E�3m��3֔p�"O���Uj4sy�L�k��'��"OJ=� Z���ēd���3j`���"Olt��%�@�iႦʂ h��2""O�P����8 vdR��R�n3h !*O������p#�רc6x�"�':�!��Z%o�VT ��<
�:���'����&�&I��� 3��i��'����B	�{�y���ܒ^~���'۰a0VKD�j�
 ����L���q�'���ZTk7$5|4@Ņ�6TR0��'����$G]��9�U�^�'�>4�'X���cf�\�2Tݞ	����'oL��K]#�D��&C���)�&�2��	j��U<k=9�$�Ш@��=�d��h �92͆ȓUD��F(J1=��u�f��E?�؆�2��|pCV�J��0J�^�V�r��,���杸>ݪŉUD�8XNv��ȓ\���6�ǄBN ��m��r|��ȓe�TY��~Pec�*DZXx��tq� Y1�T�W��b�*�0���\�x�҄O�
z?��z�̉�X6� �ȓ<Xข1��0��7C!.�椆�k�(�I�BF(m	����5���ȓo�T`Icm C7�0��]�5�>d��2d�H���!��`a�JM�M�"���H1�̀���#��I��ވL�d�ȓZ�s(�U�Y���" �P���;%�� 2�U�|0�a����񢕄ȓo��% ֨M��� ��bZ�a���ȓJ[L ��(�$q�(Y3�^�*��m�ȓ0�x�J֣�a����t�>`����Z�>�;b��6�N�bd���p ��ȓYU>)��U�04;T�ҲQQ���9,����|B��.\v:W#\O��e ��\���
��T
�o �db�,�)T=��ȓ�Ni� )�,YP����?^�'�����׎>X��1��f�O�(͈B�v���A���z�0���'LԥA!�Io�t{Q@�1O�6А���v�с��O�q��!�u�g�	�?TU�I�Yf�l� z�B�������\�`7+J	v���`�/c�$��Et�����r�p5�T��:���F��U9b�?��h�9,��h+P�O5nX����|�)�g�2d�<�J��2?��pF�0D��� A�+(*�1����	����f��DYq�Q��&l�w��7z�l�pE���(��4J�h�Q ��ހ@Uzd�u"O&e:��I�&A!qL �%o �"���$u�� ��Q�4r�Q)W�&a2ׯ�&I9�{�C�3�����9(�(��'�0��<����)�$��G�1=�${��@'n,q�h!RhZ|��U�X�"Q�y�"0��Eg��Lj"왑A�3C�T��.�3�*<�@)Q=�I�7*U9HN�)�#�6dl�rE����9KN�=kA�k������J�z܊��Yy�'���&Ko�O8�ч���vu�CM��B���)�a�,��Pk;�MY�n^�g,����J���!r��ϻ"Z䘉��\�HM�F�I�;�%NYʽᐞ>!����u'f#]��V�,^���ŉ.�bB���1K!f=�ℍ
W�䰢��"U�9�t����'��\�� �*���ř0 N�d��4Z����5�0N�(8��.Gb D1�I? ,B��
�S�(�C�5�F�Aʓj�0X%�Q�g3`��<��Oƈ*E�ĨL]�=
� �ǀ ��ys̏5Xu��+5�[c������P)��5��Q`-^�2h����ϖu�PT�����)[wR&<�%K:®����E%K���[%BP�ʓ�$�f/���]�!�t�_��B�'�԰��N� .�T<ZF�V2')�0¨�o�5��jĠdp+�&���S/�����D�߹X1���d#��.,�@J��5��õ#�<L0��I�U�tM�'n9Y2���D�Yy��9~�����wN��X���-#, �Z�o�U��L1wDڎ!3\�Z"��/`�xE(MsE��0bc�/''��'�޴x�g�;x���R�$E<`\��4r���ǭ�%MtTJ�S�����?5� ��iP�Q��33����;D班UQ\�2Ǭ�^����Gr��J��q���еX����s�4X����]Opz�:�lI�}{�t;a�f�����-VԐ	�ƭ<y�f]�2��L�6g�h_�c�����Y,SҘ�O��<5#�i��k�GW�/O����΁T;\ ��a�'yv�D���Xݴ�>��JK��ͼ� �մ㨰����?��8Ѣ�I�	}He�A.��)�S�M�*ւ�� ���矙$R���A�*kǒPاE�Hh����M[��R���l�~]^`��FJ�Kٲ�K���
��t�EĔMa����]��ល7l8	��&ݕHD�ܙ�̂ �#�#(g�}�N:�<� ���3f.=�"��OK���Ӭ�"�3&R�>Y�`AM�
|Ҝ��b޹Rxc�#�����`̻*���'_:` ���5�~�����T�0 �RA��{�'�*GԌQ7 ��dE9Vx�����sj}�ǠA�RC��#gY	/MĨ�@֖{ t ���&�r&O�"�&)�6H�m��	�@�Q�m�	ݒ��C�%P���X��$�˧s��T{��T3���(�l�0b��@��1sZ�qc�މ��%6k�w��HK����|:��_1f�����aB�B�P8�����) �(��0i]�'.8�ß�"���:�H"�S�}�Fi4AFH��9"�ě#1֐0���уI�`%��B��bN�-B��H����1]#�zFdڠ7ۆ�7�x��t?D��Ò�p���I�z2��i���:=$U*���B����M+`�N�|Q�R+2�v�sF+p��RA��FD������!Q�P��GY.�(d;Ԅ�*Y�8b�`+��X�X�>��'}��W�;rEP�C$L�'161
m�	x����:E�,lj�C��uڬ�����tHF��� <,R�mJ�z�� �;4Lqa'�ǝO8���I�EܓI�����"��<z2��g�>C�@�<�&)F � !�@����s/�a�:B͇�J�l@!>�*i�0��Y���ہ%Ev 
��P��̩��'r���7ǎl@t�B�"͡5E�e�#��6GJ�)����/�4�D�>o�D3Ԥ0oGz�P��"3N���8�P�h��p�C��<y���F�2�B ]��
�;L,��G�]h�6�P��46�4��6g$N����>V��`[jR)i�h�t��K�������mv���DA�sV2L�2A��D�O�my�eB�(� � ��h{���A�p^ d��-@����FD"�U��J��tF�����Y�BB�	�vT ��ω3�|� �q$��G�+������9� ��M;�D4l��A5"�l�;XȬ�P�I��e��4!e��?�i���
qܺ��mG�;L�a勇Wo�����g��Z�#D [�D 5�/��AHo"0X(�K�Sf���J<i'+/"�Ic�H�}u�(�����'�b���d�o�Y""Ofd=�.׊Z� ���@ՙv̡Aaˌ�d�.��Ы*N��@���p`��2,O�3��u!��˦"�����Oa���U�GȬD��	W��8֭O��@�T�
�(��� E�g�����XT�(�܇R����R
�*�E}�e�c|�u8����^�(���Z�,i��_���+E"շ,$����4��=*1. 8V(RE��B��3�^#��%"��'<��XJk�����#4.��S`�"�t�|Cv��6�E|	꼻�˻".*��'D��~>��`˺'%:ĺ�&RVÆ�㡌��8�x�dm��j$�!��	>�(��!�%KѦ�� &��Tƈȳ,�.�ēp�ݻ'N�V��,��S6�!�-�<y�2�JU
��>�4	A���p�͋WN+R�� �㋓�0�%i'͑�$�����R�V�f��c�˓�KMZsf���鞩O����E�
�(O����/ǑYth0�2�
�3h�c���M+X{%P�/�����1&nԍۤ �4P1��H5f��'���h@�@T��s�FFQ@d�5��%6�ƐB��N�'�����GBYPD����'2�֌r���>�4�� ��y0p���6�8���'R�] 8\�w�Bk�m;a���Hp4��Š�z>d�K���2���G�+\����H»w:����LM�:��ӂ�i8YP�Nv��y��tP䰫��Іr�` q7��q�(���8|=A�T���S�9+��1��A�Ms(tHq@X�5�b���2*�L�dG� ��{co�x�I�"�꽋��X�=V�0K���G��q��_9��	�#��UZ��	d�M�&�����)ز?_�5��@�����.{����j�"vQ�U���r����Z�����\�J"=)g�΋T��a�So���t #��R���;���F���	ǳT�P*\�Ul(�@�Ę�r0oZ��F����A�DL�(SC��t ��Y��O �9"B5'`4#=��;Y��1$�
 ��(s�!4��{�U1 �x�rl	?+{,��F�X��B=C2L�( ����炩i
�}kphT3%�p�2�,�=-p8��& �6��$̏�.�Fm1·�3}�1q�3:y��%�)n*��x��� C81��NUС���]4o�8[bd�<)W��Pg��Ӵ)�3'ln8�N�_��x�L�!3b��E���OЈO��Zv�MK����k�����ʨc,� i�ߝ_3�A���>"���"�b̐O�����Xm���[��
)c(���gl�f�f�PF�W�L>8!���y�X�y��'�lX2���GLW�&6&x���*������PpjaybCB.v|��iʛg5�qg� 4&|m�yX<EIc��O���r���5�D��zŉ�ӅO�D0@��DQ�7�J����[..�D�3�F�
K�q���pc���+
�'�|�t �HT\ȡ�8��l��bL�O�$����dكkK�!�p�OI��zp���v	h��٬>�d3�'f����Wی����L5v��Z F��zH��-=�Lc�.�.b8�q��1?i�M��+݋|�Zl[Q�S�F*�&ܥm���ꄴ�0�y��ɗ���"����H�3�ӈ*��MI ɚ)�����$:54��,ߕ���B�
���\�c�
-��a����.��Y�I����� �'|/�i�@* ?�a{��Ż,@]�tC�I�&���dU�Y�0�� ��M>�}�4�ӹ[IX��eHS�p<���c�N��fK)�SdZ��� ���gD'37�Д�	�h:H�������X��}$b� h ��A����+�AA�,���c�F�5�|�2 �ő0wϺ�6HK�;2���7�C_{��k>�ئ� ����� �n��<��$�\@�R�Q� ���O�^�I�'��d�:.�
4v�X9�!3��Yq*D�a�ҭXS'L�cdm(��X��F,FN�?])��J�HeP=�� �	d��"��
6����D�>�c%f��L���Q�P邙#|�f�ŚIU�P
#Os=�IZ<xL�q���
���ć
�2��ѫ�
�zRn��Y���V(��	�l��t)!a�kJ	��E�� {�t�΍�Aˆ���R"+�'I�o��h��Ӧ(����N�<:�h�qNK���x�i
0�U��ޓe�ް �ߌKX8��I6p?�	!֭�����d�ýX˄H��^g�ʜh�I�NP6��5L�6r�"�
�*��f��*��1N�Q��Xpb�e�)K�	�� N��8r]%��ik��!\���!N�Bq��j�5 ? )�EGɲ*=�d(U��yC���#Yu�'�V���B�8K9�l
e�S�/����H�X�T
@�Wb5K'�]qx@�B�)ƔN�
t��%�uҁ���1ᤘh6�6B��Trs�A4C��"�.�c��Ms�
̤5D����&_�Lpf��%4��E@اG�t1RE�Bj�5�㏫^�QT�A�#R�x(�f�� ?�� ��F�@I�e3k�:U�Q���b�vɻD�3�E�'�M����P4�}�tƍC�lܫrnѫR�Dk��7Jb��0���=)����%6P0�Y����F�z���NЩ�E��*!� �3���!jĹ�bő�p�
̇�	�=1 � �n\�-�~��� _�Gԉ�A
� OnA�� YxT���Z�-rD�i��ٱ�F�O3����ꑡJ`a�v�^�	YiT�ʒbB 4�	jw���.��k (Stn[�P�eÀ+�UTLxh ���C���@E�7�ƌ:0A4^�Q�G�o3�Qwg��!!C�ܗ{��U�V�߅��<a@%\;s���Ϊd������ Y؁k� ͌_b�����	8H6�"�E�u���uFO�`�����R�Qʽt�C�*�(����[�Z�88�r�ϯ��?DÈ#w>���gMYB���)�-c�TIR�B}֬�e���:�"�M�#v:�0�\K��HQ�/f�DQz⧂7 &	K�LY�v�X�`mݨ/����	�g�8�{Tb�1m�RYIDl���Mx3��qutY	�*�ZDZM��z�$g�D�*����H4�i8C&�spzyY�"�9~"iA� S�&\���a�R�G��'O�Py�ߧF��sW�%) 
@jW�
�p1�Ej$�	9u)�`� ��I��� D�� ����/�1("U�t�Y�Bqb�2l=\O�{���+^D�	��!f�\��^;4M̉���#��="j"q��3D /TR�aB��#c�^2����c�Թ&^@!���R&.5�!��~�'���!U��W�O��yKc&�&���"vf�[��
�(�52k�1qB�	�eg]��,�!P�zas���$����f�_��,ReHW�6c��)��Q�-M����[K�@R�dIR�y��$j�ҧ��P$j����$�%Q@��yu��+n@ʈs�.[,`p�H@J
�N����V��s���`�W���\VHEk�&9�(O�5k���9O�: piJ�B^`m�:OΕ�D� �� 9�e&?��;Fb��K�($p�I�GTrq�S�ݲb&����08DH��x����X����V���G��L�q�7�C�����g�-R��U3p�� Wٺ�A�)ΟG�P��$�@�?J�
�"���)��KyܫáA�Uܴ�"��A�D��t��?>r��6fg��l"<Zne��( ��'T��Ki��83AX`�dg�����BFnI�t�j�$�al���P�պb�μ��.ǩuK��b&�����;`�ޔ�dΆ�sA��λ 6���FR=�¥!����c�e*0C�j0��g��Z6�o�����?�@�"߳:�,1�aG^N��ts�CS11���07�ܐVF�DJ4r2"-cCkȎp[�!�dK��XW�34���$����L��P��d$	�#���!��8|�T e`݃NJ�pRA��F��wL�V��$��!���d9~�@m24	�3���i�tXL�rf�N�Fφ�rY`��i�;.�|�P�� �W��mۣ��1"mz�s�Q8l�=W����0BUҠI���E������9ch03t���u
�mH�,N9]�%�&G�B&Q3��̘��8
�bY�4��UzCB0�� 5��u*��Ѷu�ܬa��
#1-�ps�$5 Y;��wm:A3Q��'= *�/7$z8�)w��6F�}ړa���\t[�grd.U;$�%9<����yw ��{/<EU��f�(�����(�H�Gb�VaR��=.t��� �$x)4I�O��a�F o8ɛܒ��P��B'){h���f�?N���IQ�ը�?��&�Hb<ͻ�n��D����P�yo�'�H�14MP�uO�9��nW�}V�4B&�ŜG�qS'䚱N�d��7�	�g�@�4-4sF���NW�z[�<Jh��G��%g$�_����
6v6X�uʝvJ����K	=0�|KW�!�		<4�`�� 'Y��H�fՔB��r�  �0�2�
F�_kPY��\.sdSC���g*��զ�@��z����2�*�J��ÌZa@E1t��7Nd�8ӵA޷g�N�����I��D@��A%��Qb��/�!;Պ�c�`b0oۧX�F5�ȲP^l��I%�p�����m�� Sq�$E2�|RM�8\�P��PB����"�O(,����9�R�\9O������'%P,t��k3+!��=}�uJR%B%��Ò�]�L��'>�ϻLr�q��Z_�^&>&�H�)�=�.� Ȓ/-�4}�"ދq�Fd�S���>����S��ēM���M�H�L �W�N�,9q��a��y ���ʄ�yq�lۢ���|���M-J�F0�7�N6-;e� ��61N�Y���1M�Xl�օ��b0^1(�ㅚ�T=����4o[�D;��D��i�f�z`fG�5�6Hj�C
Hl�X���|��q)gå2v��q d��gZ�(��Ä'3_�3qkO�PǶ�ǁR�L����3��4R�;�Z�h��pÌ��[�_����46Z���۹m��P��K�x�؁oD�����L ?��X*�<�W�71��b")�z���/k�O>��J*�h���I>M��y�{�D����{p)Q,XE�ԧ�1^�D�ڣj�ZN�[1g��j~.�%*�+<��eo��y)� �f��|b�սy����E�Z�93�)�Vţ���X�^h��'�AE��O�0�O�6+�b8ʵ�W-X�,�b�B�`h�B�]�|ц� 憊'I(��'F�k�:7�И��D�t�>������J
!'a^�`����]!��=�`IF?*��s�~�  c`�\̈��e�"u����T"O�  �X�dG%PѤ�@�oK�fq�PkD�I5F&�P���(:JU� �*m��� ��ˉl�.B�ɚ*v�0l��&�u��KU��tB䉈?ph�p����Y~N}����7'�`B��.524����+&��+�*�	!
�C�əI#n�"CE�$���P�L�C�	�,/� �,�2*�,r�l��:<FB�I.��Ũ�M��Q�����K�yBB�I�M$Ԥ�G��26�Q3�ˈx �B�	x ٣M� ���U��L'*B�,��h�l�
�0A��H>Y�B��%#ê�YG���Kn�K"S
�C�.l�ؓ�A�ђ<r׫�7[�C��2��)��!r@�[1��n �C�I��2 ��Kn쐒�'łB�	��y��LW�:�L�D�ȟ-7�C�	�Cr�!bw�l�$hb�H� mSbC�I5/����	g)�hH#�$�.B��8<�(�,��:Z��i���q�B䉌j�n�3�Z�n"�1��P\��C�?��ĹU�Q�g�h�� �Ca�C��X���ª��c�^I��L��C�	�ḫ�PN̂	uDBQ�Q�"�C�<
��y���*2��3/�B�	o*%��eͿv��xak�/qRC�	�d�PHy�M���#+��B�	�p�!�B�W��KeG�<��C䉽����!"�;Zz<��̂�i�tC䉻	Q�1�7M	((} �5A�2xۼC���ЗCP�n�:��r� 'b�B䉜"��a��*@Etbu��c�xB䉧!Fu���	*![��ѱ��>�DB�I�:���0"��a1��I®�!
.B�	"n(x��Y+��#D��zd�B�	8���r�ߢ�|�x$üe�C䉜`q�̀�a9�.��4%�2BC�I�7����"A"NJ�[7�
&(�B�	�iG4y�t�0,�^�Ҩ�,��B�I4V�=�Q�
�ewʀQjĥ_�TC�ɲ*��cT
��K��b�C�� �B�l7~+&@��xln�[֯ndB�I7qF�,ɳڌ
��"g��K�C�I�<j��d��<Hį-5l�C�ɺ`Z�K�G���5���	 '
�C䉣a���	�n���#�mNB�I�sA(�vΙ!;G��5@V*^��C�ɦV���XC�Ҕf�N5ӆ"�(ƸC�I dXz ,_ �\=���F&Jΰ��$C(Vͺx����>Aa�[̸豒 	$#j��1IUO�<YDH�(� �A�G�#��)���8�O)��/A�C| 2�a4��Е�bG�L�@���������ȓ 4.�A�L�!G�rm�R��r���#C��6�z�'�ܙ�4�>�3��H�X�c`�B(AN�]�vm�<���d�$z�,P0�cL&J�x ᨏ�[D����l��P>�x�DO��������?��H,�?z���jCnD�x�B	�7a�l���ǩ	&�yſi#̘Bģ�)@DWG%}�T$��'��\�W����ř�A��"�p�Or��cc��sO�%���h�ˏ�i�	O������� L48��c�K!�d�V�LE"r+>#b1����w%.) ɕ�&���0֣k�,i �bS V�HM*b;�1O����c��E�B]��ˆ�xxF�'�FU��F6zl�^tXs!P����Q� ÞDyFn��0Q��]^5�'�t1�%.�2C����e���RE�L<Y���j"f��)�&��Is�US�2��Bרl���r��P�!�@���e�	��RR�X]�Q�p�e��3!�?�
j�I��xs�ՆWd��aM�,S�|@�$
	�12TM ��]3�p�Z��GĦ�'Wf���f�� \�S)Ct4�[��r���k��Ŏ:�4Ygc�p�$#���]�7W"\iSk�8bx�5"�fU�m\X(���7�V�;��أBk\m���D�4P2|)�kT9a|��c1i� v��-�Jmqp��Ea�$��S3�JY��.}H'd	���GZXyv�QP̅%>/�D��ؘ{��<�&�&-�L��&m�����h�n��m�>�ț�s���ZP	.���0Q��U`��Uh�:^��u8�l0?9#P��ܺ�)���0��c�Ѱq�R�� �١$����e^L4��H&�@�:��C�w��K��Sy��:w�U;0oXId ����w��-ʂ\�z~���n��l��u����)P�������M���FJ_I��=Ң%�~ZힷQ��T��^= ��A8a��92fe1y��uCQ�U��3v�X��?�7@�_?�%Ɂ�`��=2.Oz�0���)"�Q��A��{�	!�� *{t�j�X�F���g���x���G+$��e�Q!D�{y��+ )||�D��v~�r�҈][� j��f7FB7��)R�2��%%�!T��˓Z�B��$B�*�F�26'��M`	�%C�^���L}�"�Z�mR���Q*䏕o������-f�(y�!�$C�Z7�C?�lm�eL�'	18u�d��@�b�������1�'R�p�Q"XE @L:���&��ϧ!�M��E���)��ݲ|ـe�G���cG��� ���KQ-
�\��y�Z<uw�(��ݾכ�aK�|����I��]B�xh�H�.[�@�c�0+���I ��R��I�o4-�B�;�3?�c��b$��0A��rr�T47�N=� ҟB6��N)$�NU[�K�j6�A����E��R*O4��D�C˾�9 �NW�Qb��҃7PL�al�����Y5I0�DJ��	���'0�>8ce�Dƴ��aŋ>]z��V�"�-��S����be+��`��k�>h��ɕx8��:���8�qc!���|���6���P��4X��UC�>?a�*m��m�VNH?
�.�x�F3ޙ��o���@h�s����V.�Jr ��"����;�O� 4�E5	.�߈�f�w��u}����Բhf}#��G~�WG߃O�R#0��7 +v0�t�2ovUC02�`���.I�h�T �ՅGmv�I�=�(��O,4r��̫����D�<���Â8b���UD/i��A�=?+��c�F��YN0��&��8'��"[�o�Ԉ��xRg��m�|��w%P�7�^�,K�@��7 �7H;DٓR�]�۸'��]d�L/R6�0���CЁ��>&�	�I�{˔l�D
�h.ȨP!�S�vÆ4�l�K���<�7,�H���Ƣ�>)����r}�1�V�B~2��G��hy�mF�X فt��U��\"f`�5Y�v�����J`��yE
̧f`Y��o۠^T�oY�1a����,\��4�ç1/2Q�3o�%AҰu��lٲ+�yI3��?�nmj��Z5̌��Ж7%"M�/���}��̙�(�Yͻ[�
�xf�̠Q���H���C4�����f]�c�� �<����[4��Rq�B�A8.�mp2i�	^�r���	�dp(f�^"�h�����)f���r�D�����өE-Q��z�i��*/Xj�ə�*�:bF*`�ܙ	�@�6H��It��**�bh���\�T`D�7�۝@�Ҥ�B�'��ћt�Dj�x��)b3�z�'�Ԁ�1�Ǎ2�Z�b��ڢr����̻Ld�8��E+g:�JG�޽H�NdB�1T�"D!@h�$�O��Òm�#��<pW��:r��=(�&�`�΁pJ�<���G	(C��oB�a�nH�$,�p�i�5��Q7,)p`YU�^=Fu��)�O>H�𤐂��ɀ�

�mtn��҂�,n�8�YÝ+�����G�(#䪖jә!;���"
�ns`أr�n�ɜ;D=���@_sf$ �R�|�#>���G�C��(�3�O� �J@J���?�b�J��֮ND��q��\�ց� ��P|Ŋ��	1A���U�]	
cay�Ϛ�!�a�|�Z9��Ƙ�y�!X�r�,��T�	�n�v�[��BG��y�@� ��f��ը!A
r��x#��Y�t��@)�)³_P�>)w�7#��=Z����S� <�A�
s�P�r ����A�vn͏^�nD�D�խ����]�j������ƕM�L����:��U��NL[�xl��+u�+M�?��`��RrZT!����� �V��˒j�놝���_ Zr�he9������X+l0�,��GX/b�|��h�$�����-�2K}��bv��<I���2�ɈKր�d��`�l�D��\�I�p �bt1:+]y3"���arP��,D$�	��B�7%<�#!��s(�Z���3? Qq3BS���E�'�3/�$!*$��kl�`{�D�Fs��b��FK<��vFO�s�F8`��D�Gw��MR��X�O@��(4��dmd`aO
�'��h �(ЌB�n$qֆF7���0"�IF��ȱ18���G�N˂j�=+�zӑm�W: ���K�'9���l�?/�j(�m�S2�#���:�|퐕!J�lm�K��F+��BV���[���f3R|��i�"K.e|��U�J8oj�c�ڙD.��j�Z� �q$J)n��
!Sْ�n_0�M�Q�
�m��Z�Lқ42��[��
�O������+�8�9�c?cg�4�A�@GТ"��a�%:��V=Ga�AD�ʠpu�@�Y�X����L?��M!dn�! ��'�l��ϓ��tJ�˻/�N �FK�~�*��@��$2\����LE m�L�wϒ8�ljJ9*�\�֡
�<�ЮY>��e�H��)8��ɑ��� `�[ӊ<�D�=�c� �P�	�s�����!�&	�0E
#M�䝈��~�u��J�$7�^��d/_�+���A��e�曫���s�#�?�,P��;3�ޘ���-�d�;�A$�!�h��n�`b��8$WP?�5���[�H�� C=t�:Y�S�߈a�h�$ ��6X�3���%8B���AT��`Å<p�.u��Ğ�e�b�	�O7��{��X�U�8�H�Cٸ��٘�i�|s3*�%js�׿��Cw�V32���F���-�-Otyc@��]��agEv"�aq.��4���v&x�����BaC@1�9�h��P!5�t��癷@x�� �N�c�=*��>@{�MCD�N
4�6�Q 5�`�S$g�5Gv��P�N��H��Ź��4� Ŝ���9@�a��zUZ����9H+	3@B y+%�ڭH���Ã�;�v�A��RC���I
70���m��GM;%�z�,MqFƖ9~Ҹ ��
6�����' �GD�q���,w�ўX�A�40`�Y ��n��1B�$<�,#�Gu¤�R`�XMP1�!�!f�|Pa�[���y�����I�wĴ��k�H˂H�m>U�v�@;s�v��[H!��(J<L[T��9q?t��e��i�����4a Ё3�Ǟ_N1��(>IQ@|{6 ]�"����A��[L(`GJ�S�.���O(���%�|��p�B�#��#>� �)A�yvJ��"BT�`�2ԓ�2m���''
*#D�8�B?\z1Æ)��zrN��b�
b�"�ӵ��O����f�u��G��3^i
��^kmN�Aۓ ���s#m��]��$���U*�5�H�Vڬ0�0�O*I�H�c�a��[!�(y��ʳ	T���ܴ|��'�"\�s,�n�HM���H!��	hfڡ��O��2M� �pkG �i��V�[4LjNx��Q_��3��#��A�ܴO]�!��T�#��"��I۴��'.���u�
� }�)Bz>�jaD�8�\fA�?G21�#8���{�pJT�ưҘO|�tRtG2V%ܜ`D%��P�e����$L�FI:!�B3DRRl�1���	,.A�d
T$1*<SE�?a���d�b.�[�O'�����g�M�ҥ16�>)����ݘf:��F&���m�"6�"�s̀-
���Y���0r1�l�p��Dj*ղ��ڜ'o�GC�zb(	����d�PH4ˑ)�8M�ŠpJ��ҵ�O* ���ФA�&A�dT@�g]&y��b�)�N�q��Ƅ_)D�BDɞ:~��}j�
M -�ēQ��ي��G5{Bޭ��ѣB<�+6��{lz\���]�=�j$�N0dH�����5xG΅�3� G6�Ę,zh(��W� ���I*��{��'�2H�X�A��,��p��)���ã�Ⱦb$�9��0x�IJ�H98R�ػ���v�~!Ч�%���Ӄe�?j6�iO>�f ��^=ll�d�L�T^2�"7
Q`��Z���Dh�n�D��� F�(���顪�Q�T	R䭁���2D�4����X9p��c�@�@�>i�l�v���'Yz%�p���l���.B�r|��3�֐�����+�6(��9Qn	��	^�|7�\�2���'�.&rp�1��=t6��フ[�hx 'e'�Ot|�Qg�2(*��w���TT��SX�K� �b�+{!��` �*9���
��3++�����P@���K�M�����1.@�Q�c��R��2
�')�ax"�ͫ�`�0@b�W�*i��k���*�pfd
q ��!Q�5I< s�bN:�x��/�
��p�>�H6R�r(�<�|�"_�+Dܐ�㨜%Œ�s��X:�����M�A7F�2s�N�+�ɘUw�����ph*=7C^��*��V����4��]A�`&l[�$E�:�LZhq�%�;<O4!��ꑫ^
%�F#�DQ����R�n���@��h9��!%]?H�$	�vJ�(T��#ۛB\���ĬSj��Be$��vU�80� ]%9O�*6�:�O�jdKF��{����V�T`�t@�6'cuɤ��w�LI�ŖN@Ts�fPJJ��g̀�R�@L�� �4#ee���(4X�q��ֱe��%r��y�axҪ�"��	#wo)2��k�-�w�]Cb74y��`UNH�Yk�A��' �|SSg�P�H�%F��~~�A{w�mX�И' "�c�_%l�~ɋ�JI't�	N��W�U;"�^Ȑ���ap\����-}�D�SB��8�hz�G�2��%�R	$���c���p����/�zU�񈉯�p=�7��uNd��SM�|%t0
�)�"{4$<j��*9B�t��BF!&��$�����pDv��y.` ����y2k��zݤ���B�,}x�����v�ўp+$�޷)�>������"�Ѕ/��)���D[�g���ӻI"n��,ʀ��-�Ve�ywv����?K¶<P�ߑh]�e�WG�|��5a�FK�:2AU�ޫm?pq��H��'i���3}�����C�P�⡚fC��y���Z1�ܶf�r�i \#oN8���G)�U#��t�)�f�R(�j�2�!�c�Q��e��/����V�1,����)��<	�eR��`p��J�[���(����VV29a�G�'"�����
t��C��H,v̳���?DE���M�=��TbF������	��Uء�NE��``�P�KC�U�QW	 \P��e� � u�d�^d�h�ĝZl�LYMHK�yȁ��%T^��U�� �e��%w|zD�D��?C����.���̉$�O����	ҿ?0��Ճ=�Tm�#	k�4�;A9�B	�s(Ն>7ޕ�ƨ�>:<��ӈT�;�JY��c�m���3�r�H�ӽiuڤ��(��(�1	��A�.��'͊�M�4;�jh�OoT�9�K��fy����G[�J:����f� ������4z���d�)d�-!�(4&d#ڞO1�ͩ&��'R��S��=�hP���5��{e��8��������j��>dZ����-M=�n 0(M# <��Kv�_�=��b��K�gH*q��/�@�V�#��ϫc���;��{�ޑ����}�X "g�^"btN��=ak,M+�F��;�>��4O�?�D�3vF7%c̸�̂;H���s�E<bj(yK2��>�,���X!;�F�+��vypB �0i�[���$�֜ˌy2��0'�¬��+�>"�����1G s���8M�*��)3L�u���:��`���]�ְjs���n�h���m5�j4�O�+6I�a�v�>��x��gޑ+�D_�Q9�:s�|��E81@�Q����&�.�+OǮi*F�k�ߒR�ӹx=rE#�b�'�h b�딚M;̬��(�U��8EgǡP�F�ᤣ�Oޕu��	Uy`4Z5��H1ތ����y��Zg�����?l.�l�h�یP����Z�ɳfB�l�z���-Xc��a%��k$�d��V�َX��A�P���R�F 8������0���E�=+�t0�)�j^t��yihYd�Iî
<X���d�/Y"�L��=-@��+c���!L��ʵ�:|ɨ��˘<1���3���,^ ���wl���C��	�%K��;�BC�~������D1C�pW��X�X>��k7BB7}������5^˒-�5#�:q.2�)#���l㖕2É/lU2Ȣ M�0�\��0�>Њ�eB��X�I��̶h圙2�ɂ/mT0̲0�����wD�I��*ע��ga@pCJ�y�`L&�6�j!͚�{�p�DE��%>	̻<U,�p���� d�; ��܃ÅS(N�e��Q)D�K�N�<T(�@��~��P�xAN0�����yi���"GP��ÀGIQ����i�& b4%J�|zuL ��Jĉ�.��FR���`�ș2���*k|	��C�$xp��h�/�_��i�2Ɩ�x:L@���d	I��x���߸��dyAȄ��d!vc�D���!���^�ypHΔf?
�X�Z��p���@u�(��G#T��ĸ���
WF����ДUEB|�HZ�M�%z����,qh�T)��G�m{"a[Ր&�Av�2`�u[� ���T)��<I��n�8�%Ėj��	Z�LXd�O��X�'�I��@�"aю0 p-h�{�G��Hg�>�nDF���7Lϖ ����ap�%��!Co��A�0�MKLN8%�4�>�O�d���4&q��äUk�Y��'l6\SB��<M��Z��(���G�? ���)�n��3$�(Uf��g%9q�0%yq�ֺ?B���$غx{�qBR�hOb�eR:D0�/9LM@!HSm��#��z�aD=<$����kJ�AXT���&�>��=���m���Ad�|-(q,B��yc��Q/y#~�1"O؍C�(״aA(-�Q�Ɓ`d�c�	�:t܅K��z��r-Ҍ8*�|#�B�=`�C�ɟQ��I��X&��凒<X��C�If���S��W*���uÑ7}�C䉩x��a�)͛;��x;�g	
�C�D��0a�]@zd�`�D8&��B�4!k��y�*�--��#A��U��B�ɊQ�TP7��+-���E.��wN�C�I<k;�����V8L�@A��	3�6B�V��;ei�.ņ��$���=�C�	U������J�d��|T���'|�B�I
���3�)S�}ٸ����(o�LB��5ZF��q�M#}�TP��"�<F��B��2�f�_'|��P'/ֲV��B�ɰM�n�#�/SK���O�1K�jB�	&[�Z��u�٥.o�h:�Jؐ
όB�I�8�e1�OO@I���򮝹j?�B�]o�2�d���5�T#A�~B䉆J8�1�\�H�p�Z��
C�I�F� �b��1�R��GB�^^XC�I
kT"����ór�b�K����C�I�.���b���-�xX�G§\��B�ɾz���cab��^�EJs�W`pRB�ɒ0�t��S0����#0�VB�ɢ]D��w�	K�!�HN�`B���ܤ����FiР+� FhB�I�}J�# j�ؼ���#.�^��W����Ha�gb�>���ŚzD� 'U�(Q@D*˧[MR�r���8�tZ-Ol1A1��0|�R�!�@DZFBJ�%B�! ��R(M��I�)��!��&K�Q?��K�Y]�jɄ�0��!��n�T���H'��q�,�l�)�'F��ak6��"s'4�)E �:�6ec�	]6fRh):gb3���:�~2��߈R~���THg]���˗�SY�'ϸH��s���h�e���h�K��y-�EO6�$��Nľ�b>��!N�X�$QJ��u\���7}�ȵH����y��^�JZ��s@%�!z�ȩ�Ҡ��<i���ȓ!Tf�j�VF	������d��g_���d��2�-"�M�e4�݇�J^�a"hL�bU�C�[^�(�ȓ=�8q�e��i��i�7/��;��U��`XP��cNƏ&}�-� �Z5(
�Ԇȓ設S ���.4a�-E����ȓ5�F��+�:��q&�Χ?�\�ȓD톄0�G�p�sF)F!q"����1��Ɉ�ɘ�Y�лi�8�x��E��ˢ-N;P/p)�e��=^6��ȓyN���D"�2:�dA���=x�h���g�L��ՅN'��5���*�1�ȓrXz� �A�J-@i`�*_�,`��_�");���Nئ\����:�8X�ȓI��:R�F�P<�䋑��#k��ąȓ^6%	M�?a�%��A��)��cd����ۃQ�@X���Y9�2��ȓn��K%���
����(*x�ȓY.\��$R�%y��ʀ���xPb��
ޝ
��}kj�
}�I��{�M��K�JL�R����Z���v�%��.�81B4��J̤oY�D�ȓg;z��� 7f&�J�I���Ї�s�����L�s�����W��݄�Ll`;E	�-�����Wb�U��S�? 6��f�5W�Z�{� Z+4(4ؙ "ODq����24�-t�W�K���H�"O�(��_�&��X0�´`����q"Op�K����P����a�����"O��(���k�8`�� h����@"O����2��q�f�ȝ)����"O2�K�G�D�9���έJs<P""O�|R#�ܬO�F-�.8e\m�3"O"���$��B��4���"O�� W�m�6 pn
�TЂ�"OP�2��>0�|�d _o}2Uɐ"O
zDХBi�� ő�4c��"O-#2�'e�Z8���	�yct��"O�q��AW�cU�� �o@PKV�С"OҠ3h��'�`���$]�d/܀��"O��J���&�h�s䂌x�X#3"O@�u�� [@I����>��U��"O�suoL���$�橗g��yU"O�s7aA�Z'R�A4K��3���p"O4]�.�/w�+I��7n�10�"OR�3F��1&IP�b��@�[WY�w"O��Q���0W�qpG�^"!���b�"OT�q�@ԙf�0�kkZ��"O,+P�ڝS 
��4-%&6]Q"O\�2�Q5H�P�Q"x0�"O�԰��G�R#.��fL�_ܪ��"O��B@-K�/���q��'3��9"O�A��J7O>.�Z��J=��u+V"O }0⥙2<cd<���Wm�diu"O%�fZ�K5P�t�̍b�����"O$�@�B0[R4�q��/h�>��"O��BU�дkY�@�E�ٙ8Ҹ$!�"O.���dՒIj��a
�D"O��vF��.�1�c%tq�$:0"ONĲ�	�L"���b�1J7�h�"O��ۑB)�ژr�a�( ,`�"O = ��D�!9p��d���8R͐R"O�y
 n�2&�{��X�f�qAS"Or(�$ѪY��`1A"��z!�M��"O��X�ț�M�\�$�
/lh"O4�s!I+	:��!�AH�0��{�"O�$(��_ >��݊�S'�X�r%"ONY�d�&c���k��oF�2�"O�8��)�1t�\x�5%H�M^�W"O�ք(��rǦT�`!0k%"Ov�S%�p�M���4#h��"O$���^�)���P�A��"O}{��m�z���ؾv�P5	7"O
���E9j���&�) n�p"O �s�Qd�f��P$D	�	!"O�]Sv�9�������-Ԑ�Y�"OD���VM V��q�C4�n�I4"O-0DIF�n�����=,���{�"O"����0	0v'<@�Hr"O4{e���t��=bW���@��j�"On0�PLθ!٤�X�'�/zr�+"OP�@�ؠ"f��TH�Z��"O�p8#�ٛ3�  ��o"�`I2B"O�9��vC&�{��E
#��ٚ "O�Lq����M��`���9|�[�"O�Z��?Jx���O�����`�h�{��N#G�����E��
�H��my����1z������$%�Ć�|�*�p�	��,t��f�]q" ��S�? ���<}&59���1�xHi�"Oz!��ܤK�v���m�?�B$�V"OXu��b���b�+R�U_�q1d"O��Xb)סr��pza��
vE\@��"O,� (T>u$t�A�bI��9"O(�� H�m�P=0�A�946d3�"O6y۳�G�}�@����v(�D��"O���@�d���Kb��#��"O�d�����<P�pvK�D��2"Oh�h��\:/���W�?�}��"Ot����:7t����B /ٸ��"O�ݪ!������*� k@͙@"OH�YR�:"_��5ώ�G
�4#"O:�#@�=�H��0�C)g�eXG"O�@��*m�]c��(��H�"O�d@��������dB������"O�����8�xH�'�E�JK���"O�!"�m�4LS�4�wl��"G�4Kb"O謁s&H�?]"���76J��T"O����Q)Y�Rhk���G2���F"OT�˧,ӴX�� #�X q0��K&"O\X�*�A%�X9��!l�y2"OZi�j�!&���kЄP�^�t&"O�I��N��d�S$Ӽk���"O���A�?_�2H#��ػ�*�2�"OD�3�I���Y���-_pr<��"O"и��éQv�E�E�Ik$a1"OphY�G_�w�J�+��� Xr��h�"O��k2�8��laS�""^�aI"O�㑈�""B��豊 YBRmS�"O�����	]`�E��,�"OR�X��b>~	;��C=Ny�ar"O��$�Na���� �  !T�]��"O4�1$M�޼x�a�-V:	�G"OH��u�Ue�^�8Fc^�L�ʦ"O0(����4(sD��8>;T��"O2��q"�'�����f��7�$�"O���6l.@��1�$�1/ -Qq"OyX�.ޓq��t�P�G�	zI��"OJ,�g�.%��QV
�%�"Oh;��ɳ]���F�Q�0�0�"O�(����s�8��� }�d9�"OPD��mX�c ���ƈ?�v���"Oz��j�%0���*�����%"OVSDؿrP<e:�Z%q�"O֐!4m�9Y��xb&bK"�.��"ON��go+T�4�6`����&"O��J̞n��`��!�06�~!�"O��AP&�ua3��,%�V"O"�p7�@���΃4q�p���"O6�j�GT1tĨ7�+D���p"Oht��M9T<n�XW�8{]d�"O���"��R��U�D0Z>�D"O6���g��]bZMr�"؅EG�i�"O~�VJ�����ͪJՄ��"O�� ����@�9Ҁūe���!"O�Zb�Y�~�8�CF�����v"OxA�5�ϦM�`�W[?~�
s"Ol]���=qJ�I���p��q�"OTU��сr��5�e�,|�8s"O~h�փ��s������N$�R"ONl{҃��}Q�N���1��"O���4+M0y� M�O�{ꄁ"On�H3bå_�@5�Fg�&�zI�s"O� ���a T>�(]F�F-Lg�DЂ"O�mucR�N3���dD�3ZL@"OR��.ӑ,���B��/�Nt��"O0���,@ ���k<��	V"OZ��T]�2(J1�°I��b�"Ot���N�I]̠�"��/��4P"O�Ya�䝡%�p+���
Ni�YQ"O��T�I#@�q2�6dd�)F"O]0%*̑A�9�aE�B��8(2"O.�{5�Z��T��fĠY�4�:g"O�|1�jv�[�&^�P��u+s"O&��E
��'"��`��&_���r"O��k&'BO�v�$���e"O*�h �R�E��q��!%��,U"O�5��Ϛ3�VL�� d�����"O�囒�Fv�@Sj����"O���4bٺ1��@_'��B"O�H��Ppy�`bC&2�ڠ-�y� �d��š��م!�s�n�r�'}�+ƎS����5�̠�(��'�ȸ)'%��Z�����M��i��,#�'��9� �&Sະ{�N4a��Q{�'�"yǥ	2����C�\����']]����V�����%� V���R�'�� ���ѲQ�� �C�:~���'۸x'��<�L�ccE�/Jn���'���!m�v���N�(��s�'��U�(��FpVE�R�Ѷv*N �
�'Qb�9��|t�"�ى���
�'��D3��Üxld�u┨d:Z�S�'t(8W��2ڴ$�3rN,��'զ�G��KgBd;/�!*�pA �'^�ؕOE[5���cܭ!�ؕ��'(DB��[c�hZfB�/M�<`��'�ʝ"�̋�E(j���P�����'�@$�!L�!&4���w��3	��2�':���$��?(zL������R�'AH
 ӤMS �9f$��|���'�zF��lt�0�Ą��t�����'Ɋ�C��1'Q�9�D��l]6e�'�4�s���=~J�C��$HZ�'~(�)s��%ErP[c���`��c�'x2�Q� �"�I�O�<[�����'p�Pd�5-�T��u#�(M��U!�'�$eكK�} ���᧐�p�u��'�"�J�)�WˎU��D��HX��'ְ���n�/2�.��"�W>/���'9l�S�@���)U�Ђ�L���'~�P�R��\uڥ�Ɖ��6�@�'���B�dI0s���;w䙽�(��'������B*D���E+O��q��'��0����<�����Aiz�"�'贡�H�j�����8&�$�	�'J21��]�.e� �s�W�.0��	�'>��J�A�Ug䀊 	Љ �>���'�{ע�z���;�O�nY��'jv`HSI������`�T���'iph���Ք5B68s׍��U��89�'f���Eߍ @0�Ɔ��9��Y�'�� ��Ǭ\��p���ҐG�:Y
�'��i�  ���   �  �  �  '  j*  �5  0A  �L  "X  hc  �m  6t  '  ��  ֍  2�  t�  ��  ��  t�  �  T�  ��  �  V�  ��  ��  )�  l�  ��  ��  =�  �  �	 F : ]! ^)  1 n7 �= �C �D  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr�	p>!��L�>P^�x�#\`yq�~�tD{���O(dG6â�ߘ<����F�N�B6��~�'.>I��]�(��d_�R>`��	&D��3$l��� ��'y��T"`/"�	�|az�H?X̴Y��ǘ^�B| �e �x�@�?	hlHG �*&���ɵ@�<A&��H�'�T)r��u����`��/T�i�'�S�č��F�P�+ 8x20��ĺ�y��Y8#N�P��1�P	�BL��'�)�s�Y�1~"AۇlX<�XAL<��8h�B��.z��s��N�@�}�'fvM$��E�d^� jSG�>l%��ρY7H03�,D�������b�]S�lZ�r�̹�'i��1�	��~=Xc@ѯMb����ėL��Մ��?�Ox��W���`�~�p�B��>eBV��H�Yw�^�]�*�x� �nN}��/!D�����^����b��WL����O�B���J�l�٧�QM�H�R�ϘB)&��$:��«z��u;!L��;-�Eaș!��5z�y���6G!���.Q��G{*��\�Ǭʓ��-W��S�ə�"O^���.ONA+F��6[� j���%|O0`� �B�v�ڍq�ڂ�x��i�ўʧ`.Z��y��V�k����=y����&j$�y���^9la��&^r�8Ql����)�O�yA�B��6-�Kd�+�j���yrj�8tE�Q���T�*�2����y� G�g�j)"q� �O>&ݚg��,�yb�D�#ˌa�E��^02}RgN���'|z#=%?�j�a�/>o��rw���b��}�S� D�DjF��$o�`t
�H��,�n��1�>��p<�R�� ��x�h�&RI�$��`�<)Ǡ]�S���C�g]wh(x�ԟ4*	�)�d�p篆%%Æa��*`��H��Es��:u��n+���ᑧ y���A�^89�`�<�0��%kwL1��9MV���&̟f��CƸǬ5�ȓ��q:��Ϭc����U�� ���԰�&]/+�d<sF��4�.��ȓ׀)��[�A���Ȕ!d�(U���Ҡ؄�P��3�ǶnO�B�I�'F!�6�@��$ZB*�!Q��B��7s���$�p��� !+ց?��B�IWL����C��sT� q� Եa�B�	�23���BK�8Uzuq1�S���C�)� j��Q/�9�1u�M�I��Xq4"O�����	_��K�	��7���"O��L kމ����-u��Z`�'A�p�<iڒA�Z��N@W���H�n�<�`kÌf(����B�"�j`�"��<Q왻Z���z�䛫b(h9`�@�v�<��4W�̅RQiQ2Ć�k��Ui�<yW!R#b�H%B�̟�`�.��M�<!@�s��@�B���$����L�<A�}��D���^F?�5�p�RK�<�3��-6�&�i&+��
��XGjAD�<��F�a�<:�B!|��aE��i�<��c]!ؼ,��&�06�ݱ��i�<10m���(C�I��8�	w/{�<�3n�'�$={a��;�\��3�	B�<a���zsҥ��F]5g��(i���v�<����~9zBd��W�.��!�o�<�擰a���N?W�t�e��f�<!4)��%9g��7iC���W�Z^�<Q7�'+�𛅏�6?:P��V�<Qt�t�T<Jb��Xd,�3"�k�<��a�?pY��Ht
�*T���Kt�Q�<Yv�H6�\xa P**�Hh#�n@T�<1�
ס�ΡS���)
ֆ�I�!�z�<AE���)4�1χ(U���p$_z�<iա@6��$�9V$0�q"�r�<Qt�]%L�4�2RF�]�jq�M�m�<�Se��\gX0���r�T$�6��p�<ɓ蝟Wp��2T�a��F�<ٖgE��(
@\��2G\�<ī�}ߖ�I�E�l�`�[PK�}�<�%��{�\t� ��>D��� w�<�c!H�Kھ|&�Up�!B�q%�C��CWx� �i���-���
�B�Lu�u�4�R�i��#Q.p�zB䉾^5k�)�T�p1�3L��>^B�	�U��a���=n(��3��i&B䉺k�����Īsx`y%o�'x��B䉦*I�ӁRZt��rD�<U5�B�I�Y�ș��#|�(
�� l�hB�	'���+ρ!AVy�N9}rhB�I5���۳Vm*�b�E~�B�I����U'Ѐh�^��-�B��_�Di:rcʸs�6DY�+T�O�C�ɩNQ$|2g��E��P�a�im�B�ɭQq����S�)���sE�9SzB�*�ع#́����;��â�NB�	&��
nLo��LXg�I2^B�	;����#�����e�KO�B�;i����55�R�Sd���xB�I�E+`�A��Z��h�'��C�I�q�Ґ����/~�Da#֬��0�rC�I-�H�(�ѾSJ�ҤJɂ$XrC�I	���w@�4�>0�BL�\�TC�ɚ@�B�� �� 1�I�K�)� B��T�@-�4OW?;7�ơCI�C䉄Bq�Abe"P�'&�	���	=fC�	3/&)9��]� (���Q�G�B�I;p�i�OӤ-�&��c��q�
C�I�4(��];y`�M`�/�8�B�I�o���3 �X�-"��G��C䉷s.`�B�S٦	9TΎ�8\B�Ie�θbu��:P0��'F7u�ZB䉃>Tb�"�ɏ%�P�āc6B�)� |��V'�4�H�P��-]�(U��"O^�3���h2j5�F��o�6hp"OL,�2��9<ct�AބM��A	�"O${)�+3�y��*��U�D8�"OJy���C�H�쨰1�
U��-��'���'�B�'��'���'���'�~�����|���ZW��tZ �'�R�'�R�'���'���'���'�jp�5*��I�x!�b�7<��'���'��'��'���'=B�'�xt �j	Amtp��@ИS8���'���'[��'��'3��'|��'���Eb֖_�x�b��ڠ-�b-Y�'[r�'TR�'���'��'���'UZ��)���pi�f�0,���'���'��'���'���'��'�\���A�SJ
hbB��,l��U�#�']��'�"�'���'b�'�2�'(�����{�f��D�;��'��'I��'��'���' ��'1�����^�p�l-X���}�Ty��'�"�' R�'fB�'y��'���'����F��
�1RN͏@�"+3�'pr�'���'TR�'2�'���'~&Y������ֿ�K"d'�'�b�'��'��'���'-��Y2c@6����P�y��tkS;5��'�b�'�"�'Z��'���'?�<�\-qD�ѕoSb�"&M3<W"�'���'��'���'�`6M�O,�J+"�I�F�]��9��L�I�*��'��T�b>�z����5H2�9+0�˩g%���R���J����O|0oy��|Γ�?)�&�$�<!ⱉíURȕ��Җ�?���{j���4��$j>a������<�N�IV၆"r-Q��F�.]�b�(�	ry��	p���w$̳+OH�����(3�@`�4^�,��<)��4�k��Ƒ:�.����®���Pg�ҡQh����O��I}���!�0��V<O� Y���>�<�2�%��B�� �5O��I��?!T@:��|J�{%> ��G(ƅZ3ƐC������D-����z!4扨-yx���'�[�p�h@�H�x�̍�?q�_����ޟ����D�2�T��#�	+!gZ���a��O^���!H����O9�?��g�O��È�^�	�#(��@t�pç�<Y,Ov��s����I�.|RL�<N��tb"Er���ݴGc(��'�b7�.�i>]�w�3iy��$jݵ=�����~�8�����	$vv�]o�D~�<�"!���_ۤ0 ��ʍ%.�aXW� O��8���'�T!��'6�i>��ǟ�����\�	�<�B�IԿ	����&З;��A�'�~6�F����$�OR�d�|���?9�B�,��òm,-h��VD�7M-�	Ɵ���w�i>��	��\8vƛ(J,p8�g�.�@���9��oZe~b�W5,"�h���?!6*��<	)O��*��{_�i�I��O�����O���O����O��D�<���i�V���'��鱓*	�{�N��':���kq�'��6�<���OD%�'�r�'�2�����f�:�f��Cd�_؉�B�i��O��M���s����߹K�S>�y��ʷYA�q���t�t�I����ԟ��ğ����Ń6A�䄃�eH�P݈I�UF��?9���?��i� ���_�,�ڴ��56��b�*ԴZ�I���0
w��AK>���?ͧ�(�ߴ������g$W�o��i��#g�1X$挞sD|�	�����O����O���^�L-��3��-t���� �O�V�1#E�l5�ʓN��ƈ@:��T�'���O�'��E��0��H	�hqDq@1	J�y��'��ꓙ?���OUR�Q#'�i2B��B���2�0Z�L�pFS#]���?1	f�'�t��I�4�	YW�MkoP#J="yx��m���h�	ßL�i>����8�'<7-.����	O�lu�EZ�{=���H�<����?),O��d�<)�Z�@��V"R� (��jW�N�����?�ԩ���M��'�����M���d	zo`��%śg.(�䭆KD�Ķ<��?Q���?���?a)��="#CU���D����\�T�C��I3��ߟ4��ɟ'?�I��Mϻd��ԩC�7v��Yxc�3[U<�J���?!O>�|*6Γ<�M��'o$�j4	E���(�pFV�tb-ڝ'�P�Q.�ӟ��P�|^��Sܟd8�nȉ@K����,ִ�,ږ�ß���ݟ4�	fyҠu���+�O8���O:d1�׿��Qb���	]��y*Ç"�������O����@���x����FBњ#l;?�4 �f���7瘝��'d��D��?1fO\�$�^���B��\H�c���?����?!��?َ�Ix>1C�
��7��}0��4C)V�J@+�O�n�}S�����<�4���y7d 7|-R��6oL�S���E�ɺ�y��'��'H��豰iU�i���	�?YÇK���HS�Ř|<��&�C��'x�	����I��t�I˟T��;4.X���']�:� W�ʳ":�'�,7���BT��$�O����b���<�'hԔ3<�"����Gla@�-��	�|�?�'�?���$z�M�m��U:FP�2�[�)M�Q���Dڜ�/O�4�dL��?Y6O�ON� !?O��M�R��m�4ga�x�3Naj����?���?���9q�=K*O<o�-y�d�S��� /N<'��}�B�eQ����M�O>���3��ן��	ߟ�!C%�L�� ]<>��� �e�	�el��<	�� ��JS�*��' �t��� ���g�#<Q(L3���=z�s8O|�D�O �d�O���O`�?Q�䬉�{D^Qk�f�8�R�9�䟤�I��|C�4���'�?y&�i��']�H����=?T:�	p�N�HR�|r�'��OQ��c�i��i�!�GI�!,⍹$@q������I�K�'��d����l���P]��07.ZU��uq��@�	ȟD�'C�7uD���O"���|27Cz5�8������@&&�T~¯�>A��?�O>�O�b�I�ˈ06�LRr�G5�İr�)�D~��p�@���4��89��I�L�Oz=����>���C�J�?P8��@��Ol�$�O����O1��˓D��v��m��QҦ���Ti����"�F��y�F�'���y�T⟐	�O���\��FTۥ�X�q�U��(��n��$�O�5�4�q�F�Ӻ�%����(�<ᷥK�
ͫ��A�]� ��FM�<�)Ot���O����O����O��'V�t�d��"�=�p��M�"ೡ�i��X;f�'b�'�Enzީ�uMS%'��Tcϯz��ɀ"�ڟT�	b�)�Ӣv_~�m�<�'��+cW�� d� N�ջD%�<9ve�
A>��P=�䓉�4���$��.���H�zc aQ������D�O����O���E.Q6:��8�I����8R� ؗ���K*�����	"��=�?�T����ߟ�$��x�g^1K�*���Y�r,"'�>)3�&VǞY F�x̧RƖ�D�8�?�!�����q%d��r�KlϦy���� ������D�O9ǂ�U95�5�;���2���\}�`uӦ�Yq��Od�DMƦ5�?�;���qJ��B�ͱVϗ ����?)��?q��1�M{�O��S���1�*"fҋX���P���8�$��f��)�$�O,��|���?	��?!�6�� 2� I��ƈS��6�\�*O~(n�Fmj���֟4�	@��.A>�a�c�����"�@́��80�T�d�	i��|����?)4�X�{ծG��>W���SFC 1pz|0UM����O�����k���O�ʓN�^8D!�, >��H��1p��?����?����|�.O*�n��u�d�I�y��@TM�z��9��J�7d���ܟD��sy��',��ӟ��iޡ��)"��5ȱ@��E����Yf@�B�iM��O����������<��'��R'pdF�&��|0t9���<	���?)���?����?�����V�P�pta˴V#t	��%�T�2�'2�r�$���:����զ]$������0��U9���f��7�4�	����'ߜ�e�iY����z����t~D�s�g���կ&���V�oy����#�Fpr��_2�ܭ�-N�u����4\�$(:��?���i[�=J0z�C�@Ж$���:��� ���O6��$��?A9��
?p������+N�a���#����0a�3\6�����Jş�h��|rE��-B��`B�%H��4đ�)��'oR�'Y���[��1۴?�N����3;R�Â�W.O��!��N�?���'�����
n}r�'Q�is+��t��ܸV�ŧP�,��'�ҏ;Y`�Ɛ��ʣ'�12�T�~
eY�zl�S�Y� ������<�/Od���O�$�O��d�Ot˧��X)��N�&��E�W�L-wٲ�(`�i}6�ۂV���	�?��HK۟���)�M�;Bs8$��ۃH��X��͑!v`L ��?�L>�'�?I�i����4�yb�32�9��Ȝ�@�<X�b����y������������O����3"P4Q�hĶ����B>�T�d�O\��O ʓa��b�b��'!M�^ަ���V"H��5/&��O�y�'^��'@�'f�f� [�� z�`��D!��O�q��E�{	6M/��	j����O4)x��\�V�TX�A�3R �"OTa�爑SBQ�PK3�zM@ ��O��	�0Ժ���Ob]o�\�Ӽ@�S�S��d#ׇ0	��q[���<9��?���#�� �4��$�2]��)��O�����iV�=��%C�Q<tJB�'d��y\�����?]�	���	��;�b\�h,M�0�ڏ`�&q�5�nyrBg�~a�&)�<�����I�Op��Y	�.g#�;�x�x���crʓ�?������|B��?�,ǵk��m[��#T�]��P%1�h9q�4���W�U����'*�'m�	
I�JQ�E���o��\@CҊ/�����Ɵ���џ��i>	�'r�6E�gAX��M�$	ri�T*�8[�^19G�T^��$U����?��]���IYy2� (} Y�r`�
RT*i�-,U�!��i��I��$)P�OS�<%?�]K������nb��i�:7"4�	^��  �g�63NQ�w�2y�V�;A�M����	Ɵ����'�����|BhW�M:���Óed�Ԋ��/6��'����4(ş}��v����h�w?��s2�&+�|��AY��x��O�O��?���?i��L�>�ʣ͔:bZ�av ҃G��1��?�)Ov)n��@A�	͟ �	b��5\	ئ�.+�>A�t�5��$x}r�'��|ʟX���Q�b�N��gT(Y����u�E����:wi߸}��i>�%�'�6�&����{� ��Sa�-\"��,W�t�I͟���b>m�'հ6��o�
10w�X2=HI��a�V�\c���O��$SǦ��?$Q���ɧ�M��CK�Z��,#���//� ���şpV&���'���҉��?���� �=)��A�72��#�O�����G8Oʓ�?���?��?�����	I?$=&����	/�MS���)��DoڣPF�a�'U����'C�6=��g
+/ 0Q"��2ު!薇�O0�D ��IލU��6�z�x g�+m5H��C�zV�9c��i������O����a�Qyb�'��]������~������>HFr�'���%���0�M�������?!��
{���%�?�|����?�/O���Y}r�'�O����� .�����3fϲ�1s<O6����V�F�ԌQ�Z���S<Y bFM���!宊�x%���E�ڵ��;��^Οp��ɟ����E���'��[��/�.5�aیr�AR�'uF7��+|�4�Y����4�h� +{�!BK�q�x�1OR���O��$?O�6�#?���Z;��)�� 
LH(V�M�A���b�J�,!�H�H>y-O���O8���O��D�O�����e`n]�q�]:�H���'�<��i�f��t�'d��'��Oerb�Y���҅K��O�<h�o�2<X��?�����ŞF�h�r���+�� �R�>!�Z������MS�O����^��~r�|_��re�N<�.py������N�����ӟ�	��Hy2�d�`�Ѵ��O,��gbQ�_zxh�γ1}H�aŢ�O6�n�M�@��	���'e��PR�ڗbȴ�bP�8� ���A0=�Ƙ�@ ,ϛo ��%�J���-��CJ�pb�����L<Se9[X�	ş(������Iğ���y��6�x6#ǯ�j$�@�˙�N��(O,����M�g>9����M{I>iR!�&y�
J�d��!޵�䓫?��|�Q�,�M#�O�T��玺�
��0gK� #�L�Q��D���#�'Z�'x�i>M�	�L�I���0PC�K� ��3d�y�a�	ǟ �'B����-�	ڟЕO� ���h�R]�����Б:�O� �'���'�ɧ���(w�2���F�.?����𯑷5�^�r����!$B7�Bgy�OU����P@Ԁ��/*c�i���'{��y��?����?��|���?�)O(�m�K��3/&u>��*f,Ђ
8���gf�ٟD����MH>��Y��	����)O?__�T���L3�ʌˤ�ٟ,���S�@o�<Q��>�	�?��'^~ V�Y;����q#I��9�'��͟��Iџ��I�	���Z{�a	�;I��(��']�7m;)1$���Ol�-�9O@�oz���n�f0�@�����x��k�ޟp��d�)�)%n��l��<�P��fcЅ��/1�[6��<q6FV�ZK���@8����d�O^�$���|�����^a"Q��,
�R�$��OX���O��^��)K<0���'b5S��� z_���E莕;b�O>��'c��'W�'	t2�%�^H�7�p8�]������ !7�|�rc>�	r�O�D�5-_$�3bo�,�:�z1�F�z!��ڠ<��X��ݰ@���+ɾDb����ş��7��O������?ͻ#�X����'?�xU�äz,�Γ�?���?1�cC-�M��OB�2)���d�<C���>V���AK֚B/�'��K�'R�ɋՂ� $\e��`�a��O �I�� ��OB�D$�ӝ�^h���Z�<��*ۭɶ���O~���Oj�O1��m��e��G��J��V�(�ޠ�0Јs��7�ky�ŕi�D�������$Ī���F���t��t-��@�`���O�d�Ond�3�r|�ʓ��i^�^%��>j���/��p��[��[1^b�m���D�<���Lg����0�'Ed8���Z�9ve�9J��(�7È$��f;O��$����X��<$����)���IF�s.�x%O�Q�r`��?I��?a��?a���O����F5["99s�ʇd	$�B�'���'��D߼��)��$��ѩO�c���8�d�W�Xɣ%��@�	�H�i>1�0��ѦY�' lt���B����O�c����d��g*���䓲�d�O��D�O��$J��������y!�G�=F ����OZ�Sڛ�Tl���'�rY>�Յݾ�©��֤b��)X*?��W�(�IΟ�'��  �|9�ӽ{�(�����dǂ� �ė�.�����A~�O,I�	��b���yR��M�=ZjI=vA.]��Z
96��'��'�ʟ��R0��<�"�i�M�EJ t,�Z(O΀���]��"�M;N>��'y�	Ο�Ò��p:pq��̊ �L���������Iw�vm��<a��|�Xt��?��'�j\���o�����Ə`���'��I����P�I��$��P����$1̵��� �����!2�7�� |Q�#���O��D�����O2��J��wΔz6O֖#���$ˊy��	��'sқ|�O��'h�P�5�i�����\�p�荒+x���PN��x��E
�� ���֓O���?��.��#�퍻O�=��D� A��?Y���?�,O0�oڈC����'Djȝ2 �����!�BT[�M �"��O�5�'@��'��'�Ʊ{���A�����K�O"���!�7�Ta�S�	F���O��FL�84��,��2��굉�O.�D�O�d�O��}���^dT�t�5���j֧�8!Y셊�W���\�Z��'��6�4�iޥ ���傑J +2h����q� �I����;M>nZt~2Ȋ<�i�g�? ��cr���.�� Jti�/$A� ��2�D�<����?����?���?�Ef֮:޾8y��%>V\I��\	��d즱���J۟��	ޟ0'?��I�w�`��EV+$@�`��
�,�O����O��O1��$;`�0/F�9�'�>��b�/F�Q�̈Q#h�<���>�H�� �䓒�䛣4�VD:�Ԭit��l�p{���?����?�'��D�릭R�J���c��E2���ʞ{`qP�e��0 ܴ��'듍?���?ٰh_1�hJ�C�	#-����eJ�um Q�ش��dK�>i((�	����:o"��*��ݳ�zX2w5O��D�O��D�O���O��?)"!� lt9��t+��; 'Kџ ��՟p �4^x`ͧ�?1��i�'ČuI��5j�y�V��
((|R�'��O�����iu�I1cs�9�͵J=��r�N�auJ8�a�ɠAc��6�$�<ͧ�?���?qQ�ڸ0�x�r�)M�9�6���?����$����agH�ԟ���\�O�h��$H���j����a�����ӭOn�D�O�O���yNp�@�_(bj�Q��^�DA��䄞mTU#� 3?ͧ5
��� &��e��ث��� $m���T�
�Ii�<����?����?)�Ş��ğ��q��$��"��ӑɌ��y�D�8 -�'�$6)�������OX�!��
2?Rx[f�S�l} ��ъ�OT��ƌ$f6:?Y��ďߞ�ryB�\q����܇#��۔u��d�<q���?���?Q���?�)�xM*�"���*�H� 5`���g�����$�埀�	۟�&?��ɞ�M�;P���a���QN�A�@��8~:���?9M>�|�5IE��M�'��m`F�8gL���
E�q�'ƈ�r����hQd�|�P��Ꟁ��"�j�f���B	I�:�Б��۟�����jC\Xy2,��`�aA���D�O�̐V䈅���o�`Z�W*�O���?	c\�����%�d��MȊ��x�g^����@Je���ɓ'%�jE ލ
�E�'M�������:��'v�!(���	�#�n	 ;�4A��'4�'�R�'c�>��I�p�NI`�C �x_T�14hRሐ��
�McQA�*��D�����?�;���?j}rd�7WI��̓�?q��?1f&��M��O�7]K��� =A�@<[S�	n���Xpkx�n�XN>Q(O��D�O��d�O��d�O]��lԵq������#��6�<1��id�\���'���'��O�үB+s�Ir%\RI�v��|�4��?I����Ş5<Dej��� rRPh�ca���x��f�8z�(�`-O
�2���?��<�d�<�(�3K�เ�E�͌ ��Ş��?���?���?�'���F���Qh�����D���r��C��|�Ta34N�̟`cش��'���?���?i��(2�!��i	���2M�>��)��4���������Ol�O��Fܷcr��礂�9���ӳ#A�y2�'|��'	��'A���U�y���ea̸��Ē���w�T���O��$O��h�Iv>9�	�M�K>)tEϵ:):�P�H��%~M��ia̓�?�*O��Z�yӮ�BW�\c�T�LX�B��.���l
�4D@�$լ�����O����O��d�)2� �E�I��<�f���*�����O�ʓF�v������'lBR>�h>z����b([4˪}D<?�wU�|�I��'������S�A<S��@�#IE�n��Y�q�+@�B��F�H/��4�*=3��&��Ox4uh��G�\Mi�̗�P��e9W.�OH�d�O�d�O1�F����ڪW�DqT�Z(0�(�s�ɭnl�s��'�Ҩ`ӄ�XR�OB�$�K�|@gK�pFN@Q��V�R���O�`��GkӦ�Ӻ�e��7��Ͽ<�$A��Mè��w�܄��u����<�,Ot�d�OH�d�O����O�˧>b�J���6x��:V�\� �iyj�ˀ�'V�')�OUr�q���<i�z��P�U�,�(�T��u�j���O\�O1�Dٺ�}��扨'9� ���ߐ),����ꖵ�l�I��Y���O>�O���?Y�0g��(��Q+\�J�V�����?	��?)OplZ}{|��ɟ���C��r�/PJ �b�)��.�ȴ�?i#U���	ʟ�&���F�4U�āѷ��q¨��B<?�/�`}���"G���'j��œ�?�3D�n��18�@	�J��S����?a��?q���?aI~�B[�|���$Z���'B����#�a>2M��Vg���T�>��'tb�'��I���7�ְ�AeX F���QI^0Di�	㟸�	��\����ϓ���L^5En�mM-+^! M4��U#���y*2�'�P�'�b�'=��'w2�'�b��\>zZ�j��QXT�KR��1�4=ތ����?����'�?!q��;Vn �R�;!?�)�v�ˏh������t�)�[Ov�p��� g%��*�[&kL�q�gP+7�"(�'C��0чޟ,�0�|�W��c�a!RO��B枥�������	������hyrhg�.��f�O~�dĜ9P.�Um�&f�*9�&7O�o�g��v�����T��ퟐ�r�XJ0����6d���{VnL3+�^%nZM~�ٲ1+�PF��w^\=�#μ3�Ԙ����JkBlj������(�	���	ğ���덺q�|�
���5�	ӱh)�?1���?��i�a(�O���h� �O���A�3;Iƌ������<(���*���O��4��Q�7&y�j�+��P� ��v���aWhUb��N�A�lp�͊��~ҟ|RU���	П���؟�*�&]	:C���3Ö�p�� �g��H��Ly�z�8��.�<�����^m�hjW��m���rW&Ǟq�ɸ��$�O���/��?��%搟b������iu/J�ZL��v �	��FA?	M>g/ �(�QDY�R�D|C��
��?���?q��?�|j,O�io�(c������4D�����BJ<�┥ΟH�I8�M���o�>���a$6��	��D����6�
H��?����M��Ond�Ǉ¼��O>�Y3���aT� �˟�V�
�'�������ܟ�IƟ�����ӽS|��oD6�Z�P��2J��4$j� ��?	����i�Ol�D�O�n�7�6C��5|�L�*rM�[A��d�O
�O�i�O��d�"R��7�}���# �2 ���C���(u�j�
b-g�,����$���6��<�'�?A"aG���%���ͣ|���A���?��?������������T��ٟ�"f M.h��W���J̾��j�o�\�I��	J��I�I+r�$�:�O
�n�j�V�I
U#S�M�d��4�Fg?�����<ː�\�����p\�	r���?����?��?�O5b�9E�'�K�2*v���q+��,�����z��$��yچ�<��iB�'(�w&&��dd@�D�0	�&ڳ�@j�'�R�'Y���]���3Ox�M�}	���'r�"44�H�ʩA�CX%v(ͣ�"���<ͧ�?y���?���?��̸E;� ��Dʆ١b��z����M;�eH�����O�"|�$�*M�0I �D�c��L�����D�O��i�ɧ�O1�9�BO'}��y�%i~���� �2}�\��O��(���?�t%2���<�Ջ"-�	�%H�i��\�(A��?q��?q���?ͧ��DW�+�V�@8`��"PN@��P@�}+2.�ğtz�4��'�@��?����?�"���;֦PQmB'?F�`,�:!��}8޴�����M��؟Ғ�����]�5{�-6�����!s���O4}����OH���O����O1�p����	 b� *p�T�S��MY�(�O����O.Uo92^I��П��Id�I/i���r�ߐTd��F�F�v��&���	������+C5o��<��^�8I9T�ڂY�r��C8��\xs,R�F��d:�����9O8�X&���[D4��c-��?u�M��ɿ�?��kП`�I��4�O$6 �U�� 4Flc6�ʞ8��O^��'wB�'7ɧ��UV�r�в�T�_�)p�Z# N^�`)Ίc46�Wly�O`T���k�܀��U�EF��UeF���EX��?����?Y�Ş��d���� E�r��jT�P$����%f8!�D���J�4��'�L��?y��4�����u���a.��?��X�F�!ڴ��dưPC<��Ot�	9�<Lb��ʬ+6�T�⡒=bz�,��L>턼Z�BJ %
iCg��/0��#�Ϧ?̴2c��3~BČ�SN�{��fC�x����4�z�@sA��v�$�ė<�P1Ѣ�A#:�#>i�O�5�P�a�h�"| 8�%ɏ:.M�X���8�~xbW��(J��xC�狊!� P!j�,`9p��ʈ0:e���G���G��iC����`�£Lh���T���8;��� Jr�jťːS)�)¢���\��ũX@�\a�b&dS�M�!zF0����T�j%�Ħ��ɟ���?՛�OD��Vc�	M�Zy`��F�:z�@�i<2�(`�'��'�3?��	�TH���@��]H��A�@պi�R�'��`\���d�O��	�\H���Ǣh%eHDJ�� ��}b��',I�')��'w�'Z�z�3�1-WK--��y�i��*[�-��ꓣ��Ox�Ok��lV� dED�l]t�)�@��	��3`t�l'���I����	qy"J�} &���	��$������m��M؇�>(O��d9���O��$�#ٖ��U/OZ؀��T<R� �[���O����O��ǂ�'>�^��h��M�Bu��c��$��(1C�i��柨%�h��柠��A�Y?�0��b �p'��yTtc�BG}�'JR�'�	
�f�#��"��-����-G|}��@&�	g8��n�ßh$����ß��$�R�	��a �T�a�,x��i���n�Ɵ���Ey��p��꧉?���bS�g�D�^�n9^IG [W���3�x�'��`E3{���|bן��hrI��W䩳gOƀ("�([�iL�`Wh
ٴ�?A��?1�')"�i��f��|&e�[�t�&��@eӮ�D�O�l
0�OȒO&�>�V�*X�AP�#T���(a�d�:�k6�����	���I�?Ѡ�O
�R������.�8�Qb	�+R ��i�x`z6�D(���Hh��>����ͅ�; ���'hٌ�M���?Y��c��)��]��'F��O���e�9���Ӆ=��ar�d���P�O����Ol�Ė�X�rh o��D���� ��{���mΟl��N����<�������p@߅T�nH�T
�pt�U���G}hʠCT�'�R�'uR]�	GZ��3K�7p�=��g%|6`��O�ʓ�?�O>q��?)"g� ��`�+�<Y,Ih��>�B�H>����?�����x��u�'"XK�=)�P���l�61-�~����?�H>����?�B� B}�A�C@�ِT��-�"q�p�ø����O���O��G�`���R?��I�CJ��;^�(�H0*�%�
�U�۴�?�J>���?1N�ĸ�� qe�T�d��K70�6@jǷi��'��ɹȈ�K|�����N��>����NЮQS��%�,�'\��'}��yZw$dYb��ĒC�ܸ 0���d��|۴���D�>4�(o���I�O��ITr~R%Ï|~$�CbL\$i���(�M�)O����Oa%>m%?7��Lz���Ŝ7v��0�*3��F�ü��6m�ON���O���NV�i>�`2MC|��8�"��U� ��P=�M����?�����S��'�b�7f��ш5��@�H����DE�6��O����O,���_�i>Y��k?q4D'2<�s�ؙT펙��iSڦ-�	F�ɭ�������a?Y��D=���Z;�]��$�ڦ}���{�T]�'��꧉�'�0�b�%b�@�㇛�p�p]�m'�$Ј$1Op�$�<��S�hm�SbN�e����c+״@:½���ɶ��$�O
��+�	�p���Z#팅y��l���T02�@lZ�'�Zb�l��Cy"�'*a��֟б��ǐ�	�(��"Ϛ��!�b�iir�'�O,�d�<a�����q�s�0w�dx���%�<�"�D�O���?y�����i�OZؙ!o�=�5�Ŋ��hJ������Ħi�?�����dP��'�Nx���(,`L`�v�1epvt�ش�?�����䚒u&lt&>���?��:'��1�ߦq���`���J�rO�˓�?1����<��*�������TRd�c҆!U���'�r+ܚ�R�'���'G�4Z��	��EKS$��y�|�Qb�5bY*6��O��oDR�DxJ|�s̖2gR�P�l�˨�z�,������,��ӟ����?՗��閲~���q��:yt��k�HE�3�x�'�(4X���I�On��7���<�>	�ã�Y�,����������8��t\�CO<�'�?���2θչ�"�=p�Z�Br�ƼT%d�k��i��'I�I ��)�|����~� �A�>�,Li�R%��۴�?IP,�����X�������ЊJwYD}3��ȁc$x�'�t�� ?)���?����䑎?��ݓ��^�/�j�c��:x���
}�	����H�IqyZw&^�BO7tC�-c��Ԇlm@�4�?�/O2���O���<��hD���i�#�`����> ����H�Q���韄�	����'�V>5�ɚK����U���dvb�#g���XUF�j�O~���O���?y�Q�����O�����V��8y�oڸi�Z�Qǫ
Ȧe�?����U�'���z���3!ײ��a�Ι�8��4�?�����kĈ��O�b�'��땧PX��UM��X�t@I��Ĩv���?	���?aa��<�N>��OVBB�޷ ����a՗�>�ڴ��ţ=���lZ� ������Ӂ����i* ��G�̸��D'�0ꢽi��'�ڔQ�'^�'�q���q@H ,�r$zJ�-�����i�X�
��q�d�d�O����0�'[�B��M��ۧa���Ǩ~!F��M��(��<�����:��ߟhE�����v�!x�$�A!��M+��?)��x�����X�ȕ'���O�8�1*�> n�(+O�m�`���i?�W�<peeo��'�?!����4`D�� T�r$�VpD�`�g�3�M���6�<�Y�Z��'�Y�S�w��a隭CW�J )�:e\	�'*@�'���'8B�'��X�dS���D�R��/;n4�R�G�l�  �Oh��?�(Oj���O���
�%��P�b��*,��N��)=��xw>O���?q���?�+O�S��E�|jUÄ�l�@Jք�`�d�'G����'��V����ԟ��ɰ����
e��������7,�� �ҍ�ߴ�?����?����ެc�X��O*"�Ǵ)1��ZFXҵ��^�d$�7�O�ʓ�?)���?-�����ܴ?��(���-O�(�l�;�oןL��By�&��b�v꧁?���C3m����GÆ�C�@�[�IƟ<�I��PZ�)s�x�Icy�Пle�V÷v�)��Iϝ��r�i���5#��Z�4�?���?y��"�i�U��"E�Dv�P��_C\H �d�R���O�2f<O����yb����J�@�C�/�5z��{���,s�F�K>z��7��O��$�O��	~}�T�����.d� Cݒ5�\�a���3�M{pJ��<a�����-����`�� )9�,H0e��;1���R��6�M#��?y����Z�H�'e�O$ͫ�@�#��℃ Q���i}�I͟D�%�~��'�?9���?��OȺ}�� v���6X�HӒ�B�^��F�'|^�9Vi�>�-O:�İ<����"�5��4��ˊ��T!���U[}"䗃�y�Z���ݟ���kyB����Ba��j�0��C������>Y(OX�D�<Q��?i�����f^ry�pk��z���Ҥ��</O����O<�$�<i!S�]N��ƀ)��-aP��8v�n$��	�yI��U�4�	Dy��'��'x8�R�'Y<A*
�7M!�qPr�P(W���r�{�B��O����OL˓|_�,yUX?��i��r���n��Hb�ju�
�Ѧ`tӸ��<����?���4͓��i�dQ�0��2)����ߗ7� ���4�?�����$K�_��]�Og��'��D���kj>��V�X\��yW��Hc�>!���?���
C����9O����o� ���ɃLa��QЬDn7�<��'�2~��'���';�ĩ�>��;�T�[�H�5`�h1�CϛV2�m�����u�l�	矤�'rq�� �A;�@��
��gG�CfD�
1�ifLͨG�pӄ���O@������'���/�f�e��0K]^�c8&�a�ܴo�&�ϓ�?/O�?��	�XF\� �^���K�-H�C* 8��4�?����?��bNz�	Ny��'%��̗�:(�L]�R��Т�*ߍPX��'���'~$�������Ot���O0�k�'�(s�n��U�J��KЦA���6��mɨO�ʓ�?A*O�������*�*�h��@���h��R�0��B}���	ܟ�	���Nyb���@X
.�C�><���BB�qg�>�,O����<���?)��k]{M(s��`%.�3n'��"��<)/O���Ov���<!����U����&<�(��cA�h���a�*��FQ����lyR�'��'a  ��'x$�R��E�����92$���`Ӯ���O��D�O�k zu �Z?��5$��	�+q�
Q�m3**��4�?�-O���O����_��$�|n�?r 8�F3h>*�Zw#Ly��6�O���<��L�M��͟��	�?�� ��7f��xE["�D�pB��)����O�$�Or=8�<OT��<!�O�`�Q�\�<!f9�gZtW��X�4���U�7�ޭoZ����	�\������t�w�����P�� �'�L`���i�B�'�R=c�'>�_���}�Ul�f��Փ�/Y�{$�A�R̦�X���M����?����zV_�ȗ'�01a	\<��%;E,�U��*a�!#W5O��ĥ<���t�'����+82L,��T<M��mr���p�D�O��DBa/F��'2��ܟ���j���H�+y��E�O�:P mnZ� �	���㒨l��'�?I��?)��k!ܽ��0k�.�ApDPk��v�'�I ��>�.OR���<����l�we�ݣ$,��P����a}BcW��y��'���'c"�'���(E��� M:��c� ����&� ��ē�?9�����?1�Kd@5�.)&�S$�V�3}< ("Y@��?����?�*O^}Y����|�d�uR)ISP�c�����n}��'�2�|��'�B�1u�D\>��͈�hܖ`F8a���-��	������'YX�Ғ�(�	��
��@3tPg%��~���irӘ�D$�d�O���F�i���5}�j�6��q	��S#kϔhP"���MK���?a,OT��[�ǟ��6L���,ĥ_9Vy�U�lw�II<����?ylN�<�L>��Ocbp8g��	V�9k�.�9��ش��d��^Ȍ�m������OV���\~A�,JD����L�>��p�[�M���?1獄�?AH>A���Ɯl���rLlR��C���M󵯚�OP���'���'�tf*�ɝlR���)o��}�&]�N#|���4F�Șϓ����O��@=�h��Q��'[��%`@D�=��6m�OH���O�q:�gY�I���\?)vM�/�H�(e�(Ʀha�.[Ҧ�$��X��x��?���?�1�I!Za��
���_��͸U�#u3��'�Ęp�4��O���*���Fp���06V�@aL�6���k�Q�X���g���'s��'�O�̥��C�*��ƈ��)"$@_5N�D�H<y��?�H>q���?�V剁ri�A��ܦ745�w� -}P �����O*���OT�����7���b̑ (�0 ��Ɉc(���W�T���X'�P���h��w�� �']��]!�����6�Z=��L�'P��'��U�|+���ħ�V�)�˜�t.u!J�_@�a�i��|��'��J0v!қ>��(շ��5H_�s]Z�ٴL��M����?)O)��(w�Sٟ�s�� eI�=0��D�AB�c0]0d�3��Fy��'��O뮜#6bAᘳ]< �0�	
��v�')"k�6��'B��'��DR���{���ӗ)�jl~ِ��|<:7��O0�K��DxJ|�%d[KFT���u�hbƞ�=9T@	8�M���?����BQU�(�O�z0Q���-!���ɓ�K��H�Gq���d7��䓺?�BK�#Y���zd̆�K�rtK4�P!��v�'��I:JѸ@�'��	� �<��ak��I�+�m���U:�I�ħ�?����?9�-� Ҡ��ě!I�N%�1- �{K�V�'��):X��[��6�2�$&Ύ��so��05���䇜,/b�'���f&0?���?������B�)[��b��-C��a ��)H-j�ӣ�Wn��T�I��?���k ,|��d@�d���1��I���<�<9��?	��?A�O
6pH�O3��ϸ�	��ҧ6i�[۴�?	��?yL>�����%f���L�o&E�T�CW�(�R�Y	��$�Od���OH�>jM|��oN�B��Α,|��<
3jZ?U��F�'Q�'�R�'ɾ-��}Rܔ$\��ZR��,axn�Y1Z��MC���?��O"��K)��O��iH#��e0oׄ8��HR�	�&��Iӟ����>���FU	Qߐ���b�lޙ7N��M#�O"1pG%|�е�O6��O���O��Ӆ��� ��c���] ޔm�������G�\#<���'IJ�Ur�B˳J�X���?р�߉�M����?������x�' (�3����xq1�
A.*����+hӚt;q�)�'�?	�A�#wMX�bq�A3��E*3����F�'-R�'E���1���OH����x���h*�DAb�X�M���o$�I�|�c�X�����I΀ ��T*�9R��'��&�hp��i�2�[�~�c���IG�i���=����Qm��:�u���>!�aWP̓�?����?��O��h�n<�<�Cv�Y�3�h�K]6�c�`�IA��ğd�I4}�l�ڧ�?
�}ӵ�W���%xf�8�I^���b�˚#F^�E�to���Xs1�^�()��"(ͱ�y�`�>S�&%H � �@�k�����'���S��ێ[汪����wW&( Ek�>������.͎$H�	��'�(�8�
@9l��mJ��ȹ����	!�a�DX%:�^�	2����i�S|Q�%BkGkH���wq(����'dc0�gV�m�A�Wй=��25i��=�m(S���P�e�3E�_��Z��7H��Ct�
 K6��rWʉ- ������?1d��C�@XrÌ	?&z�k���wYJ�S@���ۘLl"L�ԥKۈ�*�����	<|�d��V��'���شr>`�V��^���`��uĆ�l���P%1�>q���'��iIs�'h2��џ,Q�7r���!�
ʐNN袃 5D�����"�D��c��)m7 "3.O��FzB�n3DAb!jôOB<܃3��?���'E��'yb$8B-N��"�'~���y7�M�&�cuʚIhDc�T 3-�X��IN�bYn���/|y��3"�|�o�y�*}��2�y�q*�3y��l��ޜ���dR�#������L>ņ�x֢Kb�	O>L�'b��?�Or� ���4퉖=J���;8�AR�_>�\B�ɼ#�J� L��4"��4GJ�%đ��'����0��j��M�,
�d�Ʈ.Ey<Q+��+H�����OF���O��;�?!����DH��(��t����)F���pfʹ]����1F?>�\�k'�'lOF}I�/D�YgM��`�,jf4d��꒔,������܌?m:I��I>������jZ����*�$��O|�d9ړ��'�N !�,2{��`<S�<��	�'/��fͯ7���f��0��y��>�)O��
��]}��'[�А�πRZ��Q& R�	��!��'j"�!e��'a�	�h+N�S��^#/����F �h2�쉯GA2(�2�ý+����I&�̹��.F%�l,j�'@�9��F�C� ��kZ�n����Ǔ2Q���t�'��1n�� w�LP�D�$6UZ�ҋy��'
$�˳�d�fxa�0�*��'��7�K�u1 ���OSS堬�"�>V�$�<I�M��A5���'��\>�R��
ԟ�*���13G�p��o��z�ퟜ�I�  �9��4������#��WՂ�s"�͏��)�N!}� ��(y ��A�-]��s�-�D �e�J~��&mY��P��2�Y��B��Իecb�'�7m�O&�?$k�+�c���/1����kd��'��V����C�p8��M�'��9*�����p����޴�?���i��k[4<�óC_�?���у ��듌?q�IR ���?����?�׿k����5tV����E�直Q��S�A�>�5��

��1�|&�|�l�nຐ"t�^�:����,"���X���#���W�q��'�$���c�VY�E�R��p�U�'"�ɭq�N�4�,�=їm� �T���N;b� ���m�<�F�E�?�i@W`[�$��\hQ �h~rA?�S�$V��3U&X�K��AX�G�	/����i0���j`��ǟ��I��@�	:�u'�'0�;���2���6KK��k	_�GT:�jC+��U� �FB5�O�L�5��^���m�?#$-Â*ƠKq����&'�O���7Q!e��T�͕+��q�Vt�"�'���'��I����?B����\���F鼹P!nO�<�"�_!]ߘ5�e��
x�X@���P̓��uy'G�:ꓥ?a��\�a�b�1�}H$ʴ�?A�Z�9����?��O^�|�&��*W�I���>A�mZ#4�G')$ l�S�#O�1q7���l�\�h�u?QѭʳTS�����s�[�N�I8�P9���Ob�$�<�c��bъ��'(�����p~̓��=��HS�}�v��a盺u�����	v<�i��`���48�H�����3YT��*�'��	,ƞY�O����|"�I��?IgH^��8�-ڈ@(���-�?��y�dE!� �.�S���*���'y��Ce�_)І�_�ft�@�O���S�\�^�$����I�#}�ꎗN�xs�m]3W�(1CQc��f��'��>U�	�h�
	��	�~�R�ԧ���0�Ɠ�% ��E`�Q!�T������HO� 1�����Y%W�V5�)�ĦU���<�I�kgbAUm��I����	��u��*
Lر*O�7t]Y�S1O��8��'��,*G, ZF�T�S 4��{�-����<���XO$��e-�C[�����<ܘ'\����S�g�'����AI� ���\��C�)� P���C�ܠP�l��������Z����n}P�&�N����8���x-�$8��?v�h�Iݟ�IƟ�^wV��'"�H�gG�x(Wܢ���R	C�̂#OD��4�Q�J�t��TC�u�� V�	�0!�тJ�:��hۑC,�40g� ���y:��'&�';��'*�O�a�.	-��q���s�B�"O�@+W.H ��Ӂ�Ra�P`D�d�x}��i>y;�ϩ!�B J���7�VqZd/:D����Y��5ؑ�ӑH~l {�6D��x�@V�S<d�K��̄1�^�(1g:D��Y�	+
�]k�I�*@ST,9D�4c�oV$ @���C�h�ay��8D��0`�_(v~<5pA�6lܙ�s 6D�Hڔ	Z�4��0aߑ
��A��6D����,`<��I] `��!��(D������>g	 I�)��t��IU 'D�ț���4����Y�d�($D�\���G����9��\�����"D�\"��1$Iu2uDC"lD��b�l%D��!��M��Xi�'p�Y@V� D� 0Eb�>s 51#�*�$Y�d�9D�@a����#�|���T�l�H-���)D�p`��>�`�; m�U���[��2D�X�U�C�Dp�Q��M�f��͐��2D��ᄅƷ|�>��D�K� ]��Zrh6D�4 ��N�}�2	�H2��H�3D� *��h�Xd{���1Ί9u*2D�� ���;Z�Y����~U���0D��1��L�g�@] �IŤgXI�4�"D��ꅨI�M QTK�.Dm�Պ�"4D�l�sdōjnBa���o|,��k0D�,BQ�
r*��(���-����,D�|��
�/o4����`��� e*D�HK�)�T ]sF�R��إ�)D��t�Q�v�ֈA��D6.��e��&D� ����r��P�G����Ub�2D���IN[Ґ)�sJ�\�8`/D�(�0��E��#'�F���,x�(D��iӭ�=��3s��i~�4�4D����C1`($aE)"l�|Xx�#3D�(�do��B/����^.��3p�$D����N�;py�-��a��h��ms!�!D���u��!n����O� z��)SQ	 D�`
��V��a�p�!m"��;1E>D�D���Ä.jRģVc�'`v�ӧ=D����bB�4S��q�EL.1n��$?D����Yp�x��y���i�e
$�y' 7�yp��Q:p�����`C��y"�ӊ1�x�9����U��D��S?�y7 Q4�� �O�n�QR`��yB���N�n��S%�Tx<%����yR��#㮉*3�ղҽ32�U��yR��6Gnޭ���v6^���C��y2`̝W2�p�U�@"Œ� 啱�ybl<,!�,B�ۊk� �˵n�"�yB�E	1cx�� ��c���2&"ʅ�yBgQ�4�(�`�&ۑ\�]ؕ'K;�yҠ�.FJ|Z�M�O�\U	_��y(M�?l�t"���@�ɹ�(G��y�(Y&��9be��Ѝ$+��yr�R5 :��FA�C���x��G�y�b�&T�{�DĮ?dP�Wϣ�yb��o��aI��	�I�&e�!��;�yN$F�3�U#F� �R��y
� ���3�O�g�<k��G12@��"O~E:d$FZ���K�O� ��H�"O��Iah�����w�@41�HD��"O�(H�A�D!"��e��O��tQ`"O�X�W/�./$=����k�t��t"O��)�P5>�$T�O�7���q"O�1Ru�W(��!�md|e�"O����#�!��,�TcvPA�"O��(�J�U[XQ��D�z@��[�>A"l�D��Ho9��i�?��rv�<#�L�|�T���ϊuj�����-����s�OM�L����|h�b�\��4AԌۄ	�N�"~nZ*�D4@C'�p� 5��3��>1�HE�<$@1��4Ě�S��B�jU��:��)����+yrߓI�dX�K0P��� ��Y��`��[���Z�+��S��$�a�G�-�Y·���L��l(]"��yǬ=D�xK����p����@����zRF;}�@�L=2]qu��/�v5�FP����~�����
T�<���8�H�h��ҵ*ߑCXa�s�ص$�ک��-���U�ֈ�}/�|	f��_��,O��z�-(�s����V�\PU*¬V�r������	�f�(��Sb=:����A�E�A�=�X��Bم+r�X��ÊŗPJ.]�D�S8�xkR�
e�t5��-�;��{�A��&��aSrGGc?�OԱ�?��t��k��4jj��C�J&C R!����frh�������O J�$�#+˘ȣ%>�Zu��Ò	��5��Z����\�~����H3A�V���Sސ�g�$-�}�%�
?p�2�i[`�� kPcO���'h�!iTk_�J������S�4�S�O�8c%��j<�qe��Ǝ��F��!r�Ȍ��g'���:��QCn~+8�1�`-#��D��=��y#'k ��1�#�_$��g22�Ce� ��9��FB�0V�lt`d_ 	��H1]w �	:!��F1�2'�W5��h�'����a3m�RHrQ��V��8���U 2 "F�Ƅ)'T����1l$���)Ψ���)B�Ȱ+ L�H���VD�>Do6�8�H�h@ "�Ȏ<!ń�A�n#ړM��!!J%PH)�;<x|�f�J�+�F@;���?&���O�Af.D���C�p��c
A�g?�5�>|�z�#☗rH1jQ�i�$0Q�3�ɦ)u$1 U���}��x�%��V�.�C�� �Fϖ}@���H�(r�f�I��<,tlؕL̴�#�OX�ڴ#�t��hCb�,��C�'m v+��8,͉�Eɕv�ny���! 7���Ǌ��xޔ]kK<Q��Y�<)���=�~r`��F��k�'r��4��c��~rHM!xY����A�^��	9�J@���4�:�7&��2��C�Oֶ�	�E2>�NO,m�
ЛD<Н��@:�{�p�d-4�p��3��6�teH��VBA�
֝9k��<�ƽy��iAG漫n�';}� Y�$!�9Yp(T�
��y�I>Yr,\H�OK��I�������&��a#\!a�.,:�yb+L!.-8` �*�`@�`�И'�v	�f��&�L!�� -Εp�4!���ێ}2C�gl��ja�-h��i�t���';�MH��IC��(à��}Y�P�rظT,�52�g�Lz ۓmU��p7G�7J�	Ӗ@��?�t�JrF��pp�@��@B��;��G�sR��'��hI����<k4٩��%qaj0ZT#E��yb��'jgX�B�A�&����rE�%,6�|�r�E	$���!�+��'��#�k�\��w&�y�Vhγp�L����а5X�q��7���c�
�B5(�V"oX9��a�~��c�8��i�'>��*P�B hd"��%扶o�acA�� ��L3w��"'`,�>�B�
Rl�B� �3�,p΂�/��T���	,�v�V�(���ӧO(:����a�^p`�V�,LO�"׭��F3D�1Ea���;�']�9+�K?�v�*ufK�sM� ӭ���D�3A��_7Uj ���)��X���@���-d!��C�8�A�)#z��ʣe���na2@��:T�P�r"�ά8R1OP�p&�ތx�&yx�4�):��[+����X� �P��'�D��"��,�@���X�\�:�٤'�X�x��<٠/�5Ux��tT�j͎t�q��̓>ER-2��>A�|�wfA5U⼄D|үY�A�vԙ#�̵/{�-��B��P���Xd	��TҒ1�࣋{y�i;!jݕt�XI!%	#I��鳓/���?I�������x��) ��9�>hI$��s}���b� Vxx��'瓶2�@9��O��C�|̓�޹j�mY�/@@�ɖ��G��q���fX�T�?E���D5�H���@Q�2rHIVC�A�NUAE��)��)��i>咖���e�杞dG<{���.O1���C-Q|���[;<�B���� H����c��d���T�'�hi
�*6�'44�p��Dh�j-K�$"<�AS>�DU�8�h��Cl(�zT�a�?�T����D�Q�C��8LЎ���-҈��i� X����hD�0�GefI!��!L$����9`����̧^�� �L�0�L��V�{H�}��?��?�����Q��=`�g�n̪��DdD��@ 6ҼD��@y���1��� Ԕ}KR�{�� �7_i���<@b@L��)� �,I�dC&w�v�a�A��,�5@D�ɴe��m����0鑗��F�M�����6�U���csÂ�ÈB䉲F��ɰ��Y#L�0X`D��z�d��-vL`@��R�(�)#KI�)rd�}Zt�R�t�0t�g��Y�$I�v��}�<9���|Zd ����r�lX��ώ�1ʣM����H��		���fhSp�n��D��J���T�C.J�"��-�.Ȉ���v�h�H�D�O�f��6ᒬH��9c��Fi��t�e�5S�rlZ�/_4f2�ʀ� �\����6犉#�6�ۓ':s�Td��:X��]cTe���	�)d~��"O�aL;8�:ɘs�ўD6F8�`�i���b۠��s�/��Q�(�Af�(�k�\�����	lD�x�"��N!�5B�DEI�mҶTO��K��Li�
X!pGD��lI�,��4Ε�BT?��2�d;����G��҈Z���(�z��קt"0���Yl�Z�,N�tP��̊Z��#�.C�u��P��L^'%�έ�ߓF�q�ś0�^��
L�8���<��\�?��ݹe�
�}pP�7�P��O����J�/P�9sU��]@8XS�'6�d��%c�\p�uc��S�si�6�X0R���ȈL�����)�<���ǡ�)\T9��l�<3��4�s"O��6GU8[;@��t�3 � )�PG�9m{D��1ݙW�8T�L���2OE��㟼���S���qT�J�3���C�*LO�9�u-ù�⍣D�M�g]\�)#ɦmm�����[#n�+�����M�R.�<:7���ɺr�Hag��j[^�#%�b��+\��X%�ݠT��)���,.�p�� ȸ�u���=\tw��6!D�124%�+�y��G��X�%� [L������P�r�M_�5�I�͔�n�,�B�C䒟<�Z�w[�`6F��
�x�)a� �1��'?�dB�/�+�Bt��˛�/��"pI7�9�!%���͘%���<���Ѝ\A���ԓWo9�$�@��$!��ͫg�N1�'���	��W%+@Z ��������'f2 ����K>:���#ɂ9z���y�/Ѳx����a*@�OU�(�̈́_J˖C,���A�'t4�&��}��7M	/ Z�� PM^1���O4���3?i��]�J9.$Ar,؏d�� 0��v�<ၤ9f������ʀ̊�Ѧ~��� �`A�i>.���I�j��g���)�KX(eF�ի�n>&�P,� C���Z/�!���:"�����6B�5H�`�!�ս!�^=B�Ɣ3 Kb�<A�ʍD��Y���0v�E�	�.m��C�0B�B�	�,'1I#��.Ű�cr�EI�8����	�Tr�fR�PG��OPK`gԷG8�����E�,)�5�Q"O,䊒F��
o���+R�\+T�[Q�Z�H�t٩��U�p>ѳ������V����#C�j���k'�0.�~��vS����l�3jv�d�>W�!�S"O,ݳv�D���<0U!M!2�av�$U6A�bp�����&��a�B9Otҥ2���?R	��"O6Ti����v��'�
�s�:<(�g[�&�h%�<+��<�R�Άv�X\ '�O(P_�1�TFe�<�hQ�T�� ��K�!SU�5���i�<qp搼�yq�@�
%��w(Bi�<)B&[OP��O��$^<B�J�I�<)�N�S� "Ąu
(3e�z�<aeI�4��q�E߂=�0��*�o�<�5�ώ	�VM3�CQ�6)PX�g�\i�<��(P����B�:a��jš P�<�6*J�t@<��%�H�0�atv�<ٖ@!�29����1T���c	o�<�$�Y�9���c�,1%�q���`�<��#cI�1)�D�'=�r���)XY�<��Γ$�n��ώ�4���K&�S`�<ar�P��vd�� [�
�� 4�B�<	�M� kO��(��H�
�svc�@�<ѣ�P($�b��"aғD ���{�<9E�̑
�px�-Г6`�	!�,T^�<9��s~�/Y�:!��̈́��B䉝V����Ч)>�l��H�a��B�)� ��#`���Q��9�� @/%輪W"OF�S!@�FnJ�f�Ɔl��"O����e-�K�'�]��"Ob�2A�Y�]6z�
h��S���t"O����G^�C�,�tǍ wXR��`"O�@zj
j���¤8C�T��"O��Ұٟ2�Ƚ��C�;=�"O��!C�Wm6aR3C[<= ����"OdQ��-�'���qL��7/b�b�"O��Ђ�]�6,���E��bs
�J�"O�H����hQ2(Sԅ�䖪)�f"O�zҌԉ'����+-v�6��D"OB�S�$@�nH4��+�Z[��;#"O�����;n\%jĈQ�uf���"O`�D� ��ɣ�0K~|��`"O�R��09zBe8�G�S�*xj�"O���O&}�%�FeX()R���"O�����>T? ք�,
�v\�t"O��A��6��a"%�$����"OR�c�Se�,I��T�V�ll��"Oxp�kQ?^��Pp]}ڼ�y�"Or ;��U�e�%�߬|�\tP�"O"D0��eP��2��YƠ�S"Oݳe����<��o���z���"O�QC����
�x���D$f{�!�t"O|�5&��\W�!p#d��;��Ua"O��[�#n�~����:��lCe"O�P�J�d��P�R�_�\ �"O*�xX���*R<y&~ �"O�����W�쩃�hD�m>
��"O4�p�P2>]��3�}��I�"OR�!�lY�$۬�6��:�� �"O��񅫎�6~�i�!�D�6>q@B"OF��ń]�J���ɤ�J�&�܅��"O�hA���r_*��@ Px�� F"ORD�G/�<P>��� hZɛ�"OXHy� дHaO�4F�h�"O<�p %�$%ʹȑ�d\F�-��"O 偅���D�95��-�Up�'�!9�Q�W��!V�e�\x�'��\+��V�\І�VY	0���'7�5��FZ`�_.Tj|@
�'Q����e=3�H{PN�\�C
�'1L��5��r~�H`FB�[�����'N]P$た\�
0Ii�P��b�'��Ñ�F2|1gН1<�|�+O6���J�!�:�`��<dKUꛐR�!�A_��Ԉ�.�.������6,�!�$]�ty88��N;|����ʧ�!�d�4wYhIaD[7?>����3�!���L�d��4�C( �H�ek�]�!�dB�M� �
S<�Ы�* !���I��	�J��)+�(p�I�F=!��<R��u� H�l�=(3h�J!����q�6+#m�� ؠ䙏x!�$F"*�D�b����N�\i���Y2�!��bI8�IeL��N�l�Z�� �!��9��@0C)F�:� o�!�$��:�@�P"�_~5" ���O�!򤑂J�b��&+	�q�nP��Щ�!��R���!e�c�88JdGQ!M!���G@^M������(�H�*g�!�DD�E"��	�nzLtP�(�Y'!�D�P��5��ŉ�bg�Ⱥ��L!�� 0�ui�"z !��Ε�{>EI�"O�P�0���;3&H3V��.xul���"O�Ds��M�4�Z٨�N��ogT|��"OȘ��.H��|���,Ua:���"OLy����k01�`���DU�q��"O,-��"F<c��܈�d�>'�J�R"O����
)�1�c-R�9� H�@"O�]�k��i�~�ƍ��W�����"O�XQ���������R����"O8����J8t��
X�xz��D"O`��bO	S�t@U'"rfV�R"O��S�aL� 2�E�.xF�e�"O0`�Ǐ�.q]�rC
SH`=B�"O�\#0 ��:�*����E�>4���L���X�ue��jp&#��H����!�!�䗱8ɪ�c�.\p���1 	9!�$
�B&9���N�R�� �0e)!��;N=}���8@n2%R��O5U!�$O@y���(Z-_�arUa�8^��φ �|��ߩ~S�K��1�B��>ctY�흊4��M��"ȩ'Y�B䉒_>�[��P5%���@s(�q	�B�	%Q���F��	H�-��%-/�B䉣P��LEa��Kל%sՊ�q+dB�3;V�S4&��*LA$��PaC�ɳ$R��? �н�V�R�	��B�&P,K`�ťM(�!kŔ�x�B�	�c%`b%�=`z��rER�Qk�B�I�D�b0�@�T�2tȲ�L�{��B�	�
��xQ�l��"�
��J���HB�I5h�n����2r�AZ��_,r�C�ɻ�B��w��>,K�qQA�&�B�	�#���q�Ħo!���v�T6	�fB�4i��}0e�N7/�NI2��p1C�IMF� t/�W@:��4��,�B䉒(���C@ͨj��0z�_5w<>C�	�j���0~�Ĩ���mp�C�i�j"�C�B���a����"Ї�O�&�3Ɗ;}�@���"�'}�ȓ�LBT�ڽ\��c�(��(fLB�ɏ<��U"�o��{���b!Ϗ�!-lB�I9GN̬8td]�h�	é41��B䉨�f���Y�+�1q@�B$GT�=�
Ó&�m��nПK̸t
�ʌ�vR0�ȓE_p��4�d	�*%�C�	�g� �r+��n��T��nl��8�I ep���ԽbW����#7��B�d��b�K�"m���P-7`.B䉲����w�ɝ>��"�� �Pa���E{J?�C�m�w��*4�]���%3��&D�8���G�mʠ�'�6y�)Q�M%D�,h���(��E@pJ׌:1~MV�&D�@�U* ������2!�09�+�>.O"�=%>�bc%���)I�酴J�8��Ĥ �O��|�,e��[�m���H��L l4��9oT5�W�1c��Z�U"u4݅�2���tI�q-�8(ק��( 9�ȓF���{��+���i_�h��чȓ�x-AAH��YK���.U�s�z-��U}֘)"��?@��Af��%y����H� 	 �,�-9}L�k&*��	F8��s������a��\s �./
���	I��!0�
={��58 !��X�C�ɺ$Ӣ�r�D�|Ҭ<��n��!�� �l��K!uG�T(�+эZ�l-��"O�j扂�qZ���L�_�2�K'"Oh�a�ʨpP�)�K��_Z1yf"O �p���%b`�,0*R��ku"O�@��ŕW�laz�!�0(ЈC"O֌��ѓ^퀍K�Fղ"� �"O��Xq�# w���ħ�Ȕh"O�)!�.��0��`PC#�� �"O�`��h�J@��
#-��w�L���"OV,�v���|1�L��&!a6"O�1`"���Mf�H P,��9���۰"O�0K�N�9`�v����!p�X�x�"O
�)�`�Ahi@lB>5��S"Oz�p&9��tJ%�YS���X"OL1���/ I�%Y��Y�B���"O�A�g�m0<���dt�|��"O��* MЂ�>�!@� 9쥢�"O�hXS�D1rO���S��a�x�b"O�
P؛��c#��T����"O��٠�"̬Y����R�F��'_^���`;&Uh�L �xҪ��
�'�����ϗ5��� ��2~�p��
�'�0��e@ MP-����tj��	�'��ɹ�A#�`���h9����':�%*�!�g.�:�@�6�q�O����T����j�	q����C��h!�3�TE#'LH4	���a�;ng!��_�/|���.ې<��]�&��:0!�Dӡp}[a��NHtay��L4K!�T=LMYԏ��<H�	kE�O�!�^�0�8e#K,N<�M2d���!�$�:�����k�H�0�07�B�K�!�d�<됉p0I4���R��ĸ��yR�]� ��r�C�}��%��ğl�<�v �	��ɐ��?.��a)�H�`�<)�C]M6�Z0'�$Jy�Q���N_�<��!l��V샫c���0Q)_Z�<��ș#T��q�b�}`b��]U�<!W�t�ZAAg��&e��|ȅ��V�<�%�\�m�"M�@�K�g^���'�U�<qs��#k��#(G�W�&5b��]�<�RK��"�^A�QB�n�V$jD�[�<�5��q�X��5���?�X��M�<F�J�!4 �G�H St0a�GEH�<Q� 7��@�wc��T��Q o�@�<�7�$���ǙQ����a@�hF�C䉸K�����W�>�v(R�S��y��+&���M(l��(�y���K3�(���J�XI��c�.�y���������$�=R�4��	=�y� �0#�
�as�ة����T��y�K[�YL�"�<L�谦)Y�y��b��ܪ����U0F���y�gZ&�=�惚�D���c/�y&�-j��z��z�L8!��В�yR�аh�Z�������^2�y"��LR��ǎ��<���c�V��y.�9Q�7K�:.�^�[F�ҹ�y2�������a���"�Ҹ��G��y"�Ľ&�H��$lC��zE2aHS�y�f��/H�`���M�ژ ġ.�y�I�/FZ �w�N$\ږ%Rd"�y�	�l��S��_f�֌C�y�L\��"���WZ*�+�$N/�y
� rPaա�=X���z�
?�Ҁ"�"Oҭ�4,ƞ8����C�l�.�"O(-��Z�l��+6��G+�XiC"O�h#��~�:V�S�<x�`�"O�Y�qmQ�,=B@�IY�fe|U�"O��!@+�2.�)�I�ad�{u"OP�(g�]!P1`u*C@&<8=Ȕ"OT� !��S�p� s"ȵNr�("Ob��+ۋ&٨E��+�$]騬��"O| ��BCw��@�N2	����"O��Qi�)�h;���y;>���"OΩX�P�;�8R�M0�U��"O�u�BQ7a�u�K"U�*b"O��B�[��}�R �-Z Z�"Ovu)�K��E�j@a�m!(l�у"O&��f"��L�LH�ČNx��"�"OL���,� Z]<�1�lG�E�5"O|1�ۆv��R�$����"O��&c�>%��s�_�p�(F"O`H8�ʖ]j1��D^�J�� "Oz-h���u�ISf�IR����"O���f�+[6�x��n���9C�"O�B��E8^��<x��r"OLH	�DN/R�&��ӂ�G��@�"OT1h��"�0) �݅�^�x"O�TRp��j�3�I��2iCs"O��+gh^8���f� k���s�"Ob	(��Ce�\I��\/ v �"OU�CN�W�^� ��/v��}�@"O��dhS�4?��h��F<�|��"O\���Zt`,rWв;�F��"O,�a�g��D�����p�dc�"OT��ǚ1&7��p �Ńtq��"O.�#��+�6��"�9{s��"ObH#`��!��x�!�ƢD�6 ��"OPb�
"9��p�������"O����i%��!��hԣ ���R"O|Ջj�0�aG˓~ �Z�"O�,��j	!Hx� �E�!{��\٧"O~��� ��0=�P��	)p���s"O.9�W��?�H��Ղбi U�$"O�db���+S��Yu�ȋa��Q�"O�L��GZ�O���R���MG�`��"OJ�v�U�!����#"K�U�j�"O���V��;1�[B"�2TLݚc"O ��$��8��|k4�$0J�y{�"O���Ԭ̋4v|P����uF�5P"O�Q�FM�5
h�m$!9���"OTY�:3r�#�
�k�D�0f"Oج�f��;��Q�Z	G�lq0"O*Q�rdW�dT*��@w���"O
��!�[���䆗*,j���"O���j�l��I5#�6U^\��"O�d�W�[�k��H1p���X|� Cg"O����g��B�0`ӏQOez���"O�h�$bJ8`��y ���-^�4b"O$���l&`��l]�Ma��{D"O���ŀi��tx6ldS`���"O���� UC	~j5��;4��R'"OZ�K!J	y_�dQ�I�T��I[v"OpĚɋ=^�j��%���~����"O@�"�Z��lr͜�c��%[�"O� 3��ޒ\`�E� l^]��9p�"OE� ��5X !�Qʒ�6�z�R@"O� T]�a�k�^-��&\�8���V"O�X�h�$S朒5�?�\��"OL�[ǀ7in��ac�Oh�k�"OtT��˝�|o|��U�U� ��"O:���Pr�&B�X�&��v"OZ�XΒ�?f�*�+s����"Ol�{eρ�)˺�sF�ϔS�2!��"O���Z�p�d�؁oWX�>x��"Opi�F#�|�\x�dP�F�T�s�"O|(JdaV+Y��0��)g||��"O�Y�R��JUp']�4ZZ|K�"O`:We@�b�ec�-d3r�u"O|�j�W�QR(]�R�f0YP�"O.���c�;Ld�9�d�O�]���"O�`�̿^I��hD-�p��Ȋ�"O� �W�5a�"}c�*ۭ�*$�v"O$b@�ڨb[��q���U����t"OP$�c&O</X1�'W�${�d#�"O\��t!W� ߄)i5,�4&מ��G"O �#J�we�����
�#$=z�"Ob�����3t�|Bi��@��D �"O�x��\0"e���+���"O�|J���$zҔћҡF<i<D"Od$�7 ʴE�rx�^pR2l"Oz��΄F�]zv/�@���� "O�D{0�87[>8CT���p�0��"O� ���ߢzN��P�W1P��"O�P3�Ο>oB)�E�ʺ@�@<P"O�0fh�5�JC��P��>�b"OTeK�Z���)����jt`�"O]��ݒ�fr�-ɪM�Y��"O���a��?�6�X�L�J�>��s"Ovmh�OC�SV��U�Z�A��%�y�լ9�±��hģN�X�Q�߬�y�\�+΅�C(N�|�n2e��'��i�r��%�<��O�#Y"j��
�'���9���+x�@D#�*@��Ѩ�'���ݓeS���Z?+Hԉ�'i�U�c�ܢZ���
�h�;\,���'���VE	�S���E`��8O� @�'�*h��� 6�����5*^ѐ�'f�M"��������w/M�XR��i�'3,���-�2~
LhDŐ]I���'���BQ�����H.QY���I�'0�e��I!y L�S�\�O��'H��V
ގ���@Ǟ�u�0���'ݠXC�$O;:5Ps!ȋ�8��e��' �����UʆdS4fЫY�|(9�'|���b�Ows�,��Y�M���q
�'�R�BE	�)�TJ!L��m�1S
�'0�Cc�%Q�ع@)V��M �'������G��ቀ/O�NYX���'$~y����k8�s��A��ih�'�d����r�hx��3>�}��'�FTCd�/ZV�jG�M(-n���'�<`J���i�>xA+�*z
�!�'<LQ���?{:�Ѩ����$wL��'����%�/�0�
�H!�hm��'�:h��L6\���ɡ�Q�?��� �'����ٶ71�b��<�T�
�'�B*�@aX���7� ��
�'o
p�E(��|�5OT8'���	�'K� #4NL $�l|���-�F]��'n� A�Ӊd��ݛ�%?_�l����� 𙡂�0��Da��R�r@q�"O��;�䇁��� �#���vDk6"O�t���g�@ �ԃ�!��a�e"O�`#E�$̙3���;���"OLa��Ie��� � �3k�4�ٴ"O.���^�MJKQ:j�XbE�4�yλ��#�� ]���)��� �y����m�G�D�N���%�؊�y��,O�t�bg	�L���,�2�y���g1�0	�ȑ�7���1CM�;�y§�=|���SJ�3{O��ӣOſ�y���T�d�U���W�i�ᐲ�y"��p�TX���%q-�)kfZ/�yQ%Vv8�1��N�dZ|a;����y"�%_ ��R��k����vfF��y�,�$��VJj.� V�Y�y���2bz�VgH\�)UFץ�y�� �q���`��hBDoŷ�y��_�u,F�@��G�Y/���
1�y�lU�2����0U$Ԁ�	��y"�;wq�����S8E�`�9�G�-�y�_
2�ր��댁l�D��!���hO\��3Q��@���8����F:џ�F���0R\Z����R��� �����hOq�ܘs�b��S#�d��[F �j�"Ola�W*|�=HE��)g�6I��"O.P&K�-�$��Ą˙s�j���"O�Ġ�m!�^��EiOYpTi�"Ot�@C�7U�:U[(�ak�y�U�'��Ⱥ����[nx��Ve	�ܬ��p�)D�x"@���6@+㣈�)u�б�-D��0�b�NdNi�Ҫ�'��xk�)ړ�0<!J���d�������!z�R�<1P �;*:���E L���qd�P�<��LȊV�����l8�9��P�<d��i����UM�I�fe�t�I�<�-8tC.0Q0Bԁ+����G�<1 �K�j��9A���;sL�+�j�p�'�ax��.OoD��Ƀ$o�8!:�#����<���G�>R��� ��6��0�ΚZ!����V0xbK�8� -�v����!��$:AD�� �h:�k�"�!m!�䗴v ��jSoB�s��!��X�Z��'�ў�>��1pw�x�H\9`��@�Q#9��7�SܧhL ��ԧ�l56ZF���g�H#��͟d��5Q�ϛ%��=E{��OȂy� �;e32�ڞ��y0M>�,c��`�Ӎ-��-�gO�V~Іȓ`X��'6��}���"?~!�ȓF�r��%�"jO� S��ڟj�
D��S��xĸP,��6��D2�k����C��$��y��;j�B�j����x��C�I#n���Y����|v̈1����?����) ?��+b[�KED���I�<����;��Y�4�{r�mS��K�<Y`O��X `�YЦ$SPnũQ�F�<�2��{KNA����0I  �m�~�<OխC�*���[�K׀�#3��}�<��UvF��$�^ AmH;C��A��0=A`� �JlB�9# _�O/���U�V{�<��q��x�l�9jv��P��z�����O0�$��N���
�nU�����'���S�%�g�p���<�(��' RYl��;<��B�Ԟ.k�%���� <��b׎ }(�(�Ý�F��q�S������|�&��CO��P+|��"A�-6�C�IN)&��P��6"��5�t�O��x����x�'�d�D��l�Q�S+�x ���x�
��z�u �R9 5r"F
�y��Ăr��9�M��*����'���y��]�wRIaf!�r�0DF2�y�i-�`jDjq�e�R��y�ƅ;Y�|������ 3��8��'Gaz� 	y��%���4 ��KAn��y�A�� :�&Ʈ) y��!9�y$�"���5���'Bz�#P썋�y2m@�B*J�C�3{x��4��yr-C T�Xӱ�Ψ�����y�g��)����e�_>o�0pbC���y�J:�0�3��LQ����T����0>1nR38���ѣݥ?N��R-]d�Ik�'����<aD��Isuj�!A8���[a�<�V��v������on`AkA�x�<�T�1|�
8�T�:K�R\�C��?J\�YB$��Q����E՟B]�C����b3C�:Dp�eC��Q� �C��/pu���!��*�q�^1Tn૎"�)��lN֎�"���#WX^B&�Y��y򏀰<�j�S�lQ#Kn<U���D0�y⏇=}�
����Ќ>� �����%�y�E��ZĴ�#me� ��װ�y���eH��t �"U}��hQ*���hOr���@+[���kakŭ(��TK�
��x~!�U,v���%	/+��hC�nF�)�!��I#�J����@����#��2O{!�DǕp	�£K�El�}�`�MI!��kH����٘Kh��Ӕ�Z!a�!�ċ'@�<}R$J3�,������!��_z��Tb�
|8�:3*���!��W�b����I�p|-Q�
��!��\C,�|yvN�U���cB�7��O����xg*Uh��:E���O�${!�đa[J�;��@�%#TJ���S!��@6��tI.��[p|:��"C�!�64�jL[��I�h�1ɖ�!���)�`Pg�_�"9H�'O�!��5I��x���v�8�c��r�'Vў�>��>Y�a��6UʚT�§8�$*�S�'�Ƒ��L��^A �Θ�o �t��	b~R�.���.��җ\ @�J��
�'��#G�� p��f0��	�'k��ImQ�=�aS��D�2<��x	�'E���/Xǂ,s��#�����'�`�0����У H#ZBQ�I>������1?v�k� K�vXF@Ƃ��+2!�G+x��z���
{AȘ�C A�,!�D�!z$�5�ƤKV���<L�!�J!�����%��DK���A�
|q!��U`�d��@j�?\B�P���!�Đ7v^T�WJ՘!Br�h�/G�!�I�Qi�焦j�lhq歁$.!����4@���V��)YWBƍ<!��L��1��Ց:{䍑�Ւh�!�C�0���t/X�Wu ��Y�!�DĚN���nmb�SO	�!�$	�gy���g��`�`���z!��Ta $��OE�p�N�BUI@��!�$Q�e�p1�g�����a�`)ȣXo!�� "�ʎM`h��lDj��@�"O��Y�LN90#Z(Ɂ,�)���Is"OZ����IUR�È�;?�d �b"O��Z�fQ�3�j�����k����B"O�
6���1����0�W8�T�p�"O\��3C/w�dʄ-·v�>�1�"O����.��P��A��'��'��6B׆��􆛜_��@�ȪB�!�Ĉ�G]�rdB�
����흄*�!��)g��I��D�������&�.�!�� �)f`�i�m�>w��mC�LO�!�G3� L�g��J����i�N�!�K2F���-�0�Rq�o��T�'�a|�E�'�<���'X92 �j�P��?�(OL���P� ��`i�iA�X
��6d�o!򄘔V3��hs���y
F��6B��3|!��D_�\J��Fz^�����Mx!�d��Y��u�vJJ�
����!��SPnm�En�0��-�6P:�!��j�$D����6�r R�횎b�џ�F��M��2��p-�<O��v�B:�y"��>��ip�+��E$4k%@՘�y'ԹBo���g��<�P�)�
ŷ�yB-Ln�R�C��A-k��TnK��y2#����!c(  ��<�'
��y"f�2-|����$�Pˆo���y�e���҉�1�Ѽ"�As����y�	ՇjR��#�#=�ƍ��ɨ��<���D4�\@���#�V�X��ǚ*F!�DV*L��0��RF�0S��,[+�y��	� JmX�&�WHf��*]*"B�I4�e�����iX(H���+'B�C��6q��qm�c����va~C��1R@��A�����p��OE��h�=��'���eZ�u|�[��Zܰ�ȓYa�S��>�h�c�FIa�Zȅȓt�>9su�B�m���5� �r�4���鶨��F�A]]��,��F��ȓ_ЮL��	\t0ؖ��'𮹆ȓc�l��3,����[@�A�Ky�!�ȓ7=��IE	j���EdF�%�0}�ȓ��-�rd�(�X��s��=�DX�ȓ���h�G����cs�<i�x����T�f�F�T�����6<N��d&^���#�����*s����ȓaP���2��9���7����qզt���c �#6NM�Q`v���$����m��镎�3����ȓT%��`�8r2s��W��%$��G{���M�v"8�;�\�>-��b�X�y���V���<x��T���y"F�T��z�㌮~�t	�$�E��y�&S�#( ���B���tɇ)�y�j]���
��;����AG(j�)��#%|LR#�϶5n��&K��j�|��ȓ!������Ի)�: ��q,XY�<�ǌ�0���@P��y�ҋ�T�<1��S�F ^�䁛�FsМ3b��w�<���߄mP��1�.F������p�I}���Oܚ���ɗ?��´�:�pQ
�'<z���Ƃ�Ϯ�Aw�^���$�
�'��5R��8.+���(� �ک�	�'|` ҖGр�,֯.�d�I>y�z^�I�V žDz��RfEI:l�p���S�? ���
 9�FPk��l3����"O�������#]t=�w�]"D!}��"O��&֞�(���Μ6n�ű�"O��Ђ���v��(����c\D�""O�Qc
$T^|X)w ��E�x���"O& Z�/߹')SRA�"6T�p�"OU��+L�oB�(���Q��"O�ɓ�%��(���!�0|����G�'����ʱ�iY�}����Y7T\B�ɵG�J�(���4����[	2B��7
�`��E�$O�q�%n�����0?��Iו6�z�pUbY1|�:�*����<a@KZ!�&���
.O�Z��v��~�<�Uo��B�(t�"��	��[cN�}�<"'V3{Ĕ�J�/=M�Лg�a�<�5�& ��l:�l͹}�l����`�<��Ŗ��!��H=�2��І�R�<9G[0)���ql�UmyfKAP�<�Ч��@r���	�B@��NZK�<!�@���䀐��	Yj�@D%�]�<!G�	y'���BgQ:�F!�*�n�<QBF,�.�el����C &�l�<AA*�,�j�`�/c�l�K2�l�<�aF#����G�"{�.���͈k�<a���@��"6���+�0����j�<��ܤ[P�J@����D��e�<�#L��M�����DЬ7�� ���`�<�BE!l���#Q�Lޒ����Y�<a���3h��c�G�-Z郔'�Y�<y��3M�!�c� OA����U�<���*��p���oV���N�<��˝9_C�ة�X�nI�y9%�M�<i�@�s�^�I�*��9$�MG�<�o[�r�,�@d�d�T@Q�Hn�<9�.��E���i0 Ô~V}	$�Rm�<��F]�S��H�sĜ;E ��*&̚k��hO�':�!J���;l��g�eI�ȓ�M`Ʀ�)�(@T��!�r	��K��|��k�h�I��Ɇ�D ؠ�ȓDI�E�J�ʅJ
��!��|�<�V�ι\�p���7�ؔYâv�<�w#�;Jz1��.4ROd�I�]r�<�+ۊ`"�=化�Rg�:3I�F�<I0b�8.�1!���N�����E�<���Ő՘��D���:p��DC�	�F��-b��ڢ,v�UkEOW�(L�B䉘?������i<����V;,e*C��	h�P�7��D~UkQđ�N@ C�'��哳���/*�T8���2:w���d$?��-^�	E�l��}��	���t�<�K�
vŎ�cal@���Pƨq�<�&��?>w�t�삁W��`�)o�<���M�w�l��Ũ(?�J֮]A�<��K�z���xg" 9JV� R�<a���v�He�!
9ȼi⧛K�<1؛x���᪛!X��a���k�<�m���(	 ���!�Fi�<) �¿�\���--�xi��Ky�<��0pkH	�*D���bNL@�<iEK�� 6<8��R#p��J�I�d�<�R�P�V�~�4�� 8_��R-a�<)ck�X}h(�6�0��X
VT�<��a20�mb��:�
�.�S�<90�3eD���U5t�����Ux�`Fx
� �)�W�ϓ{?D��`�݅)ٸHW"Oj���L6_&� WC��*�vtI"Obe���y�� ����q��jC"O�Y����Аj�D~�t���.�S�)�b�6{�Ԯ8���G[�{=!��-v'��i�� ���1%��5O!�dߟH�
�A����[fEL2!�$� �$0�ƃ�:�t��d�!��Ob�=���ukƢڨQ�>Ts"��4_\V<�"O,=k-�T��d!	A�W�!k3"O��C�B��E�g�;@�~���"O�����H����MJ�"�SC"O�)%���W��|�7FE#��RD"O��D��[��� ���k��@�F�z>)��`R�r�
P�r�_�i'����Ĺ<�+O ��7�&�J�bOC L@a��p�8��"O`1ƃJ�E��x°�U�<n�b"OJ���DD$���&�/Hk�,��"O����
��\�-����f��KG"OBI
�7v �M�񯙿
c�mb�"OTP%��
�����JK�h1"O� qwjİ&r�Vj_��
�����Oأ=�'X�x�0ԉʌb��Ԛ%H�6d�L��Pa~U��J�?��zχ2M���ȓ%��e��'��Y��P�߮3f8؆�?�\��bʄhGN'G�D�ȓ\~��$$:�y�Q�D>\`�ȓu�@P�"h	�{���3�J���l�ȓ�T�a�׏S�TY�んu. �ȓ��M+3 �-/��MC�ꀕ;���ȓ/�2��������sEm�i�✄ȓM�e�T朅1D,AS �%v����ȓ4�4�����0q�+��!=X�لȓՂW\�!��=�� �<O�x�P"OLa@ ������`ƅS? D��"O$�@�HZ�0+��-(��"O�qb�/$�vD�&����D8�"OX��U	��E�.���
�����"O&�KtC��u��(q���z>��E"O`�{�����ʅk��g�P�"O1��M�c�N����7-hL<�'"O)@r%LY��p2 'ϖM]���q"Ov���C��O�D�[��P+LS�dI2"O�|�!� ]s��y"*�%�>��"OJ�Y�S~�X�`@#G]��0��'��	�6�����Q+bp�$L�4C�	:�v�bi[�W������FdC�I4_��@����)hX��.O�DB�	1#_�ѩ����J� �B?H�8B��*.��eR�b�r����f��(�"B�	+Xk q���ڷo!�B�ɚ}o`ȊW��(�İ�$�\RivB�	A<z����	 '��d,��O�C�	O�8����՛D[�FF�`��C���%���{%�8�|��"O��O��a@FXaB�P��p= �"O:�r�Г:8�z�M�;��ʲ"OL���k���Z���S�;�HH t"O`�cb,U{JQ1��h~@QQ�"O�� 4ĝ[�q�L�k��c"O�mj�̕
N�ՠ�JH�,�J�Jd"O6��s�]�|�:��ށ�tt`�"O�@�TH�02�IuGK�N�z�"OT@hb!�4'��M*�-�Qj�H�"O�  �r@�P=�|��5Ɯ�S{��a�"OH��古P�,�4@]�A�da"O>�HD�c�u��Wx����"O�iX&@��	�غ%,C�Bd�'"O��(�Œ.�@����1+���Z�"O`P闇 ��/�/�TY�"O��X���E��̈:�.Q�"Oȵ�0C�7�6AF��l.��(C"O��!g(�M�6��!h��H�1"O8QѓҒy�L ���Һe�Җ0�y�ŝ�b�B82gb�	@hZ������y2�I�o��EI�ď.Mdc���y�%Od�}Ycˈ%��DQ0���y"E��5�0=hu#�O	�tSd$���y�۴>w�M�F�E�vh�S.״�y��?w'�4:�i��:��8��)^�yB�,{�`	�$̎�1��$��f��yRG�#��L��$�te�ä�����!�OL�H�%��T�Z�:�`G2pq^���"O����K:�$�QW�Ę`"%p1"OB���u��X:�-E�NL�$��"O~\h@�4F�t��FT� V5�"O"�@��%%T�Eo
�U��'|�cF�D�[ ��k�	�R����'5d``��uQ� ǂЌF��)�'v��JU����&Ը���'�R��
�' <��SF���(֫P�1B�
�'.��7�(O~T�ȥ��*+�L8)	�'���*pȉ�.��Aش`� p�h�	�'? [��,I�f��qX�� @	�'�l�эNL����AĠt���'�He��C@q�3Kքp�R���'�H�3�/�-,�}�[�lY�-y
�'�X�h� ø�����Nxr	p��y�@��<ҕ�C�=*���[aDI��?��'���F����,���Ƙ
L�0��'�Z����K�_~�XYQ���|Q0b�'S��)Y�?��e��,=�NA�'�p8�I14������*�T���'qx�Q�Um��H@�E��� u0�':���eV�Xࠨ�b	�(1��'(f�2��FĂ5zu��*R|f44"O�����;tV�z�HL�I��"OH��!IK0��	S�N0.<:�I�"O�(Y	ͭO\�3��G�rz���"O�|���ÆcZV<2�D%\�H���"O�y��@M?u�]�t�+}.�˂"O�2��R�"�X��vbI�s��Z�"O���5�������DBk��R���D6�O �;�Eu;B\�g��G��a�1"O��y�HW�dU�e�4%�����'�p�e*W*��B�D�V�9�'^~d���<�=�1FN�B�y�L�edPi�A�;�ވ:��P
�y�	T�M�
����N�:c���Q&�y��?��!�i��+��I"�4��'Jaz�(P�}� ��eω#�xs����y���Z�B�D�i��lZ�(G+�yr.�.p�v #W$װY�R�3c�O��y� Ҥ1��q�P�Ь(ب�r�c6�yB�S�efACǉ�P�l(����y���B��4Q�HH�H�ƭK��ݫ�yjkh�� ^u�x�0J�y�U;��%�2g��ӇF���y
� �U)��-wy���T����"O\
E�6*���I�*�>[e�U��"O�X!6LЁJ�&������{"Ov	�Fg~F����A;;�����"O"�[��?S����&I�]'��"O�hI�R����bfF�l� Bd"OP�C�\�&q�h�#U�z�Q"O�5z�/�0{f���fc�<-�ꍂ"Op�
�G% nd�#T85[��4"Or(��ʓ@� ,٠a@I����r"O����#�;Q��x�31-����S"O(��Aa�q��mT����o"O���#סK�^`�&cD9%�� $"O\�(wI�2J�xl���O�b�C"O��B"-u#J�
u�L�L���1W"OL�[�O9�lڒA�C��0��"O���.L1SنB ��y�D�Ä"O�E+���.n�T �a^��b@#"O���M��z$�����8q�D���"O�!�DL�}���R�-
�>���˦"O�@1VeE�7(j�����/;��"O>���l�Τ�����$<h7"OM�ӊ��25��:�U5��D��"OH	�rlF+g�x���?Qڌ��""O"p�Eꑍo�P%��aײX]d���"O�V���/�Ea��@X�B�"O��R㩋� � 8�).,-��5"O� �d��0r 1�Ph�$^$L�"O��p�I�&�v$�I��`��E��"O��*1�\�
���*y�z�cU"O��fF�i9�ybP���2����"O�����e�4�+�^����c�"O� 1�Ō
<�P��DUx��+"O��bV�DrB�1��)�9y҂ �"O�̪uk���I���&#f�dp"OL(��nS<j@+d'�4����"O2�93��o���p�����5;�"OnT �L�d���W#���W��_�<�HS�"�9<�E �-�S�<��=>҈4���܃DЮ9Xc'Q�<9�n�$w�$@�T�CV`3�^d�<YS�bj��1��.:��T��G_�<)��X+[�ro�)-����!�B�<���+�e{�ʋ#}�KUHOi�<�`�?30Kd�
�xt��(i�<yf�Q<`�ѧ�P(~7td��K�<g#�?b�H������ � �-�]x�8�'���"c��5�
1�`׳[�|��
�'ۮ��D�'L��r@M�6F1
��	�'s�p���Y75��h�į@�8z�z
�'M��D`�+c,�aHܧ4h
�'6R亳e0$����\t����';>�$S�Y��A��.<u�BP��'|<)�e'J5g�n�2�Q�j[b 

�'�*������֠��D���&��
�'��*�c����K���c%Д3
�'����g�,-�QfGA7' *
�'2�!pV<H��9���	v;	�'\�9k�A�6�.y{5�W&����'���A�?&�$49�ۚ���'�(��������;���'���	eU�f������-��"O��3F�V$dn�ȦCΫ\n�#q"OZx��'�z"�?\�@�"O� �x��S�Mt�R(��j��D2"O����Ι.w;Z	���(~V4�W"OB)r�gM}�FQY��S� VR�X�"Ob�xŇ��b�����D�Dd@*�O`�T��G�6A1U��,^�:�xT��OPB���&��PփRA��m^�C��4x2%RP_�'�����2�JC�IQO*xQ��:����d�~4ZB�I�k�(��o"$i�AӦ!��R�<B��&E�|pb��T�m�&a2A�+ �&B�ɋw����^� 
%�U�$-0B�I�~�RA�P��%Rl.��ՊJ��<�&�D{���+�����g�Z�1��,�C���yo�����j�"�p�3�Q)�y��?nb�hEc�#h���B�W��y�삽R�� &B�;a�~�9�bݘ�y���ff��W���*�x��T�1�y"!͔S� )�G6kE��Th���y�	 G�T0R��j^�i�5.��y�'�:m쨱�h�N�KD���y�J�Z��U��@����)3ɘ�y"Ϛ+B*,�bT���%�r,
��y"�X�q;������� ť�y��V�c~����Q1l�(BPKC��yU@�*y�1G�Z�x�����y���H�����d�e����5�y�l�(bX`9�'V4��('#�-�y��8B�0�K�R���B��y��3�0-����*\��	��y���gk�E����k��g<�y���2K��x�'ò�f� �AǼ�y���D?hqG�U\�,H��G2�yB�@�+9 �cd��a�تvBօ�y�WM�ޜɴ��_�xI!q���y��ŎI��˷h�?DCN�Y�j��y���S�t vd�$�b��+�y�����$-��~�#��^��y��͚��c�>	&�C"KW)�y��H� ���FQ�hR	0"�̉�y�j]�6J�x°�X6���y����y���1]�o�$�t� ��	#�y2��;^��}�Fď3<�6D����y��;�.9�e?.6huP0	�y�!	BnF6�0aEH����Yi�!��\h�=��l�[)�]�"�	b�!��>g�v�d/3.�Xa��&�'|!���e���x2���n�`�"�p!�Ǳņ��J�W���	v��Wb!���f��iЕ�N]S�b�a:wU!�D x��8jV� J�1c�`[�H!���7�F�;V�G=jE��)s��:�!�d�t���z����  n��F�W5�!�$A�\5�=�pƻN���m�js!򤁲0K�� !��c�#j�	=�!�����`��DM�N�Rw��	!��.�p�EY�z��8w*B�	�:E�9���"Df�� ��:L�B�	$@ P�I�<}�l)��1�C�I�b�0b#�+�8��A��F�C�>'Bi�a�@)%t|S�$'z!��D�F�BMCDS�	3�A�����&�!� s�\���(��1���®+�!�D�g��bV�!l �.��O:!��'6�J�hքS2*B�a��.H�!�� �d��.0w�\�{�Ù[$Hã"O��[�Nߝ2��`З�W�A$�'"Oe��.��K�"e��Ce� )�"O�p��ߔf~@$���֨K��}��"O�"�k�qRΥb���O����"O�!�1�X-N�ȡ�4k�(�"O�R�`ڪY��m�q�F%�"Oz�z_)n�KBb�H�r�+��t�<aPa�3r~j��1�3d}V��[�<	v�ɓ��e�%"�1�`I����<i3�����2fB�!��d��Jq�<�&@N�~sfQ�#� ~�J���/�C�<@�R�l�Sw땢U��9�uz�<�S\����ǝ���Ш_�<�"惲8D���h�p2\����Ea�<1sL\&J@�B`/D �!�/�s�<Q�֖dz$13'�'3����.Ll�<�+�4�4Pb�c҉cAE�#Ym�<iw-�2��͠3+[�`b�#2�~�<�d�;'D�D"܀W���Ox�<�� ���q��LQ| �"�MHt�<��@M�d"}� _y81�VCBo�<��G�{�N(AC� �D0���i�<���[��d]	n"tBE�l�<a��Zx�1!���w��l�eÆs�<Y� :R�ְbE�/c�Ƞ� �q�<I�C	��1 �%�?;�����DMo�<�A톽nh{T��#|���
�g�<	Q.�<b'�)�	�&TD�y��	d�<�UfL�A��	���C#��@U�<���Ӏ,3p0�A�ӥ#��հ4N�R�<97��f�:T�֋ӇG����f(�Q�<���|�<Qѡē�t}f�%�S�<IEɃ/9V�02b�0u:�z��R�<A�iD�НX��Q(K� �@CTE�<I�o�O���;�&P ㎜H#�w�<	d��@G:l���E�l�Cchv�<�#V�4&&�22�R"�"�"!��q�<!�(��%��\A��/m �)�b��l�<�t["6��њ �@)Z �]�4�\M�<I���Ӿ���K�	/�+C%�J�<�BMM:>�tA���"������]�<�W�#��j0�&^|r9Z`O�X�<9��Q"
�VD`Q��$G�F��o�L�<a���@��h�U���QP� F�<QVe�-���#�Q F:�P�A�<afk��,��:�AB�U�v鐵`�y�<)��ȍG߾�;Mɶ<U�]���q�<�� -	��R�F\��J`�U$Jq�<9\N���c����`ĂF��!�$�2c_Lx�$�����у*�!��Ro��	���+�-х���p�!�DG�F�(�dS�8	�}1�=�!���N�Mj��90��i ���!�D�sN^$yB�Z4Z~e#D�:�!��W�jp�"�(O���+��Z�>~!�$�;<�Bȥ.��"g豢T�N/A�!��?d��j C[�d�颴"�V�!��ϋ���r'�`F*t�c���!�=
.�1b98�ؘ����lu!�DO'p�� ��mߝF�E��Q�pg!�d��h%�Ԙ=a ���AO!��R�
������xARX)�/!��ث_:$9��a�;0X��ĕ�j!�� L5;�cW/|�C���>0�P"O0R���-aӦ)��e:�:"O��@T,��e�J	Xp&��d�RQڠ"O�����VÒ�S�n÷�"r$"O��� �����l��,�*�"O��ԥônL�A{�m�	f��H�"O��7�p �ݸ��_�Ph�:�"O�SF��bąH� ��[I��8�"O6�b$�:]� Y�͂�$2����"O85 ���%��h�`L_4_,���"O��	D��fHW�IjJ�)�*O.�I�k]���eO��)�'.�hǆ�7����
���B�'~��t"-?0��B�H$
2�Q�'2B�@1'��B�:���d$��
�'frY�v�G�$d�X$';Vg��A�'�68H��KK.���]�H���
�'��BǂӌP���Ίt�؅R
�'6(X�#��-T�a�#Ѵo���
�'��ՑtmOr��ˀ,Ѓ\��H
�'��tZ�h�R�Cp��"(
.<b	�'>0��d߅$Y�t;!�~t���'ͤ�Ӳ(����Yj#��͛�'�\<rEL�? Yk���@xd�'��azЎ^�d��,X"_�� �'Kp�A`�E�8��ɸĒ�
�'�0Y�d
G!������ݳo��k�'_ Ax�B��t� �&�Ǥ7/�m3�';H�����;W���o�_�9z�'|=���A�F�
�8�=�	�'�R-Jt�5�
ȹ��p@�:�'�^����6O���)�Z���'1��{���-�`�SR��!R!��'ᄄ
��Dmnv���dS�'h�8�'������% K�6d	2�0��'�!PA�Π;���,��r-~dY�'��y��&M�2!D�[ŧ�=v9����'h�x#7��(<�|h�΋#n2z�*	�'���rSN�'�������e ���'z��"���k���(��ʊd����'���Z�)܂V��<���6c�jA��'eB`��)�Z�|�r��֊�x�'䔽j�NR�M�z�3��/���y�'���hQ.Y@�Ӳ�͑,�8�'��@p�������+Y1V���i
�'��5�⬜S��5֍P:b	��'�P1�\l��[�,W�Eb��',��V�S�wM�LJ�bǝD��I��'�6��cZ�s"��NΥ<�q*�'����%a��psL%���G�=ޚAQ�'* ڇޣgz(p���B&3����'�݀�B]�:V\��4�@�0P�0�'�@`���6Y�&�"[f����'��$��K�c�Z�Y3��)T^�$C�'C�b��� >ڍ�bV?,����'�x��#��Q+��+b�&0�j���'լ��b�IS��x�Vi�#� $��'B�(\u�:@I��٪"�hi��'N8�R2��]X(���$F�`�'ȡ���.��w˓ HT:�'��1�Ǌn��!k��N:z��q��'
��gIL2%������@�"a$%��'9N\�RBV.q���g��p�'O�`h�S�M�hp�v� e��b��� 	�g)�&���N/��q�"O�5J�b�%#���E�D/m�J���"O8�� #EM�~�kT��8O�N�۷"Oh4�GrrcŪ�1�|C�"O��3��pbԩ 1�L�]�X�H�"O
`�C�&J��6�5�8���"O�ݨ`�s�T˷�ݥQW�Mr"O�Țp��;���3,`�@�"O�y� '?�h�щ��R&ى�"O-��� �8���@Q(_5�^��"Oĸ��a߿x){��]-H}�"O�PQ����;�
���Y =����"O:	i�j��x��!���RR�v�P&"O`hHܪM@��r��h�"OL$8�æ}L��2�@�_�m�#"O֝���I."(��E�A8sY.��"O�,{@/��ձE��
V��z�"O0u�R�-BC�aI�� 9Q�e"Oց;`#W.����%W��;B"O�����s�ԕX�H�B<d �"O֩���� )����M<*�p�G"O�Yɰ膩 �@���G�$Dыp"O��eGۂDĐ������>\���"O�if��f�z4���w�`�"Ojx�B	%(I���h�
 g"O˶&>d��[����E)I�y� Ͽ
���[5��Y,F�h����y�T,<]l�sg�7F�(Ŕ/�y"�	�)�	�	T� �g햩�y�m�#x::��(�`��c�O\��yA�_F��@����T�ʭb�Ɂ�y2c�	�N���!��\�CfFP&�y*�=�� ����?~��pɅAƼ�y�IUr�0C�m�Ic���܏�y⃂ �Bd���u�`$�`��y���!��d���q�ؘ0�.���Py�� �|p�D�X�~~R�;�EK\�<�E�T�H�p�cVs7�ȈY�<�F̛�3�,�#�J��2C!�\�<AK��V�H\@�H��o�RA�@��[�<��I��2���.K'\G��c'�Zl�<��C��(�ʌ��CO$Bye�q�<�ь�6I�!ie$,���y��B�<p�Q��R�D�I^֝��E͹!�!��>��"k�,u.���'�^$<�!�䍖?��Q�ɜs!"��"�P1!�� �̉`�B&�8���!�4c�!�dD�Y��1���̫����*�#>O!�d\#X�$(��v�X/�	0!�P�-��L	TC#V�M�!��P@!�$ޙiY܉i�7 Fv�bw)s!�$.?D��2Ŕ!4
x`����!��2.<�w�S�@��1��A<�!�$��hb�����N�lά��C'�!�$��5U7ʃ�s,ۂk:�!��J�o+���6!Ƨt�q�#ߢ�!�d��K��Uj�Ybl��@�8x!��,1YG��p'��'�N!�$�0B�dDq��3�ts@j��^�!�G	����&3r[�(T,!򤜀Y��#PHV�Jyn�8�s!��ݜab�4����m�^` ��S!��0%D����"$Up!�R��H!��>�(���C�+���b��>]!�� �	�G��R/���3jX�;(N�9e"O�\3�(�TlC�� ���(��i+ў"~n�	:"]
�g�=�Ȝ� K��?_F�OP����(b�lJp�[�$k�d2�,¯���^�� )0#C0�X@�I9uD�8��5�.�S�'T;�L��h�!�P�u� gBԅ�e�L5H䩞�6ǜQS�+t��Q�On���ˇK����93�\��"O�2��ec(c��ƨX0��`"O�q/�R�J�W��	?(֍k��'��	6 �"D���
-|����YqB�I�&>Lб�^�*�(+�O�g�BC䉔� |�DL�b%���'杗V��B�	�eP3 ��	���!�+?
�dB�I�)-^���)��drs�KR��G{J?%�2c�/�@%�ͼ+yH��g�j�=E�ܴ��@��S/(p�qw��X���D{��'3�ؓdO��QAn
?/�a+�O�����X"��mݹ`H=����	W+�	�<�J�ЦOq�j��"
�2 Ҩ9@�.��J��7�'i�!��؇dl<��{@�V$�D�MH�	Ex��)T�r�R���� ���P�DY�=�a}>iC�C�Q�p�ްf'��(Ɇs�g��rD�C[���iƲ����f���'h֐G�tcv��yu�P4���L��!�p�A�4D� *H#	�Z̲���-}$�P���T;�4��SF{@�;fIؑxR ۟<f�|*�c ��y��{��ѹ��U
j 
��3���y"�'=0A �O$PcPd2�I8*4p%q�'mڌ�R�*��k���*�����'m�(�P��=\�&��f�O�"�li��'>%���N+�!�ך.6�)P�'���a�/�<ƙ��O�z���L<�r�"|OU)� d`�L ����DH���Q�O�U"�c;S_�	�e�]-u�  	�'B���g� x�B�L5����O���D�4D)�6����	!#<!+A�C��y�"$�z��G�$l��D��yB"�3�����gdv��Ə��x��'�IZ�N�2-�&��Lʂޜ���'�a��ȩm�)���.춨���N��y2iLO�2h8@���<MA����yb��/�� c��	"��wI���y�nΥ#����FT�O;&�/W���'�az�n��`J�9�, BV+�N���<��k�*#��<C�Ӱ�*l�$��@
�B�ɣ.Ԥ,Z�hf�=5st�@!LO�X�>`�Wr���Z��Y�q�� 3',��<���&"˪EksLP`�jYZ4��y�<�U���(���a���Ф�V��t�<���2f�(����4H�9	ap�<��c[�C�,��W��0������k̓�MKS��>IO|J˟�m�!�����D#��?���q2������'cʽѥO��D)fx0��2Z9P�6&2�S��?�&j��c�! �N]D��"'ȅX�<�(ΕkT�E9��؃�|yz�	�?���'���`cT�Y�uNU�͟�L��� � 9��ۋR!����F�"���ȓyl��2�J0Q��Tj��ٰ�B����O�'�Z`3�K\����j1�$Xz�N��3��'����E
�i��\`U%I�O�K�t�Ik�����>�6�ϡU^VP)�'Q�:�ّ��o�<�!�4�0!*���<��ᱠ�7؈OH����(D��ɲ��ԕ5@`'%M1!�� p}z�C:*��p� ٦sH���%"O&i��U�I*(-c�\kB�����Oe���i�Of���@Cn� � ի߰w%ȥx��x�We�����̅Q��Ӑ�|��Z��-� �=���'o�S��?K&"U���Ucb��@h?+.�C�	���r�G5^��)�-�% �P�,�S<��}�pd
�M՘@��D��Z�xQ����Q�<9%��I[�x�HȦIx�����c�<YU��*k���AɞyM"I���J̓J̑��'�H� ��R�B���l�"ap�q�+"�Dܖ�0<a���MVB=��� eߑ��J�͙�<�L>!*O?%���1����BK�_-�x᳥=D�����.Z4���bLK��J��0?��O�Ósl$rG�M$r��"�ߑR��p�ȓ*����G!4Q�4C��H�<�;�4s��oDC����q�:�M��y��X�]��!�#&�8:�R����e��D�>��!1���fV������az��=	\\��?)V��d̮F�!��1�g��z/�9��$ma��"O��Чm��*�R��R0̔�"O���
®�@�{��V�t�5He"O�u��HGWwd�qw&^(g ��6"O,��[M<���� w�(��"O`�t�r�:Q�r��vO���0"O��b2�-e�pm�*]>�H�"O0(��H��L�&	���	~=0P�"O��r�;�8���E
�:-4�"O�Y��1FL�<I+E0E���"O���B�Ƹ4�b� H�`����"OFU�A�V���dȚ(���P�"Op,��. �q�$��1	�L�c�"O0�2
G�z(`��0�����"Ox����m�`4���  �^E�!"OD Ys�ԗF��5:�A,Z�ne�7"O���� J�;��4����*�z��'Nў"~ZЏ�y�ɢ��

k�O-�y�Y�">�b��S!_lTS��@�ybDPn>�+���eϚ���"���0>iM>�dn��-J��q6��/i��H��^�<1���?)d@`Ri�)`���@֨K��hO�1E{��Y*T�kbg��k�Z1��+����m6Uis��5!���W���{� ���$;�O:�PCg]DRڅc�,̏e�t�(�O���&_^����f�3e;d�"D���,�R��R$�t�S`�!D���W���!Y� �wj��/�ȱ2	�''�܁��� C��!���$�C��hO?���5v��S#��5@\� ��<��ضT�<�t�O�,�	��NV{�<y�UC��<1�BJ$��u��5T�X��ث٢a��-&�|���:D�`���{�������Tlf��i&D�����\(2�`

Z�t���8D��S� �@߼�I��l�BV�:D����A�;pZ��dȉ�C������7D���%�N����wd޹rD�4D���q�G�b#~���N߹}��1��M(D�`� nO�`�d��-�{�l�� '&D�̐�!<e.hb"V
U�h��4�6D��1�"�:b3�AT�y��\*g�(D�l`�`ӧ��|eb�m�R,S�*O�]I��0y����Ǒ�Ȣ@�"Ob��RL��NVi�էK�1�\@YP"O� Z�2޴bz������o�^鈲�'��/���9�G҅@Y8�$ �27N��ȓn������ ��5�C!��l�$�ȓfy���rJ#"��F�$|MB%�ȓM��`W�;4��kš�
��1\L)zr�\+J~�y��!E�cȶQ�ȓN9.Qq�Ƶ�d�W �#|(X�ȓx�蕸���3�2����$4t�t�ȓu�x|�'Ý n?�h`w$7�i��yGj<3���.vH��v	ʞ?+�ԇȓF�F�SݺV®u�� +�1���T��u@�(r�͕�[�]�ȓL���@��s�I˓��
j��ŇȓC�Z�J@a[*�J��� Uin4��l��Au�$<�-�@F�{�rU�ȓ	���@U4O���%G3�ȓ0��pQ��2y��U��l۾�m��F���(Q"��(��=��l+�h��p��|��)Eh��:�l[$��@��v�d�##���X0�D*��Ԣ3}Ω��V.8 NJ�������Q�i�ȓ9�.D�s�FZ�4�F!��jk`������ʦ�Ė{8�A�D/[�4U���Y���g�n�Vcؠd:\9�ȓY�Ju��cٓ-���B�����b�(0����!A�H�p��1�K�<D��9�F���K�/�$��C��J�<�T�>Vf��ad�*�<�k�A�`�<�&,8'����.	��ࠀ��^�<A���%*2�#r�� �)X�V�jąȓ������KL*�!���L1�`�ȓ%�ֽp���$Nvyat%�,{�*�ȓ:�D���d� �Q�mơ�ȓN,�KE�H�<�0�"*�|�ȓ�α&ߟh�t�p�@ԟ!8Ҡ�鉷M�~��
�fNH�n#�Z]�i?Pn8C6ဗj�FC�	�xT
��􏛑<�D�X �ŗ,kC���`6�V�I(�C����B�Id�Z�`�#d ��^���C�I	�!B)�6&&أ��<<2B�	1$�T�����\��̂�e��C䉕/��iuH_� $�1��>	�C�I9Pv�:�U�I(x����0DzC�I�=�"Vܪbep�K֣�a�B�I��T��X[��2fiԅ:��C�	��F��M�>E��:�cH�'��C�	��lX$H� �)$�ʬj�zB�ɐ z�hp���=Ghd���F
nDB��-�&"`F��l0�3��+ �ZB�0�$��H��p�����i�n|C�ɹ.w������0p>��Q��V�8[NC�I�h�Ѣ�=Y<��!AmT�UZZC�3=�5��F?�F���s�6C�	�!���[�g�8���[Q�Ԥ	�C�	�&u��*�E�H���x����b#�B��1�A�0�V9X��d�%e]=x�B�	�]V=J��ѕ�p �M،L��B�	!Pu�yP���f�ba`t��U�pB�I{��� +�M�z9�U�̞$;<B�"���g�P	�2AK1o7�C�	+.�3�nD�>Q*�@��8��C�	#txص��=%'��Xr��
]'�C�� ��YH%N�8,r��C��C�I�v�^I:���bU�]p�	y74B�)�  {�!J/)B|�!�XTR�0w"O�XTG͋#7d�HR�+]^�G"OhAP�.�7 uz�H!� ���%"O.��
Q��e�1) Y�f�z�"O&��7��0a�9xC��ɪ��c"Oij�D @��[�!�'I�8P�"O6�(�K�!?�ě��]-���5"O�����6%&�����i�P+�"O��oͮ2��q���K�GX0�F"O���<w����Ɓ	*p^b�QW"O"\Pw(ͦJ�Q�� �Qd�S�"OؽFk�4�恊��W�'F A��"O\�"�f�2��I���$$��"O�!a5��$k{�$��Z�O�Qz"O$����*"h��qԎW����I�"O@ XG�Ø�0���+����"O�P����ݶe*d�Ӧp��h�"Oz�C�.M��;Q��('0HI��"O�h�� Z�:bb�Q���X� �u"OJ��/��h�`��E����E�"O&-�4���0��4����.i�>�sQ"OBTx�c_�>8PZ��ګxd�Q�"OHd�u�ܗc�4��Ao�B�� �6"Op��Q�۸1O
���N�1��}ʔ"O�*�N���r�{��ʬ�Z��'"O �����]�H�cю�}�<ms"ONX����h͚��*L$�!��I�8|���%��TT-9��]�oq҇�X�[U�|���<��U��JȕD%ƥ0�6'�B䉦#W ��-~8:�f�+z�On�x��`�(4A��d�#f&����K�i�x	�G��<F�|2�_4{)��H�!5���`�;9�v�H�b�on� B�[�J���	��䨲�qD@@xP��).V�<A�������rM�pGFL``�
���i��]����F�ή�˵N� !�d#o��!I��K���@�왿�9�&��"f�X�t�f̖��	��o�Q>�����II�邬Y��Eʆ�E�Lf!�1(ƮI�ж�YzT�#LВHp,X�aӦx@�#L�A��T�Ʌ������'����b�.`���#3h�@�r=*
�i�5(�5z���+]k����$u���h�-�-C�ܩ�V�]�O�xͅ�	�E�z95,C�um~y�0�Z.?h�<�C�@�n)i���venY�Nڟ,;n�R\ws�D� -�_@ĩ�Mnf�M��'WNcB��� �zWʌ����wń2 �ӑ耮t������|PB(S8���$�!U�P @t��6J50)�"O�%�3N»>��<C�+f�-RT���9�4�Ӄ�"r4��R&�� @>��vd��=9掐�H�<2�A���"mx���6bۭa�Yc��P�]�<�DLW���*ƮY�B�ջU.I�I,� -Wz�z���qh��tnκ-�,� Ř���O���+��vx��A�,Ϊ	[B���K���@�:f�\���aR}t���Iu~d�s����Js��h���wI|y �j<bb`<�'���c�˂�Sg�-cÃا=ML `��{�'e@��V�։I�8PR��C�2��'�J\��f����zB�B*F�l C�W!O��1�faH� :6�:���1�r	�d�߲m�,rb�ª���P'r��y�����FLU�Y��z�ʊ�9��D(j���?y�ثk��8�q.�3�5Iv��>��Iq���%B��[�`�>�c�MP�!�8����}�'{��� �0H�O� ��Wj�g��(���ɇC�dj�H�=W8�ӕ�Q��Q���#j_���"�9%V��#��ĸ-�v%��)}�sB�<��Z�r*�Tx��.扯_�T	X6/�<KK��A���Qʓ]� �G�1MlR0��/S���e��dr����zם�t�,��Ã��z4H5{��ѽi���ɟj�ہ��W�az�ě1@������I Zj�Z#pD�9;4�J6�,�� ��2+�h!D�C����-�V�!�9#ن	�c�3���B*�������t��@;�#����]�q�Bpo;2c�P����]�uA��(��s����z8j ��L�q
�r�O����CA/b�N=��]�T�#2E	5�d���ɤtJFu:��	�'�f��E��	P�(P����$09������1m̥��Bo�mJ#�I*}Ҁ1�V��P�,RCF��&�(�"�p�ɓ(�R|)��3A{`ʓUKDQ�� �������r�4Z��Vl�	1Dsl8�Yw�51��lB(V�d�a��<��I�'�z}h����<� |!r�V'&n���F.AV؄mא#lqA�F�J�d�����K�r"���$	ƮG�S�<qt��0t�T�[���n?�� ��%F�~b)Q c�L�LU�0y6��s&B �۠nϞ��0�BPy2��U�V*�D��|[�lZ;]��a�?kT����M�Y�џ4,36�����ͫ�ħ_�l8���I�|�����
�'���%/�$�����M��?�`�f�cG�s���ə'^�����)����Q�*�<i�/�<���1}��)�'S�j�Þ�(�I�gD_*d��Эu0��A~A���剷J,�:��W|x���N�pq�L���2Ǧ+���&?���G�sKZ&
��q&���y:�0H��,�Չ�[��|��V|Nm�ǃC(x���bG�X;e�U'x�'F�H��%	r,���)_�Zv�+��J0�AsaE1v-џ�	�	�\�>q�p����;?�|���*��C�M%�M{��׎!0�Lh�^~���isf�1 �)Z�ؠ93b��0h�)Olq[#f�;X�H��|�2"��$;P�%iG-Wk.%�0�r~2�X��LZp�'s�1�1惭8>U�`�\��@Bc'=}�aܸ)�5�����O`j'���:0��Y#V�}*��X8�p�
�/�6!`�g��l���͉4��a9�cC�Hr����� �OV�Xd��`D�<���&Y,�t��ɭFm�邤�R��O�b�i0�V?��4�&��{$�	�'��ZA"G�G\�[���>����O�$��lY+O~�O>�+A%ȵa��Uc�ԁ,.F�g(D����u��(W��9l�ᓤ�&�I6b��A�Q�'�*�p�&�GL\�9�͞>	΀�	�'@Zt)!eѶO$����bD�� �'{�Ǭ�v�L0���?��M�'bP��,F9
.4���V�e��d�'a�1�0o_2�s�KW�X����'����
.H�@�d�78Ɗ��	�'-���E�P"D�.�af+1欀�	�'���h"��\��@�s�$ �"O�8��R*���`�,P��"O�m���6R��˄�ƥqֺ��"O���A�8VXT ���!<S|�Y�"O*�:u�Z)%L��T�Āy3"O���7��+D�\� `�-P���"OF=�)D��H��V�9�>H��"O��kP��MC��� c�8چ��#"OX ���,Bp�"�".�R1G"O�D��H04f6a��)qs��@�"ON):2#�3@n<���݌SP�d�"O�u�6��*a��5{�-ٯp^p�"O����oA�1'F��@^*D�P!P"O>�H��^�S,H=����>Ա�4"O~$����/~"��fƂ�E�< �"O��SaI�K,°ڄX�I��(ܾ�6��i��Y�\c�H�6�� �P�H���	4�-D�k�OַV�k�F.��5��ͱ7�bqsH�g��|��]�tʷ�GI����V��<	�/O;�d-1e��!����>s�r7�i����'�~�!��D�X��QٕzI�]Ys�Y/C��)��(��F 2\���('�ߵ�H���H��Q�0�z�Z�E)oj�<�"O��!���u6�e�I,gL��1�Q���{'����j��A9�q��'J*��%�@�
��%�"#@�+�d	p�'K.���R<=3��fE�����a"K��"ٓ�C�mA\��1+�h��|*�*��R7��Qǆ7H��`E�>O���-�>?�i"'��*)�6[� Ǆ'��[e�=�x"3PwE!򤖏I0�R.\�T'P)3 \��	�q^X�xńM�qwf]�e����G�$O�)8�� "qO�f����W��y��
�}�&��è��A0S����gOC9:�B@���[�"mI~��y"��c"���@�Ӗ�>��FG��?�^'`>$L��Q�o�,�p
 �6�`6��FAɀ��A	ӓ/0��7�E�Cs��A��3Wj�G§ށ���"��a�t��Ċ|j5Ȥ*Q'L�Q��Al(�Z�"O8��Sb҂
�fx��$���<��^�p���ړx�\��ʸ������g�π ��a
�>DΖ=q�$�h��Tx�"O����J��߬l�5��N�ĳ�
މ�0��m�'Y#��`>.��O"1OB�I1AWb�ۄ![v����'{F�aQ�Y-�����ȍ+y�Ȱ��C!dy����J�=�Ș�)̻i<az2i�&��}�r�7|˒D���-�0<Ivo�� ߬�V�˽#`�����g�,���I��2LD�һw�I���`��#͆�+�u#ӏ2P+H��'V��f�`�N�0A Uz��D��l��7�~�K!���ty��D��y҃U9f�P��!�){fV���?
5L����$+ �D�RK�ᓈ�L>)���j�����ʹ)f���H�F(<�ō��p�i��J��=����Pg�|�	��[��=�D�P`GL��w��?r��K�OCX��j��}��5r�(�����+��b eJ�ju2Y�*ݾ�y� u�"EA�=>���D� ��'<:���$��
DD�dD��r�	."\R�-_��y��V'[s�P�Cl������Dt�%���\ܓ:Α>�^�`��2���q�:�ӱ�\�|z ��\w����͇F����c,�:_�L��ȓN\���2 ԋ��5�ɘ}����m�T٪��؞cAq�h��������!I��эlǮܰgj�}5
���ڜ��w���]�6T �J�<�j��ȓM������M�=pL�&��݆�XH8!s�#�$-h�(��A$) ��\8��0�&L�}�)emU� ����IN�{!GG=#��Y�HI�3HB����bգ�!�%�����: ����)�9�� Ͼ82��7C�h��V^he�U��1	P�Q"r�W��Xd�ȓ!��	��G��!$'L%iż9�ȓ� ��Y�;��6�T�OV2\��'V�=�`)�54�j���i3C�J�X�'a<� ʎ���
 �
���'���3�X��u�
����!�'I�\�Ձ]�MC``4\+��[�'�c��Ho����	j��
	�'f\e�X����̎xe����'�,{s�U
K5	a��вogQ�	�'��!2ֿ1�~�c�lۨc�.���'��tjP ��X�.�!3�ޫ^��8@�'�v���M�*ffNt�CN�Snd��'�B��e�>Ev�sl����I�'Q|p��4$k`9���X�F5����'�ruq�`[
�h�Q�.��7j�y��'\��i�ρz�^8s#V))U*�'���s��]<,� j'�·$g�Ԣ�'�� �d��>����6��WC���'��q���Iv��LiX�'S�@Ys�!y!�U#]"D� 4
�'.V��,�氱�4l��Nk����'��҉��L���H�6�Th�'#���dזj�R�J���7��U��'�v�ʇ�Km`|S�iH�g�`�'� @F�1�d
�(�Mk �a�'�t���ֶwn��@�ν,��p�'�8���H�'D�@g��v�#
�'YlE{0��>. 0d��3
!�`
�'@p��
�H�T��4a�� �8��'�4Q�0%T�k�Аrԋ[.�Z9��'���DN�-F.�+VfU�J�'Ԛ� 	�Am΁��k9�	`�'��nJ;���C0�J�<��ݘ�'���Ǭ;�Pp[C��2����'�r<s��j��`�"��2�
��� �A�
�qIZ��G
��'AL���"O�����MR\5�P;
Nh��"O<�����/MƬոdF�J)d�h"O�t[bgʀ I"��`�-+�x�"OX-xP) � _�X�@dU�7@�w"O��	�2�yh��W;�@��"Oޘ��e�>&��c��F+*��`�F"O��)g�3�ne��%�Hc^�8�"O���E�*����'��9q"O�5 _iW��q����P��jP~�<a��˦cX�$�2��mqo�t�<� �	/%U���g����#�_q�<)�
�5/�;Ą�f��)P�/G�<�G�I�\y�́a�4�cA�<Y�Ɖ#2��I &䝴0:Q:��|�<iA"̫}�A���7��l�΀x�<�'�čn���z`/�@S��	e�|�<���RK�,:(��� �D�<����T�\[�H?�\� �B�<Y�*@�sI����ǻjr� p��U�<!B�ObA�֨_�F���h��L�<y�!	Р�hх��l�v�<7��0�,�J,ax�3�n�<I0��*�|lsnD_���{#Dr�<9c�"����+/hRT��L@n�<��O��?v8 �4d-ǀ[��So�<���\1F�Ll�k��x�ıå�HA�<��X�u�gd�*u�D ӑF�C�<�&W�V�87&mv�c�&�S�<!̉�pT�H��n��2�l���J�<y$�Ϧzr&�����N0�ݠ�Z|�<I'��`����C9�t)�� ����ppH��9J:�$�"~F�6鬉a����X����=�yr�y*��Z$�*?Z4��L����T�"�^MЁ"A���<�1' 	d�����l+#�U2�o�t8���	>^�`�9bC)H��ɱ�MȘdta��H�1�2��ēAd�YC2��*O}�9���"�b�Fy��En�q��+M��vd9s٫5s2�8��#x��C�"O�DMԌ ��`�7DZ���Jġ�c�P�h�O�zD�-����2�W&t��M�r�I"LvxvmI�y�a��z(8*�Ń�r����P�~ba��+��PP#�.�ayѦA���0�$�%fC���#_'�p>a��H�z��u ��*�]bUdL�T��ԯ4l~��	�'H}��ϛ]�pp1�A)1o>a���M@U�AΙ^�tb?ɐ!�ھ���C
��`b��3D�tiS]�E�- �\ �C��<M�u� R�T�
*O?�d������Д=�T�H�l	�Z !���N��d@���z���+~9�O�-��4�j���` *W�h�ɠ�`Ϳ:�@ܳd�'�DԣDM��K�4�H���(�L	X���z�<Ћ�"Oh�������{4n��mK�Qk �'�H����37�V����$x�T.�
ynD�I�;B�XX���5��k���`��U����,*��F|�&qYC�&�(��O���ia�	_�BըeL�Q�r�ON��D
,a����$�r��Ac`�T�h���H���]5�{��F�,��!�h��s��O��	��D覽��#�8�x`� ��c�G,��ڳ��"w�J�҆��E�\K�"���<J�JĪo�~�j�@�A"�x�񮊡p�Z���4���f�9Z��D/2Z\���?%B6i��Ǵƣ?aQ��H���p�E.� @xKv�	3CL�"������ �
�{6GQ�3;��pbI��y�Dp��8�C�j��c�ЂŔ�mMr��PE�>�{��<ف�Bt��pk4�ݾ. �HQ����$TGk�@���� kݑC�T��b���8��������Ҡ��c�d�Y��'7X:��Y0�#���8D��A�"�E��]q�#��`Z�3d-,;@,���?�ݠl�,`鱂P�($Z�8��Z�0� �5�[i��
*#N�T�.X?h37
�'�S�g Dn���×�s�P�(BAO9fzZ)84�K�^;`WZ�4�4Js�7� f�@��4�I)�!��$|@�W�	��d���*H��A��(Z?�m�2�o����<Ǌ�1
�(G���F�ќTE���W\�L��6T��B�>�%-��2f' I�`�w�ބ<˓`(I�ߟxZ6��D�x�3�l���E�O�%
`����6)�҉O�:�2<���*���6O� �c� mS.�b��!<O4��DE,�<JR�ݐM7E��%���"1�A�%V�����J_(��l��.���u�Ij��넭G�nk�-�S�E,/4p#�lF>�p?��o����MYw�O0h�|m���@k�$@Y�tG���X�d� $A�bU�!����#�ħBʲ�#s5D�@#�F M�u���U�'�V!�X>�&>*wi�pW]q�gA'z\��"�N�!p�Rc��Q0q`��O�	\�AU��Qȟ�d�>��y�AƝN�~��L�6.��uH(}�Մ�2��S�O7� �C�_�,�J}h����pX2�'��-���U���� H',O���.�Ew٩���7faR��k��C5h
���`/��4m֝�;AF�1�柄d+X�q�z|�Y�b/2j�����}����+T�D^xQh�&'���1�S�,�N�[L>��/�Z�dE���O��a5�
<�H�Cf{e��e�'�WƎ��c��2a���<1�e�O��p��g�#q'B��ig������u�Ds�O?7R�<�ʽ9�+�>i���Gg�?��I/n+�f�KH�S�O��!׾�E(��1�Z����g~B �.g`�p�'.NPPn�8i��ı�K%_<�1��$}BmǖO�`����O�Ģ�� ��S��"CPv	��Q�]dZ(�
��+�1���D$\rDȱd��.$T��[d�Q�'2\d�e$�O�9Y �V��A�!eT�1jB2��� Z`�EXw)ƕP�O�d�,0�P��U�V��tMi�'u��1��+<���*��:7pX�O����v&l�O>հ J)`�҉�J��gr�d�;D��p)F9S�&a��)Ȱ7  ��+7�Mȅ�'��y���Pw:)��� ��p�'�Vt���5��L $qZ�l��'dv���KT%?H0Bѣ�_�hQ(�'�J�;P)
c�|l��GD�~�P�'���� ���1|���Dƭ�%%�W�<��
�(X�}iSL#0��iS$��y�<A�^�>4c4,����a�I�x�<��섚\\��YS�Ԗj���Jh�<6"�H|��a!��in�E8���N�<���:�,�����<�D��`A�<)Qըh����`���.��D�B�<1��ܫ/|�9�!�5oSfx�q�x�<�F��LZ��E�D/�6��AL�{�<�WξA����Ɨy�f���"�}�<)���C ��K���E��{@�y�<!�C9E�xr��[u���f�r�<��($�:Y�_�EZ�j{�<��;,� ��;"4%J���X�<1�O�>������A�:4H1"�	Y�<I�� 
r����l�z`=Z�gNW�<�&F�rd��h��:y�b�Q,�S�<1�i	�F�Se��4}�����@O�<�t'J�:]x�ǰd�DuɄ�P�<At���fN�+��׭Dp�l�ƫ�k�<Ib��B�(���+31p����x�<�&bH���"ή:��MB&�B�<y��_3v`n�t��.iL��z�H[x�<f�#y"&�B!L9��|�<���ޭX�%3����l4z�y�<Q�%]�Ɣ v)R���\����v�<Q�]>ob��GG�x�.�ǃ
q�<A��J�z�3����N����7kXi�<��ٶ�����$2��(A��i�<Q� �[����Z�j� _r�<��'��ҹi��!#P1����m�<�F�3ڹ�6�հvA4XK��d�<0/44��`3�
p�z��A��f�<���4�b ��&�vD����J�<� ��
G��!ip Y�s8�'e���N�KX�h�b씎!���0�L��;�d��F�$lO���%�ԭp�*��#k�dḊR{�=��@V�$�NB�����sI�
8���	�#T���� �A�_�h��V�o[<� �L3�4x5��1J�C�-��D��-�39Fx� 瓝𚨀R�M6j�6�'�-E�,O�P��1H��U�䃁�wt��0"OȌj���j:Ȝ�g�ѭC���C�L(tx�|�f��}�a|"!��c��M��+>k�0��T�G��p=�/�6
�*=؁�x�9t#F&x�N�B@�Yu�Z�� a%D�T{��Z�5<~��х�X�ٱG-��ܸc��F�?�#2�U5Q��8!�u��� 4g.D�@��+�ʂ�����2�x���6
��y�l(}b�B���`:z� 0DX�v`x�B�Q	S�!��z!Y�P鱴��9���A�_b��U��JZa|�̜�K�l��L��Uʳ���=)�)�4H|޵�'Q���5hKz1dL��g�"�¥�	�'��a���-�%��-O�^�q���\+7, �G�d���'\���bƖ4�|3!��!�y�H�������* �M�y�*߅H�!��A�v��Bc�L�<ٰ
�4=������O��qI���}�<����+9�R���,G�S��а�]z�<�D��!"�\��L�[��0Ɔr�<a��>l�	j��ޥ5[��P�)�s�<ycOZ�[	�e����)?��p���g�<�TmG�~���CρAɮ|HN�k�<)��&v,�AV�@�G�j�c&�	{�<a�JR>lTU2i(Φ)��oPq�<�R�
�V=�bGDROĔ���g�<���`�j0Q' �#"R��t`�E�<i��D����J& �D]��NAA�<I�	�l��-y`��&�����d�x�<	"�X9*1A� :Z8�Q+Ʃ�o�<Q嬘�/LdY�alL5~yڭ��N�h�<IW�`op4����7���D�R�<A�&	~�
�`G-�0 ���T,�u�<y�s���;��Ev�s�<�A`_�v�B�i0�P:(��Ӧ&
`�<qď�5G�j�q4��8N6np�`.�G�<���O5�B�PA��ED�פA�<9ue�9�@d�ҫ�4��ax��U�<�u�$�j���*���"�Q��4!0��G�L�f�-T">I���6i�	�k�W�  ׄ'D�T�!��x\�uc@ꐳ9)���Dg)D��i�!:��	[���/�-"sH#D�أ��˷%�
��c�x]F���g4D��A�F�(g.���d�(iZBIS!.5D�B��=�V��5�V�Q�EY�5D���D���;�p��%o�`���>q@��W��H�<EcC�T�M��hBg��X�,��imJ���R��@(O���T��DI�W��7m�(h
���'%U�]�M����z6����oӦ�"�����ԧ���	-vm"u�AF���q��e{r瑦R�"~*2��I۴����R�@:6휖"B\�Ey��	ƻ"���AI�1�@��_�zTQ�P�W�O���3!$��B<���gQ�7^-X�{��[���'C�b�'���b�!��U.1�O��ڋ��i>a>V4��g�)|l�u2'�����5�hOq�����r$|��E��t�A��1U�b�>�O'dc>a0 ����)���=}O8A*��4?�CO#{��t�D�/}�𩈣s.Y`g�ϟ'���hL:5��f�������$P: ��)�p���8t�\&c<�y0��S�L�G�^C&�a:6�s��8u�{>U��O��~4�۱�̥mE�3Q�X�&��W3O�X�F������	[�@���mI-1^z)�o��s߲a��hJh���kY�������� |�bR���Q���]�Ƶ�3�'Čĉ�.�_�S�O]�\�ə|���1���,!(N�����5>���|���.u�`m�<Z��hC����(����{���Ipa�DL?,�ر`�`O'h|�z�̉���i~�r��)�)k�.��R'�L9@�)`D�9�PB�I\M�x�!GB X`�l��FCBB�ɫ8^�:)��pW�m��^�lB�	=�P�B~�������b)B�I�aqrk�G�>[N|��T/�)P��C�	!�F���l��0�'��_G�C�I�e�$�¨�<����É5JjB�	�C�Ҕc�g�>��t`�R�B�	}���'ŏ)��5�ņ��c`B�	�{ǘ�ٵ.J%B��1���\~*B�I:m���W��O�h���_,PC�I�%֨ɐ��D�<@(s#'�3/"C�	kB`��H;,�$��	cUC�	~<���r�E
?�P�aQA�|N�B�I%N�<\@C�O=p�zm���=e0xB�	:p� 5SgNӥ/��<�q�Z'{�0C�_��}Ad
iF��w�Y�?8*C�ɣ*H����*�J�8�&>@5�C�I�_TQ`Gȓ�Z���Rӂg��B�	T���e���,���,]�OtC�I9~���h��C����T0DC��zJԉWΑ�H���b�;J�@C�I>#D���H[��"Se��e�RC��T!<�5K�^����vՆB�?{�9�� �4r0��*U��B�	��0�"c�|��A'J�&VrB䉒F�I3K�I�j�jpe@0sddB�	���躅	3~�L�q���}S�B䉫wY�Hr*߉k�6d�m�1ѴB�I"g��K���"u��{b�Z:6<hC�I����n"��]�1�vfC��t{���W�ʎ$`�QqE��,4C䉯F�P�Q���pi�p��?�LC��&-�` �Mϊ1�4٘���y�.C䉟^-6�@�įq;u #��dIC�ɍY(��0�9O� J�ˋ��B䉪]_T�p�� Wm���q�(B�	�H�S!��[��a�4o�(B�	� �x	���	i�0 ��6q��C�	�0�<�+�J��7��� 1j0fB�0�t� ��5R{�ݫ��P.}MC�-"�B�)[�ta��b&.��B䉺4Q��Z>1�R���[�|N�B�	�@=�@+���1XH%����?wj�B�	3�ޑ��N�J����/��B�I�\�B0�<P����g��B�	%�l���ɾ �n<����1O��B�RE��A��T�mJh�4�̬w�bB䉘E��e���_�6�"tÅ@L�C��2\��Aq��>Zjf�o�|C�I�L
"�jq#8���)c̪	KFC��''BF,IǠͼ'�z!��\g-C�<G��9�$Q�v.��� \��B䉸*�����X5� P��M[�_q�C�	�H�T1�H�@�� xT���d��B�ɪJ����%e;aoL�rW. �y`B�I�ӡIW  ��P��X|�C�	�d�0��c� �g�`���ͣM{B��sHI;�J1�T�*���qi B�	2a�^���/�!7H* �u�yC�)� �yR0�/d�ܥÂ�m �!�V"O��R"_j�&���'Șz�%؂"O�P����S�"���f��.e)A"O����g41t�I�rE�h�nTAp"O T$JӦ9�2���#��X��"O���H>u2� N�T�T�[�"O:��d�^�!X:�Yf�ɀ9�P� �"O ١����%2�����r-R�r�"O�yB����N��#hԴ^����G"O��Sm&`:�b����H�"OXMW�E",�sg̉�U��@��"O6%�%e�(^,��`
K�H���%"OV�IPB��@�4lkd��1����"Ox���K(2�`�ڕ��JV�`�g"O���󈄫#r��gk],n��5"O��#�in<X˂���*���H�"O�I��_=<��aJ��G>@���"O�LYrI[�#޸�qe��71��98�"O�<��%�[�D��eЖ? z�"On�#r�F�hH�Y��^34<��"O(к�lZ]�Xq���Ĉ�6��s"OԬ`W��0 tH�BE�J�F"O�8����%<�z���12jļ�q"O@À�ƤiU�.�1,2� �"O����ѯ%m�BV5I�y��"O�	��c�/f_����8A��z�"O�H����*"+�9P�"���t �"O.�����E
�9bF"I� Y�V"O���*@�LƖ��!��zW(�{�"O��x��c~�����0c�l5�"O ����v����C�X,�1"O���Q�)I8�X��-5�4Ń@"O���5G�o�ųe�u�j�"ONXv�״_K��;��D�:h��Y�"OB8�6 ȷ)s��"�(�iN�j"OV�Y�S�I")e�̉o\mC�"O��� �0\���T���:8�/�!��B� vЁ#��(����!��a�tp��O�0�ά����8�!�T��:,˂L��	R�I�!�$���<���@%h�HDФ(װz�!��*��)��̐Z��cQ�ё@'!��Ê|��L*Ā�7b֌�Q����/!���)~�ˀ�Q�0k�>!!�x�����C�I�RA"P/F!�zKnl"�}$ъ6����!�$�14#��X�!'8b	ru�P/C!�$=
T�x;j�6Q0|��ߩB�!�߱��90��.}��|A�4�Py�E���x1�N��=z�z@Ԝ�y҃
9\����ǎ�1Ҧ}�m��yr� 3J���fލ&�%����*�y�+,� \�%�$�:q؅�
�yRQ��	�L1~Ezu ��yb+ػ�2��T@�p��4�I�y2�P1m�P*�G�r�YBT���y�I ,?����8Yu�@�C+�y"�@ �U�"�$XZE����Py"��,lF�#�E�Y�������S�<�d�N#!BH�EK�5��e��@�M�<9���]��β��X��K�<Ɇ���W�Fux�l@+6����O�~�<�DNY.`��ő�f	�K�z��I�y�<gH�B��9�,:j��YrH�L�<� �����((°b���#Z7�I6"O>=h��
Y�!3WjY 1>�x�"O���E��:�4�G�!Z'$e5"O���φa�&E���!�m	�*OF|�n�T��%)���K�\X�'A�ʧJ�%)8Ȱ�Ƒ&4~��'�����W�`|������Q�'��x;�@�l����g'�	
��d�	�'�l��ЃZ�V��4'�6���S�'bh�!�ț`x�I6+Q�0�����'�q�+Ee�� z]V(;�'����J'5���lo	���'�`%��X�ڔ��Ya�����'����`j������
T��� �'< yk���:	#DD"�K�0��
�'0�u��$�K�H��B�M(�o@M�<�wb�	Z�dd!��6]�*��T��H�<�4��B)��g�	;Zk5�Ec�|�<��B�T��P�s�C8�Z���Q�<��$KA:�Ȓ֊~�X\	���N�<����p�=*�Q���|� *VL�<�7ˉ�9`�S���Q�O�<a%)�'r�
�aٛa�r�E�<a�搐)x�1J^�%V�II7̀Z�<)�I�k4>`3%�Tp��� d��R�<A"�M��x'��R]B@iqiBY�<�p��9W��a#���|&�}�s�U�<�c�AD�%�b
�+�� �MT�<A"��*��#���#9�l�k �.T��K(k��X�ժЛ_G�Aڶ�(D��p������ӑ˜p�]I��%D��Z�`E�~ia;��=R����Q�#D��ZcfY���;�!�	v���s�"D��S�* <K����JM2�hj�#D�hy�g�u8xͰ��	+u��e�?D�����."�&��B$ǔ�y2�=D��!g@G�Eon!�׻2�PH&����yrG�0��D(f�ը~������yB��c����'
�R�)��X��y��˟��� ���L�}aa���y�`T�b�*$sR�Ĥ"yִ
1���y��4:��h+���I��I��J��ybnH�¥
�;E��ݪGƑ��y�#Q0�S

�{@p���0�yc0%ṑL8_����i��y��uE4*ޔ�s����y� �*`��d��-HLQ$%�.�yRk_wk��S2b�̄�ق���yB�:�xd���򈫂�y"#�i�`$��O9|����&R��ybܺ6�Ќ����,��X��喷�yRi��R�p��8n5L��r���yR�I�q,�$��Q3p�@��J��y��8x��dyV�ȝ<(��Ф��y��Ʉb �BRiH�58������y"i�����k��0�q�/A��y�G>�͐��[(�5���E�y�ㄧs�:I�v��Od���ʟ�y2��-�D��@��I���(�*��y��"^b����؁luĠ�	��yg�D���C�ǘa��!:�	T:�y�f&|�@A�F�Mz�ލ�y��+eR�m�.� $y"dT�y�%�|��Õ8Q؄�q�!�y
� ���/�F�b�2�ʃ�O�a"Oj�Bb�!M��$��k.pֱc�"O���,�%F�`1�� �Rk��"O��N6al��S'�Rbj����"Or���B+K%H��BFU:�j#"O\`QA�3k@q���!oҔ�"O�m"���p/�]iZ5V�!"OX�j"C����E7H�
���"O�b�	   �