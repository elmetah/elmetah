MPQ    ��    h�  h                                                                                 �J=���������L-O\v�!��=���E�[���d���'����M��8��%��L�=�l�i���2[,��*��B�p�83�w0��S\,H���2`��8�:M(<��:��v�T���{�x����p�������?��}�_"Lk��y3&hGYT=�u�
+Rsq,�)Q�\.��O�|+(Lz�ٓ8Ęi��Ez�����a�h�p�@�xۆ!�HV��| �1S6���$�'|�,X��s�1K��M�E��^��ӿi���4,>�'����MRC+�G?��́\�Dgf��X9�
H(AB��^Ȥ� ��^�9$��,�m����a�TC�0�g�	J��%�ɕ�s4���>ʞ+M2Kl�Z����(*�L#�x��:T"�L��u�y�x� A�R��!26w����Ak��Q��}�Ȫ�t��,��Q��
�P�2��.���1�;�ۢQ��?}��#.j�����n��@Ә��u�\r�M��(���8�ai6v:A�.�oЩ��C�1�P��n+a��22w-җ����_=Y�sxd��^b�żzߏ�Ul������!�__H����p,/�rt�6%����K�UЊ
�N~���P��C$�k|w�F�c���\ܭ'^#��v�ܭe�h<�pm:�8�RϪ��s�Շ��`c��p�΀rp>FLH�gJ�	v�E�����)�&�������6�|��O8��	J8\�6˴6il6�;si����_��V���*���l��_�y;����E��H��{ >�."���'�8q?�D��^��鰖�fX���a=@'�?���4��D��Us� A�]al��SY�j�m�DǗ7�����Gb��* ���f����ԭR�GI� 1X5B:�y4nY�0At�N�?���#ez/�d`x3�&0�=w5kVĘ���J3g�G���j ����g4:Ke��K���o]��#����_!SXK0~k��݆�F8���N{C����3��E��_��<i���4=�!ڸ}A˜�y�2b��*�:��c�ú�H��Lе]q�nתc�>]�q������rS�IxK����	S@K�g֜~$��M�;���`��`~��mkt:)�r"����̀�;��ቛ�4��p�H�'���0ڂ���5��цW�'�^���������+E���E\V��ɔCr��Z�nrK����T��:�L��PJ��bۤ΂����|s������6Xv=OZ���N���,ͣ��{69������X�!Ry/_��.b��lA����+FF�%y�>���@+$�ex"�:N#|$�o��K&���SX#[03,�2S^V�1��ڈԐ�J��)�(�h2ԁ�fc�7_�h8DGϜ��"��QM��m~�h#&�!<t6T�sG�ߨ#Z��re- 0������
�ߦ���WY��Jhb��HT�~
7�@�>��O�cm޿��URbt����v?)�?ENXb��j��1ri��,����#���zJ_�?����J���^@�1No�@�a���H�V���,��ը�֭��zq��jL-Ln3��L�������Z�=�I��#��V>1��.��t�"����ߧ��4޺�sm���	��\��xl�.0UI���cՍw��k`�=�R̈�9$Gf����ف@���s]�����i���>���Y~�.��%E������z�^�v�w���E<P��W���-nWqO�����";
Q�n4jf˕�����''.~�l�����+�\lm�Z���ra�I�ާg<��y��p���$�lh[�>j����빷FT�u&�FȠ��uߠ�-;G�uoF�+>۱�|ܘ��rV�{-�w���S�4��2��J��Y�χ��j[���Gf�h�ڎ@H��B
$��9��������n|�ζ�j�x�j��nG&G@�4.Tw~���.��a���}�P��F
�-�"�F�d]��W��39 ��&0�@���=La���{ii{�x�x�7���1�P���B�����,P
������9�B�UQ�R�B���8������<�I�/B�K�ܴZz5Rgn�9�u�1���W�Ai[:PX�j���Nf^(!З�-�f���9ƃnS��J\���� "�$oh-�vm��W����<����;�y���
2��I��>D*��w�}�zP_�V(	���]>ap= C(es�9������vUT��h4��DrS��Ö=_f��O���C#�6`��o����K
����W��K��yDU��<�\�� ��~�j���l�K�����vq8�9�����p�o�i�8ݾKla)�j(@��z��&D�d���V��G���x`��z)�H-@J5�b��؂jqVwf(��o���#\���}Nt���I�-־f�G�EQ�HqD&}wB���Z5�D���Y���_k��S����x�l�P}[R�v|�[�p��K�'.[��en߈��F����WH	&Rd�M��Ng/>���qϡ*���u���� 2��XtX#�gN��C8���4�P�`�(���*��ݭ�,y���\�G���M�`�"�MN/%,	���<k��w��$Y�I��Wet{?����_�
=�L��?ϵ�Ԓ*j�a(�e* �o�iY�p�PQ�\a`��q�:�:v;��8d���-�EY֬|_��l��*�o��!U��=�̤DC�ׄ5�uy $�S�Xڨ�wH�B=`	 �����8)э;Y�)ʣ-8�%Ƕ6�5N�l!��ȃ_���l}��3��^YAD�ަ��f��#H^�o��pѢW-���1�����蜁�#]�d
؀H�@����Qe�b�o��w��:c&1� ��[��,�����v��� "�:�H��T��qg|v/z߈��s�%ԟx_ǁ�#��h����ʚ��u.���v=�&�-Y�诇�fF)k���
�q��3����z�^-�h�rO�j�v�0ߩ�I��+��Tk�Ro/5j�v��>�"\�{�6��~ۈ��`�Яbؖ#�zk�k������>ZN=�Fs!�ۇ�6��g6�6h�tڭ̻t�N﷋���ם��,h �*�lB�3>�sQ~wˈSW�Ţyc`�E\8'V:�ƃ�щ�����A�v"���opM����$?\�M�x�L�9h�ȩ&cv\Y�K�u���m�����,�n\i��O|��+#F�zO8�(������
ũ:?a��p���=f�|JhH�E뻗)�A���I$L|u)*���1���M����y�c�N�h��ؽ4g��'5t��R��EP��>���t����9U 3H�x��7^#�� Iz�T���ze�H����׻T�0q�b�	�%c坴��?�����y�m�A��bP���S*����32��U�0����u��2�b� ��X����6�!���Hk�c�֖�ƍԯF�,Ov�����rN�D���\v���ˢ,�y�z)׾"��2\T���m�C����הFM�8��r����v5)��� �d��C�[U����n~ܬm��ȑ톂v��O�.j�dиpbv~z�{��/j��*����!ں�:���pG/Nr�Í%�J���{�%��NyP��G�������Vw;QuFq��3[�H$^0!��<� ��<�F�:>�QR�sƔ���h3�c��s�)?�p�ςH�(J�u�߸����V �&Ŷľ镀����8O�)B�hl\1��Ѫ#6°i��=�3�2��1�*u��l��g_I�9;�6j���HK�� YtZ"7�"�Mqz�瀏v���X��бXJ�e�|��'3��^��4���bؠn�5A��]�H�nYC��28H�xD�72����db�� �����p�f���-	�I R�XКn�t��n�z0��4�i3���� ��C��kPd�;��!gFT5& }ĳ��o��"µ8��#��i
:��<�'[Њa�Ҟ>��`�!��70��S�F�(���?{^��J�A�lg]� �<�mN��̕�|q$8ĩ� Tǚ�;����u[��õYK5���pk��/3��D`]��=�#@�jM�D��z�!�w��S[�9��p~��f��Z�EP��Y�ɻ���Q�4tUīr�����̻Q������^��#��@�ܶR�&>#5�`���X��S^�/>�h�>�A9�+`jd����V��~����qnm��\Ƚs��L��J�x�b���	-��%�rs����j�E�\?�X���Zv)�g�<�#ر64�v�_聐�8m�!_*<N.=��l|��Į��FAHByQY`���b$��"���:��|_��o6:�K!�D�1�X��0N42�i��{�j�_���J��G�^��h�OہVJ7�I���D��՜o ��,Q�&�m�9��B������T��xGOSl#U��r��0h�^
.���Z(Y��*h��j�CT~e(@��m������ޚ���T�t8@� �)\�E	 ���	9Ҭ�����,#�p����+Jw�� ��ߙ?╁��9�1��@@v�6��[�Vt0�����J��Qƨ�U����oL	����*�n�K� �u4��n����Z�l(����c"6�������"�"�m�kE	O��u�s��.�H��c����eƎx���$�1���z��^���]Մ�f��㲚�I������$� O���;e�5g������}E�E�)��`�pbn,:��Ȥ�t;%��;f���<J��3�~�W̱S\,��	�\�OuZ�r<� ��Z���ӃtWA��NQ���hv��j����n���&�	�F���������b��o�[Z>�܊|pԫ[�V�|��!8�@34p�2< Jg`^�
�CC�[��{����h���@cGB�u��/��4��אwx5���x��t�K�G���`�TMW��Au.� �aYGP}�UP�@
t�"��d�|&W��34M%����@K8�X����͟�6i��xJt��2��6)�P�����|H�>O�s,��(��}} ܦ9�dWU%;�]τ�f��Ԗ�<.\/�˴�jEZh��`Z�T����q�2�A�9�P�v��� fuy9(�S�H��x4�^����V\��k�FZx-~�q�
>������dH̒�6�u��+2W���֠'�YV�Ll�}�����K(�w���I>�i� �L�s��k�p��Q� ���4�W,�?�0��$�������KzH�b��quOߖ,���o
N=QȨ��fA����Upa�� ]�~�����'
K
m/�p1vLh�t��%�k����}�yYl|��j�lk��Z�]���	ٓm��L���x{�dz�ry-�|ɝ��ӱVr�u�a�l�Y�w#w�<x��NO���ҕ��ȩ?f����skU���DA�B}Z�Z���*�p%\k��׺Sӻxd�P�o�R\_����_ɰ�]�.VƯ���∓�����W�*]&Z��d8�a��{�>ۤ�q*I&����͝k�2s�>t���g�yC3��b�PN~�(���*�݈1�y�� ��F�B�H�'K�`�[��h�_/��R�l�<�%ݔ4�b�I�e/������C
��LY"?jvT�f�jyI(@$ �>�nx�KT[Q� �`�%B�5�v�C[8b=�����և��mFlCjN�j^�!�4=���̿�6�Rt��PX�$'��Z�r}�B�4B :s�4�ڳc{��)iP8q�B�1�Nl*q��z����+��hp�)D|�&ƾ1w�~r2{�w���Y�����1������@��S�_��;-�[����ye�u�3VTZ%Ď5|�&�\\�ʙa[�i����լ�����)�t��U ��,.t|���zZ:H�N߉��t?���_]��b�ElD��N�k�=Ĥ��h`��Jv�fA������,�z3�i��O^�a���v~�{�4v���_�T�eR���j�X��m�� �{�[��$ֱ�WFv`�jybSt ���|�C�>Uq֡����UsQ�g�^6C9}tC��V�N�e�l�,�p;*�,3Blӄ���wf�vSR~?�cQ`q)(8B�g:C���6���+;�D��q�Ů8δpA���j�?��I��lLፌ���X&^��Y
z�ur���["\�\�\�O��+`�z�lp8����7;��ńɐa:�pMͩ�"m���KH�U?���'����$�{
|F��ٳ�18BMD[�ܔ�p��
��4�A'��9�pR��h�j
���:HO�X9���H^���}�^~� +�o���~E��#���4nATy���]	U	 >�%!*��MS�y�F�T�V�m���+�����*P�����m�ppg�B*�u�{��� w����O�6-�#��Yk4�2��=|�~�����,�-��]I�$J��ǅ���#�1�'��T��`�Y!R��o��n �(��N�R�sM����S?4��2�v01Q䰱�yaC�e�F�n�'��¨cq��}I��!���Hd��Jb�V2z���#�*uZ��=�����j�pbO�rj��%��������U�Nt�e�AW��!��a�w���FL���nTt��;9^dڑ,����q<=y:��*R�\������Cc�²���p�y}H�	gJ�����Lՙ7v���&��$�i��[�F�_�O.y���\<K/�lS6�E.iK̅��CMV���*P��l<_䖒;��܊�pTH<l t."��j�ݯ�q�ξ�*�}���8[�Xn�˗7c'�M��9�4?[��z�i�&Ar\�]�O���`�Y#��D=~7͔�Q}bz� `�'�[��Y6���I;��Xk��o,�n�0�A#���`�5�gμ�G���d�5��R��5�h��FM�@�����s��P�뜋<:�����Х����؅;��!�0�� ��@�F�$q�4{yթ�ŧۦG�5��}t<7�>�؄���(��f��N�(�q��������bFð�	�{*�+��J��Y�M]v���^�cHÆ?���ծ�2<Sv�?�]]0~�!�����j���r���p�Ձtp�r[�˕�������b�����&���׀�\󂡧�5�����^�]G�^��1������#+{�j����VuVؔ��l�AAnh�]�.�L�r7Jx�b��ؤD�l����s�#��Ū~���X���Z��{��W鸾T�6/��κ���Κs���_��2.rl��=�I�+F<#y��T�X,�$2��"r*:��|�p�oь1KJZ�l��X�%0i\2I���VGN�PU�'�����(Zh��ۜi7U�o��LD��p�
I��Q�m�E�����������T��2G��g#P�[rڽ0#�.G�
��ؽ���Y��h����>�j~�9 @�����y��u<�v�tө����x)b�_E��I��g�'�����w,^:��H���QJ�i�s��C��o��Z�1Ŀ@���ҎCV���t�a���o���b�0���-L�h��(e�N�K������?��ٓ'̺��3�����"���N�?���n����m	Y	�\q����ntJ.�[��e��c���~X��YM��C�$}��x"�7�F�Og�Z#�_H���[�AK�d)��y��W���������+���E���W^^�2n!���_��;@��d	�f�>~�$���]`~�ȱ��͡��\�Q�Z�1*r�����{��K΃o��&9P��	�h��<jxIm�@�-]Mȫ�F�,)�+��a�&}��o<7u>�'|Rů�F��V۝��-b>���473 2�E�JBV�E����[˺`��]hLh�@~�B �����6���D�r/ضZwxk����G��l��T���7�.碒a��}]B4Ԗ�
�^"u\d�NXW'273/����@��s
d�_�z�i�x��z�-�c��@P}�W��,ܾ�Ne,ƺ��0m���N9C��Uǲg�xC�.O/���S<i?/x&���Z�4��x��o�3�'+��`A�7nP�<��y�f��(����c���:�9�o��\1���!��'-9��%D5�vtg��\��ѐ��Έ2����Z�t��ǀ�}����(?~�����>�� ��Ys��`��,r�,Ӝ�Y��4:��:���x,����ڽ��$��=쬪��1	8��R0
���c힠��oUK����} �U!~���f,���dGK%
	��q!v'�4��hUK�<�f�Q�CX�4�Wl�6j����U�Z� ��'�>��u�=ɟx�J�zI�-�uT��W�ظ[
Vm~�	�	�#�4���KN*1����c��f����α��GD\�B~�UZ�@�YЏ��k�(���D�x�tP��?R�ŭ��;��ᣰ�'.Q�3���N1��(W-=&5��dsHL���>�lq�B�PD{)���gm2N�Tt�3fg��C.�/���	P	��(ؖd*�q�c�iy�(��RQ='Z��h�`�$�Ӄ�Y/ӈ�G?�<��������ID�ce����h��U4v
�wL���?W$�Z�jԼV(�� ��_�õ&�Q��`+qJ�0B"v��8�˺�P�;t
�b>W<�l� ��e�!�Y=����<��̓c�+W$b�R����m�B�({ ��i�9���.����)@N�8V�,��Nh�S,�>��2��b�宅���D�^ƹ��ټF6{��ꩢM�p����7�d�B����ձ��#v�v�t�7�e� *n\e����0�=&��7�E�[*�������,�Z6X�0���Ѱ˔��d%|�
�z�"�)�����Ƿ���vi�HY}� .���G2����=�Pg٣�H��>f<͘�m����G 3�Mޏ�)�^�ki�� ��jmvyj�����š7�T�4rRetBj�Zˬ�\��X�{�Ө�M���;`%�b�q���̱�gZ��l�>P�����T�QCal�^g
�,6��t~`��ɈN��v9g�c�E,� �*���BG؄��Tw��SMW���IE`,-x8],�:�c7�l���'���B�lJ����p��Q��`?Rra
�Le�J�?&Y4�Ye�(u-�8�=��gⳒ\��bO�`�+��z�8NR����X��_x�au�p��'��2s/H=����5]���oB$�|����ԃ�1\�M�~ܯ�%�D`k��4ݾ�'k��3RT��x��Y����Z�9�6�H�lƻ�x^ٴ� ��?��|��0���X��o$;T��X:�	[�%�|:�� o�����/ݳ�.��+��ȼ*�^��ߏ��.�½�u],�)ی I��@6�N}�HˠkO=��Y
n�Y^�%�),�Ӟ�����a�%���ی�d9�������Ì��J����:
ky��w0� �y��9-Mh|��,��2Ǻv+Y�?؂�ڋWC��6�n���㺏�p��x<i�p�eդ�dC�blOz��C�0��������pw?�%�p}��r�* %{�����#�[+�NoB0���r�t�I�Yw1N�F'���m^�~|f^�����{��W�<3S;:4e/R`eV�$����j	c��-���poC<H�JZ�� r�r6����&�j��(�@���K"O��b��\w�ϴ��6���i�ZZ��Ҝh-�+*+��lJQ$_��;��V�2H�� �ة"-�^ոdq�ʀ���jݖ��X�c�˲�')���l-4M�d��=2d��A�1<]����i���Ig�ފDxj`7h�B�2�bՌ� ���#�M�\@y��TvIv8X��j؞nj?�0rص���E���Η�@+D�d1#
�5���5�#���»H~�ع���2Y�[���:\�	�|`���ɊҔ�]�i�!��0O�g��M�FIa�,6.{���@��"�i<��ƾ�\�2 \�)Ӝ6h��T�������Q+ë��}���沨eJ��u]Q9����)�b?�:b�0����S��-��P�~�tK���C{������q'w��8St�Z�r�W�����1ć�RSU�������X�A�#��1�5�]��73x���c^��a��Ѹ��+����xb�VP������+inc����O���DL��J��2b�⿤�5�[�s눡� ����>7X�rYZlw�m��L��Y��6*Ȁ�'Ԑ����o�_ ��.�sl����?F7�yҝ$M="�rj:��|�{�ol��KL���XT@�0���2���1���kِ����I��uhc��۷��7�V_�9/D������r	Q^�mE������������T3+�G���#Krv�0ޚ�IP`
$佌�9YA'gh31�9��~k�@Ezx���\�i��P���tn3���LO)��E���.�ҢY}��b,��9��?��'J-��p�k�#�|����1��@� ����V*uI/������GW�I���L?3i��F	$,��㬫TC���7´�d)s��R����N"���	�Q��uú�ޫmZ��	�Ռ-��i().A��� #c&�m�������9ȴ$)����ْ���
��0�(���ɚ��=�|�o���9��d��.⸫����"�s��E�[���O�4n6@`Q��)%;[U���#�f����_gi����~��_�	�3�\�\�s�Z�Wr�Є�����8��j��ҁC��U_h��gj���Hlc�h��F.�F��?ކSn�p��|�o�2|>l��|��c��VV��s���ĥ�6T4R�22�LJl����yh[��a�X�h_�@��B{x�ʐ�F;��~}m���-�x&���ܝ�G�|�G�T�̄�ҾX.�D�a�}O��:k
jD\"P+dA~W�k3*��7�e@�G����w^�Uai,�Ex����(�}��wwP8!��)Q����)�,����|	���9�	�U�`��y��W����<�#v/����Z�<��^��;o�XХ�u�AV�P)"f���f+�p(R��~.P�n!M�X�G+\�(���5�w-�f�@j��]��u�B�lL�	�!2�F�L4�ȏ��B��}�f�Z�(ڤ⦸��>r� t��s�ͽ�f�n�B)ܔ.�4�Z{�5a`�ӐAn�j�����A�g�1����������
<�h_��ņ��$�U&���S# ��r~�T��؝j�K@Ǫ�f��v(:����]�a���z(���Z�l��dj����kp�ĕ)��5e7�	/�f���x��Iz�?�-�;���:�S{Vh:e��F�ϯ�#��n+�N��H������f�|��)��y@XDwXEB�zZ����K�I��]k�z��	�hx�BP���RR�h�PQ�!�r��.L�3�vC�	^��!(W~O�&H�d��J��>�T�q��}�4D�aե2)ۚt	�ogvBC)]��yP�$(��*֐�>��y7싈�{�8�G�ݥv`K�Ӟ�;/�֪�"��<�ʔH?Y��I�_*e�vm�T�Ђ�
�6�Lϴ ?�W�n�j/PA(��  ��ځ;�ƀQU��`�܊�+!pvL��8�U��#\�X��=xe�+�ly���`��!f�}=G�1���U�H���vm$��)?'�hGBN=� ����TB�ک8t��V�){S�8���'��N�ʜ�ί���~��mL�`2��*/D��Nƴ'��4'��0���W¢�����1��rQ��G�7ujرd#��Tʲ���e��5������+��&B���@�[EB���{��x�ĕ5/�AP�,�����z|�8�zP�'�b�P��R�j�ȭ��o̰���`��a'&=z���κ耳�f7Ϲ��.���i3�Qu�E�^��ќ#��;�vt7)��.%�\/�T�#�R�Fj�|��6���	�{�kL��侈�+%`#�bI�]�ű�l�y��>K��WZN�Q��{�g�6� t�Ӫ̌�?N�ᭁ�&?�$,��d*xs�B"<M�$lnw��SHP'�b�`�PL8x�:9b��G��br�z�g���4p~~�3WD?�`�<�wLW���^&TïY�6}u�1�wf����\{�OM��+��z`�8	�Q$18(�:Ga�Q�p����L7H����|C=����$��=|F�0��s�1��iM�����ڿ�n�_�4z'k���R���3K�96��0�h�5�R9�H�K*ƶi�^4�� z�������t<���ӄ����T���S��	���%��δ���o;�
�;��r��ج*�,�d�U��M�8Mhu8�Fd� �������6���]�kj4�����4��`̔, �h�ߡ�����u�����'�#�����+Ƭ׏���Ide������m��H�rMCN���9���{lv&���tЕ�qC7�~�<In��N�Ӫ��?�sO���F��_C*d!�Wb�g�zx��A9��`j����1��R��Yp��#r`�%Vcb�7��� INj���X��/�^�w��F�_����ݫ^,��⶛�Q�	<N�%:�^`R;���_�96c� �::np*-�H,�J�[>�p�ޙ����'D�&�t��eA�Ѵ���W�O$xu��\��c��/6���i��K���$`�*��l�� _�;������1H|1� ���"���Փ9�q+�	�`} �	չ���.X{y��ͱ�'�t����4�3 ?_ҜA(']M/��!s�Va�	�D��7j�3�b0�� ��M�>3H��Fȭ�*�I��bX�d��e��nŊA0-�죺}S�+X��rf�f��d�F��yWW�5We����6��ڳ��G��M4�/�:�*@�7-���-���N��?�!?a�0�F��z�F�-,�+{�Sr׻쳦���K�q<m;��TH��'i�Q�Ě�Ⲗ�o�&T�����æB�F�СT���B��O>�],
��YC;���5��P���S���Sdt~���9�.�;��(�̟�傼�t�U�r�ي��J�l���cɛ���ܥr�Q�-	�����5o6��r'���@^����y���r��+�}P��VWV+>'�/������n^s���c���L˾J�!bt������k%s���{�����X�mZ���G��b���P6%��pv-�D�U��_�\ .���l-����F29ybh��Η�$h��"�v:oM�|�fo�K��"�=X�0��2?L���e�ơ�]���צo�h�����7K[y��D3Zc�@��Q���m �B��[����r�Tnw�G n#FU�r�\0��fdyr
�Q;�g�zY|~�h�V�4ܬ~v��@ �S��ߧ��+*�Aot	݌��)�)q�E:�A�I�]�<��|^,���A����ØJ�<�+y��0�������1:�)@G�@��T�V�G���ŋjW���;��К�V�~L���݄�)�||k����5YL�B���i�r��ؾ"G�~����! �v�m5�0	 o<�W��d�#.������cA&e����K�tl�$�TC�і'��y����ՄK<v�Uqǚ���ܷVhϚ6H�-F���f���⋀��E�:W�Ͳ5�P�nk}�%e�Ո�;v�ɗZ^�ft2���,��7~����d���j�\ص�Z}1r���5k����eX^��m��eh��Zjn�.#Lֹ����pZF�82�ᨳ��p����o2No>G>|�q��|4V�?.��B˥q�*4mh2���J��͌���-B[��~��SBh�u@��B�)���q����)�zHh�ѶLx�1F��v�Gy"��T��٬m�N.��aj�3}�{�
��
��"+b�dIS�W]�w3%�g��!?@|���H��	��0C ig��xb��#Q4�G��P�c��D���v��_�,<�+�f�����9��U=.����$���e�<�V/�;��Zyo�>
w𥫒��a��XpAU�rP�'����xf���(�ڛ�����k�����O�\g���r��g-�qV�[�	�lg�Ҩ�0}/�(��L�2h���.
ȪH�ʽ	M}^J�K�#(u���>�" /{�s����Kמ�Х�Ϙ�4pW�0F��.�)�ɔ�꒼�ɪ�j?�"u��g"J����
_���D�����eZOU��H�� .E|~������X��K[���R�vݷ��%_��V�\����-�ݪ�l͉{jov�F�~�пͷ��Z�@��]Iנ� Jx̐�zVT-�!��Nz/���Vc�r<$��v%#�P���N�2��:���f�#附��4�-D���Bt��Z�}�����A�ak�쌺d�x��P�kR͔�_7W�\F5���.G������+�<�yW���&�ٸd��]��yP>�\�q;�ٍ�	_K�b�2tDĭg�U;C$0��s=(P��(�&*��|���yr�ψ�Ʈ3C�8t`nӹ�/����D�<W����=I��pe`
��3_�K� 
otYL
�?;x���j��(q � ;��U;ߵܮ�Q��`ah�& �v�~x8P��>�1]��]�:�l���[\�!���=,������B�ᴼ$���ĠA�c�lB�q� kR%�o�	�$��@�)�x18B�E�"L�N*�E��V��XS_�;�.�JZ�DM��ƯRP���/���䢢C/��\q���H��Tg��us���l�4�����{ezֱ���+�A�&_	&��o����[`�Q��t}�f�І��������f���]2t|��z�Z��A�ԋ)��c��6���۰vڈ�V�܃�=U��6�f2�6�#qO�]A�3�ut��X�^�y*�^X�ֽ�vo$:�E�S�G�T�2�R[9�jj���q7s��.�{#��5�����2`>��b��8n�WX��l>F��ֲ<���~	�`g ��6Ԡ�t�f��'��N�/�,4w���T,Ԁ�*�FB�~2�_
�w7_RSCi��t�'`���8��q:���"�`���k���b�I�Dp9MQ�N�O?H�FL�J2����&Or�Yőu�������b��\U:TO荰+n�z�8�8����Ͷ�7
�6&a��p�Lj���H�DT������a�{$8�u|�[c�ʃH1.Mu����b��:k�:,&4S_e'�R��ɧR
����Ts?꫉���m9A�H/��Ʊ^^�_Z 5�������g���n�����TJg#�N�		�%O���&���-��HYa�aEX۾X*a�?����
�³�u���b HP���v6>�p��
k�� �O6�v�ԛ��,�����sZ��}�04�휊�;Ģ�	��f���*�����	��+�Y�-�6,%��^DM@��gD�hP�v!	
����P�CRD����fnr1*�Y�4�u�n���&ٮ�!�d<M�bb�]zSL�||F��닎�D�&�Ę���p�o;r�#%1VZ�r?�Б6	Ne��泚*���'C�w'˿F�8�� �ܴ]	^
���=�[�5�<i�7:*x�Rצ��e���!=c�ز�x�p�6H8mJ��n�K�����&��l�z�:��I���O�'4P$�\�Y�=�6��ii\cw��Z�;��Z�*�l�;1_��-;~v܊OPH7�� ż�"#K�n.�qf}���`R�I��X6�i��t'���ʋ�4ðs��"$Z("A�<<]��������F�T]D7�}��T�b�� �J'�Y�J�Rm#�� fI�V!X<=1�`��n �n0�eǣ�+���ɥ�MD��Ndg�\��g��,5�����±�_ڎ1�$���d덱�:�V�������Ҋ����6�!z3r0�������F���-{�¢�6?��.䆵�<����l��$��l���5�qB��a<@��á%���W�\�ݨ��Ԫ�&�]	��M�����0�H潖�c&�S����Η�~k��t���[z��}?�'8�=`�t�p�r�4��\Ļ�I���U��H��7iͨ�;�HƂ�5J/ѭ;h�.�T^��u��ye�-`�+�n/�nkV↔j���a��nYMY�nX�_ROL�J�6}bO`^�������s�n��*�H��X��Zb���AI�S�h���`6 ����妐�J�ٳ{_R�.���lh���%�F-ty����}�$�7�"��N:J�c|K�Po�DDK�Ú}�(X��0��]2�׉��י��ː� 0�˹�ʙ-h�~Z��b7��bTe�Dn���ۂL	�VQ��m�y���B���#Mn�T��G�a�#A�r,M�0T����
�޽B��Y���hi�W�/�~�-@���
[~����0|��t�����&q)skE����d�$Ҙ>G�Wki,�����|��J�]�+��K��� ����1u(�@�?�����V�9��!ދ/_w�=hZ��x���<�Lu(������Fw7EW���$��<M�j,/}e��0��+"�Bp�B� 섺��m��	;(�c8j�_�:.�U����c\܄������̯06$N�6��U��H���D^�f���5��Ir��%5�5����h�߸!z]��G�iãE�9�����6�n�6IȐ�;�#|�ո�fO�Ӥ���.�5~�d�����t6\��Z���r�Zɴp[n�n��`C��7�͐�jh�j�S�K�����|��F�� �<Y�����̝o��N>"�|x'��PV���>�Q�,n�4�<2(y�J�������e4[�>���h}��@ϕbBq�.��r㑼�H��Jc)�k��x���prG����O�T9����.��a�@}��8%�6
`�"�ud���W�>L3 A˂�m@7ׯ����Ei�	�x�Ft�Ɇ��F�P��\�_��ut���,w3���u�'�9T.iU���ɣ.�Ȍ�@6`<��/I���� Z�<"�����;��_ߥ�[�A��P_M���9fᚨ(Ȣ5����d���ʓS��O\*�� ���-j �v0�琼҃���#�#m���2�#��G3�ř��8~#}9Nh�8i(Ru��?�>(� ��s&��\����
#�4ު�+K�鉹^�-�+ӳ�7䷪����]
A�_7�{b
��KȔ�L�����qUܴ|�s
 ��=~�1�w�e�֖Kv�F�\�v�g5�`
l�'�W_��0SX�e�Yl�qzj�ZR�!��vR�k@v��p5⸙Ƞn|ex�cOz���-�'<ɉ;�؉��V^��ͷ��E]R#�sd�N��2���48tf��t��D���D���BZ|cӜ�~���_�k�~���X�xP�P �RH�":>M��(�RDV.Bz��,�M��WnWt�%&Ƌ�d$���UU>Ǆpq�&V��z�:W2�t�t�gUU�C#n�ΏP:5�()64*�4����y��g�#1G.�����`�>{���/�=�����<����~���)IU�7e� �N���X
JҢLE�v?ָ$���j���(,_[ V������fQ��4`���!?�v}8�˫Y���O��$jFl�N�VF�!f=�� �+��>rS��$7�_"��^�OB�& &2�؊��ڟ����J$)�8݄!���Ny��]�������X�|�셪'D�TWƪ����[g����K��G�7�q��%��)��
��+���'F���d-�w�SeU�/Q�\�!@i&�����[{(��[��A�����)Sמd;���|��|��/zF@������ƥ�ǈg���{��Y���13���T�W m=0��T��pxf-3�~�P���3�ۏ; J^t0s���b�q��vj1ǩ�g���~�T�a{R�KqjE լ���)s"{z�gʐsL�C�d`Y1b?*�{G�� .���>A=��?�����eg{@V6�Xt/��¹5N֝f��a����,�p.*n:�B�ᇄ���w��S>������`]��8�]�:/�����l�ؐ����]����
p�;��iÃ?�S���BL�'�RE&JAiYvsfu^,����Rs�\��O�T�+
%z�8 �j�'WX��D8a&8p����a�C �HnԸ�k���<=0$s��||�-�ųf1m5M0P� �5ڵ z���4�_�'<Z��ćReie�A��o�^�&������9|��H�/Ƭ՚^��/ �-����@�j�V��)� �T�D<�I�>	l?�%
P��Z�eH����+�2���V۹p*�����S���(��.�u�����[ ����+k6��y��k��U��/��1w���,V���e�r)���z6�2���Тsp!�*��Ňó��+ ��ϲ�QG�>!�M�Q��?��E�v�*P���Cm8�2�0nM�5��c}�/d�i�c������dW�b���z.nȼ��O��� ���3ځ���VKp�;rV�%i�����,l�N`�x��ƨ��B�w��pF��l�Zy��O�~^tؑ������2<�Ur:��FR�?W��鸇o-�c}�����p�`HS�wJvD��&�(�#�;�]�&��<��W�G���O��+�\(�h����6��ui���1��r�uu�*�}Ll��U_P	�;yV��g.�H�� ��"�fC�IC�q��$��̣��
�����X����
'�OW��K&4�ky�iE�U��A�q�]��Q���p�L���nD)]�79�}��b�M� L���t�U�ͳ��t6�I'(tX�5��[�.n{�<0�\F�����![��(�M�x�d���Z���5�H��:kK�,~B�i��_��*���S�:m�M��&��V���t��M�!�%#0 �l��4�FZ&4]�2{�Q[ױ�����7����<�d�Ĥv�CF �1 ��v���L����D��"�)Ü(]�D���Y���ŪE/�]� x�J`sqrĆ+l�AK��_�S�Kh�I�h~F]k���`LA���Sɂ����#�tܫ�rӈ�7������#�����-�LȨ��[�c5���g5%H.��o���u�^��Y�/�ϸ�9:+�V��V᥶�����nTG���:,���L9��J��Db*��0`I�,oJs�w��1|c��\X�,Z�v?p[���e�*�6��&u@�����_�g~.�b0l�^�ĵ��F(��y���D�u$��
"�3�:%�|�]�o=PK"J��ksX��j0�<�25�X���=�<n�>F����%��h��x��`7A�v/+7D�<��v+�F'Qo�mv ~�
8'��(��T�o$GVu�#<Cmr���0���+o
�Jν�lY��h4��*`_~,��@vP��%hv��:��q�?.t?�0��C�)��E�&J�t�a~�2݄,J/�w!��wsPJ>�C��J�f,���d��f1��@}�߾��iV;L�`:�Jt_� E��@����LSZ��`5���-����q�+@:�E���3�����ӻJ�"����:���;��lj�m��H	vX�8=�Zn.R�h�Q��cw�̿�$Z�_�����$�b��4٣֘�;Ϊ����K��`���-����m�a�Ê��܎	��u���E^X{�C����xsn�4lq.-�K�L;����P3�f*�����R�~�WбY�͍��\��Zs��r��3��k'�	��[NҒ"͐� �h���jd�D�k��
1�V7F�īޗ�^�MҮ�$^o(�>��;|>�7Բ�eV�a����X��9d4��2�jJ�m�1�oJ�>[���i
�h83@���B����[�ґ�!��i�^K����xW���-�KGҳ�TtB ���B.��a N,}I5�@�8
�z�"�/	d�רW�ؘ3��H��@�ζ��|����f,i�f�xQK��au���[PiIQ�zO�6���,��2��k��G9��U�)���h�1D��<U/��l��Z/*�������I�y~@A�pGP���ݝ�f<�(���ϟ��߼�ƥaj�A@\�ڂ��WF#(-%�#���~�b���^���7;=?w��IV2��}� ��
kʳF}r��ׂ(��¦���>�(� ���s,�E���잘No�E��4��v�&p���}��]��F��2��>�옿�ߝ���vRK
���O�y����[%@U���3L d��~}�7��o��;�K��@�׳Ov�7+�����ЎR�f���� �"lzaj
f�����FLK�މ�����
:�)�xW�z�"-bMT����$�]VY.��(S�� d##��d߯�N�����4�ϫf��<�:����$D�S�Bjx�ZW����u��w>sk�0ҺJ�x90P�qR��!e3��*���a.=�Ƈ8��:�6�r��W�v6&�]�d_������>�̣q�m�<O7�?��W2��t���g�tUC6��)GP��(D�	*����ϸ�y��S����)�8���`|����R/����ʲ<�̕���o;I�X~e֑@�i�7�A.�
%P|L� �?qU�j�j@��(罄 q�VK�����Q`�ߜ�~�v]�L8ƲY�te'���Γ�C��lJ;*�QP�!wc*=x�m�F�ʹ�◒+$N�����Yf�B_:` �1�إ�Q�h�]tf),#,8x���l�N�H9܃�2�N~���P����D��oƥ��E&"5�+_��9�ѺQJ�#������\��惰�;��de0�Z�2ain�A�&S���q4[���~a���6�F���?�0��9���S|��z��B��#��B-�#������r:��t�'l��Ҝ�=@�ُd
�Q�;f(�E�ٓ2�Ӻ�33���^O��Ԝ����ve^Щ�3�ō��T��RQ~�j ���瑆���-{u����jÈ�s�`tMCb��&�б����J�Z>< B�ha��=:�؊�g��6�0mtj��]�tN�+����O��,
�o*�M�B�dM�զswm��S9�e�*k
`|�8�XK:�0����z�K�oX���op�J�ㄩ�?>��ͭ0LФ��&E0 Y�A�u�Z�����N�\��O;.+��zqj8:%5&&����s:aa�pT%g�{{Ն�D�H)�!�9'�| ��$��!|����!1ȄM�@��g��0�����4��'ׁ���#R��d��MFꡪ����9�#He�uƧ��^E�e �~���\u���j�[=�T�BM�D>o	�,%�+��0�/����ʛ4��si���l۴�*�E蕺���f�©�u�/�L	 ~���r�6�'e�4҃k�!��E|.����r�,�׮�w2��zV����M����JI�N���܌��`1L����v�����;�l
��Mԃ��z!	��Yv9������C�����,�n(�q���4j�
�dHڹ�]�Ր<�dr�GbXq�z	����b��1�.��3��ܬʘ��p��"r�x�%盚��;����qN[�3�i��`�]yGw�-F��˄����^ H��P����=<���: �R�ȷ��*�
YQcx�s�KU�p[��HnO0J����^3�����&�Ri�0΀��9<�O���W\c�ٴs�I6��i씅|�)��@��*��l6��_�u8;tV>��-�H��= � *"���$x�qܟ �1����շ����X�z��h' {��+�49Gӌ�vP4�A9Ǽ]~�L�
�����jJ�DdCs7Ը�x��bA΂ Bf���h�H��Ol�Ib[XrN��VȖn�,�0^si��l����u�d�q��Q�hz�5��|�UD�§zq�D)����Ź���:��$�hSH�,�Ҁ�����!�7�0�>�����F�R�U<{ ��,D���`���<>)پ��w�L�tל����Ж�'<���l���×K�WǶ��]��q��W�]�X�������&ZL���ٷ�S�����^�~!@V����F����b��ȑ��t��r�r���)\��U���0x��Oc�D�V�~{p���5 ��#�(�dQ&^�)z������3�+�Ňd�rV�����l�bynOa�$���;�LT�JwUxb^��k��� s�\, �����X3��ZXalK�ͩ�aw�ţH6��΁$��u`�x�_��._G�l��*�P�F#J]ys�ە��E$���"w�c: �|��!o�	4Kh��3qX@Cv0�y2�N�-R�w��.�T��q����hO��#�J7��
ZD��%���!Q�jmm1��%�3�~F8p{TcG�#7�r�9�0�!���Y
�	���Y-D�h����%�B~�p�@1-?�@��t�,޼~��|tڙ6� ))��Ek��ԚdKҎ�A�o�,��7��r{�J��J\�2��v��w�[J1��@�þ�m�V�~1�ڋe��3���w(`���L�����2��g�6[����c� 2��!z�:i�Ӷ��"X3���IøV�f��ؼm��,	����Y(�U8�.������c��<���Ȏ:���%�$��Ŧ�3������w�������;Q��h$K�k���+��]��Ù�3��_BE9���~���!�xn���b�h�;�qy��͞f�]�K<��d�~��رu���H�R\)<�Z�l�r^dδ���!}�Vy���A�+h�j�����TE�Ȳ�iF��2��hĠ3��o�`�>�}�|y��M�rV�"F��ߥ�%�4��2�6J�N�l ��6a[�6��Kh�y7@aBg���6�q�2~��KM�Y���!G:x���H�lG�.��gT��Ѭ>9A.��a{��}�[�
V"�"�ƌd�I�W.�]3���f�@����9������Zi�x�oh� �X�=P$�iÕy|k���A,�#�7����9
��UnWD��M�╹���E�<���/���^�Z�7�o����m�枥T�PA`P��F�ض�f���(>
x��ZN�Z�ƀO3��\8���������-�} ��B���C'�9J.��z�����2y ��8�����G�.Ǵ}�"��p(Fh��>��~ `��sG�B�RꙞs=�܀��4AẶ!���?b|Z���a�ޒ-Y8���}�Ӕ��88ڻqb
p�	�
�ʠNW�ֺ�U����� ���~xǦ-�؉�uK���R�Yvn'q���R5R�M����8���Ol�0j��΂��āB�������2@�n�+��(xjuz�Y�-=�����ؿ�.VTj��}����#�~ZqSNq���4��j?�f��@���0�eGFD�<�B�Z2{�7�y�=�k��u[Dx�uYP:��R>;��	�M6����.8���t�������d�Wj�&|Od�����&>�4sqLծ������yM�@2���t��g��vCiD����P��(_@�*��ݪ �y#9��Yf $ݖ�I۬`7���
 �/�$l����<���48IIAEe����@Z��+
 ��L�Y?����Gj��,(�<R �*��'ӵm)QAz�`2˽�� v��V8�����U��*�֩�$~(?l�^�Lz�!���=3���a�u�4���r1K$�+��a�T[�B�Ι �Q]���Aڕb��8��)g��8���,cN/ӹ݃�i��à��E�����Dd@Ơ����n�G'�FL����(���r�^�J�%w� P��7؝�����0�m@�eW��[���x�b&���,��[������ˆ��!ā:�_侞��w���V9|31Iz<��p�S�<�EǾ�ڣ��+�	����T�B*�MY�=�D��+���Wf#��4U�����3N��1.^*�Ԝo����v`�U�V ��HN�T( *R���j�C,�"o.�_\�{p��F�Z��v4`���b5E,������ښ>7��ã������rgq��6e('t�����N�N�ُ�=`�
�Z,%��*d�8B����]wP�S4tȢ��`��8�s�:%���)5�N�ј���S^O�Z�upjy�㟯c?������LC'-�Qi&@?Y,0Pu�XM*|��)�&\8uO�A�+ �z�$	8�i�A��8Ŧ�,a�:�p�(�v ņ���H�S��T�-	'����$�ڕ|�����sw1#�:M����6�ګ�5�˺-4�^'r��|R~��������,��W�9�n�H V�Ƣ��^�O� f�ޓ��`�žE�_����T`V�?�	" �%�'J�K t�[Ձ�v��
�K�2�ۯ�*r�8�PA�����$�u��P�j ˦���	6On����k�j���蜖�	�L�,�l�˩��(��a��h)��.�)�(�����L��}��88���Ș�)#�4M��鵮	�9�$v@}zЁ�CC���(z�n�ݬ
t Oi�_��7P}�Kzd���b�	�z䝱�-_�������7�]�̼�p��rL\�%����#�7�b7NV�����8�xDw���FnҺ��˞܅��^�;��N�\�=q�<��_:���R�qȔKRP���/cs\���kptH��0Jl����c�����^�&����g�����T�O���\��>��I6�cim�#�7��@^k
�*r��lq��_�";ovY�MmHh�� ��"��8���q��̛�����Z9WXg��9&�'�k�[+�4tB�����K��A�<]9��+B�B3�E��D�I�7o��sw�b�n� ��������à}�*�I�*�X���Qn1��0�0�&���p�ީqR�0d8}��g��p�5C� �p=��"���չ�$n`��~��:#���#���G����rK�]ێ!+ja0V�s��ntF�<�,J{�dק���iԙ�7^<�Z��t���Uײ����
�ղ������X`lÒ���i�ЍK���;��]��&������U�!h������0RSLm�?�~�B��%Nc�l�~�n�8��n(t�r�oh��Ȱ�X�C�Y抛����Hs������������5�ل�^8��L�^������^M�+}��hV�������2�YnJ��u���Lo��J�b�U��Tp�b�Os�aE��րy�4XN�Z�k%&里���`� 6�����Ӑ0�*�$_��.:L0l���mF�yΑP���Y$��|"�T�:�L�|��os�K��Ꚏ�)X��0��2+:��x�ց�����[��G��*�h
2A�>|<77'��D�9��ܧ�Q%�m��I�@�h���� �TZ�UG���#2��r=��0��_�]�
�Ñ��=�Yh~h:�&� d�~�A	@�)��[p�ޗ��-�tuô����)��wE&cԵ��	��� �,����*��m�xJ�r?���Y���6��1&��@��_��`�V���֚�������~�R0B�B�LF��ɼ#�^ph_s�2UĪ!�����'.0���>9ӱ<X"��D��i�q�bg�m�\�	��4�+�P�(.pt��|c��Կv�c����`=?$Ca��R�Y�B��A����}�AC���ܣS�����e�y��R�N|�ڱ�E�_��U�[�n�~K'����G&;�HėF�Df����������~�7}��7��U\D��ZirPr9��!�5�?yȃQ���HW����h3��jZ��ù���M�tF�Е�M>��óK5�o�t>���|�J����wV��O��]1�4�eY2��Jd�C���4�ϛ[���A�h��@ �B�/&�5��m�ޠ�P�T��|��x����c�G�����T�0w�٧�.�Na�0�}�nBvOu
��"�} d5܉W�k�3߂��@h�E/r��͜
�iS��x�����&��l?P߮�ð�Q�,{�p��,(�	�Ҫ}ݰ�9e�U)�	�S#�b���=<�cw/�8}�LZ�d�*����1�	��/$�AA��P0~k���df�C=(�m_�6"��`�[]Hn��\ӛ�����	i-�l�����X͞�Ҳi��s�3��ǥ2��C��TG�Mlʩ�o}�87v2(�Ef����>9� Ιsb����	��NL�ܻ��4�w���f]o�|@���ʪ_�]�����ԏ�l��
���ŭ?�#�o�Qp�Um���4l ���~s���jD�DgKK�X��͔/vI7��w��HQ��A��ݖ�l9��j �n��քļX��<y���ÿ��J���O�x8�z�!-�4�:?��Z/VOƧ���ڰvѱ#4	��R�NL��o+����f|�����u� ,D�E�B`��Z7��r���[�k|�Ќkx��fPU|{R��d�СH�ɰ#��.3Qz�=�����R��C|W���&Wa\d�7r�&��>���q�\����˳����2pK�t0e�g&PC�I��FfPkθ(z�*yP%݅h�y^�(��0!�О��*`�x��%�?/��*�i�h<C��O�� SIfI�eL���˄�7�
۫�L��N?�:����j�8(]�� ��yAa'�H��Q|��`���\{v8!8<�������Aք�\��yl���G��!-VS=�>��|%Bʯ��M�Z$ĥ20g\�Op�B�� W������}v�()�Mw8�
F��N������7I�D)d��Z��6[#D��ƛ>f����]�aY��/1K�Ȱ���u���1����<5s�X�c����;fe���!R�d{��q&	_����e[�q��t���ҥ�ļ���V��'���/�IM�|N�z��ےK���w��Y2C�����j���bX[�]� ��5�=����d�|�f����6��I��3iF���6�^�Ja:�B��v[W��,���TC�MRGC�j�p�]l�� {kC�ʡ��t��`�!`b���as�C�����>2�y��u�5�g���6@@1t���̓�{Nǧn������$,@�*��sBi�(�Kûw�5	S/'���`��.8��E:�:u펗񉉬��FvN�Ȯ�ep%���?4���L~[>��$D&;nBY�>eu�2E�o��k�\Aw(OTh+���z'^�8��\��u�Ł1aׄ�p�(b�q�0�T�H�C��o����K��*�$$0|M���j1~�Mag�Q�.�&���4? '13�u�Rv8������m�K��|��9-�JH�(�Ɲ�y^�4� !���,����U_� /��	�T��W�: �	}:%;Cs�f�����`�Q��EV���'�۪D*�������-CIT�u�*�D� ��m��`�6��Y��k�ӥ�;uW�{%+ԇ�,'냮��z�}��Q���}E���~�e��R��ז�ų��y,���EFZ��hݚ�(M�G^��[����v�4ad�<�C�,;���n��y�E,@���Z����bB�؅d��%bN�kz�e�h�d�g�ҋz*ڒQ����p��r�_z%�a��^����̺NQ��|��֫��/�wE�FI�9��� �p^�O���W���o?<�w:�R�:���6*�@Fcn;����pѝ�H��yJ�)���0���B�.5�&��־��xܑ�ot�O�%����\ق���7�6�؂i�����
��*M{Sl��<_!��;j��x�H#�' 1["W5��A�qR�T�g��������X"Ư�T�}'!'�6K�4�]��:m)F��A�ѽ]�2o�F�:꽎 �CD�o57
t�n�b�.f }����B��>G	�8I�[�X��u�L��n��e0� ��A$����ιʋ�͎d�آ���w�@5��HċV?ӳ���hl�����y��:~1s��c�b��v�X�8RM!f��0�Q���;�Fk��$\{6���"�d�D���rj�<ts��O�T�Z��ؤ⚅���ݵ�M���ϡÍ��,�HYe��J�� ]s(���Y�B����R��O�=S3�˯��B~�e|�`̒�&�y�vɓ��)/t-=runj�Ȗ�̓����w���aꣶy��6:��g���	�5�R�љ̹��h�^�'o�@s����+8s|�Z�Vr�&�V����O�nE�U�ڦ�K�L�W�Jm�#b��ܤ�����s͆��Bi�4=�Xi=�ZN�ji��?�ָ�<�6�B�7�͐��E�W_hF.q�lT?�Ć��F��y)��uT�$���"m�:�|7_CoO�K�S��۔X��0&�42�EM�Sˁ�"�d�Y�O�6��hŭ��Yo67�}��<PDZ��G�K�9BQ��^m��%�[r��ti����T���G'pl#-��r��	0@%��&
�e����Y��h�o��~=3@�F��v$9j�T�r��h��t���Z�)߾&E���Ђ�҄�l���7,���H߃�h��JOa��6o�j��mm�$�1a�@N����s�VLC��X苛s��)
ζ-Xt�}	�L���Ě�F��#��M�ɪ�
��ַi^6�p4�Ӭ�"�6�kє��Xi��m|ڥ	'MX��F�K �.cc���{�c�����*���e̛��$�5���Pٴ�7�l+)�ҡ3���1��؜�ޢ�ϡ�����\��f�i�r�UA=E�t���5 �W��n�S��+��|G�;�?���bvf��'�����!~�׽�+�M;��\_��Z䗆r\\����˃L/Aң!L��ZhN��jՇ�j�ƹ����WF��ި3��~T0:�o��>���|�� ԃHuV�����m�]4�*2��J?�Ɍ�"u��[����z�qhi�,@; B]�{������Π�t�O�޶��x�:K�~��GyGqi?T%��t6F.İ�a1�1}z;c���
L�/"rTddp�hWdeO353�Y�~@#v�0������w��i�>�x"��
��daP������a���K�y,c�C�mz��sy9��|U��5xZ�*3����<7�/� cxZ�Z@�n���,�����
��A|��P�#���HfM�(��ʛ 1��Px��6����\n����W�y-V{����Z��vB������R��붧2/�����1��$�v}��ru�(|,���g�>��r ��Bs}Vv�HI8�){&���4wd���������㔗�)�#N�:lM�I�t�n�ݻg�
&8HȀ�ؠ>R0��E�UH�o4J 5�u~nݸ����,eK��ߧH��v$g�L�#�:ݎC7���(��Q_�lTR�j{H����������v���t;�$��Z+�xS�z|��-�~��u�����VJB��9�ذ18o#OG+PT�N'�ڌ�w���*fwF��K{��
�Do|B���Z�N����H��kw�+�rx<OXPp��R4J�������P��*T...cƘM�k����B�W`��&2��d����X>�d�q��m��YC2K(2tk��g���C/�:VP&�(��:*���`�y���9���`�!��@`�/x���Dl<~v��`s�)YI�qSe͸��v���/
��iL1l?B�v��MjQd�(�� �6G����#tQ���`h���1vn��8�/���7��S��_�d�f�l���B.=!���=��̗�v�*p��(�Z$�_.�h��J��BpW �A��l�ڋ���)�;8Iw��	[N���IoM�Ra�߿�Ӯ��.�q+�DT�	Ɩ	��VE�Sؤ|����:������P��[t���"�����i�3ղcW�e�L��2v��&d�<�wR[�tv��4<��ۧ���,����S_�-��d�|i�z2F�&fmԲ֓���㣪�Q�ŕi��%�x��C2�=����@��"k�f{��7��3�
��'~�^�K���sj��=�vV�ԩY>ž� T^^�R�ծj��ì�������{f�����/ܔ`Żjb+�;~�!�C>-	0�y�k�nCV)��gg"b6x�t'��.dCN)��V1��XS,[q�*ZH�BD�>���w>;#S*Ɓ�;��`I�8
�:�)�i%>������IF^�iap�6���?��^^�L���� �&6��Y�l:uJ,`�I�5�N�\|֯O�+��lz���8kShw���\��a�p%��l���qlHZSt������C�d�$_��|�I����1�2�M�a�l�|ڡ6��d#4z�	'����`R�d�p�ۄ���םWW�9hehH6ZƘ-'^V:G �0��GU��V!��Tn���TQ�P�5�	�@%�~ ��f�Q�K�,�����h�@ۥ V*(>��Ʈp�H����VuZ���I Om���6[��eg�k]�Ƕ!^�Va��7},^��m���.���-)���3�	�;��K��ss�1�׋���� ���*k�Meٴ�+)G�oWv���k����C�v��un�!F���;�N�Ua���G��U1d�Abɚ�z�Mۼ����Ji�u����d��B��p:�JrB�%x�����9И�SNL�M�z8��?��:�w���F$.I�F��ܻ�F^񃘑~���6<�m�:��$R]#���:��ۛ�ci:�\��p�G�H��
Jb����k~�C��+�&�P�A�;�3-�@�Ou#�w\��D��6�mi#)B��p~%�1a�*(e�l統_�{�;ed����H�� L�o"�<�յ�zq��̀�K���R�.�Xݛ��o 4'�Q���~4�ٌ�GA��AJ��]����aN�8
���D�D7���iٷbR� 8�#��������͗I��XCX��Gxn��0�w��\r����ΔV�)�dn� ����y��5��TĦ���0��Ռ�K�R�E��t�:ْ������}&���҅��!�.p0�[��(FFƗEI<r{QΎם�_�8<��L<7$���$�c���՜�z� )X������_�Ètrh����"�\�1�n]N��6��ݜG�������
��SN��5yc~�����j6�>�t�z�����r�tH�sr��x�������ο�g|��| ����u"����ys�5���Ԁ�5�^��C�������+Sćձ;VM����J��h�"n@o��5`>��L��J��b��T��g���5s���MJ��X��Z��;���z�$����6�ZΒ�琦�_`3_}��.��l���!k�F{Vy����0�N$
)"��}:�w|rJ�o���K����DA`Xq�0Ao2!q��.�/�(���tP��覑+;h�I�t�87-�?��#D�����u�Q�<�mb���vpJ��*"��T��WG�)#(�@r�90����
�����UY�)Thpn���~�D@b�/�����-��M���t�v����):��E�����A��*���,6$�㳣�cSJ�� �����o��Z˕��1�{@�=����QV���L6U����B�����LTL|=ο������Ьh5���'±�S��B�Jmӧ�"i���&�C�����X�HmWx:	b��j{z�F�S.�v �=��c�J}�l��� �����$U�@�������'5����1�7�����/���<^ګ�H�/p���!����A����E��/����Yn�Hݿ��7g;W�<]4f����k��5E~��������y�\z�Z_�hr�⾴���u���G�o��L�r7WhixjPE+��Vȃ�F�\��I6�9yU�po��>i�w|*w��jV�%;��t�Ө4�2���J�ߌ�I�`Y[��|����h$�@V�B�����Vp��Rr���Jgb�2��xC���-�G��D�CT`�>��L.�2ca���}5(h�7R
��""MK�d�`;W�~|3����X@���K�h��R.Fi�x��K�I30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�/ڜ4�{^�{]�$Ht�E/Z}1TWZ�i�ˀ���9��Z6$�x���<�������5~��ߣ�L�8�6Z�^��3�B��˞� �Z�>~� Bc�wz�荏�`�ر1�y������P��v���cz���Q�ا���@�j�{��T�,2)��2{#��X�jEǁwNրv�t-+ ���2���)D���?&Ìw��K �ڀ�-���9E���YW�%����e�1�8�3��c��<G��Y>i���9+��=��in3�4�S�@���`�����j�@��I�`�39�Ǹbн�>D,:t��N��@wReb�T�
�1�掚l�A{��K��ү�!��'���^g}h�2�+����1�V"5K�AO���9�����sǑ9MܐxZ:"��?�_�=�h���G�9��eХVN�Ѩ��vdv&r���C|�7��|`D����S,!ع�9�P!0d��-s?�n��T`BY���4�זQB��ǝ�����-�M�����6��v���>���m���zh@��k�5�"z5G��GԊ+��Y�%[�Y�5���¢�>$��׹:���������n����#@�ᶻ�&�������2�T��8���ln� -S�ɀV�ß����[��i��;��/�@x���9,��I)�x�(�mF�A4�}��Z��i���";�'��#����ZQ�=g��fKc�o���C��"��ևB�4���;g|�t�pbo���t�6Q�+1> 
+zI���
`T|K�!�_�}1�����7��uI\�_��LVL���r#�A�$U�n��t�p��������0�Y-�+��#��*��$}u���4,�Y��e>�u%0���U���3,!�w(��kҾ��8-�[t��/&|Ώ�v���$XBn̊����z�3�4�q;.P"�0|B0_��I�܇�A)�<h**5����r���r=l��H�v�;Uԍ">�nJ�Ğ��q����փeu_|�Ë7���>>�HD#a��P��Boq�گ�9��0��E��B�	��e�J�"N����j���*�S�����q:�Ӓ�e�*�L�7��6D��?���M2��z�W#4���;���-L�ȵm�Aw?s�Dޝ���кT�P��5�L
W��V��ސf˽����E=��EQ^�ar��Äj���0���1;O��b�����N�׋ B�Q�d`���dxS��ET�M�x�(\d%>� �y+%�������{�Z5�;����Cg���x�.kT�h�W��x"(��yZ���;:l�@c�̴��;�طç*f���#��c8�J9�]�8B�0Z���YK�<F��%�+!�go%ki��F���S��9�Ħ�[��\ȵ���T� � ,9�?3mh��	)�)[c������ib�l��5�*v��ph����`��ܘY�.�h�գc��5��4e����l��2ǐ��¨��'��nԤ�s��b���=Ua
��ºa�D٠+�w��WC����*���ص�7�߉�v�V�}�<�Q�.�,�3Qu:L��s���߻v�Pc[��ňy�D�JO�`�q][��$>�H�_D%~��-ܝ##5�y�����I���b��9����* �t^~��ub�"o�9n��wj�����*4s��6(<�4��W�����Aޕw�}|�,��Q�`����p$�)�e&��m�J�g�y?F��Q'ŝ��N#��ͤ+�d�,EY����Âv�6m@{��8�>+Vu��}]}PG�<�����F���8n��]8vbʟcw)��ْR�s������9��t� �uƦ�k�U`ʅ�/���$� �$Cz|���1"��p�x�䗥q1�~lp\1r�%��z�Dg��S{��)�~6�i]l�F38��~��l���-��B�
�PΓv�n�+�IF�~�+��UXd-�wU���?�A�U���=�����]����Xm�M��h��}��4~2)k�������aj���m���2���?l��>Z�3G��|�hb��&_�V�]��T�9�uj�eGҖKLζ�C�V���!�^��9��T�X��|Ǣ�w����`s�n��'Mr!"i�fi����]0r����)������ځ6�3����ߟ;/��쩚����+v�M�a)Gu��cD�-!�\r-�Y��"�G���b��CE���>y��[��������`���L0w�bvd��EPztZ�?P�,G.ݦ����5�F�/�@M䅉0�J$w3����a���N)�W-����[w?ZۉGr�;��[�'ڢ#�c9��dH�n�u�3M"(2GZ0�p�a'��c����ّ��r�Ot/6�=Y"!~c�Mp�2�}�|���ar�I��8P��_=�΁o��<�s���Ø�Y?��V/�d�+�{�c�$��`ES��Օ�{��i:��������~{B$nb��5b�J�i��~5P��b\��26~�à��B���B�c�~��~q�qc�뙐�����,��U�y�$�{��P��^�܇ҽ��IN�u��K$G��
$je�k�x�R2�@~V�N�1Qji�lw�O�v�"ѝ� 䴼2}�~�&5PDU �c�2��d�o�~W��Q����T'�ćY��VIG0���d1:��������D��q�G��Y�U�0o�+�{S��83�k'4%@���˄� �yl��|@=���Ǟ�3��S��'ʅ�>�DP���Z&N�	�@�fe� 7ҮW�1�!����{�5��ӷ�ߩ�B�K��2bhBϰ��.���`����K�RP���0�#S����>9�C�x~�������z?�BZ�������e��N�Q~�(�P�W"�Sʵ�;5hqR���v�;�WN��y3��`�k�)����FeIv��� ���8���^u��������ZͲ� :h�יՇJĨq�&�uZ�:���G�v�F`%�O��F�I.D�"gǇw�.�x]y\�2{}���O!RTN���t��n�L)�g��-�r\���o��N�;͒f"�'_E��)=8Yn�x��_Rz42��p�ی��S����Ȥ$=磍W\h����_ڈ�U�?�1�ݎ��M'
�a5O抢�֭,}�j�H�K��ݹ����$�h�j���9���M8O�jO�+�?J�|�������I���d��%��t%S	h�}H�����RH���k�Ji�A�V0��5�;:uI�$��7���Jc>�a�p�kȚ�l�Po�ބ�0�6O��x��q�N�k��/��S�k�l|IV�E�E��Y�x)�i�[֠
+ȁi�0�z��2�E� 6
�v�ps�ٵg7�4�����ʱ�7(H��s4�M�8,9	&MA����$��q�������)º��,CR3ѫ�����X�N�4�)��W��>Z(N��Y�Jnz�X���q���kf/F��Bҷ�h��:�s�y����OX L*%��9�ћ�I<��a"�������r4[2�(��:~�<(խDJ�r����(~=#��(�z3�:�+��!�L�w��_JT�������3�]�Ԍ�cٞ���NLaQ�"��>���D9�0�&Cs9���	�iO*6�a�r�<!f3-o�9)t;�v�<����>��vr� ��[��NHR��}5e;T\7��C��IL�|�O<bV#�H��!m��Yڭ/^9�����Y����2-�w���Eo����|^p�j6�7/Iv��e�S���guJq����1aA�M��yt���ي7j�A(ա��r�td�ml�LV5ۻ�?�2�^�5��i��w��Ė��;�`V�ʥ;��Wh:���a<��ŞQ���U�(ہ�c��2�e}���6�Ӱ'�~� [RB��c��lV
�/��X�H}��B�xO&�/NVh�W[��ب!�
��)o��[ݞ��R�d��Ѕv��W`˓\n���H~�/�1	L9�*kdi��	��p��L�:>S��+���1H��vQ��閂���NX���Lv���0�7~�\�r���)l������]y�����&�J��=�؀��b	l�r(�cSe��\��� �����
�s����@��rr�)(��}�#7
v�Vw��Ŀ���Ć����PA���_yZ\��� T�q1r^'{~=y��&�i�C&���ރXBk[�S�.O;sG[{t!�&@��H��8��dW�xp�8�U!+�s�U���g��T�̈́S�M��J�˱��Vb�)
p�u7qb���S�I.EM�n��%�6/��'NGn���?���\?B�����f�	��4v �Ul�'#g�,���yL�H�A������&4&���ƨ�ޥ'�0�W5 �+=/�YBF&��J�	R�۰?xܮ����_�s�������<��-V��+$�� �`8�q-�jk��N����=���Oh֎jz���bJB�l#��GWmzA���k�ù��o;D��B�b����T{���K�����L>�,W3�����O�/ �֤i1�*A�؜�Av��.�W�F��B.gW�SUi(;+�8��;�ʰ�W�?C��D����v��X-���K'7�APWzM�#"C����&�h�[]MT4�n�� ^ F>PE�2u�{��A�SY���Y���e���c?�������� �xx��j���9����[�|�CK%� ����g�g�PI�m6���y�s���3�g&x�JPu���u�S^��K�L����[�"��y��"�H��,/�+$^� �C	��p�\����C�=�Y�;��+U0������̂υ���r�^��`�~lJ�����s�� �zN��JF��Wk��V<��_���0�f	Gw+� $��� Ғlt<Í�'3_���d~j/������ɴ9|,$���l�� ��.������^�i(�'���9CZ ~��#�j�@g#�uf�=�m}�)�Aغ�8�{�� 6;�������Sz"e"�7$�#����.5�� �5�E{QȲ?���c#zY�e[k.��)���W�b�� �]�s��H�ߋz�P3�ȕ���+��(�S���bn��/f��$��{X��o�I�Bb`�ԅ�yCv�feUEA�w.�iI�-�~��׉�4�sh�)��=�{�|hsE.�W��@X�_�H�͢)aY�{��� ����-�͌M`�U:�^�g�8�s����c�9�y���LAR��ǢU]8'�'��&u�3/U˄�ݒ&�e$GLx��0������<���]�P�/��-4��⁽>���	�k�J9O<��a�gn�οa	�n��PX��E��	fN�_"ۇ�4Z�:�O�e�.�'�$OE{���eΟǀo�ԅӑU�L� �h@ |5�.��5�}�/�	��b�$�鬂�H�X1�J��K+�5Ľ:`v���:��}Y�9����\�|J��@�DV\����'��b	�ř���\��aW���iN(t|�q41�2����d�gI�)X6�#n`�k�M_�~q��C�$#�C�@�eE�KY+Le���'��*�����/��XL^�����K���^R���Ļ\�+�%���f��X�m�}�
�{!I_O���a����%�Av��6�����m�)�g7�J!��wo-�V�+W�c
7�X�-�����5g8EFQ�Ր�9��Q�j�o��|\�� Is�r��},Rjf�������ٸ�q�����*R�ڳҦ��f��KGGx�N��E�5�3��a��M�s/8�
�'!�V���jkΞ5G��`Y���}R����ռ1�}?���7�E|UR�a�_��o^��g����(fߴVŭ%,ь��\�Ht1�>�B�g�Vl~b�����³A�(��OtNoukQt E�Z�Z��t�//pDA.����������p�Z"K��~&z�[S��-�g�O_�(�o��ҽ�E���4�m��,�����@6��\(��M�oQ�~�E�n�zwc����r���Q�Ǽ:�&*�:��Pw�^�z?]�͋���+u3}��@Gv�>�G�7�d�4O�!+\~`����ܚ�jTS(��4^�Y1n傉M��/6^Y��⏩���9�{e���z�X�A��gj6����5H�4�gʨM�R��1�O�����Zc��։�7�:]e�a��@��������"��V����v�=]]~,"��/_g.�'Q7LCL��	�ꅷ�OF��kԿ�Q60D�&e�[�71H1<[�R�=n�U��J���n�Db�r�:��ƶ��d��9>�O�i0-V����b�=���������L8� ϴy���ַ����7Gp8�!=�b�O��ŊD��������*�A�O��!�R1��3>Fm��A�مj�fg���($��b dtR�"�.�rda&���
���9͇�{�����p�90&`�y'��:�L��9c�Qr'�><�����*ygئy.P�� �OKt9�c<	S�T/�Ɇ��켇�E7rk`1گ@}�SY�N؆���;1d؇�- �un*3`/�Å�8�JOQo�4�&���	-�ep�vu��\��ͫ�����hv���n�JE����k����5��Ut@�19YU�%�fVN�tI������&�����ٲU�t�n@W��0�'�c�F&�"���2�.'��$��Pnl�~S��P��-��1[�H��iDY����@Es I����%@Eֺ���.P��
�wZ�:4��g1"��4�v͕���Z��g��_fش�o v����"H��OV�4�F�ӈ�|����o�Gtn�`��P: 8�I2a
^�|8�!K+)����!�k167ɻI	�ǎ5��C�,��A#�[N$"4"�/��}|�2(Y�0СѸ8�#��4�s�uDVL49�L����>���0��cUgT�­!��3��1�k߿��2�¨�T�����C��XEǊ^��}?��T�;{�����[@�vJw�T�X)L�=h7�p�_r[r8��_�@�_�Xv��.U�^�>Yş��x�(������R��	m�d4'��>P#n��P��co��I�ǥP9��m�]�P�]ݯ�ݜ�e�
��o��}e�3	*V�R�h��{\ӟT�e�_�*#��7�=�6��h?3�X�}{�N�W0`��n���L͕JmY��?���D��T�o����=�jڂ�L�����<5޽�����x�nhJ�~��{^*������ju�V�]N��v���͘��骸�I���] /?����>7�x |�E�&Z̊��}�r� ͺ�%pq����t�HT�Z��;��L����h�I.��@m���(\�dZ�$�H��l����>��u��e�Χ9̬q�F�-�8ȡ�
�B=����uY��)F?|/%�ؔ�o2Ё�����S��?�Q��[�I\\���ZI���v �+?c{rh�	�+�[����n���	l�5�zv�*�h��\�-��	�`Y�����h��p�5�e��gv��i��v;n������x�'����Q�s��|�=�EC&���a�8q�釾a�g�v�
�<\a�0
S��$*vy�D׊L���T>.�Q� ��:��à�5ě��v-b[�&�&Ǭ�]���M�q�X@�Q�vH��L����:]�Р����л� �8�	b������*yK����~[b2��o�? n�~w�'�hw�*��}�ɬ1<Wl-ۤ�P�{f@�ΒUw�c3|N8��yheL�Qu�go�]�z)��IL�:PK��}�?S�QԶ��a��#�ഢZ��+�dw,_l�p�#Ï#��㻽��8�"َ��+�RE����}�#�<�o�v��F�f8[�q]�����)̫l��K�s�I�X�lWk�ak����ߘRk`�ޒ����1���̉9CǗ����+�ߥ�R�d��1]��pi�B��Esz]��u��U�~c�]9��F�� �������SB�/��
��k��Ŀ����F$�+��XX�8w��à,�A��Y�$��jR�X�e��ǘm�釮�w��j�g���]2VS֑���	���mF��2}?Y��>���G
���5����_
�����Y�bT�l�u�b*G�8�L�ᙰ���)�'!�O�↠DT|(�	���\zŧ�;�۠�4�!϶�f�����r#���̅m�N�&�G�%�@����1���;��ߥ�'5j�5Q܀��^Md��T�h�LV+(�Y-.�q�O�s���bb$�CRcճ��1V���B�;o��|0Dw�b����R�tA<\6:�(W�3�D����t�#@Za�ݲJqk���Pa.�mNVp�-�O��f�wL�����Έ�.[����/�cfH�d���k��@D(���G�;p�u� c�*b�ޟ���at<�=XF~��p��{�
���"�a?N��f<�"&t=�a$���.� ֨=��� ��.09/�W��{�H�$و�E� ��Hq�i��������Ʋ�]�$[���¶��w����8�~�y8��
P��|6��ÍJ�B�po�o�3�K��~��c�P�9�����BI�y�Χ˨�P�'h�F3ܔ��k�&�·�8'��Vk�j����Ecm2:��c������j�r�w��\v4�p��^ ��D2��3ѸD�㰲2�/_��lM��&�V��J@�Y��I,��AE�DKn�ꪝ�3��Q47���6��6�K@1ݹ@����Y8I3�����m�G?D���f�3N
	�@m�`e,mҀ��1Zi�b�j{�)���[������i��?��a�hT����:�PW���gK�5z�����i�����9C�x�|�Z�O\�^��@BA���/e��N"寺���)O�e���a�O�Dw
�M�
N��3g7$`�Jq;t��!�I������ �ӑ��l���Uu�����ਬ�DA�::���kO�N}u�R:���G#�7F�N�OvS�"��z�gY*n�����\��}���O�OT`�9�ƺ0� �)XQ�?6{\Vu%}�� H
ͤ ɶy[��'7)�Gn�2�@5:zƱ���ԇ�m��'�!�v/���o�R���YKU�|�v��`u+_~�\�5�I΢c�]>�j9ۀKI��݋�c�
Nܯ�5,�v�(��8aDj�Gv�ј7|g���ځěX������^���o	��(Haܼ�Ŏ.RZ�Ľ�Liy��V�c5��KUb��	�d�����cc������k�8vlʨE19&X��0�mcO��Fx�2�w�ks��㝊����|�l�E�.Ά1\�x{YS���
��Yi������I�[E���
�k��
�k7	K��	����7�B��\��_��,��MӀ�V�$��q$�1|���(:�䙇,�M��=]h�S+:�1j����x���)qH>l�N�O��J�E���!��0�%�dVk��a�A��%���G��0Ӕ�wX2Bb%ٮp�c^��Q^�s�0�
wvj�=r���:~�:�k��B}�Qr�k9գ~�P�����.�:*���L���qݬ���L��/GҌ#����Jrga�{�"�V:�ܩ�9rB�&�L nY�[X]O��a_OT�N��3�o�ˬ�;}l�<Y����o� va�H����+�;&,��复d�L\�v!}*V&~�H
��mVX���9�e�Cp탚գ Jډ]�� 5�棭��[�|p���c���紗
�S�1���������x�����&A4">xɭ(V�I�#��{¡K
�F�m~1�V���Tտ����4���	X�����H�M(hV��;�)�h�1��vװ+}�Q�4�'��()��_sP�ĳ�}�RA�Ht�y�ղnBik����
'r���*}a�B�q�OxʅN��W-�(غSK
/B�o�ݭ��=d� ���W2�9\��h���E�B�y1�΃�#d�b�	+7��"��LTZ�"{]��1�vch.�x�T� ��o����yO�	e���b#V��hw'��A���u]�I��W��{qq&���Y0�=�1���*	~{�rz S��*�.ʩ�m۷?5���k�n�@)��rj(׻�"��z@#I��̨�O�bV�[.N��VX]P�-~�xZn:d�R�q�F�^�B�=�v�&.nA�Րw��"�ޕ�1k�l2����sՆt*�i&���ڀ�8w�\W��j��ĝ!��^sz�`��iŦ�P��v�M�yI������Υ�u��S�qt�P�=�9���Ml���bw����' ר����z?����)���4ȥ�U���'��6,�$y��N�ӆ�����(Հ4Z��٣y��z��98㎩e �w5��F8ӜnR�K�ۂ�������s�]#�T9U�N8r�ah���ф��xJ`J�-���읱˵��O�!�g��h��zřs�ڦ\Bq��#|ŵ��zS���UC��A�9V�|B1[?�\#TMM�]�d�W�ؽ-H����є���"! DK�i��*Sw^���XAPl.lw�X9�����W:�i��ʮJ�!;��!����C\w�Dǿ���/���A�i8'Ir�P����sC�a��8�����TƧ ���^2�lP�8u��3�nAsA�CQ��O��?T7����5�\�YQi�ҢixZ����U�7�R�[�W@-%���w"��y�zIĚ�$i��b�����U��iF����u��^�|���w����T͡��"���*S�=��^�C���p_�4��3I�`�EYZ9���:0������*�^���qK�Ƅ�6^���7J����!(5�7H�ďzJX��W��'V�b�_����B���Yzw��$��A�2�l�e�v{?_aaZd�Ʇ�bB�t�9N�m��Q'l=!g���qi��yƻܒ'��9k�~�*����Ҟ�_��$��ƿc��8�،v9��� ��w�n�z`���e��et�$gF��9�.G�L F'Em.�5���~z�G*[��{��P��\��������E4`H�oz#�}ߕ�/����+ő^ԥ��Bb�Ǻ!���aL�^X5]��*�br���׏�y��f�*ES��.�I֏�姡���!�s����n!�{�u�|z��.�ihLn@*��_�����l)�{q �� �
��.�U1X�y�f��h�y+c��yԶ�➷I�]�U/��N'8/&�/'7��xs��G�*������!<��9]�q/��4�u���e/	Y"��\��<�x����Α1��18V��d���Uh	���N��g��g*Z{7��!Mj�@N��v�q{L���7��ǒ���&�������hR��5��(��R�����o5��V]��t.��j�mJ%�+."˽�Z������X����x��nW�JJ�Q����\�|�9iu�����+����@�s�M�Bp�(M3qs2��ݤ���I��6��������P_`�rq�d��6R�Ci������K+��Lw���yn)㼚O�	/��X����K2�K���p�}��`�\ R�%g��f.�[X��}��p�MKIq�$��/��n�\%Z���.�:����J7�9���\Uٲx/������c$�1{-H���f�NJuQ�Dq���#�ܚ��x�g����ŞD�C}>t0fI"�X��يJ&���h<�*�ʳ�����f�VK��$x���W����;}a 	-�E��8��&B�����<�ΰ�;����^��R�-8�紳x ���S>R_��^�͒gk��� 1�MWd,��n�-t�����?�g��%l�>Թ�6"����A�c��6�tU���"FT:�l���D'/�
A �<�w��~��@.��4������_u�����a�M(�
��d������m�,!c����6���(#�CM�紺P�ν��̝c?���D����x����Ƹ���#P�/��̗�_�~���"31��ܒxd�����	Y��F�'!}��`��{���jf�+�L�Ʌ����l�>� �(���4�	}�<qB^7�O�I~N2N�W�:=؄��
96�o]Zug�滰-6d
҅R�W��\J}5��L�茿�1e׸�� �dŵ�	u���q`�Cܾ,�:���1��]v-�8X���32��N��0��Px���zГA��sH7-}����#�ɐ���]����t��8[&���c�H=�JY�L�H	H��r��S�d�z��.ַI0b�����@�l|rt�5�.ބj#�"̲UJ��h����uĠ.2�PI��RZ8P��\΂q���^��9=Ua�&8���V�)�&�_�k����
1�s�x�t���&�� $�,8�W�O*��gJ!��s���L�ŰL�/�BM[�j���ʀ��J�$�˃q>s�Gp��%��M�í�����'�8��Ѫ�|(?]0�A'���4҆/U��('�k,g��y�4��!�+���4d<m��%�
x�%��9���FR�Ӧ�R����܊L����s����m����k������U��`*�-��!���ɵ ���k��qEs�P�zO�$٤,B{��#�� ���FzT�(�C���9�˱B H�B;������Tע=�'�g�a=8�wFH���|��z��� �^�i�Vr*�Ŝ۟�AR��.�(S".����W`��i�Z�w;1�3&ZC�uD�����D�4��,��'ԈP�|y��o�C�
�'`��-+T�V�^��<P��u�p����A{�5�Z�������~���P�?%/��\��x�������M;��'k[��Ea�%d�F�fF�C�IB�n*��z�����Ø6�&�W�	u���^�4t�(1�Y͔��&�ծ�"�]3�/Bu��%^�C���p�K�}�9�j�AY�1��Hݘ0a���u��t����N�3�@���Z$'J�ѩ�l�2+��V�s�N0J"��Wǡ�V��_^���!
¹ywO�$RV����9lкN��q._� (dZ�$�-~𾡹9�����WLl�kT�(�ݮTt���'a�9�ɛ~�Z�~����2������?�Ȟ��!$F��3�F�ݔT��I^9���]5;�@;vщ�c�J�<���E>a�a�N׹�-'�^Hw-�؉��#Ω�[?n�ڐ
c�Rd�<��J>�!��(���G��pqD}��c8Vd�Gz絠�t�=\�~�9p�J�k��:?|a��y�'}���=�֢����|a����\�c^����/�<��� �{��%$�EA� ��B�?�ihc��ۤ��fh��}$��[�#:ɶ����u~cM�ߵVL�6�O��Bŀ���o��i~���c��}�:���a�؃ƒy����)�Pf)S�|~�u�ålW����yUI��alj����u2�XqDդ���jj���w ��v����| R2�.f�a$D�v�Ѿ��I�ϭ]�,(����y�	q��Y�������¨1(v��a��3g���s�G�NJY�����j�+��ު�R13j�14�Bu�I�r�b�'���Y�@k�-�;�3�)����|����D>N�B<�Nf!;@I��et��\`[1]@=�>r�{�2�l��A]���+8�9{���h�{"��h����B��eK$�~��p%����E���9�{xl$k�6إ��;i�:1����:���WebU�N�'�����<i���=xrVT7�S���N�N3Ô	`�S��¨���I�fn�\�f ��6�լv� u���XX/���E͠��:��C�~�h4���u��1:�eG���FN2�OR��~I-r�g�[8��	���\��q}��O���T�N��L"�\��)4�����\2����w���0� ���U	�)�%�nS@��q�z"i]���0���I������R�������c����B��a�U�X��<B���85�5=9�?���Cj�bK����g�͢fR���ų��L��c�8�j}e��-r�|C޳{��w+�R��q=���	�*+H�Q����R� �ę�PiվZV޿x5�1��7��@�|�U~cloj�^1.kv��l&O#���i�0��YO�lx�2���zkOY�?�f��	|7��Eb����lJxWuÝI}*
�L@i`��Ҩn����CEu,�
!A�B*�j���ˠk�Q��g�7�R�8mq���,g&�M/P�2�j$yмq����3�~�|�@~#,q��љȎ�/.��d�|Խ�����V�>�sG�+�JM�ӯTԌ߆@p�kT�Q�=�R�VB�h���g}�p��X�,B%��M�O���m`�ωv��:s���r��іd:������I�rK���~+,���׬�/P:䗁�n�L�E��ͯ�ƭ�{�}��a�H���~>�,�a���";�唸��9�U~&�5|�k�7��O"#a;ܲ���3[���'\�;Y�<cOe��:�dl� [}!ߖH��H�kvn;�h�Lxx�@�ML��x�A_V��OH�%wm�?T�[\�9=�c�j���
������Yh���9��0��7w�p��?��7�H�s"SP����:�8���T� ��A5��~��ɉA������o;ԡrT�"��m�3pVc�L������+�����[��J�r����ƨV��;�·h��G�[㷰u�Q�r�F;({c��;�� �C}r����
��U����BE枡S��
��F�}=��B�OT��ND5W	h��ƃ
 (oo^ �R�B~�d�l؅dd�Wh�\�ƫ����螵�1�����d���	�z����ը��������!1��v��t
ׂ��0��!`\�z0	�՜'��]���������u⋐� ]�w��@]�W��&7�T5�=��˪��	���rV[�S#��
�تj��ζ���JJ�@��rFx���nǐ#��̄��� �˿7�q�2����P/듙Tw�Zʾ��.�qR^չl=��y&
��1겙{�;���k����~�s�g\t���&n�U6v8Sc8W ���f�!��sV0��'��ł�p�A�M�6��9i���^�Uh�qпA��O�7@TMH�U��S���'����c�;���?0�.�̋w��4�A�U�:'ѫ�,���yze�/�{b���46�V��,$�V�o��2䎅�@�y^qYF��s�x׵R����^ ������#Ys�u�0�������=X�ݼ^ۧ�a`�!�-�|����#�rpw���m�C�T�-�z�r�6u)BMB.#�����zz�6��2���f��c{�#�B ���T)�2�&��3$���Ə�o��/���}�� �XLiߒ�*�Kh��8�Ad�<.H>����px�Wr�i�Ȧ��@x;�{F�EˋC8Z�D#�N��9Z�F˙~Z�'�~:P�y`�xCi`�Ȕ�(��CT"����-^���Ps�0u��B�J\hA���!����ц�yPY��I������xpl��q����.^[l��3,j%v��Su���|�I�=∀П��p�I=y�]̩8mP��:$uBd!^�$�:ɮѫg�)���%�"�0�����»^�_C��Ip;�@��Ǹ<�Y�t����0�2����������M ���f�����lY�Jd�ɩS.u��h\��`�J��xW�.YV*��_��e��T&�_w��$��|Î��l����Ҋ_=\�d�@��Ԅ
����9*���Sv�l췺}
�z��@l�Ɨ�'sʈ9��~�w�t;�.�;���vUƛ�/���h����xL d���ʥ�<�Q����ePy�$�w��b�t.�� "+3Ei쐲�t
r~z��"[Yg���~�^ZP���!�3��!��H=|�z�zh��7p��\=+!�^ԁ,���ǖ�I�r�z(i�X�b����bΖ�Գ��y1;�f��!E���.�/���硦��}sxs�	M��d{dP�|ֹN.�kQ�@w@|%_4�J��{)O:�{M��  �1�[(0�;�U�5��O1������RW��y0%x�z�Rù}�U�y��'���&c�o/f@�K�U��c1G:<V����#��<�d�]�[!/`Nx4iwz�늏����	5{�ʸ><<���U���m�Э�zY�~�^�3�E	��$NP�۵�!Z�����ϗ�,��R7{�~j�z����Ս�C�P�Α�h�(a5�dL�#�N��~��w����,V�P�����J�+�?��d���h��'W{�Tb��	QJ&����[M\� ������B�Ň񘗙���).���(b�`q�K2���G�k;�S7'��Rrᫌiƌ��>�oF#��P:<ko�H�s�19Ɇq�	��>��[�i�=#e,�v��3U�)'�_@*�r1�~���s_��AVe_�I*O��7�+Z6�q?�י��0�����W\�~C�	HLyoRm���?L��D�iX��+����QڮيL����:�i�W��ɦ�)�v��P�^V���}|�j��
�	=�*�覢u/���������� ��I�Ս���sxLJ�E7���զ́�W��U yD4%�0��|j!�t��ZN�,;�I�͜ ��9qҟǾ�!l4���(�E�Z�m7�tlh����{����Ց'��吤��
/����8�����BiǷ��+�Y�YF��_%�V�:T�o^8f�E�X���hSm�>�}h�[s�\��,y���� ���?��2h�3\	��[<Zw���Z����l>�5G1�v��h8�HtL��#�Y�n;p���u5J]��n�og��)M��Ȑֹ���kD'�@�����s;_(�=ǽ���z�a��s�dFi�39h���w"ƚ�h����.��*�v%��׶��骻�.�
��u":���L����iZv��[�.��˧�(���_�q������H��e>P��f,&�|����+�g!��d��b_>���l*%����g�Ab^3oo��n�J
wC�)��-k*MW����<�9�з߄'ج��9Pwh��|zZ��%��E��Q!��.Y��	�c)=�>��f��ހ�?^�Q��}���*#�*G��R�+���,>Y$���ûX2���C�<,8��ٺ��+/�P�f]}iO�<�P"W(FE�;8�]�u�xZ�)�}K�8c�s-'����ʘ_�y1�.o��D{z`�@ҒH�E�]6��x(�C��얰�W ��Q���IR1	�ap���~�Xz8={�`[��$�~��]e�FLd���J[������ۄ#
��	�O��$8�Fг�+܊�X�Vw�x��ظA�0r�����XT������m78�����q��s�2�������[m�7�2C�)?"">7�G�?9�a�i��v�_6��^J���Tv�3u#�G��(L�;�\�U�!Lb���T(�0�5�;�P�x��c��N`�!{� f��/�$�rO�(�x��z����7�l�-�Z��|Jp%p�S0}��N�$KM֌�l�ռ"!:�M�54-ZE������ʚb�K�C~�_e˚]n0�l`�gB����0p�Cb����~��t��V�����1��_��t*��H �)@�V׉�M�J�[��_F!aZoBN�V-�u�3Rwx�3���δ�[����[��cE�dADf�CZ�l�(he�G��pw�8H3^ccP���J���lth#v=��~��/p��X�6�de��ak���읫N�c==��DԮ,1��|���v3����/7��xQ:{�T�$�EȆ�@�t��iSH(�&'��62b��հ$����ж#N�� �~N�� ���5�6����9��B�u�1��w��~�W=cݥ��击��X����y��?�T�fP�/w�����ӥ� ��s;��h����zj>Y��qU�2�)_��L���j�w��v`�1�5< �G�2��_�_jOD����FԌ�H3�(��W�g�J W��O7#�YT������1�Ǒ����W$��u�G��<Y;�����*+9�E��?x3�^V4�*��ȧ˽E���#��r@��&��3��и^ޅ�TpD����Z�Nq�@�:ae?�҇�d1�Av�)�{?��H�L,K�B�v�9����h;�]��VD���ǬS1K/0��S\�C�p1�쐼}9
u�x�����g����(��Wl�g���e�g�NՋc�ac���F��yV����!�ܛ~mO�4zEN�7 3�`0����H�-n9IŐo�� � ~�)흄!����u2���cn��r�kM�:A!���K����_-uuY�:'�^Gj�F��O}�5�	��]@�g �"i�=��q\c�}}��DO�KTG(��W�>)����q�\��L.�'�͋��@�G:J)��n^²��4�z�m����߶4D��'���G���ő�y��ɇZ��ݣU���j���$d���n@5�F�j��%�oj �6K��F{�qeܯ:/��N���H�8H�}jh`�xa[|$i���������Y�m�	��-H\V�L�R�� �yEi���V	�Q5�����@���ǐ�`"�cה��)�k��+l� ������0;{O�Rx,���Uakz����쟽��c|�OEh����x�����
oi�#�ғ�p���E l 
,M	������Ep��{�7aU,��'}����,�7mM��]��$�q�Բ��E��)'ºKi,�	(�d�!�Z���g^}�:�1���>�9G˖��J�����"����+�_k��N����a����u.�2�ӛ��X[0%���
M�������Q8���
r�$�!�1:�x9a�p��k�rV<���~�q��ׄ(:�V��$LI�������1!#�F���6���
��ٷ��{�aw�"F�M�#p79��&+�c��"��Oc�aa�n�����3��߲�rR;��v<�D^��YRӯ� -,��H�`�6(j;-�����'�+
�L$>���V�|�HQ�um}�چB�9�g��
�W�A�P�����)�gW*����bX$p����*m��oA��5S[\� �m�����q�A����ɛE�4;ϊ�����Kʡ=$�M�Vme�VN#[����ɋ����ee�}���
�4�lV�4;0��h��t�fȂ�r��Q����.^(��&���k6�}*d������V���!Bp�%��PQ
�Q�M�}�vAB��hO��DN�YW4+dء��
�9[o�պd�ۻM��d@���/�9W9&�\gJS������GP1bk/�4%d=�	R:���3ݏ��aD�1�;�v�u�:�{/
'E&�F��e�� ewА/*���j�z�����됤"V]���D$j�ӄ&B�'�E=�`ߪɛ�	e�:rA<nSR!>��-�uv޷�ks�ðV�u�@;ir1��b�6�
�#�!���}�˘ſb)�Ľ�!�0PzZ��4tZ�1̙�qֳ)^ U&=r�f&��|9�&�T��A�k�����zBs �gtp&Yx����8�)W+����V�!�s�����N��mK����MXeɎDm����������q[�c�#����@M�g�`Í�U��''E��Fp�ܛ�?{t0�>*��F 4=�U�;�'�-,�J@ye��z�}8��4��9��0nƁp�� U��p_�djK.�F�Nb��HrR�91ۉ�.ܧ
��RvsQ9�� ����������B�`1��-�f��D�������讯��sz�z����>B8��##+/��@z�79�eU&�|�f�H�=�B�p{���TԳ������(�TA�Ԏ���a�h^ �Еi�&*���<A/Q�.s�? ��[N�W�vUi��/��� ;CO��Cc��D�������ۑy�)�}'��P��A���zC����Q�t�PTmR�SƸ^���P�Cu�p��u�2A����(��3�c�>�sc�|
��.��$�x�8��3g� F��F�[w�����%A��~���`��Iܺψ��<�wj��T� X���7��{�u���^�J	���:�VF�4n��[;"͑���$�+^��CBׯp��p�w���HY��`�Ź�0~O���e
��̅��@���c�}e	�7r.J��©ޥ�������K�@J�OW�V��p_��W�)'^�NwdP$O��Ù�-l����G_h�ndwn7��c����9��Y�^q�lWwH�Q���W����Ƃ��'���9�P�~&��R���j�f�Z�Ɔ�b�������)\ ώ���űg��L9�e;�$���M�.�K� �8�E4����(��zr�,[����H�&�i������و��L�<H�p�z� ��<{Ќ4	�+,���S�i
����>����X��b���bٳ���y�ƈf��gE:>�.�+��f C�Q���k�sK�7!{�P|a��.�"4�԰@���_?�:�fRe)�{x�B �"��F������U��:�����1h���f�y����e��HpU����5'c��&.��/.W��֙���KjG�!��x��.^;<<J}]��./�:84��7��-����	�����}<V��� �Θ��G��iP��~��	w�N[�� �MZ���(�H�'Tg�=P}{���y������mk�6���n�h9��5�8��n%O���	���Q���}+d�{���Q�Jɕ�+իG���h��t�:uЎ��T�5�UB�J,�=�\Oq��ok�����R&���g��Z��	��(�D�q� #2o����$I�f�6�cIg�����7_p8q�q��F�C�@V�+�K2��L^���@;��c <3�/$oSX�y��r�K����Ws4���\�n%�m�f��YX[�}ɺp�T:NIXY����̓[j%�4��. ����&���@.�C
����f`uĄ��c��O+!-oQK�m��1!�Q�m���٪��'��v��{B�KX}%�f"�����XP�]����*���������f��VKDWx)fЗ��R���aG4��L4�8�f	��ď3Y���U���*;7��R�Լ��<���J������%=Rs6�_9+�^�fBgrfe衑�<��8�,*e��8�t�yȕ��g��lw����iS�=v6A8d�#HPt�Ä.�M@��S��&/hM�A�q%�r���gl���o�Η�3��Y�������b($��ɋ8����A^mԤ�,�����6
q�(j	�M����W0��V��,�c����k�Mf��`V8�������Ppxu���O�H�?�3�0���i\�����]�-!D#v`.`��5��j�o�ܓुPZn�xjM�d/6w)�@�?�l�a���{����3Z�����$6��U��HT�8gC�Ő�N1@�+�_?�S����f�p��]����l� �?�N"��D�rX��<�vm�]i�"�]D/�6�.d��7%]��^�ꞫQO|��25��_QDYSed��7
+p<T�m�7:�ȎU��-/��>D����fO�֟b+� ��R����?� ^V��M}3bp�뷏��螮�0���B��e�-�}�"��dk�Ojp1��=�z���	��?���8�[:N������RJ�}3w�:�vP��R����l��X����2- ]��R烷g'�d�:�mf�HZ��@ x�s�����NK0_�*y��_:rUe��z;Q+2�>��09�f5gA��y��h�y$�K�J��S�pT��{���%��?p�7�LN`���ٶS2����g�։,d�3-y�|n�m!`Ȕz�׊��#=QeT�M,����-��r�|"��v����{[���{�̺P���/���k����5�L�MU�[�Yn ˘����\��lS8�_������m�DnYɹ�iQ����&\
��<|o29�Ի�F��n�GS6���\bW�R�����i��ƻâ�@>X�b��	',�~.��3[u��8L�î�Z����5s"��Ȧ����:Z0�g^Y�f�Y�o����	N�"a�ԇ��]4����z�|w�m�IL2o�L�tg<����v P��I�*�
��|�j�!"r�|��y�ք��7g�Ib�����4����S#��$��֘�u��P*��:�0i7�q��#�&G�l\$u]v4r���$B>V �07��U Fk0�!�V����k���> ��!�zϵO���1�ʛ*Xr��,*����}�:��;��$�˓v��O��M�)e�hpC���|r��#�����o�v�xBU�]> 7ɟ
x��w�2�p\���{�S�=�����>7.#�w�P�bo7�*�`qY9V���6���
���$�J�3e�d|��\�qh���n*�4�K����t���pek*���7}6�_�?w��v���g�vWi�J�xe�Vk�Lf��m�u?y^D�k��.� �dVR�����L��m�ޖ9f��@��+���$�+�^���jC�j.���6Qt���������T��Q� �@����^�ax�yE�Lx����.���^ fE`%)Oa��ZQ�A��Z�2;	�G�I?p���p��\G��Ǩ���(U��Z:_���>l0�)\������;�j� �n8J�c�`B�Ն���Y��%Fl�%����Z�ok����E��SZ;�
{�[��\���s���ׇ� 2��?ܣ�h�E�	oV�[i�8��eD��>�lK��5�@iv]��h%���� ���A�Y�R����ѣ��5�t���pC\�wC��߁8��Q�.�'
	�ԪP�sk:��Y=�͗���XTa���q����_]��Lt��*��	�����-v�`����H�W?�.X�N����:W��y5�ĔAdvF�[������?���q�y%�*% H�'��>h�s��)y�?��T~t���b��W�~��*��j�НD�b�#�os�inG�wp���a|�*�_��G<�z����o���.w��/|G&'ɒ�R��Q�L�{CF��):)��wk�6�3'���3|?�Q-W��ڙ�#��ԢA�+É,"މw���Ÿ�<��A!8�o�G��+\@6���}��<;E���F�y#8�"�]~�zʥԜ)�=���+s:��L���=&�� �ֻ��q�F`�})�����j��%NC@����%���~ָ�]�1v�p�۹+Sz���M=��DU~<��]2H�F�tv��hM�r�%��c݋�P
@QƓ|�f���BF=��+�e@XjIwK���A\�T�����C�q�z��Mm��ԮTkw�M��zJ�2/���{�O�(�*rCm�.�2�_{?�w�>�J�G����.�2� ��_C�mk�Ҡ�Tc�xu�j�G�7vL�5�ɲ��b��!�����vT&|��E��}$�Š�b��m~�!(�Ef/���wQ�r�T���.�GH��`�M�y1�����e<�]ﯩ�7������i�M}�I�r��i�������a-牍�(���fba�C��o�����(��Ydl���n��h0=��b�Zǋ�t`q�q�������ʯ��F��k��@��a�6,jJ���L��a�j�N/�!-����\w����MW����[������ic?�}d�7��]�y�(��G �$pd_�ըAc�:�����C�tu�=_�L~)��pr�h��<w��$a8B:��X�[�v=���59�1��� .^Ș�}��G��/D���%�{G�3$ri�E������A7�i�EΨ3���>}�Dx-$���{S��P鯕��"~�V�\��T66DN��&=�Be���H�3�D/�~��c��L��N��J����� y9�!ˁۄP������͗�ķ��;���+��jk� �>ͧ2S�w�bs�7-j/1iwx}Uv� {�D� �<�2IU�l��D[���)��E���V���[����c��D<6Y���Y�!�1���ⵐ��F�F>�Gd,Y�[��5h+&5�QTN3��4����j����P�2���@ÿ �A3�-��LGm�?W�D����UN��@���e�| Ҵ<�1�����^{L�?��aҙ���/�lޑ���Vh�6�.�9�Vd� =�K|���@�BL��K�]�9w�hx�q������U]I��'=�E*E��8�41���-B-����ʱYȅ�F/e%~��~�No"6���!Ƽ�QS�iQ�At�[�"Y\�օJl�D� ���?Sjh��o	��s[�����F�Ƨ�lu)5�;.v�	�h|���:���QY�������`35�B�WE}��z���S��R���'�0�A��s╢lx�=��B3����a���(���wO��W��f}Z�,��� �����avieq�zo���՟.��1�:�'Ð?Nċ�v�[���88�M��=-q�c��AV1H}{T���*b��{޶��Ы��(׶b��W�u�*i��q
���
b""]oʌ�n~�.w�p��X�z*� ���><G��۔*"�k�=��m�w��s|>���i��	Qe&��Oh�Mŝ)�N�r��*�2�Ģ[?CX�Q���Q-�#���J�#+�}k,���`́�ֳ�����;8��a�~T�+s[{��&�}�(�<�Ef��F	x8K�]��}ʼ�)��Ӓ|@"s�r9���\fd�QX���6߈;�`�	����q�!@���jnC����ړ�lߕf��T��1M��pYE��2z�K}�BR�E��~S��])�!F�M4�{\ƹ	c��C!b�pl
wHp��}O��GF�d+� �X[�w�����$A��.�1��H���
m{����6�Z�ű�2F��rI����L���m6�+2��?I>��G��%t���o�_����q��Iz�T��8u�}^G�YL�L���X���!����v/=Tl��������ŗL®��$+!��f�l���'ir����X�>}�7�J�0�������ܪ`�,L� ��%�I��;uMT��D��� �����@5-�՚?S��?)b�X'CB�գӠ�!����o�+:2�ۥO04�Lb���B�t�a�LuJ�	Eo�#C`�����Rd��@Jq���iJa����])aoMNFy�-vvfwkw<7�����x�>[����7�cVA�d�v�`{�0��(��G�-3p�o;Xc�����Ͼht,m�=�8�~���pɿK�����a/E�V9��c=�2��@��"�@�-�֘������/��Bܼ�g{�'�$�E�E�[e�L<8H�i�uM���q�z����,�$K;�ɲٶg^���� ~���M�y}�6����}�wB����_E�;N�~Ό�c����)���6�2��yp�f˘�qP�Ν��܄M�[.��V��(�J�F��j�uN�5��2*g�S�ݥ�J�j��w�\Fv$ˇ�UW �pJ2��×#�;D�~|�1�������gx�ܰ����:�$�-Y�V���X�bΔ1��&��������+G���YnW�m�=+}/����3يG4�BA�A�ˁ;0���\�-@;��D��3��;�C����hDM=�11N5[@���e����1��E�m��{�c����s߆3���x��Ph�p�����m����K�2�����yd�m�T�9NҬx{��%&1��G^��R�+��<�e���N�/�%�5�������<��,�±���F�N%��3Ҟ7`t��fb��q��I�ࠛ�h� B�����o��~�uvu)�'�`�7��/!:�m♒�!k:�#,�u�'�:�{�G�tF��mO�K�� 3���g�B������m\�h�}uڲO>�9Tf�����k;�)#�Y�j�\�I�t�kv��OѶ�H���)��n"�s�˯�z�}Z(�;�x�曒M��A&g����9Eб=I��5��F�UC.{��+��I���5̋��+*�u�jDYjK�޽�V,��5C�E�k�a�Y�Ұg8(fj��V�<#|2�K�5�&?��ု�7˼1�%	�$�H̑����R����H�idn�VMa}5^_�`qaF���/���$]c($���k�#�lu��<#���0�O˪�xp*�b��k�����m���E|F�LEQb��\	rx�ޝ؉�
H�i�(���d���\Edj
��M�,V�9T�B��Λ�'A7%]�'*ǃ�C",�@M��d�i#$���q(zn�����m-��8�, ���(2�������%!����Y���|>�����E�J�����=�����ob�kcJ�,�Q�%��%Q��$~��:nX��-%䕲��&{��&��`����U�prQLN�媍:�-%FG��[r�Ĥ~�8�Eoٴ&:�(�}:L��@�b֔u�x�
Ȝ�z@a�ά���l}��a�"�"
���g/&9]y�&`�9���f��O'u�a*���y3
�+���;ț�<�q����s^R JSd�dH/�����o;qN���yX�o�-L�^���VQ��H�P�mA�����9���NTe�;�Kڴɥ�&%��?�pgz�n>tFi��b�GS���D�Ǩ���8c�D��A?�ހ�(�xq�t�7�#c�俎���m)�IV��U������̑ڛ���C�ƣ�|��"V&�;�z�h��2�*�����Qo��r��(ʞ�j�f�/@�}al��sUd�{՝8bB�ro����
2x�U��},��B��O�IN�r�Wx�?�e�F
:#Jo~���)���d�����܀W}��\+����X���1��5�NK�dF,�	�2{����U�-���]>1�5v�������?�hkP��[������f�ԅ������+�S��i��h�]֖F��F-K&3��
=j�d�x�	)N�r�9�SǗ�� ��9�8��j���տ��^@�#Aru��&!��]l�#t�9�3�I�����ā�6rP>�.�C��Z�`����1q��g^D="=6��&9'��@kZ�jJ����4k8����Esd��tՓ&��=E��8B�W��f|!��sűm�vGű\k�P�LM�׻�(?�3�O��<מ�qNL�H8��F�;M7��$/m����'k=먲G[� ��??��삤{�F	f4SX�U���'@*�,H�qy��q�>�#Q�j�S��4��0َ8I��p6��]z��@��(�,`��Fc��'l&R��i�͜x�k��� xRsՙ����y6d��+��l��K�`�
]-����d̵a/�z����^S�2z�Kم=2B|P#� [���z~�������@�O���#˧B<�̧�FYTFH��Ɯ�x����I踔~N��D^ ���iΪ*~a&�\A�p�.���Ax���VW��/i�_V�u�;��7�ԯ�C��JDrB�����U_�mp�'tR�P4ǐ�
�C��������T1�%�h�^]�(P"[ouoS��|A\���n����P��H�B��Qe�D^��Mx�M���|N�r��[;�~�62%p������$=0I ����4ѻ����D�������`u��^��B�Ix�њ���h��V��"�Mo��%/��@^��C��p*����̸��AYE2��	�V0B�-�㾥��oӅ<�Ư����w��5hJ�5��jN3���w�6��n?J��%WHt�V��_/T��o���[w(��$�E��]�plQ~`�a�x_�ȸd;;ʱ���߽F9���" �l�{�Ld���ݏE����'�3s9�~�Ӡ�w���>&�<��.T���&֭�W�.���| ���YS�?��"e�:$��Q�.rf6 ѫ.E����\SY�)z�=[h����)�-`\�?������ǐ"�H�ѵz.z�� �x�,+�&?�0+��-�G�+q���W'2X�����_b�Zd�b%y�.xf+-DE��?.�
�*�h��f��L��sE�g�Y#�{Ӵh|%��.��@�<_SB���b)�k�{�^� O��͊#܌Ji�U׸y��0��P�
�d�ZV6uyՑ⩫���} U��;Hʩ'�9�&�BF/r�䰚��	�sGI����j���L<�ݵ]j�y/Ϯ�4��0�����	${ʇ<<�D"��4c����������s�B|�	�{TNP��dz,Zf�1�l.;��X�����{����x{ǽL`�
@�ҽI�=�h�3C5�o�2������F�|�?�BA7���E��ҸJ;�+��ؽף#��{��~f�����ýe�%JU���y\�{v�d»�?5
�:Y�����"�M<C(q� q�
2�ET�AyIy�6���+H
��s)_�I`qP���a�,C����F�KvIL"�k����'^H�I/�M�X)1��6�K/�)�T��\�P�%2��fY�#X���}��^�� I~���g�����%%SP��S���{��Al���ʀ�'��I*Js�ȵ�cGCoo�--3}����+�M�Q�2G��e���;暬�Yc��}+)���}��"fT�Q�ò��U��*���*���磻���Af�P�K�Gxm����o��Da�곐�s8���Mo��S-m������n`�I9ZR�g��y�$�s��s���[�R75�_}A^�&�g���eR�<��:O,n��˙�	tU��S
g�B�l;���Gf���A|��Nwtࢌ�[� ����O��/,WZA˳І6��c���+����8߻]�ۮ@�X�N�������(h�Y�O�b�����m�,�%$�L�~6�g(��rMv�ɺ���yd��c����^�}6ǤE�ƣ���W��P4Q\�����&H��&3\���]}��]1�T����s�!��`����y��j��������/nQ7M�E�6�"V��"��.���a�{B�y���'�2���ef�6/�*MxH�Hg���/��1����,q��S�|�4ى]&��0C�] <���"�я���������:]��"\��/<>�.(��7iE�rOt��)OC�X��4��>D���e(;�7N�<^>�{G��RO�ҫu�D?�\�*G���RصăX��"?�L�+��V�P�㑐Lb4wT�����[`���i�I���Ս8����fᙙ(k��TG�p���=����L��'z��|1����^��镈R�� 3;PAźΖ�i�C�O�鶟�2j !�R^�+q;d��o11ݬ�}Y������W���sh0#��y�n[:6�Ѭ�1Q�A^>5��CA�⏵g�oyˀ��=��KQ�����S5&#T�I�&����z\���7L�g`32��Sv���C���d��-�s`nEHw`ȋ��&��g hQ�⺑a����-8}��@�����4���D�1��?�|�I�A�k�c&�kC�m���5Q��q�� �Y�=��c����B�0��^w-�#�Ԧ��2�1n�
��-��� �& �����\2��j��)���¾nɌ�S����c��9�%:Ni����@����-�͘]������M���?�b(Z����r��"_���%��Zۦ�g���fU��o=��͆�"��N�L)"49y-��tR|�3w�foڀRt+����D� �>I���
�Wp|¦!�aw(�)폺���2�7��SI�x��r� _ǚ�)#�."$�jp��=��zV��-L�Q�y0����5�#	gD�0��u�q�46z��7�>+s0{U�}��t�!��	��Yk������������Ιj$��X��p�P�^[�~U�;�٭��6?   W   Ĵ���	��Z�BtIJ$�� 3��H��R�
O�ظ2�>�k�����4�?Q7�-0�" +�|f��+�ᅑ t���fӊ�nZ�?��R���'q�V:O����6(�Y��FR�hzy��'��*��ܴL�qO� ��Z�M3Dc�e߄��w �Y|��ya_E~��<}��l����d�U#���gښ��%�<�C�߉��H�"-�jU�H=��Dq�L� )R?#�<!�#�J}2m�6!��'
B1u�(X��=��t�#�C��.O�)k�-G1O�t'� �~��;�T�&d�>���7nS���A�H#<i7("��B�nAۗ�5�ޡ����	4�O�!y���?�4��	�	X6�����F�0	Dx"g�Y�'�p�'>�=6��e#���r�Qc!T@cO� :��	7@qO��xB X,�h���Q���:��i��Dx��~�'3�=�Gd��pR�s���K�ޡ������'�zEx�P~���w��a96Þ�K�$�z�ߓ��ǌ�ON�`���²H!9&J�y�.dZ�b�+�.�Dx��z�'�R%�	�Y>��� �I	J���k�!w�nb�h�P�	��'f��Z	{zq��L�h�W?Iѧ=)O�Ւ�'�����dd�ڥ�0K@(����u#�*3�i�F�Q��ǃ	�uW�O���oK; B�X1Ɇ�1���"\����Oҧ(h�O�|!w�T��'&6�����t-�d��f��gz�useH93!�Dy��DT�O`�1�"ĄH�@�`���H�0"O�#�  �                                                                                                                                                                                                                                                                                                                                                                                                                                                             �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  ��   �  �  �  �  7*  �5  �@  �K  vW  �b  �m  )w  �}  �  &�  l�  ��   �  D�  ��  �  ~�  ��  (�  q�  ��  C�  ��  ��  �  {�  ��   `	 �  F# �, �5 <= zC �I yN  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C�x,�]���O_�!aH�+dmP��u�U�8'|1j�'xe"����=����⋋w��Lӎ��'�� `p��+U�4���@[$#Q�@�'���3g���>��C㛃�<��'�h0�W+ �X�j���=��r�'���wi����1T�,�@���'Zn��dڞ?�N H������ZK>Y��)�Smb� �G���t,%h�k�"O~@J��2�\Y�rχ�Vr�(�"Oz�X��<ɔ<�E��c[F`���']�I-��<!F�����mJ�v�ܔ��'�aҀG��#.F78EdY��̛(��?1�'$ �Bh��e6TkB��H�8�'����ޗE�&�#_�?�ɫ��Dʜ�h��t��P�{��∑�[g�����Oz�����[��cW"&={t� ���r@azR1OP�Z�O�|�SO�p%�9�ͫt�S6"Od���+I�$L�h��C�G�����Z��t�E���G/P��9�ī�����AdQ��x�Ԟ2���v号@st(��֌I�B�IH�j%�Q�P,xs. !�kV�Q?�#?	ܴ���	��˧v�`�GC��`��CA( ���J��� �s&.qp�lڋZ&��Gy2�-�S�4�@�l�S��~���/�<�yb(�#	���  >�R�`��	�y�#X>Zb�*͟�:�D`�a̚��yb�[0���q�C@(�H,�SΩ�yR�'�zi��@�97�AC�ʚ4(dT�3�{RK�M���g9~��3"�u�@`[+��Or�)�����d*эJ�%�h�Ey2�|��
��B�4T#f��+w���[�BC�<�K�%!i$Xa�g�)�&�����$A���?!�'��S��O2��FƗ�*��IV���R��'��dE�D�8�K^�k�F,��٪:u!�7/ :0Ђ�](-e��SA��"^Iax��	 m"\qC����&�<40<B�I#MD�!��
���`.�$�"�=����0����� Yn�4� �O�ĺ�G�y,D*Dv���G�F�P(q��'%ўb>�8�hܧ&U�!H�֩,�̥ˤ�.D�2-��_���B��K�z��'#+�	L؞� R��7f��x�f��wh�^�*x�6"ON�T��=%�ݘvf�P���9O&�{��E� ���?t��x����3�@��ȓ"H��ٳn��.� bHW;Jx͇ȓr7l� �N���^ip�a:%zZ�ȓh��H$���n�fYX��ǲ�ȩ�ȓT����*��"X<TЧ��-D��ȓw�t���)r�)(�h��m�ĄȓAAƤR���
��R�K!/���ȓ ��2���4��� ����j�ȓO���#�e�~����؃d2��ȓq�|+�˂!�$���J�8P<C�	-��1�A�+L�$#sU:��C�	>ii0�RF�C�%Š�ٔ�-z�C䉶W5b\���7f�qX�ʍ='��C��;T��<C���O?\0+�A3 ��C�!1�>�`�J�1Pt����vìB��6�f9ᕡ�5_H��V��+�B�	^�;w��V�D���(B��2L��<2$
�� ��AJ'�O�$:B�I,��LC���p�t�����C�	�>E�㩋"rTF5�c��.)��C�3�-	���<�a��,�1[�\C�I�USZ��Y�MT� 	�0~�C�	�f��Y�cI�u��	3ݜR.
C�I+�Aʁ,&	���q��/k=�B�	J^�� �μ(t���aK,�B��F�����`��3,4����y�NB�	>ڝdGO0^}�G�ŵf�B䉻~�@D�>=�@a�@��a�C�	?k�����,	�h-QDo�q�C�I�e����ߊ)pL��G�<ĠC�I�(�V�c%�M:)#���d[�,C�	�J��-�2 4]*q��ș>C䉙r�ʸ����	t�1B"���B��%i�����	�D]�s+�)w��B�	�L��(IA,T(L_r��g�Z$�B�ɕ1�����T62�X� ƍ�ӸB��4*��jF+���g�r�B�I�rȀ���,Q�x�
A ��>U�XB�I�U3t��X�
L���*UPB䉴?��B�?p`�pf�A��"OTX�0'�9�&�"�	��A�ʘ��"O$j㮇v����h����nY(�y���0 `*S��F��Aq&�yb��k���4ê?�4�Z���0�y�KjFK�9��)��3�y�Y�4Bt����R�A��C��yb�Չ�V���F�?g't��R&���y����ph�RƯ,`Öa@©��y����hٴ�:eC^�Zu��"h(�y�Jɣ��Z�O�$NR�BBꗊ�y��(l�	Vd�r�<i1����y�E�2�©�UoGm��A�#�y�$�4����!�X|�$"Т��yR �bH�����,Rp̵@���y�k���c���[%�}��lċ�y�.,l��$��͍Q�~x�q�
��y���X�@ʚE�TY�A�W��y�h@w�f�m�$GlSTFG4�yr�J�4k8�8ǋ�A;F!��m���yrN9��� &U02�������y�h��v8���P��&@da&c�0�y�ϝx��y�VΒ�$�9�0i-�y
� ���G��I��D�1��%N��f"O�HAgN8$h`X�$�����7"OZ ��V+
�6��`#�%x��U� "O��ۣ���]�-S�A�I��"OP%��nC�Z�3U�z�����'���'Q��'��'���'pr�'�����$�V�q� �����':B�',B�'^"�'�B�'��'4X0r-�xZj,�W�N%1�'�r�'>�'��'l2�'���'��`��,(ސ�!gB����U�'.2�'=R�'�"�'���'���'#�����]�a��,��"G07�.� ��'g�'���'���'���'���'i����'@q����NQ"�(�p�'H��'<��'���'P�'{��'F��H����'t�*�Ô�� C��'8��'��'���'\�'���'<�0�8&Wl(��ɏt�X�r�'`��'���'���'��'���',nEQ0��1R��q�Ψ4�hݩ$�'H��'���'���'R��'�r�'pS􃏑+� ����Qp�R����'���'���'��'!��'�'��i:�3X�z�3�W�l�Ĕp��'^��'���'���'�R�'�B�'PtL��E���y�J�+Ypijr�'aR�'���'�B�'���'S��'o�]��+�\�QkO}��u�'��'���'0B�'B�d~Ӟ���Oȱ�hL�wBajS�
�\'�}14��\y��'��)�3?��i��ГF�D�^4���	��/�7V͢��'�6m'�i>�	����� ��d�P�į]ӈ�zÆN�X�	(*�pn�}~�1�$���t�I
�,,Ap,�&~��\��6I1O��$�<���)����q�A^2r�܀2�.256�m�>hijc����p��y�Aڔ ���(��S�CҀ�SFE!_�';�D�>�|"��N6�M��'i�
0$GA	|�����=a?�DJ�'O��G�����i>���;*B �A�l[.͜���H�(;.�	[yҞ|�|�RA����
���#F��`�"�Xq(\�6��⟰ѬOl���O�	f}��ړ~������C��������O:%(�˹)�1�:! �)�0�$�}������Y� �<Y��<4������O?�	�#���� ߦ$F��27�P�|�8扆�M[Tl�|~�k�6���A����j����)A.YG<�����Iߟ� V	Wئ��'q�)��?a�v��}G��`�K�K
��Y�̕B�'�)�3扫Y���b2�$&8���ąG�0�8�P`��/ŘM��'�b�i�?İ�ĥ�\� �A���r�,��'5�'�ɧ�O���'�_�vqkS�ؘ`T�ӅP�x�Qh�^�P���CV��i�IRy�_�y�9��R?\M����b��'_��'��O3�I�M�2&1�?Ag	� ��<���	�U#�샵�-�?9$�ip�O4�'Q����*��!^��Qu�,l������Y��oZs~b��*Ni���'�O`��н�ni�ę�$�@�¦�K��y��'��'2��'���ɔf�E��hd� ��u�{F���O~��W��a��G�iy��l�d�O�܈���*Qavi�a�$t�8�V ,���O6�4�v�0Br���17b�A�l:O,�`G0c���[QI�O����r�	gy��4k�\�e��"������ǚM��48�4v�[���?Y�����|�f������Gd��ⶁ؞!W�	 ����O��$6��?iA�G��>�<؋���/Y}�C��$>D��%�ަ��/O�	G/�~�|�&=�9��ȗ�L��Ra8q2�'�r�'+���^�h)ش@.����6l.
U�B#y�9e"L�`�n�����p[ٴ��'Qh��?y�i۟xD2�
#h]�S\QP$��?��B�8�ٴ�����z�'����4hs�5.��8F#�=,\�Cy��'�r�'<��'�[>�����	�aZ��Ɂ�\�ɆA&�M�D��?)��?qM~b�ƛ�w򂡛��H
& \8bHD4B��@�'�'җ|��ԏ�	]h�<O���7�^�^}A���3�Y�>O���~r�|�Y�����D��G� ZW\5���v�0���ϟt��Ο@�	yy�s�4йQh�O��f�3"θ! �� ��Q+Ĭ$�I���$�O��$����Lɦ�s�&A�<�$$�h���-M��E���	zېc>}���'ѐq�I�i�ʐ�E�˵e���H�f�lI�	� �	ğL�Ix�O�RF�s0��1e*X)���Q#�7Mi o���K���Oh�]��	�?�;��
b�'�x�؁=�p�Γ�?q���?)5�+�M��O��t���j��C�n�*a�֠Ӄ�&����(C:�O.��|z���?i��?1��]��1���]�"02�k��^6���/O]o��>���	��,�Il�S��๳/�!k�a�Vf�o.i#�-G=���O �;��	_�T^(p�a�0�@�1m� !)̬���b*�˓@�0���j�O���M>�+OV��b�j�0�R�s���ن��O`���Od�D�O�<T�ir�)���';V���k����Ǖx�HC$�'C67m?�$�Oz�'�"�y�H޲d� �h\#uԘ��_7�z��İi����~=�|��ܟ����� ���4TB(вDfL%�t���6O���O����O6�d�O�?���/*B�����18cY)��
ߟ���ߟ���4cS�Qͧ�?�G�i��'R&Md���DK��ZFfߦ(k�����|B�'+�O�h��i��ɔIg��w*��p�Bn-9D� ��~�"�@G�Oy�O�B�'#R�4GJ��
7CU!a�;k��z r�'s剠�M���ݣ�?���?�-�q�e#��0C�gLfa#7�����O��D�O�O���t���Q�^ O���\�_���H�ρ�A��Q��hy�O�f�ɓ��'C�ّ�2P$�\�0��n�b��f�'H�'����O��I�M�`AD-=��9���	i� ��[�R�$����?ae�i��OB��'�"mw�V-;7���%�XS��	�e���'%��Ӹiy�I�U��1���M ��=Cv'_:x����cb��b��<���?i��?����?I)����b�KZ<��LD }~�lI妩�e�˟������%?��I��M�;u�T�6�
,Vo`��l˶I�,�����?!M>�|�����M�'�ĥA��7y@�Y�n ��*�@�'M�ɓ��]E?YL>y*O�)�OF	��A�+��XCSH�K> ��Rj�O����O*�ĥ<�w�i�"`!d�'*�'�b���I�(zD��8�(q�t���b}��'K|���^��� ���?I�����ղ��$R5�lwakӴc>!� �O��d�Bt�������,�w�A'.���$�O,�D�OL�D.ڧ�?	���e��V�2n�)�VHZ�?�W�'��%���?aq�i��O�0�@Š+G-R�V1�a�\��O2�$�OH��DaӶ�Ӻ#c���R��_�T�� ���+�~�Ӳ+�VEh�Or˓�?i��?Q���?1�s^Эs���$Du�"SA>:��/O��l�s� �����	R�����A��$ul���d��d�|Ys�<��d�O���*��)H�0��&ځ|w��J�
\T=b��eӶ�<l,e�衟@'���'	rS4㓭mߔEXe�ݲ}��-2�'��'�����P���4:Shi��1����O@�nW\���Ǒ�*���O�V�d}b�'5�w�>��&년W�����	�_����7�S<Q��ƙ��C�_�Nf����a���]ʵM�$��JR4`%���x�H�I���Iӟ��������d��k�����O���M����?����?1��i�n���O�"�j��O���4k��Ay��]� 4�8��.���O��4�J\I7i���>�D����(d�iJ2�Q��MPr �����D�&����4�*��OT��\9R�{2���.�T�#��̮e�\���O��*��fdWR�'�2V>cK.x���t��/N�(i)�'k���I��D�O�$6��?Q��/�]���Db�"I��Ys�M�/��	P�	���.O�iJ��~��|�ȟ?KQ�lq�VC�9Y��ac�'Z2�'&���d���.��Q����4B楑����C$��W5�rs�����զ�&���	!����O� aS%��P��r`딱4'�Y�#L�O��$Ж"�87�b���	U�����OcN�7���1&K@)����	&�|�Γ��$"|O"%X�l˱9�\��.[���7iTɦM���ݟ��IޟP��׶�y���/�*`q�N	�n)�� �HB�'�ɧ�O�Vq�T�i��� 8�@m���������H:}~�D�'������O���?��6��##��Y��Ų�Iޫ|������?)���?�)O6�lZ7�`a��͟��	}�UA����Ԉ����[���?نZ����Ο�$�`9Gi�b�*R� D#R"��s !?��G�h���W��Ņn���䀎�?1"�؂+�<P�G�L��Y�%.��?���?���?a��9�xq���z����K�#�`��O��m�((�"`�I��4���?�;;FI� &�>b�Ȁ��d�+G| 8��?!��
شX�.u	ݴ��䃓q�4���O"<�れ.(������b��9�|�X�D�Iٟ �����Ɵ�X��d��)&BK9=��1��)EGyb%}�Ztc,�<���䧌?A���0Hz���R��'o��E0�e�r��I��x�	Q�)擏n�pWZ�J�]3�̩4�@�Q�=C�f
�<���H���If�IeyB�O�u��d�B0d�Y9��J U!2�'}�'��O��� �Mc����?�vF[�sֶ��a�F�iV�d�ab�%�?1��i;�O�Y�'sB�'��A�W��$�ԯPȱAsE�F��p�i���Q�yy��Ocq���K}��8���
C����Fe�j�$�O���O��$�O���8�S�@�%�qm��6���@
<(�Ƚ�I�h�	��M��FS�|b��mr���|2�7���z�(�8�P$P���j��'L������ΌZɛ&��2�ō�xEV�i!V�Os�݁�C](e#����'b�$�������'�b�'b���%��#9r|@��ژZ��P��'��P��2�4w������?������1�Z$��A��ʎ�w��I!����O��%��?�"�o�v��D���P�EWR])�CW,"��$�F��Ԧ�j+O�)6�~B�|�D�v&(��eĐ[5lE�t�ϳ>��'��'���4W�,aشN����\%��B�`� @�T��g��?Y�T���DC}��'��a�0*�!�l 5`W�D��M�7�'�H	G@����֝�!�p�өD��)� �����%Y�5��"$s���4OD��?1���?A��?q����i"^zpM@w^!�����ْ1�n0c�,̗'�����'@�6=�"��P�Zs������.[�Y`�'�O ��:��)��H7�i���������	���C,m�\�b��p����H�ry�O8�%lu�=p�@
�rJixbd���b�'*�'`�	�Ms�n���?���?��.�!Uv�a��C�.��踷C�$��'zH��?a����h����l�|_�0�0'�;�'���`�$Z��v �����e�ܟ(��'v�aq�a״e*�l�Ǔ3
[zP���'<�'S�'T�>���/+2P�0F��dc�y񭟬=���I��M��`
��?��I�f�4�Vp��fƳ{��pƬ��`�l�y�=O����O���� ��6M+?!&�]�\cX�S�-���sO�(�>�5�۽6�A%� �����'���'���'ٸ�+Ӈ��h��9�`IY:h`�R\�j�4)�dEC(O��$6���O�9��j��2���:�E�d��}��dHt}B�'��O1����>�V�Q�N�?3nV H3k�]!J��3�E��ͬ& n� ��M�Ob˓]r=���լZ��M ���;l p�
���?���?���|
(OX�o�s�p����ЫV���k�X��OQ�CTx���M;��>!���?��8����J'�®Σ-D�5q�G��M[�O���䏟�(���N�3g(�m�U�ٺ ���h�(ˌ0����O���O2���O>�$0�S1i����N S��k�L�G�����������M� +��|��Z����|d�j�hҶ�G$6�|�f���:D�'�b������]o����E�Z�̠3��F�h���#�i3���0�'�h�&�������'�B�'�,�;2d�
�Z��Ц���2�'
�\��ٴAC�I(O��d�|rw�h}���fL�_2h0�$�(���؟8�	v�)
��Լ���J��#�D�� C &�Ӄ��
y�0��D'�ƟH(`�|�ɅR.n}ʄ͜�+J�������'���'����R��ش�By��?
=�TЯ�52�@<ȓ��'�?���A����A}��'p�Q���?��2G'c|;��'��gC�8�V���*�)G��d�~�Qj�#	|�(��\��ȪG���<�)O,�$�OH���O2�D�O��'�\H�w�D�W���e�&zjF�@�i�,h���'���'(�O���n��NѕbL�r��t��vf��b��d�O��O1��r�v�T�I0}ʒq�d��0LdH�Ԥ�1%��牗I,�Tӄ�'G�=&�X�'���'=.e[�cѲ�°1ƃ�{��d"��'��'RY��8�4)�z����?���R��,�+��\vp �s <sE��M>��LZ�Iϟ��I_�	�-�B������x0�g�3+��b)R7�[ ��V ��ӷ�~��'\t���DB1��e`��A�y)t��	�'Xh܉��D��Cʀ>t��-@Q�'(6��Jv@�$�O��lZG�Ӽ3 -J� p
���J�xL����<	���?��|lnE@�4�����L;������fB]�lQ��3!�0I�&�B�S����d�O���OV���OL�d�B�<I��PN����ei��=$˓[!��fΠK�b�'nB��T�'��%� kī[L�h1E文HF��c�>a��?QH>�|�O��9��k1��6C�1"�	�^�d(�!�J���Ą'ybVѫ��.�X�OP˓)dXD#B����@�X�`=�y:���?���?Q��|�.O*�n��M�>Y�	�zm�Wd�ط�D�'3̵�I5�M+I>1��Uo��韄�i���}"�2-R�~����Z h\�,o�m~��k�>�����'ڿ;�ן@�<p% �5(�ujT��<���?����?���?���?F?LT�,�'X��N�]D��'���uӨE��+�<1b�i�'�&8�"����G�G
7�� �ǟ|B�'��O�f��p�i��ɿ	�ɻ�)�`Jjuy�.�u�v��k
8+���"�ļ<����?9���?i��>	H�Q)q��&���X�	��?I���$��-K�K�ʟ��џ��O���1��.W����v�
�<���O���'�B�'ɧ���V
J#/�/��Q�SbL"z[a����7�V7m8?�',W���p�I"4&����A-V�|��'��x�j$��џ��	����)�Spy��hӒ�z�G��K&DE3KC�	���y�#�o}�ʓM��F��Bl}��'=<����^Zk�T��A�m9�����'(R��Ln�������֟#Q�)�<)%��64 ��cE"�8�R�Z�<Q+O:��O&��O����O8�'�����(L�l��L%/N`� �i��u�@<2��'%��\y��f���[�?L�0B�ԃVZd�6E����d=�i>�����c�ƍ��ϓr�a�(^q���FE�H��ϓ�R��5G�O�N>�-O��d�O>ĨяK�M��� 	J�e(�����O��D�O��D�<A��iB��$�'�'�D�fPgd�D����y�0��|2�'���?!����|M�m����-C`Y{f!L;T����'Y���F
�"�{��dK����{��'�T�ԃ�-�d�Յ�L|��"d�'#��'Cb�'��>����BY�UYc�]UbF�O'1�H��I��M#s��#�?���]��v�4Ａg�Ls��<P�e��%r(p0O�$�O��d��WN7�<?�b��K �3� �[C�?3�(!3�ɢtYdɐ�E=�ĩ<ͧ�?I���?���?�G�g�|ykFl"PEp��c���������0�Gޟh�I�$'?a�ɦ���N�>�\��W,X��O���:�)�S�r:A��A%BPԉxqOA;�tuJ�,��-2q�'���5i	�p�T�|rY���mہX��Y�D�t�H������ݟd�	��Iy��x��a�@.�OR��F@�N4;���0�r̘��O�m�I��x�	؟d����R%��?&<�Gn⢜��M�Y���nZk~R��44�P��O|�O���]>{*&}�e�I�+x@/I�y��'XB�'�B�'��)� �Z��ռ`?�%�Q�[������OD�Z٦��Ugr>����M�N>y� �f��% �n��TȘ�P��ѝ���?Q��|�ݔ�MK�O(�D�^&N4��
�=7� c���!8]������R�O���|���?i���E�Α.Sm�s�	;PgH�����?Q/O$-m��� ��	����Ih��iG4b��9�Iо@N�Hç"S��y�'�:��?�����S���iېԙ��.+p A�]�+.���cΔ���*3T�擋8T���B�	�f୨#�ْ'NZ�#� @K.,�	Ο����L�)�wy"�`�0�*@��(z�d���fl�D�:/��d�OF�m�T�Wj�	Ɵ�X���l�T���
�!�И�gKOsy�j"l������FHE���D�Ky�)��9��V�}dJ���ݞ�y�]����I�\��`�%�Aǘ��� x�l��4XP����?A����O�:6=�vE�b/Y-`��2Ci҈f����b�OR�D)�󩜤YJ�6�c�I��M�3�V��0�έf�X���}��8iE-	��D-���<Y���?�f�_�hX8�I�X,4�����?����?������ͦE{��M�x����p'anV�UX��O�
�L�QQ�D��|5�	�T�Iw�h�F j���h"��y҃Ǡk�����hu�]o�hq�|�e)�O|qY��4Ln��A�=R�"��ď'Na������?����?1��h������#�� �=����cʀ�'��d�����Gڟ�	��M���w$��Ï�Lp��yu�D%R���1�'��'����Iz�F����3R������;%Z|K`a5p�nT{�%��IZH8Ö|�U����ȟ|�	ڟX�I֟�W���0:�@���U��tr��CyR�`��U�G'�O�d�Ol����E?/�lKuI�O�0P�o�$"8���'���'�ɧ�O���c
�TrlI���3[?�q��B�	���Gy�Ø1yp*8�	
U�'t�H���@@�

f�1�ݫN4��$�ڦ�1c�Ɵ�&�"D
��A�m� 
���3����(��4��'���?1��?QF�[��I�E)� ���@2�[
" ��ݴ��DɤC)�����~������Q%K��4���YJ�B	%�ȅY6��O���O
�D�O�$=���%̎0�q�D�t���i��N;�y���P��/�M�ׅ �|B�J��&�|*�>x�NQ��m9C���p��*��'Qr��$�O9n��V���](x$�(ÀoԀ$R�ԁ��%$���B�J�$H��|S�h��ğ��	ǟ�p9�#�@�A��AEi��k)������?�(O�l�H��Iğ���w���Ы֔5ҔȠ4�	a�ME�����W}��'�B�|ʟ�0�����Mt�-��"k�PP)��	�F_,� ���-����|"p��O���I>�j%�x�@Q`�h��1�0# ��?��?����?�|�/O�0n�#�M�R#�+J�Ș�狔E)�0ğ��	-�Mۊ�c�>a�+���Q6s�II#O�.��]����?YT��MS�O|T��-�8ĸO�.q��O�2:��ݡ1��ng0d3�'������	�������,����G�@����ͭA���NN�(6���=����O��D9���O��nz�A$l�:`�v�)T,��!Y��ܟ(�	]�)擨&^��n��<�@����H�g`�=?���A����<a�I�4|P�Ir�~y�O8�CZ,j�Ё�4%��YICBz���'�r�'`�I��M�&ђ�?	���?�
�h�\!�N)�0NY�B�>�����'�=c%$K%4%��R2�z���OHP٤���脋G)�I��?�g�O�J#G�,נ�hÊ4>���30"O���K�X��\Q��"D�R��Ł�O�$o�=t�6��	ʟ0�۴���y��εE[��z�e�?Q�6�����y��'9��'��jֲi��i�e�ѯ��?u[4e�u�3&ц6�j-+�'���Ɵ�Iʟ���柠�ɘfjBE� �ȶp��P�#���~����'�7��,��d�O���;�I�O�m8�'M�\%���ϊ$St]�� A}��'�R�|��d,��:������Ã�_�����iP�˓TDP����&�,�'^6��F`6h��mi�J��~��8U�'.��'������S����4␘��I�ԕ� ���A����E�̂T�*p���J��&��`}��')r�'������:&���6A,c�#sa�_w�����A@�L�+n�����t��T�ޟ����\�W� �S�;O��$�O��$�ON���O��?U:�ŅT���!�;]�J���x���d��4f���Χ�?Yнi��'��,8\ή��g�؊8��l��|b�'&�O4(��v�i��I/�n� �`����!z�8c�'S�c�"uCN&�~�|W����� ��П`�T@դ8���j�@"�4�j埄��{y�c�������O����O�˧!V%��^�B����f�;�e̓�?��[�t��֟�'��?�ڵ��ǉ�����`��q)%��U�S� ��4'V�i>U��O>�O$`K�,��AT Q0C�_K���4"�O��$�O ��O1����� �*��@*���
u�0r�%&bPZ��'R/bӸ��q�O���=%�� Q�Gѝ$��	"�J�%`��$�OҼ�2�b�"�Ӻ���S�Z"ʣ<� ���@�x���x`��<�(O����O����O��d�O��'z�b�x�,�,y��Lȇ�ȾI���0v�i��'���'��O��a}��N�3|��u��s�ԍ��L�p����Oj�O1�(�f�gӆ�	�H�)�"�@0�"�K� \��ɂ/���OF�O��|���iv"�k��O�w� ��6FIa�����?i���?,O�\lZ	/������p�	�5�P�C��#��(��.�_f�'�������O��d0���b�9�f�6kF̜���̒x��� m���c�&H�%��'?�s��'����7~����Q��~!vxZ��Ƽ)�C�	�!��Ɓ�ZFNlKw΃n�P���.�M�2�	�?���~>�6�4��)���ǳ�$=c� �y��0��9O��D�O�d�w��6�!?9�f֨4ͮ�ӛ"נ�"�ڻ
S�k#�]A�J�$���''�'��'��'"�Q�����
e��uu��k�S����4O�8����?9���O�L 5�5U���ϐm�4��%�>i���?!L>�|�'�ɡ[Z(�����q�!ݰ��æ����͇Y�^�I�JS�OZ�z����Xd`	��R�+ ��3��?���?)��|"*O� mZ=���	<�:�"Ė�ȩ�g�����	�Mۊ/�>�����D�#�(b��"(�~�;��ǣ&�*��&�j�j���X��(㟀�O~��; ����4E�3d���ɤ@�Q�D���?q���?)��?����O�N)r�B	k<�7�-����'*�'�7���$��	�O�lZD�ɟAW�h�DL�&�tI�G�Kƴ�%�t�I����3�� nZS~�gP!��r�A�3P�P� )9�MI���h?�J>�-O���O��$�O6h2V'_�if�z����HV�[�/�O��$�<��i�J䣣�'s��'��ӯ5���a�^�2rJ�8��ܝ|���ҫO����Oh�O�ӄa�j8� �\�.! ��'$~�E���'
����e�Py�O�,��	;R	�'E́�F�^<`KD�R$^���3�'%��'kr�O!���M���� (��c$͝\G.�r��2C��D���?���i��Od�'�R�Q�@�~4�ԯ��~�I�o�H5r�'�*DH�i����c,�#2�	�$�@ SrA��9:8�ȳ$ϧ4��D�<���?i���?9��?!+�֍��>o*2�"��ʰ47ڱ�-��	UhEgyb�'��OWff��E���i'�^�,�a�+?�d"�)��)�0\oZ�<�t���8"2�	��^��$ �C�<�#��T���dM������OB����L�b�J8nm��c�B�����O��D�OL�W�����?��?A4"�[�hWiO�
fZy�%痦��'7���?����na��	�B\,I�eiVeW�Y��T�'9�lʢ�uƛf�2���~��'d�؋��+��%"E����'b�'b�'M�>��	<gĜغ�ڠ�n�Ht‪lx�����M������?Y��>ћF�4�b��$���ƌ�v*��8Nd�)�:O��d�O��
;c֎6-6?9�"�`@�I�����ғ��|vـT���E��I>�,O��OZ�D�O>��O�h���O:�cv��Q)�lq�n�<y��i��B��'2�'��O~	�#y4��"j!8�R���h~��?����S�'h~,`׊[4^~�X�a�P���ݐx9x��ʚx~r+Y�!�p$�	7q��'��I?~1��i�sUb����/���	Ɵ��I��`�i>�'׮7R����љm����Ї���r'�? ������?�w[�p�	Uy�X�a���bnRz�HD`Q�!���3�ip�I�EÆ F�O:��&?%��
pL�Q2���)b���5��4���I�d��ʟ(�Iٟ0��s�'��i�_�N&�ܯ�@2 ��a%�O��$�Oje�I$7W�	�O �lZn̓XyD�Y�l��Z�{r-�%O�'�8�����S+��mp~�.VQ=�Q��E�I��� ��O=�y�bt?�O>I)O����O����O���̢�.E�M$��m�B��O��d�<�v�i-~��"�'���'��S�BAp �@�/OV�b�##����ş�O����O*�O�ӛU
q���&I���T)T����Y��P�d�ċxy�Op�E��-b��'����-��"�bWDT3r�'���'5R���Oa��7�MC�
L�B�ޡrq����*mT*� Ȁ1���?Q�i��O��'`�ɒ7OW�dR"'	S�ƌ�u*ߍ���'5B|�6�i����&��� �O)�'{�H��v ٛu�.<�D��D�,�̓��$�O|�D�O����O^���|2�_�SSB�qԡ���P��򛶠R>��	�$?	����Mϻ`r�i����Fq���7 �5s��	���?)L>�|����1�M���� "hs��="D�!�O]?� �y�4O�""��~�|�Z��A�܁`M��x �Kq�^*(o�|���M�3땸�?���?y3��2L�y�FD:\
�� W3��'Z>��?����q��-Å��rP�	!��?v��$�' ���C��ba��ѵ��D�J֟��%�'�4P��Ƞ�`m�S$��q�@����'�B�'��'A�>q�	 NF���OU�h����Q�!H5�	�M�!�?�?q����6�4�0�����\?�;4��>���A:Op�d�O��$S. ��6�1?�����y�'�:Yp�]4����ƬM7s�X�%�:�$�<���?q���?����?⦈�]w����I2bz���I^���@����5&�ٟD����$?M�I�(�b�zw�݊/�� wjՄm�s�OV��O"�O1�Is�ʊ�F�|��E�,!K��3���%S�R;�ξ<R�O���^�dYL��lƎ�"���4'��%���m(|��	�c��Q�ƅ^���p�C��HI�fK�'���IF�Y@� ZD�	_�h$���ɛj�XI�3����*"`��ε���5H/��C�·��dT�j�Vx9��	�jhX!a@�#[AV�v膐Mg�d�@��Cf�40fi�7	%q���I���p�$�Im��)3C^�p)¯�wp�q�o�)5]��A5�D�,�BC�
�"�୑-�0@Ĝq!V'�:B���R����Y��ITU(�l��V��(9�b+�*u�Y��'�`��GG�6>n��K�huM��j���D�O`��*�d�Ob�Y2Ww|���H>`�d�l�"���Ki���?����?A+OlTJ�-�D���'?L���Η-�������7Xj�k��l���9�$�O��
�N�R����=Z�̸s�LAy�x�@w�����O˓Go<���Z?	�	ޟ���&Tl2݃�M�<Qdf] -��L���N<����?Aw.�"�?�L>��OĊ�w�F�	\�7(��	�v�ܴ��d�	mȴ��O���Of�)�<�1_e�jEB��fވK��Z�I�,n�����`�"<�~���ڜО���(�p�i3	Aݦ]1%% �M+��?I���BVW�̗'�民�٫D�2���C�R�'r�ba�h4��D�'�?)�L�+ )�q��(�(e�q�ߵ$'��';�'D����>�)O�D���*0�	$� �"���1uO�i�a$���y��`$����������'n��*;ln�c�65M���efӎ���8\-���'U�I���%���:�dp���L4:�; �S-����
��I>���?����$C4r� y{V+�9W`��1�������eKw}R[����^�	����I�>��1!F�WK�H��r���AB���7�R��柸������'�l8�~>�A�.� �T�x )	�-�,��i��˓�?�M>���?�����?y�f��:��@�F21�Τ`r��'8b�'R�S���5+�5����O�"�R7��� v�E-�܀c@��ƦE�I_�͟@�ɯs2ʵ�=9���*�<��@� �|��%�̦�����'�yA�j�~��?	��2���R&l�|ltc+T��"m���x"�'.B������|џ�<'ϑ�e�r<��̛f�8"e�i��It9܀)�4�?9��?	�'T��i�-�kL�JC��j�:%'��0�h�r�D�O���$�IKܧC�R��+����+��;B�lZ�X�pE�ܴ�?���?���l���Qy���.8�h�:���P�V�	�+�7�,o���(���X4���5.��cY�Y��D�$�KҸi�2�'0�Ǉaj����	��(��U��[!�=N�h�I"
͉9&�nZZ�ɐ$):�9L|����?���v�b3��.�\1�@�|.�d���imB�۝"�O��OZ�O�2�zlp#C�
�İ�W�Y4O�'9"]���I՟���tyBՏ9Q �b���#S8��玓3/𘑓k0���O��D7�į<��/s��"�F�Fc�٣�a֓?Q�9l��`�'���'��Q��a�����/ɒ7&��"�'�P5i��D�O���)�d�<�'�?�PSM�5�� �^=ީ �Y�c��I؟���П�'x}IQ�'�Tcbh��޵�<�(�Ċ&��qo�ӟ�'������'{�'kkx�1/� �Xp�e��%i't�mǟ�IKy�,�#5�:�����k�=+��Űì��Ps�
:�'9�Iǟ���V�s�� ����-V��I��0PIZ6m�<Qv�2-S�V��~�����p e�>�lUR��,h>�5*�aӠʓ�?����O��M{���;�rP�פ��	�B@������Q����Ο<��?%�����q�q��O�#���l
\&l4[�OZ���)�'G��5�vE�q�&�A� ����8�i���'��T4��)J�fL�GR�� ���b���N�O$��~���~"!�{ʕ�RC;YDcԈ^�MÛ'@4lh/O���O$�O���#(��K�&�7��D�`��2b�l�	Gyb�'d$e�t��*}�n��=��ۆN��Iv������Ij��?A�'� ��JV�9�"ʛ�%��)޴?����'L��'C�Q���q^&����L%i��5p�"_�8/,�zTJK���$�O ���O��?	(�N��4Ye���p��R=�馏��2�'{��'H�P�$PǏ���'f��5���I�/rA�p劋T���s��i�R�'��۟ȗO1B�~��hݎ�!�)M�@����c��A�I^y��'��A�^>����<�s�� N`J�@�$��M�$�X38R�����x��'q剽{��"<��/�K4��3AX`��ڸZ�Ulqy2�0x�7mYE���'C�i<?�l��~��`����.޾��b��Ʀ)�Iן8�	���٨�����i�TڳE�j�N,��%�">�(H��4rL�`�i��'�B�O�O�Ҟ'�n�H���}P<0W�&)A��m͟ ����d$���<)��/���dA��A�j��w%eζ�SR�i�"�'��O��}��O�I�OB��%ZЌx��b�56�r@�㈮��6��O^�O�����O��ɯudD%�V�>V��	���%7Mn�����<��X?�?)#J����9Pd��+�u˂mȣ'߉'�4��ON���O���<�rk[�f�@���ɥ2 X�o!�M���'��'&�'�iݵ��I�36v`R��*26�9Pdӈ�d#�d�O��?�R���d׮@M*-��EŝuSr��r����M���?����'7�IjI�6�F&9V݈�ί"�t�a�b�f���ԟ��	�4�'!T����<�	��X}�!N�3mN����b�*Ҁ�oZ�&������'���Tq��ԋd�*CC���m�����	byb� zB>�2���kL�$�*�t��~�m��iN%n�'3�Iҟ�Io�s���$~
J�锬ЏY&��à�v�b��?�Ѐӟ�?)��?���*O�n�*'�B��4��_�D�Gjڛ����'��ɀ-, #<%>���`�6#]`�C�hY>9 bl�E�w�̰�tD�̦��	ʟT���?���O@ʓ#�i��+�%-�@u��kJ; �L�e�iH��1�'��I��@����4R1���#����˔� M��:��i��'�G ]_듣��O���0,�\٘�-�'�:Aj�F��,�6��O����O0Q�0O�S���	̟8sMS���'�Jt<�9D�)�M��b�U)�^���'�b[���i��(4�]�+�:�ӥ����};S��>� �[�<�-O����O�$�<���:`�z(@�2p2�́;��ÑZ���'�R����������j�0��!����ի�i��D3C@m�ȕ'Zr�'��O3:����l>�[6mV�+aN����l�2�;�mӶ˓�?�-O���O0�$����۬S��i����FF�T��+տwP�H�'���'�"V��1�H-��I�O�ik�e�iՊe��ɛ/,̡c��Ѧ���uyr�'<2�'�l��O�iϼ@4�Yk)/L. ��ϵ�M���?Y.O|�	�E�b�4�'I��OU e�@V@\��cEʃN���� I�>	���?	��~ڌ����9O"�S�.zX�����K������\��; L��Ms��?���j U�֝8e�����
D}�C!ތC��7M�O��$Ð#|��O �$�O��>���H��@1��g��b9\��~�ʕ h٦��I̟��I�?�9�Or�Z*��r�A�3(GĬp�,ϻ��PX��i��S�'*RR�4����y���J/��m;ŊC;�f���i�'�b��vv�����O�I (�[4��AV�aS�i��=lH�	ϟd9w�x��'�?Q���?	@�[2q��#F� ���V�v�'Sb${DG�>�)Od��<����������B'�lC�m�g}B�R.��$�O����O����<�����0��_��5c%����+�^�ؖ'kb_���I럨��Lk`�0�m,'1*6Aŭu�J�ے l���I�8�	�t��[yr��$�擈ER�C�K�%ޔ%#�fZ.k�~6��<������Ov���O ��'R]3dcct���*��C����n�>����?	���d�9T8�(�O�rcմ?�Ei$�[��x�fZ_|"7M�O�˓�?����?�4���<qK������&��R�"|�ūgJk����O�˓gBܐ�\?1��������f�B�Q���'u���//l�aӮO��O|�$[;��|�������:��=sdl<`��M����M�*Otq�5�U�e�	ן8���?U�O�.�J�ā��j^�T�Uc�W���V�'���yR�'�"�'�q���`)��Q���)�>�jtyַii���Jj�|���O��$런D�'�	K�`<�En�ikŚ��:��@8�4N/������O)bO�"�����7{v]���N�6��O��D�O"\A&��U}U���Ii?9@�Є=S�dh#ɩP{�-9 EB�	��Uy�����yʟ���OD��ЄR�����# �C%�:���nڟ�땠����<9����$�Ok�^�]���zv+&At<�r�S�
��I���I֟P�I����	ߟ`�'��AY$c�)v���{f$�a,��{`OSE��듦���O���?i��?��JFLDXIVǆU�z��v�Dd����?A���?����?i.OaS��|2/P9*�E�G�,81ڌ�Ѕ���%�'�W� ���H�ɤ2���I�r-��g�G�l��tcH�L���
�4�?	���?�����I7P�O�B�]�5b�9æ �*�^a ��P8]:���'��I�����\y`nh���M�7nT��)x�+o�b�//�|6��O��$�<Y���%��O���O�rIi��7[u�l�䨑V8���G�%���Or�DU2fp���.���?9땈��X��|bE� ��0���d�˓��`A�ifL��?	�'jg�	 ��)i�	]�
y)�B	�\_�7�O��d��h�P��+�D;�S�&g2�+�P�oSԨ9E��k��7M�)I��nZ����	���ē�?�� ���'b� ��hRE�c�f����i,,|��'��'��.�$�$�� ���؝#z2���gڪ�F5lZ���	������'"��O�,jƛn1�V�C���[2�i��'�ސ`�d>���O���O��q��˃F��X�C��#�$�瀍��a�	��t(*H<����?�L>��:�������["�(Oʘ�'u���'�ҟD��ПH�'�����x",r���~H !uʂ�8�c���m��ߟ�ɀq*��E����6�	pDd������'RR�':T�0�cD��d�ܐ~4@	#�ÒPz�A�@l������OT�0���OV��ªmmX��H�4��3M�	z�\z��Z�B=�'$�'-Z����X:�ħ"´A���ɄG�����ۻVp,r��i��|��'�2�66�>ɗ��g�d!bcշ3���k�gYӦM�	矤�'��K!��'�?i��>D�8�ykJ� L�
u���C�xr�'��$۫�yr�|�֟y��GH4�=�b
�n����is��_(,D�ߴ`��Sڟ��S���d�%H��Dp�O�0�����3���'����O��>� �i�/s��*��S7|D1��m��,��Yݦ��Iߟl�	�?��K<ͧV�0�:�O�bV�����ʝb1�I�0S�X��Aya&ҧ�?�+��aj��ߝG�\��$�Ұ�&�'h��'>@���'�V>}�IO?A@D� 1�g�P&wUR!@���{���9H|���?1��uN�C�(°�����V�Z&v�3�i���pO��'�B�>�7� 9�Pw�٪R��!P���m}�
���'���'���'tL9gN|!����X�R!23cZ'M/8){�U����͟8�	S��͟<��3�(�w)W�ļ��f�J�N_�n�(��?����?�-O���EM�|2�e� 4sL�'�T���
h}"�';��|2�':rE�������\�@�S�_�	;��^���	⟴��ϟh�'ВX�5�+�	S���c�K�y�̓v���9�n�8%��I蟠a��'�I�od�0�qGڒT��aA蒄$$7��O����<RN�7FE�O���Ot�|���hfT����	�ɘ#,�d�On�$��A���'%|P���C�ThC��I	Hq��n�Oyb�ըl�L6��m���'.�D�$?S������.������������� ��?�S�"���Ԇ�W6�'��?Ln�x��X�4�?����?��'~��'�P�yD�����6��+��- 7�Q�K�"|�J,��F�)A�ʢ��.L�	��i�2�'Z.ӱa��O��$�Od�	�mlm���	/U	Z�`Dm�*b�H���%�Iҟ��ϟ��0�$U�2 ��?���H�"��0�'-P ��/�	ӟt%��0Į�AthK)�~�h�YN&��.��<!��?����~��ʷ�0s��0�u#�;bP�����a����$�	e��� �	<7ԥ"��O��ΑjB �
pL,t��	9�ڟ��䟠�'2.�P�z>����%���el��:�H��>���?qM>��?YR��]}� ։J��Ȅ���s��Ϻ���O��$�O���&�����D�R(2�D�r��1%6�!��7�z7m�ON�O6�D�ORl����+ n\S@�#E���G�S ��V�'5����,#t͕��,�I������?Ap�F�ޔ��b�>d���5��3�ē�?�+O����i�M�����ki�P#�(�!��­NC��^�ċ��2�M5T?��I�?�H�O�������t�R撹�6e�C�i0��'����F�%�u����9t�(�ٴ)w�ـ��i���'��O�O�D	�D�ZA���1����i�p�P�o�;*��#<E���'� ����'h��a�Y!��dpP+`�8�d�OX��!N��#�)�On�	sN\J7̒_�b���q�J-ˎ�d�V�����	ڟ�9�	љw����\H�91��M3��^n����O`�Ok̕�$B����&<��b�;���������Iky ��A�6R�0��)؜l"�Cp�=�$�O���>��O��	�k��@�����jmI���Q
c�H�I˟���^yrkM�Q��7u qS���:p�� k҉N�hB6��?���䓍?����r�':�²o� }���K��+l�s�O|���OZ�d�<��H��	*�O������|�8��Ω4NdX����� ���O�$�� �O��@�R4L.���#�8$� $�i4��'0�'I ���'�R�'#��O�Y�Q��3	����%&Q'DRA>��OL�+`�GxZw���j�B������/K��|�ڴ���Ym�Tn֟��Iٟx�S.���ư�ŀG�H����ϼ`��M�T�x��'�ў �OF�I�dZ�x����0<�	c��i�Z�ô�'>��'/�O��I^��ɬ:k����"B-��c���y*�'I��Ex���'X⹢�A�:�6���㈾��@��mӦ���Or�$�E>��D*�	�O��I5q���`�@�o$#��]�>�.���dZ�SΟ8��ܟ|j�L����ᰖLE S�ʉ����M�� ���S�x��'!��|Z� `9(��R�$Z���%��-�E^�!'6�	����ٟ,�'����1D]DԢтd���>5y�O���Od�D�OP�Of�d�O���0��Z,��w,؟8 ��Ѩ0A1O����O����O���G���$��sݒ	q�Hu|(6�ڳJ��PnZӟ�	؟'��IXy�h�Mc�W�w�朩�냼��!Äh�[}��'$B�'z��(P%r݋�����W8�bY�����K�1PV�ymZ̟T�IS��?�{�Bѝc��%c̈^�݋J��M[��?��?�4b������O�������c/m?���CA��`Sfu�@@a����Ȗ'��� ���&�C0J��C&�������xR�C
R�52
�PF�=����x����c����D��=A�e���ŌI4ҁ˖E3=��%���5,x� t��fE�A3#]�2a��AZk�!�G9)Έ�HR�;fqXqp�.4;�NL
@hD�L	茂U }�Z�Ұiơ
�~D+��-R)��&+"��J�jA�X1�lB�y22��w���-���\�t�~�K�8_�x`�fy��R��h�	�|�I��u��'��,^Up���/R���&e�Za����-"D#�V I7�����hOz��pk�a��� K��@�@��qo��@`ը̀<�*A%�X0+��퉃l�Ɯ��sYy�aN�by��I�<�4���OȢ=9+OVԫtkܭ\���ӄ,�kl��H�"O�lr�
X�"2���J*)�")�� Y���)�<ٕ&@+�F�v���*b�+gr𰣅
U}q"�'�"�'����'��:�P�F"m8y!�<9���#ٰa�s�Yw}�Q�p�=<O8Q�@�gN����T�̬���Y�#���Х_�]�
�F) <O����'�"�X��4�J�i�+NP�ў@F2�H�dz��n`{N�GU1�y�
' �5(�)X�+>��n͝�y�>�(O`hr�[˦e��̟|�O�p�Ԥ��Z�:U�qnΔk�:���!^�JA��'�b.K�x(]��T>��
k'^�+�"�Z�n1���*�)kdh:6�SP�R��״]$�fV!5\�<�AÅȟ�������I`�D�̺n����w�S,y&:D���E����s�d���l��u ��ݦa��4� � �O��$����»%+f|��m\7&M�@x%,`�`��'�M���?	-���!1�O��$�O��(W���V%��)��,'��`�NB��V���2��E��\ןʧ��?ɓn	�c5�U�5���A{n���F�<�T,�U�T�n5��0�a'F���'��Ayg��@��= �%��rY�53�)��w���'Y��H"|�I<P2��"i
�~�BE˂���c������X����L��}�#N[�?$<uCQ	����"<���)�D`Ҍ~<-Ig+F��u���7�?!�i2�4�q�O��?9���?����OT���7���ID�{.�p�/G�p;���v@�}�k+=��i1֪G;���ͯ�~��Ƭ��>!2��C92�����(�4T���ׇ�?	����?)���?�gy�T>�Ɉ+�wD�~�Z�q�م	.rC�ɲ
�����,[�nD�)��W"�P���?Ք'H�+��bӨ��6(�(Ҏ�V(;���O����O�d7hY����O��*��+/�"�ban��H�P�	��u~]��1!�F����[�_�������i�Ȭ"qʍ� �`�$E�E�-(�
,�BmX�ї:L�0#��I I�����O��!	�pS\R�
2x�2�	>�d�O��i*�)S-��Q`v��EV�CA�ՊA2!�D�4%�rQ�i͘5�9�����2 ��o}R�)�Ӕ+X�0Z���L2^C�����VB䉨	)� :���={�:�R�0�tB䉓k��A�G���t�rH�/[
`�C��*}����p��+24J��,ZLF�C�I�9�P�)@�DH���b�E�`.�B䉭AhbE�C��8*W��[J�B�I:0J�p&I��&�M0����BxB�I:o�-�%�8Z7��z���5_�\B��9U��|��A���K��^�n�C�	���	p��R`�P�ݍ=5�B�I��(����ر��%��f��B�	%\�ъB��(�d��d̝�k��B��"�e(�W[�u�3 �BB�Ɇ0��٫�@S�I����b�9�C�x�̠A0-�TA��ʫV~B�I${����6�ۦ
��9���Ǳ!RLB�I��]�с���}�v.�+��B�)� $�� ��j�t��u��,XH@��"OXM	$cױ1'�C�������"O��S1��r�V���e�0P����w"O�k��!�z\�bE�+�f�Q&"OD�sSB�3)����Pj�b��L�6"OF��v�*&;��$J^+Ӷɫ�"O����PQW��[��V
@�J�ٲ"O8�t �z�p���%!�\��"OF���S�a���w*�C�T�U"O*=�Є�.ml"D�2i� )����"O�L(bBmf�ZTƈx�z�)�"O֭c�A(w�����$7�`A��"O\\8�"ݼk�*�0��E�ԥ��"OQ�B�0{��(�U��W��s�"O�찖�Y=��jrm�&fG��;3"O� �D�G p�Ԓ���{bDx��"Oҙ��!Z0=@$x:��@�p�$@i�"OȨ�+�N�k3�=b,�b"Oι���Ӝ�� ��A�h6�@�"O�X�Х��A�,��OA�xNr��'"O4q9v/��BY#��D�pe:�"Ot�F�1�佢 ��=Z�4�b1"O i`�&�,!�Y�tm 7J|Au"O�)�ԡ������5��}���ps"O$A���1b}2�l��c��	r�"OZ%�D�]�t���C&�=7�i��"O��N�C�b���zٰ=J�"OH9c"]���q��-jШ�:�"O6(a�g�5)�xX�E���.�q�"O�3�b�qn� �0�E�4��T3u"OH���+ۗa��T�%���4M��"O����߷:Q��o�+��X8�"OFY�T%
8�xmO�}�f��"Oj�!ԠPFv`Y��(dq��Q"Oڑ��*W�0s��f���]�����"Oذ�'
��F�0����/(�Q�"OnL��k¨Q���ʲh�4q
�m@�"Oĳ�ş�:���نʁ),�:��"O0�� �IFFu��ʇ�y��BA"O�ĉ���73>��p�JܸJ�P�p"O�Lڣ�1��-r�
 Q{|!��"O��hQ^:c�BH�B	Ƈ���{5"Ol9#��S�+�j�V�X�~�l̹�"O�6͍6+c.Ԛ��N�9�d��2"O��3��HT ��� X�l5�R"OpAB��T�qb�%�Fe�*s���8"OB�qa�!=��հa��+��ģ%"Ol��Ϙ�+��X�5C8M���P�"OLD�4d]�2E�������t�z""OZE�F#��W�
k��E��"O�ّ�TK:�$��ɡk�j-)E"O�|A�BQ+S�𠸰hN���`C"OFx��ʎ�U���Ʀײ	e��C0"Of\S�O��h*�1)�f�8Gd��	d"O^i�GC�'���#��]!mIm�"OA�$��4I�\xǥ�'�BP�"O��3���<]SV��g/S�ƨ9 �'k�<@��'�q:�D/	RHp�1�Û6���'(ji����S{~���οK!�u�v�K81e�">	�Oҽ�h��!hR�&��-
��;p�\�J֕>�1�=A�CڂZB�j^�\cPf�b/\��%eQe��1���F�&1)���]���Eӟ�S�&�ͬ1N��1ӳ��&���f�D"'Rp�ȓ�ơ�6oP��� B�z>:�A�<��P�JA������	��B��� ��,Z��y�;x�upu��0.4��GG��4E��ŵC��n��}�*T�#�4\;�� �� �.	��훂 N�(d8 ��h: m2��DȜi��ŊF� zv�	?I���>I�Ҏ
<����*�r8sg��C?�T�=d��Q��˙K̜%	be_<kŞ�Bdl�O�����Q� vKC�ҏO�<��a(D� ��}�L��t$.�����z&�����U7t')���=3�	�a��9�uBu�2z������:�����U?�p�9D��.[4H�8"�,ϰf�P�` $d��}�h$U�D��HK ZNl���4�Q
����P��^���XpB�� ��y�M[�`�ܠ�,9���J0t�Ɏ>�b�#c �y:�%j4�|X#=��bW?;�̐�5�]h�4�Mjl���O�&Q�F�bdՎ6j�Q��$$le	P�j��>��0�DJ�V�'!N=GƝ�р"G Z�\ڨ!�0��x[2��tȡ�"��< Aʅ�u�*Ȅ�:�L�5RIф@§{�|��c��"�U[�)�4��~��Ȯ}Fe�`Đ\<��Cѫ�<y���mL�ZA���W�|1�cO�Y��'T=ɑ�wT��"I:n\����E�b�	�<���z��7Qվ@��lQ�63�cg��5����'�*���#+K��D��*ߠaj��R�y�R����ϺY���-&����XJB��p&@�*�����$>��iDAX�x���O꟤JQ�)r�%A#B
��˶�21Y6UH���d�H�N�4P�"��'2p�!ԇN!E"�D���^0C8`9�'��P *]�(�T7��C�p�#���K�[W��1jE�N6����L\�4X�d�qM?s)FU��k^)zF�$	�;��I\���e�{��S����[:���@	Xض��牁_*(�@�A|P���k�3\���CS�����-��I�a{b�?�$qąV�pO��Z��ĈA�m���X��hOBP��+�c���q�b�( ��"%75�h�&C�,�(PG��0#����&4�-Wd	��KC e��n�2�ޅ���I{�b�2{�@��8r�dd���##&��=kH �cgDV&Np�Hy�j�;7@��2N�	2�<�(�'[�9�J�!;��7-��g]d� i�g\R�1`O�B䑟��r�\D�:u�QA����$��jG��B@�B�^�d�:)ܢ
�����|�8�1 ��5$D1b��֞z�\l�Ӏ3lO������Ip
\�ѹ`*R,>g�
c�ע+��|�U�`j
��z,��c��쁘��Ӿ
j�iVD�/y�h����O>��{m5�6�J�:Ҥӧ��Z�~Z���jڿO��c�O� ~,N|k�C�'r���(���O�R<�a�G� >�N}i�K�2R�	� N���ѺJ�n-�$���B��L���bHG���B�	ЩY� 5XS�͏��es(Oޭ0ElO7c�Ԙ㠣E=�&L�B�'D�u1�D�N�Z�QmҴlDެ2�y�'LΌr���'Kx͒b��f�45PEc�8*X�@��.i6�Mb�EC#�FL�'�2O`d�6��f&�x���� Zt��CV/S��%����+[��)�b����'^�d��(iT*9`a֮�D���l����ē�J��.�^�37C\�.Q�L�Tm3�Ru���D7;�V%��M���"�fPHy"&S�h�&@�����):\�v*��F�Z7b��B�r$��t�xYG�c݊�%�@ ��,�a���A<��f�Y�c�n���)�>�T���#�ryr��8s@���túXbR�ȑ��']��Ң�R�����' ���PM��#OA p5J7ME�%.���P��z��J��W�8���_6���=3p�uA��7�>`�Ah�O��1�+|O�����_}��1/+ �s�hl�b���B��d �
џ1� ���xBZ��n���T*��#��cb�?9����N&� (U�Y�'�K2�X^�h������'���u�LΠ"�F���ہ\m\��J������c	�<Z�y���:\�x�g�!t�H����q��fa|��l��k�f�R��#�x�<Q��+c��y2�G.1Jfȸ�f�H̓D����̏�`d�� +;�u�O�9Z@�A_?I@���AO�y#��� �����N�<�	QҚ<!Dl�zw����n�J�$��3Dv��s/ɼ��<q�L**Bd�	��5K"lr�cm?&k_�w��Xؔi�Yx8B" u�'\Ɉ�Â;Q�@ɪ�f\"z�OL���o˰?�������1�D�i���hu�-�Ǡ
�~0JXX�D�[�R��4S���&(��ԛ�쎚$�P�#��/M��h�ŝ>��O�$�
�'6"\
Fk`�H�@͠k-P��teC�+2��=����5Y�X0X�T"D�\i�JEE�+��Ez#m}.8�S�A4W42O�|0���A?��Y�����y5EqA+�9k��a�D�U羍�#�è^�ҝ�C?6���Rq�˘x�8��1"�Ix�\�t'5�Υ+�o��x�yBn��(P�.\�y �����32c.l��� g�ۋ{ǚ;�z���G�6$"�BՋA��yr�$~��͒� �2&��m�C�(>�N`����eF�_��M���ޝW���g�Dݼk�O��pH��h�瀸X�=2co�\������=	��`���C�6�Xu�>'����:D��x0a��Q߉'<�h�D��i}bp�d$ʲM\ps$->gF�E}R'5MN��D�2C�"�3�d\�|BU�^9#�1rVg=��)�k�`}B���z�(��	Ĥ�x2MÛ7�<�k �3X���ɑmΜ�ga^9Q���� fډO��9�Q��?��#O 8w���ǄC�vކ8��'D����
�I�(��7���F�r�G	/����4�c���bC�ʦe��ʚK��O2��;R�^�H�%T/Zx��q�����+�i��:S
��������&�HO?i� �� 
��I�j=�2�ҵP��1�"OtH1TBV�� ��/Z%1�`"O�P���Q��X��'5W���[�"O��0��Y=�8�Q��![��m�d"O��� �<� 5���M�h�D��"OJt(fҽ2�нcD��(h"OTx b<ڵa�!�LT�"O�(# �r2��d
[.G9~�0"O��S�\ki�7Iu!����"OBDx$�N/�6�3��I+@�X�%"O4���CK���j'OM�3��):�"O [���..���cN�=�jq��"O���&ʪf �ś% �~���"ODM�S�
�4j
hc&�>C�h�"O���&�,D���fͮQ��+"O���$�$3� ��FR�Qꆔ�"O�PrJS�lpΰH c$՚h�"OQ���RO�&qw���{��� 3"O�9����1R�j�qV럠|���"O��⤂�h����G�݄!l"I�q"O<(�TB�P�܀�I�8s��1f"Orx�@j,L#^�S(�h��A"O�����,�~��g1b� �"O(l9�`�(A�	
��#[^�*�"O,�	�Kܔ~MH q%�5m�RF"O��E��r"�����Qj�U��"O
��0{>�����C�"M��"OdX��ȝA�$���F>�mIE"ON�(p�N��U+�'��Q&b�("O��(�hI�Ԯ�ca���6 L8'"O*@���~R��ED"f�R	1�"O� @��] ���0%�Q��"O�ʲj^�<<�#J����k@"O��k�A\�Q������G�:T(�"O�����6�*�
9�8ز1"OFu�#��'o� ��S`\�Y�!Zg"O���D���su�]?���H�2\��#�xF�tkn�"��!�ȓ3T*Lc�'��4cDC�<0<�=��%��`㒉� �	#���6j^�4��/7.��#O4��-b�E44�|�ȓ7�x9#��7?�����T�!�<��ȓVA������;?���+��\�D؇ȓlB��G�:2d�C�"�F���ȓ]��9;cH�� �9�qh�Ai2@��`�e[F9J��%�S�!�a�ȓ+�X���h	 ����gg��A��Ňȓcߞ�(�(H�~������
-U�0��B�p�C��� {���s
�����tǢ��C�H���ĳg�Q Ee�ȓ0n�Ը�l�~�*�cf�;#EȆȓqö����ߖ I`�֋��n#�Ć�l��EB%��9 #(T	w ߣT�����`:d��6�,q�,R�֎�ȓ�&Xҡ��R*U��R�BT�y����!3&��n��J�
~�L��ȓ p5QуK�O�D\�

��4��<�:< ���<^9��{d���S���ȓ-&�����
�SUMMS0~��4���
E�A4G�Fp{A��)l8i���.r�OR�!Tl��3@B��<�ȓV�,���]�a�ЬP��EJф�g�����B	�6�N]��-H)��~�,�`DD�A,�$�����d��S�? ��� �m'jA����<7�$���"O�D:B���dS�V�y�.��"O�z�M>C��<
reO�|���	"O��y ���YN������3��9��"Oɸ��؃w����LX�8b�Ӑ"O��ؤ��:z ���ȃ2�����"O*ey%d�Q[��"тy/ ��6"O���+�x����A��D��"O,�c����%�P�ϞQ,��0"OlY���l
�]ۗML�ThAK�"O�!�F��4i�eH�Q��`�"O�SP/��\L�fL٢�z)�"O�չ3�^�ޡ����T�ƙ�g"O"ق��_45� ���\(y��1p"O܄��$��u0b�A�h�3j�,�f"Of%t.P?[�%�%GN�88(0"O�Y*p�ƞo��fE�	�C"O�t�t�ۉVÂā6挽 �hh)c"OB"SE�o�d����.8�D@Rg"Ot�H�IB�h��8IN�(��"O�a+��G�"d�L���S:\J����"O�U�BE�1;�ܠ���	S�����"Oj�ZB�B�J���"#/B��jqZ�"O DЄ$���y�NF��|��"O�\H��ʋz#&�#.^U}F�0"Ob�yW@�02F�#��,pS`QZ�"O��X�l��x�d���L��|Qh�9�"O�isbhU�1��"�Q_|c"O�p`��RG����J�L\E�G"O�U����<�z���8 ��E"O4� �'B���pc�BaIw"O�H1w+��O
`���I���s"O4���葵8��r��:R�\��"O�ͱ�¦T�f�	��U=��ur�"O� ��*�8\7��0��9��@�`"Ov����=�<���I����4"Oؤ:%^�V����6NV�l��	��"O���g/F��`Cu�7;P �a�"O�,+c�Bo0bu:��;E�H0"O�A���s�n,��ݭg�򙘢"O�@J�딋>'��kg
T45~=�s"O6�gdA<j���i�hiY�"O��:����3�<��r	��4�n���"O
uK�c�
p)$sC&H�8z��v"OvЃ���dj��H��jZv�F"O�L胊�,�� w�H^$�"O|}���At����q�ڱ��bE�yB́�k]Fk�l�(<����i��ȓ#@&Y��v�Nؑ7�L�h�ڠ�ȓX����(D/w}�PZ�e��(�lq��O�z4��h^"tz�<�ƥ�^��|��LW���p@o����o��zv�$�ȓg��9J'sҘh�n��d�>��v�.Ԡ�.^�i���f�CD�t�ȓA����2��t�f9���A� 
9�ȓTpt$�U��1m��Wl��t���iy��c`E�YG�Y�i^�k_����8
��hR�0��fB�%�(��)�DJ�OO�C�,��/��,fr|�ȓj$]��ߒP)�L�XC��F��:\�흱=�z�H4bؙ!hC�	�y�#��K;>ZL���Vv�C�*R>���'̯I�<�1sk֢�\C�I_n�I�o �BT�7�ћbZC�)� ���Q.1�N`[���y��"O�=PA�{�t�i$&��8
��"O�5A�F�6B�ݲe惹b�p��"O�*%�x�b�0`��V��y2*�#{Dp ��1�:��ğ��yb�P8������i�)�(M+�yb*ٔj+,�85@�
s4(1�e �yB����й�d��Yu ��y��{��%���ʼkV�9�C�(D���/ԛ���F&�~��4��l0D��㪗��@��$� ����
e�/D�<�@@�'�̩҆�>A�d���,D���+��2L΂l4l94�&D��@V`M6n28��M�/w�A��#D��8�&H7t�
��݄ao̵���#D���㚬N@a)�?\:��d�'D��zw��=�{�A����� D��f�ȣq| p�����Ok���V=D��!g��,z t0&O����s@�9D�(r�o g4dl����X��4D���!��a����Vq�Q�c�0D��Rr �t��h"g/h�ĬB�/D��:�B�v�(�?p�*�"D��B0�4�t�u�m[v�k��5LOL㟼�0�Ʒ�8�w��-R:hs��4D��s�S�0��` }���# D�D	4o�1(^�}�"c�j��)P��>D�p���^<s�f,�)a�;�IK���r�4~���B� �L�2�aD�;D��Ѝəl�p�۵��B���"&$D�@����~wX:�D�R�x��?D��#��Ʉ3k�Uӄ��?:�V̻�e?D���+Һ����j.O� ��Qn��ą�ɭx�PWd�?	�:�� BLB�ɊI:Pd;a�?N�BX� �]�}B䉇O2��fH��:�����ŢQs֣?	��Ʉ�7[X��rN�i<��qq`C0w�!�,�Z&BPΰ�4I@�k$!�d��%4b}sg�2n�4K��,?�џ(E��).J%��QT�Z�z�b��cض�y�c�4r%��/�r*��9���yb"�
���i' R
iHx]H�Dȇ�y�+�.v�r���e_w�! �*Y4�yFǆ���:��ޓ�"���
M*�yB�A�B��Et���B}��Cq�Է�y�)_4��<[��D���I �
�y����d����$̟�P)$$��ƈ��yB'�+_��Tʅ)�6=�q�Ѧ��y"IN�v��sn�-V�qq�ܾ�y2EáY�t5�%J\2 4�i�_��y⩀�nNh����5��KS�T�y��� \`�J
ťv���G��y��M��6�Qs#�\v�[����y�Ɵ�'#bh���#Z��2��Σ�y���>�f�аC�"Yvx(��c��yrb<[-<<Q�Ƨ��i��dR&�y��k��� ��W�H  �Γ�y��_;.����p�_�A@X���ƌ,�y�O�p h�ik��0�s-K��yr&_�+�ŀ�`���cI��yrNЏ9@"��r#«\þ
����y⠛8[:���J�(Pټ��BH(�y�#ƾ	���Q!�� ���Ң���y%�d��!a�G+^v�zK
��y
� ��H �P?uÖc1D���5"O���5-պ1��*#X�q3��Y�"O�<c%@�j�@Ly���9��"O~�Af)�1�<Bȼ.hx�B"O��Z#ʓH���P��4�x�"O:�x��Y���XC�/l����"O�J�K��������t�b�x�"O�e�����#W�l�� \ {�����"O� ���<� �s����8���`�"OR������P���խs�����"Op���Ǆ9��Qbo�!��T��"Oj�B�� =f+�c��H%N�x���"O���re��#v@Y���&W���t"O*��q���,�8�n,D���ɡ"OT�u�>jP�EB���95�����"O�x�6(A�d��QA�a�8,��"O�"'k����� ��3��q�"O�ݹF�рT���S	+G���J!"OB�1��r��	:�H�u�R<�0"OD���m�3����r�H���"OTP�Q���9����(��E"O"�0���6�z@V�- b�=C�"O)au��i:(P�dI*�H:p"O�ӣ�ӲA�^谄�[���["O�`[W�V�C���w�
f�L�G"OL��� @�P�$�*RD��,FZ"O�QjvHB�7@bl�7#D�k@]��"O��T�H,/z${�AFs-�A�s"O����-Z�X�p�D
&r��T"O�Y����'=\����Ȗ}D ��"O�`���� ���I�"R�YI	�'ˤ̃@ IY�D��"��}
�'�W�ám�����_�Tp��'�r��%A��'Ӛ��,MM��z	�'��d�T���z�"g�(>$��Y	�'b\�/��F�X���O:6�ֵ	�'I`�R�+)&IұQ�E�1�$`��'��0b 9 F�X+ �ʖ0�tj�'�����ιe��T@��+�����' ,�H��rČ��.�F�'{��.�'Wy��1��)-���'RBD�3��33�F��E!��IA�t�'�č�ӊ��s��X��jCH"��'� 4��bqN��A)X�:����'6�1AL�Щq�Ѻ+�bH�'�0w��\�����Q(��\��'i@�Cdş.�HH�7�C�M��y��'ޚ�@�)U�Д�(tz�Lp�'O:r�*�9����lm�d�
�'��Q�7Ʌ[U��%�C6z�h�
�'iXU����ޅ�C,�F�J���'MV�x��OH��a��LA�8l�	�'��`	��Кu�� '�}�CF�y�e3,�i��t�C��yreU7?����*j(ÄV��yR+��u�E�o��r�����y�.SIIk�*S��$Y"g��y�JK�'���Ѣ���w���!�6�y��À|9��^5v� ��B�y��^(�pȐ���!�uE�<�y""�	
�X����7��E-���y�.@�m��� �n����C�'�y����P�Q�U3 �~����,�yrE�-V��pU�v�U� �-�y
� 0qb��/5���qMA83�Bݑ�"O����T�&����3=�0ѩ�"O�py�8Ov�}�/V#E�v�8""O��8eN�,v�<IZe!;2�@MY�"O8		�
�N�� gI��P�!"O6�� J�(�D�pd@$�,��"O���Fi��X/��s�)`�z$��"O���E�r![AD4����!"Of��S�W���H!c��Q�L]˳"O2���`� CX�"���4<yT�)�"OvI�`�G�9�����ǙC^U�a"O�*�fM/�=�6b�F�L0S�"O؄�`�\�O�����@"O�@1���E_�TҶ�̓D޾UQ�"ON��e蛐�*�Շ���p"O���\6L��˔�	�Bs�r"O2l򁣃!J�v�:�ieT�u�W"O�X��邡g�.p��n�>iQ�8��"O��(u
R0r���µ%����"O�T�I+b'э �ms�"O��B�*>�ۇ�����"O$�h���-0�Q	F����U"O��1%�>��R��60�*�B�"Oy��N�%9�tS�'ݫ~����"O�[��C)me.��p�ƲF����@"O4��5�Y�:~�`%�.<�1U"O��S�E.��=Q��<[�D\��"O�:3BIz̍	5�]b���:W"O�$�I��"b@=b��@�Z����U"OV�B0晭9MV��m�4gь<07"O�T9��ԂS<n�k��,��C5"O $��BZ+ŀ%��� {���'"O�%�ટ�#k"TC��9V~LY�"O +.K�J(� "&�`�0��"OT���&N�8ЦY��C�	�j��"O��y�JQ�F����V�6����"O���G =OPH��JENG"O|<�����A��c�GA� �"O�����6#�p�RI�"b���"One8�E�rCr���!J�rE��"Od�!'i�'輥P���4P�m:`"O��CK	�b��\�W��(9�X�"OV�R`�{֜�jR�F�37�ي1"O ��,�4bz�����"OVMX��^e�ɡ���7�ځ�"OBܠ`j�1v��Bt'܊trbM�'"O�hZ��`ʜE*u�!h<���"O:uS���j1P�A�tR��"OD�2Q+�g�0L�`�T��]i�"OLY!��3'�(4���\�j���"Oʥ9���(;jN �F?d��I�2"OD�8�.��|>(���*�&�s�"O��)��WB���C;>��EQ�"O *V��8/�F���d��-Q�"O&���.��@RD�P�h�"O����a��)�ΝȐC��R<x "O�`!.���X�	� �X4"O��#ᢜ�������v��,ۓ"O��itnVLz���&~B�d��"O�PZs왑
l�+�L}/lQ��"O���c%�y��h0('l��hR"Oҁ#��z7�}*aF����( "OԤ��$� J�4��g��4��A"O$RC�"R�떆�ony��"O� �����\�-3L�"���E[r(��"O�ݺg�o�Hm��fJ�Y�)D"O(\�cKԠa�pg�?SKF�!�"O2t�w[9�����V+��X"O�|��+AR"��u�(c�� �"Op��b�Z�F�V���OK,T�B�"OЙ���w�0��0!@�&L��P�"O�,���.D6� ���:d�t��c"O��@��mA���b@�9��!p"O�p� �C~ ��D��9�e"O�L����Dͺ]"�&
��k "O ���Y
5�|��>0���"Ol�;`oU�FbH�`�J'S�q[r"OP�9���R'�e��bA2a�H�"O}���#��=�Q![�e%�,�f"OX����*>�Hl�pO\�Mf��Ȅ"Oh r�	�5@yڕ@�<a֜��"O� �9"d8(f��p�*U	"OP
�쀣;�R�{� �.� ��"O$��q�=e�j�sb�L�t
D�"O؅����8�. �V �
w�5�g"Oļ���6yN4ኤ�
1�H�X&"O�X�/��M�VL9��Dy�,Ҧ"O�)��ku����'QM����U"O���ː<=#b8`@G@QA�P"Or(Ƨ���4`��D�!p� ��"O��8���>eu���ć���Q�"O�ܻ�L �<��bM�	Kt"O:X`S��q���U���2����"O҈�l��FBʠ�g�*c˘Pq�"O2�`@��8w��-P����*�4\z�"OP�V�P
n�$�b��"9��!"O�3��ukL$�&�B�^��"O��!0��;A��%,S ��8(b"O�D2u�ۘ��@R2+˜�.B�"O:��R��w� ,�U	�o�4��$"Ox����7%�(uڃ&����P"O0l�A-�>\��1�L�i����"OeH1�F 5�k�D�4���!�"O�X�r��_ �)��U����K�"O�ń�>���Si�= �ڄ�"Oz��ʇZ�`@�V�B�*��ESV"O�,8��EQ}��W�ߦB����6"O��FnRDɒ�E$�L�ض"O( ��%C����X���1"O���3+�\�ᴄߴf�й6"O*D �[}J� ���:ei��A "O�=��l\�%��	�׬[�c>�A"O�ՓG�
�%g(ty#�2}�d�"ONIdg�N,jT�A�
k���'0�'�b�����[� <�#�b�^����3��a������89��E룬�Ϯl�� -D�@�dD�
�. 2��7E��<��+D��K��*��8D䛄9snH�a�*D����&�I%DY �\�s'#D�q�"N���p��	�HH�O$D�(q�/^�Z���G�%+��$�R@(D��xeD
A@�b�ퟗe�x8��%�����l��l�8o�6���mC�[	�y�"OX�Q����)Z�/��{R =D"O�)�T,K {6e�!oE4/=���"O�0[��é9Nl3Ȓ49�hq"O����AV�sP�՚A��Ȅ��"O�lb/T�,�d����>�>��U�'�ў"~�� �U1�ӿK�n��#��"<n� �"O�a�t�1cj�ؑ�$�>9H�&"O��D�3�J����hr��"O��ځ�C�/.���[�	�����"Opѡ�J?<RTRc�`��(�"O,x��ğ�!�b�i�B�xn.]i�V�`'�����25�iS��8�L�WiH0}�d��5��q���,p� I�2��Wkz��&6D���ǝ!hO�U�U�<Glx��'5D��1�.�������ʫ^`b��e	3D�Lb�H�	�]��[6�6���=D�(j�kS�;��Q���{�V�i�b:D�ܘ%�ɑ[�A�2ʇ@���� .D� S�OL�H�xy'�Ks����#�,D��R(�C���A
Ǣz|)R&?��'�Oz�kG�]�+� ���l	<_w�(1""O�1����'G�$J��Q�b�%�b"Ob�KP̒�k������1�j�Q�"Ol$b�B4?�F�[��	n#�}��"O25KSg���"0���y���D"O�!ro�5�ƸҲʥQ�*�c��'�!��̱6pq{B%O<��H��g��'Tў�e~b�S!q�؈ #
�� 9��	��y�d��q��|�(
�Q*���y2��#5��آ揊���]�L'�y�Ǖ�p��-
soǤ>��2c�0�y�#Ǩ;������:}R���ҵ�y�ǘW(�9���6�>j�-	��y"��y᲍{RbR�8�t�I����y��è�f�AS��D�ޥc�%��y�G� �����cӦA�`�5�i�!�A %�|�@���(l����!�$Q�4|���3kH�qPz��\�U�!�=t¼��j��F�_Z1!���2�ృ�lE�Na@��p�4
!�DI��ބ���
 n�d�ݯ2!��ΏL����kj仇�]^!�t��o�EK�80��P�u����W"O���g�<���1�#ګs8$��"O&\�E�c���V+$H��"O�L��d�`�F��1 ���g"O���Ab� E*V� /re��i�Z�`G{��i���k�#4z�V};��K*��}"��ĺ$����Ȩ�
X��3-/D������+6
�D��x��+D��B��M2sI���%ҭ~2$�ņ+D�����Ӥ:WLȸ��� �*D��*�եs �AI�$T|��	ho)D�qӢ��*]���Q�W�(D�0�V��'<b������?���H��'D�4*�j:4����e�=h���xqn$D�k��8o��,9�'zר�r��=D���햵<�U��/��h�6D��31��X��M#F ��H�h�1ړ�0<�Յпr�>ݹ'�U"k�� ��jV�<�V�=1(�Y@'׃P��lp2��\�<	��E-��YDKM ����JNcy�'��qYc��+%
5�D�JP�����'�ep����(���mP�t�A
�'������4��r+OoYཡ�'��$����:nDʢ\�m�t�(�':��z2�D�y��(#L�P�<
�'�(%+�$�d�V���ނ|����'�ў�|�b�Ͼ-}>��%��r�� J�/O�<� ,�2FcK�z�b��w`��\\���"OF�Q��N)��l��\�(!|�""OI����_gɱ@n΅K�F�k�"OD���e�@<zE��l�;z�d0���'#�[(>P�)�r�߫=��ܙ�iE"8��O���ҝ�dT�E��!����G
�e�!�dS�)�.�qee^yh9ʡ�̲n��	A��(�R#�)b<
	���-\����Q! D�$�T�W7�~l��(�5��A�>D�(S�E�6v#t@ �bL�?�a�+"D���$�+O{��pC�,�"Yk!� D�l
v�@�E��ԃ0�H�)i��Z6k8ړ�0<���ۋ��m�B���"��n�]���O�~�8gI	I�j��'�mv
ar
�'��E�ŉ9fy���A
ļ7vf�	�'�<��N__>��;�� �~}2h��'��= �H�!7��h�u/?z�*�
�'|H�0�.�BVyV��j����'AD��-V1O��4�0�S{�J1ˊ2�'x<��%\��d� `C�"Z#6 ��'s abщ˙Z��5��c�j���'(0D�'@!@t�-F�.�q�'0	R�џ � 8T�Vo�e+�'��ly�"'f {㭍&=���K�'��!���nt~��QH�0�\`�'J��ڲ���$E��OF �"O���DЛ*�C���A!�Y���',�|cZ�e�z� �"$*(<��E,D��C�EB�8x��LP�C�MB��+D� ���>&O������5g��uA�)D���dHʀ`��A��əaI��7�$D���u�WP��#[7���Ĭ!D��
�L^_.J���&^4�V�)ړ�0<�pJřF�hy[��C�iĶ��&�HS�<A����C�zP�E �j��E�Հ�U�<a�FU���I��V�Aځ�Z>bB�	3H�v�W��gi�Q���i,B�ɫSH��1�Q maŢ��@�B�I�	�Q�YT�В��c���D>�S�O�T��p9��)��M�:0��r"O�$� .�(As���k��n'�TC�'�ў��D�'}F�A]uk�������BEZ�'[�]83�o;⡈��ʃu|�9��'��Ti#�$x�I�#M��:Ȓ"�'����.�����-�!`�4&�E�<�t)\z�(�׎	4�mH�@�g�'�axOS*!Bژc�!�67 ����V�y!�6'/h#�N/�|蒤����y�L��k�j Y��R�(f��2��A�Py�@֚	FBP�g�.�~I�P�`�<��Ɔ,M���X+A=m���`"T������>9�6e!�+^�y/84{��&D���#+�[�6U2QjP\G�,��a�<���z�PaF�<�����N�?;v0��	���с[1�~9y��B�:`]G{B�'ў�_�e��Q1��h2��bi�Y�<Q��T:�MɑE�w�0�����W�<��iZ�AVġ*���Z�<���>�p<2�F+Jr��T��k�<��!U?U\@@c,�&dƲy�Fk�\�'�?]��l	�6�p퐬��hzo?D�H�UgIH`zx�6��7�\i�`N?�OJ�5v� ���E�H|����C�	�cg�CC`ӎP��=����p@�C�)� ⨲'Ɖ�C��Xq��L*8�}��"O����<M[��. �hQ"O�-{�Ø*5�Jd0�)L'3H�I�"O@�0��n�P�Q�<~�ȣt"O���ψ3(zȴ�F6jB�'^1O��7ʛ�|��Q������,ZQ�'�ў"~�n��q�Z8��߄���0�K��yB�H�nUxy�|�Pk�$@�y�JX'TDI ���73jHSRb���y��8X�@��ԁ�5;��C��ڞ�yRh3v ��b�J�&�t}����yRʐ�^}Ρ:Q��,!ɦ�{�4��>��O@(k�1i�Xk��y4�i�q"O8����LJ ���e��`B؝�C"Or�0���A0�<��+U0�Z�"O�s!*ˎT!�d�Q⚮Z�%#�"Oh$z�c��mB�aR�W�����Z>YH�(E�g��HԂE����!(D�$��m��2\Q'"XFxh#��%D� �w����r�)�#��}m��J)D����B$Ea�]��&��	��%�1 ;D�H����Y��"�.T�$���a�7D�0I���9�z�ر�8fR� B(4D�P1LV�6���Gd�&�"�X��1D� ��)DjX��E¾W����g1�� �O�(S/X�,��q��n?hl����OBP���9����*��v���$�3D���3�U�~K�,�f�~�>@��H0D��hVD�;i�Z�i��/�f}�a�!D� ��K�m:�L�R�{#�,D����4�Y�t�W�-C�=�r�>�������R�}�B(�5�@�7F0r�l��/�!�$V7
�b��H;Ȉ
�͊� u!��4]�� ׌)x�J!����1�!�X,v�L%��o��)��^
f�!�$�#��$#_Fy���(�7\�!�d^DD�a� i`�����"F!�$�L�L%˔��*mc�YF�L�<!�$�|��`*�cMPDZT�� 2.!�V=GЬQ�B+O=$��U�v	S0" !�$ڼ,��P��
!	㢙��O4V�!���5���2�
p*:��/G�!�dW�l��I��۟'r�Cԣ�4}!�]�gZ98��V^h��
!#� Zc!��.eg��2��Ӕ[Pi�q�B�oR!�$�"�1�g��(,>�I)W�хL�!���5A�L����\�(�eb����sK!�d�9`Dd�##ț�U	90@�M6!�dH�q��3 O
�AA�	@!�U>�h�p�M�=$!3���'!�D_�p2���4�� �U"Dl_�X>!�d@:�dCPdG�{F\q5�Y=8�O��=����qu'V�h�Nc�"�T�}�s"O<ܲ��3�&�8fℋ|�����"OhdY�AT�gW��x �Տm�E"O Q�ACڞx �؃�՘BJ 2�"OX@sQ��$aa���Ԫߔ'	�}G"ONt� ��
#TĘ�&����y�W"O�͠���0$h����6t�"O䌹��vo~p�Rb�u�q"O��@ ƚ	+��l;t R�$�0��"O�U�'�!I���OY�V4F]˲"Oh|i#�Jn���`ь 2{"O�0��m�D�Ƒ��n�u	
��"O� �4{d�����Cd��qX�A�#"OR'��i�X�d��Lpe�`"O�%�$��p��D8v��:��͈�"O���pAU��Zt�2�׬D�H![�"O�,���FXP����Z'�L}C4"O�PCRJ�u�Y`���X9r"O:F�(u@H�PiE{Z�Yt"O�p"��94���e��+m��F"O<�*0�ݕe�(�c�>U��
�"O�� �Kw5���#A�]T�%YD"O��SW���� �a��_�,��R"O�q�*�5@~��;��چa�m0"O���1�=f���e�ĝn�&�r4"O����<Y�PqP�+=w�t(G"O���w)KZ�3�+6"��"O�Tʵ	
e�"��Wd�!���A"O��V)��oi>X÷�Z�M���"O4AQgf/��}��,D�k�	�_�<!!�*Ybr���M����W�B^�<)�����w+H�����F�@�<�6	RWEXm � 9��)�R�<i�)�eL[@��h�q`R�Oz�<�2a�$}a��;��B�t;�̘�(�ny�)�'u��Q3J�*Y&S�k
J&�u�ȓs�|��'MF*SB:���V!gL��'�~��w��G�@�4	X9{� ��c��H饁T+�4�)udď	�$�ȓX���
·+oZ0׏ՉQ��ȓR�h���L�F�#��B�R�l݄�#���Q��.KЖ���Dp\8@��jRX�Bg����D[֋��F�V���.^<!p'T5So���HD=C�R��4
��'?&L�q�A&�y>��ȓVE��������eΣr�l��&"O�|"a�¢F�[wE �8�SB"O$�Ci��xhj�cϜj;B�0"Odq��i_.P���ja�@,Z�[d"O�S!��$m'� z�.
|�t(�"Oh���S�1�G=}�|"�"O��p�&��vPU97�H?8=$�:�"O�ࣦ��Q®�a�O:j��%a�"O�ف��^P�X�E�7jZ�P"O�X`�oE�O}8����Oo�Eb�"O ��� 	<^lq���_,*n���"OzX�6-�|,��cj@�N�`��"O>m�2.�Z2����ޛ0��aA"O�s�⏯Q��L��f�\��"O"���P��lQR�]�Ė�{`"OH�'�8�|��2Ǒ�G����"O�hz��UM��E���14D9�'"O�m��
�$d3�(i�+P$� �Ӡ�'�1O��w��4K�%1��N�e7Xq�D"OH-[�!G�Xq�Q�U��!J'���"Or�Z��O h�q�LO� ���Q�"O8�E�P
z-uX��̠%H�<ˢ"O@Ԣ��J��PJ0F:P���"OH0�"M{�X1�",�5V��!"O��!���Qf�Y�KS>Ov�SE"O�Ś6CW��(� �?8,śt"OR0�`� �f[�� �n�g#�5�G"O�Y��4HyL0�.�h{���"OZ��������a�K�jt
!�a"O�	���j���î�|Y6���"O��)�J��D<!/i8b�!����y
� �)��M_]pw.��"���Hv"O��ӓ�3`�~�q0�=�Q��"O�a!�HW32ښm�e,bybm�"O�"�*��%�a����\k��q"O| ȴ�őhm�CDK�PPC"O�EZ`��OM�Mi�b]2:8�"OPMK��3a�`��F�$)N:$��"O
�p�9Iئ�3�D�yb��`"O��0�h����s�Ɍ�T��at"O|�0o�1-�R,r�jP9!P���"O�}A�`�"-ɈDhc�ϒ>R��E"O�TP�<Y�<PDcK�3�����"O��cF�̲s�	� ��0�@""O���s�3q��]� ���P��u�"O�{RO/w���*@ K���K�"O�{a��*]$��"�n�(�jI[�d3LO@q�f_9L�Ц�-j�D;�"O�P��E�VSr�֚B@9"O��ӎ��#fyh2,̞*���"O�D�v)��v�����)2L�3�"Ob	�r�1 �aJ�	�	4,��Е"O��5H �85����ۑ=>�#C"OR���8z�eK��If� �	T"O��Ԁ��JF���܍.]�I[V"O
��iX �:#��7T6��ɰ"O�	�v�͟S+zE�߾P�I86"O09�r*�-�
X�g��0f�H!�"O�q�����C��thqAP:|R�X��"O���$��킣m-[5d���"O>�p���1qB�:Q��:Q'���"O����ċXPDK��D�g�$�� "O�8ɧ �$ ���m�>=^h)`"O����V�Jq*'?b�R"OJ��'兯C0v�;��+1����!"O�����ȑ5�X�k!��*�ę�e"Or����!i���h�N[ƌ��"Or&��))$|��th�!+N���"O�IbC�A+5����UB�Q3v��V"O�dzQmT;;��)+�g	 �!�G"O�q�q�p���E��FZ��R"O�(Q fA>�Fl9�d��.��p��"O��P- �\��*�G���1f"O���EŵM�nb�����O:���ApL����H��i�j�]T!�Z"g���J��H:@
"$�a����!�+Ϥ���(��RhEa��>�!�$�Dʰ8�յy+Є>E�0*�'�2�ؓ�Ӓt;`�Q B�GF
���'��HWGW�O�$q7(E�C8"��'�����@� L��c��@��̺�'��-�E���9�l�+/iBU:�'��RMP'�.Ӳǉ>&��l��'�6�`�#�i��=cg��U9�Z�'�0�vo8�ؕ��5���'A�QnG)^̅�E%D�����
�';������ s�5����1C�'{jp�B,A�2�r�䗘��a��'�z�X���,Y-���Ɠv��M��'��<
F��m@
l��̄��	�'�� ¨�:%�ɚ�F�QF���'S���K�n�%
�"��M^TI�'b"�3է�6�> ���\�I{h���'L�9��Z-��P��O0v���'@�+��j�$YgޱH�@P��� n��2aܗvӊ<�bc_?�p�%"O&q� E�0�d���J,L��	��"O�Zf+7�>1�o�KK,+$"O�i(e�X�oO��[�-�L��<{�"O� T`�(��%��̴+�|��6"O���s皪z��'�U�p4�"Ot�I`+� i��z0E�S��hЄ�z>�u��{��ʡ��!;�x��#�O���O����˵E7$DhcCY%x]�!�RZt!�䇾�A��A�w ���DC!�Đ$t��Y�.
� 
1C@!�SrTTݢ��&�½8��H]6!�#t�BƩ~���r`͵����ȓb�@��B�A�P*���IҳG��)�ȓ��)��o���N���
�\X�Ib<�v�V!5���� �2+_:4��h�p�<��m4r%Ɓx�B�l�����X�<I�j�!I�����
K(z$ ����K�<�R��,`�A!��(8��bZN�<PM΍
kV@� ����\�J��@I�<���M+�Uz�"�e�p�p�b@Kx���'EN�1���.R�FD�$ d��[��?		�S�����k�([��{W�+ �� ��x<���25�CC��v�T�ȓk��1��>�d�9�@��1D�L�ȓy�lX �-V�'��u� ��<0�*��ȓ$⠼E�[��ࢆ._�<ߖ��b�z��=%�(qB��;s�hi'�0�'��>��~~V�Q��1"�lqb��8��B䉣�t,w���H@��M��lC�I_y�ɓ�_���%���F�I�NB�I�
�J��A�:!]�}� �^
��C�I�jѺt��|���1��q�B䉲Q'�8#��߽H�ȀK7��6%RB�ɂ6*lIFgV<Xz����L�C6(B�	LK8���%�+*"���wdB�	�N]�d�T|ޜ;E��.-�*B�I�v��nY|��$���$��C�ɭ2Z�
#̋9XB"y�QJ�,�B�	&R��Ӧ��HY�,r	�B䉧s*乴�F3hǮ��s�[ vC䉸u�IeLǠmz´�W�[�m7B�I#p@��c���
lS� E�)g�`��ȓ	T�+�cV�Q�����D$
gpD��V�D5Xg�Y(/���c�R�����R���{q`�5�u闀E�]c$�ȓx��Y �',(yt9	#��n�4�ȓ5F�5)fb�<ֈp��jY*���[x�-�r[�p8L���Gŗ�T��ȓ:Ơ����=%�0�3`_(U���	p<�r���[�n��6�:1����Z�<�d"��%����B�J=~���J�k�T�<aٞe�H1��5Q��qІSv�<��i���s��X�pTFą|�<�G�2K� �9��7C9
��cAJw�<)�G�Ych�pN�2]-P)�`��Y�<y�	=?`!ʲ�6ӆ,��(�ן���W����� �T���ȣ8pb�����u���� -�srg@!R�.M�ȓC�lh�NN-Ll���u�D��ȓb �)c���"����#ER�mV�ȓ_L(��7�T�x��h�^�ZȦ]�ȓQb&����B��v S�1�L���)���r��U�f���AC��`-��	ҟ��	�<� ���E&\�� :��̱V)Mi�"O"�j�m�=��O��[	B��&"O�eʶ�M.+PL�B卄!��
P"O�5�#�$���T��jU&� �"O�H�BS�2���b/C�EP�< �"O��f�Ã4V������%X$1�"Ol(b��X��*6�\'-R��'��	�<	�(�=����HV�Aeʱr��v�<a��ˡ �Ƥb��
*x�`�hq�<��lO�~�V�:�"��?�bX��d�j�<���]�L�C F��)�8��ǅ�l�<a$�P�A�٢�3��<x��Vf�<q�e�2Ux+w�Ҹ*�򁳐i_�<�q��n�6`��5��H�� U��d�I�ϓ6�F�(�DO @�r�nKK�9�ȓW�*U9�AǛe�"U����YX���F��PA���Ѐ��o� .tV-��!6���c�@����#I�L�~���bSd�Q��9_pH(U���x⁆ȓX1DRP�N�<�%��n$|���|���k�55��ӧ�B�T�jx��s�,�Cfꂟr�r����I>;���ȓ?PIaSL�T��-��HK[L���@����������i��E�ȓj=�����X� Śȫ��D������S�ۓ@��X2�@"Pq>���o@�]xV��8m6E���� \��@�ȓ����̇{ �L!�E´��ȓ#��C�A�)@����2�<��J���,�;aU�	@��8��q��!��p�(��\�|�����7R �lE{b�'=��*�A	Ǧ<sӪ�u��;�'�:<`��f���i�"�p�C
�'����⎓>r:��SL��r�ͣ	�'�$t��)���j�@�� �kX��Q�'�X4�<FxF���`C�j�x���BT�dD�������T��5�`�8v���hOZ��D�%��(u���p �"�8=��Oj�3O�Y�#9Ѵt�.�	6zU@�"O���6k!Ʊ�2�U
"�j�"O��R�F�[�&���B؉d��"O8��`��3�����&P"^\�\Q�"O.EJ�X5~�d�3%啜D&��A"Or(@�"6`0XR�� ��"�In��S2Ώ�.\���F(`l��5D�3�aNW:�dZ�R�#5D��yD�S�/�X�n�<�HE!��2D���Mk�v��a16YB�l1D�xB�" ��i!�b�.}lI�Ɗ0D��@�m�9V�$hc!��}`A��,D�������
��6Ԍ5�<��+ D��ɗ�T�J���ҥ��"7�ftqǀ D�0�э��izm�e�O�o��l:�J2D����O?���D��s��l�ā0D������|49�fV*R�^�{Ej+D��e��1&y���Œ�"�`�*D��C$�]T�E�#�[�a�����+D���En�>
�(�Z�Ԍ<Ϟ8�'�<D��R�&W$iJMb��^P&�0�V�6D�ț1��:a�H���j[�nt��5D�Ps�Pv�c(�1U��&�lB�	>T�dY�0`��h8�tAwB�C�ɸx ,�`2a֎&�jػ�o�>E�C�ɝS`peⒸ��� ��XD�C�)� ���RBC^��1�&��K�:K0"O~��"�ShpF�9 �Ly��"O�UA��[�CY�]�k�S�*-"�"O�a�H�1)�����5,�n1a�"O4�0��6Nn1a���Ru�	�S"Oڐ:�CLWF\�ꡈC�"t�( "O~X��� y�"�q'Դ!O�!R�"O  �cI�.6��ؠE��a5Z�0�"Oй�$�9H�P�&%U�]ȩ
"O���/X�`-�q21D
��q�"O���� �{� �D�J�y� ٸT"O>����}c�|s�͓/�J�"OTrP��MJ�ձӫ�8~7*@!1"O�h���	r�z��3�C�,���"O>=2��^*&A��k�9'�Lz"OD�3�lU�K\n��`
3'����"O$ܠU`�$?E8XBe)ܳ=>\aB"O(!r�U�{��s���;0����"O�+�j�ip�t�g�M�$t �E"O�P�$/�"���4��.�A-!�$�/�6�X�)ڥT�
�C�/�|!���X����6���>ӘL�FM5!�$��0�4өD���|%!��U2a��ȉ5Gܑ��T�b(VH!�DU>���E��=�Й�G׫e�!򄞜_ݺ!HK( �̹�'�]/!�d�sذ�!���*�Ȩ��
�S!������\R�g\�E�hhY�'m1���G��)�ˎ#kvt�	�'���S�N) �ly���_0.`0�'�:�Λ�u:����߮ehz<h�'���rE� "^�!G�HZ��<B�'s\���-U�T�G�E�Nj�3�'i�p��DuPV�̊}���
�'��7�ӏ:�
��V�Gq�L���'���Kҕ6��(F40`1B�'�i;POA-%��{��ɉ��̀�'d�d��
W
���/��tr�'-�M���hwbH��܃
�n�9�'F��I�e�@������'F��`�Z�'�`d���S�{�H���'�~�I0O�l��a;ƃ,y+h���'���SM��$��&_��}J�'��J)S�xR%�ė �P�x�2�'j��3�*	o�p�@�υDaҌ��'>�M�B��="�p����H)"����'��	q�ʔ�He`�7	Xo�XX�'�.t�u�_s�]+�J�Q����	�'}zmS5BC#[& �C�H7�,`	�'K6��K��g���b��B*���'�|HZ�@�@ܙ�qCY�f4�F"OA8��ۿDg*9�'���eP����"OX�y7g�a�pT� ,
B<�a�2"O�2J � ����3MG�%kf"O��1���6x��X��jS=%7T��$"O<����0{Hx&j�)px�v"O�Q� ��L挀���h"�""OF�ۓ�I KI,�3�W�l`xR#"OR}T
�O��l����Ou��1s"O�y#i]�_x��9��	91�)!�"Oܴ���
4C\<�w�A�x�v$�q"O,�{0��P\��;�n�5i^�f"O@G/��.P���B�0��QC�"O����`��7�h]��G&x���"O� �@S�y��5p��L|��%��"O>u:������h3"S�:�2m�S"O�<���PL�B5�c) �;t"O:e���!��R`@� @v���"O�P6K��t�|�{3"<�G"O��s6��f�L@M�10���"O� � �d�Ѣ3�3�JbO,xCb�%�d�)�B�+'Zn�"�m2D�L�1'�J9a��Q/J�TX�`.D���ר��W䖕�R�R�����b*D���"'ȝ92芴D�f��C�&D� �#GT%/�@�3��(���
WE&D�x�6B7EmxE�1��Jv���Cd7D�l�&'Y�s�`����}%���5�"D� g���(&���S�tP�J?D�D:�.�y�������$(��	+D��m*@Ҋ�ؖ�E�
Yi��,D�x鴣�q��9`ǃ�hd�йb*D���IN: ��"��>>����.,D�����o�$�祜�D 8+W�(D��xS$V�F���'��N��}rso&D���E/�V?�}�u�
7=	Xcm*D����MCu\�"啺;$���j)D��3&�ǎf�0���a�en��G�;D���r.901~��� G)sV!J�c$D�hq�%VK|���o�a�D��#D���5=h��X�R�I����$D��8w��C��dV'&k����Q�-D��0�'�^պ}�F���<'ޝ` ,+D�܁�ڴ]��*Q��0gr��X�,(D�F�U0N,B7	��QH4 �&D�H1D-��S]�h�2� Y�2�2pL$D�\Q2@,)��X�R�[�.����	!D��iΚ�Z�vL��CY�zZ�Y�s�)D��A���&u��B蕆i���S�+D� �`܏}����sʒ�V��!a�)D�8�d�AF}�9�+�G��h�E2D���GS>%�e�R�'Y ��$	4D�0�Uh��q� ��6�Cf9$�$f1D�`����7m�M���n��4�b�0D��U�U�|pY�V�H���q�0D�H�� �/$k\��W�=���f"*D��(�U�d��lzã���Z�f(D�lY��	B'PH� M�-x\tq@`9D�|k�\6Dr�ᱢ�FL9#B6D�l@�-��Ȑ�K��ʗ0҄i��4D�0s�� �u�C1]��D�v� D��+"JϪn�H=��H�g����&<D��qaHl�Ԣ#oĶ*�J�Z�/D�l�
K�����g��O�X\��+D���'Z/(��!�L���~d9�)D�d���Y�yV�a-e�|�[�*O�\�@(5�"-�f.7���W"O��� &Q��m	�k'>��"O^lA5�
I�zdqVE��=n�p"O�ūR�̬B9n-�W�=[д��"OX�Z#�Ίlh"i�di�7!���F"OX'�ݵc�����i��Hs�"O� ��nT5O�Z��a���Kr"O���B�ԧYH�i��f���p"OZ��Т�-Z�>����]-�xX�"O
����5�B�Z�G T��k`"O� ���>���1G_�'���S`"O�LЖH�;g����u& ����"O� �p��Ҏ)z-��oԡ� "O
���iJ�d����X8$�v�"O�S�J�'����@�"�.Q��"Or�B�`ۿ)�J�V`�(�8U"O���F�-v��|pv$ܲ���8�"O~����Ń���F�Ǉ�L�2�"O^%�+J1@���t$�=���2�"Oz0��>I���IG߁.��Y��"O�ec�e�
'�E�� ��|����"O~aa���B����eK�4�p�1F"O�@���,;��p�wd��8��X��"O x�7��.�.��Q���9�bՠ�"O�Ad�
cغm����2��xA"O�-y3HR���E�K51��$c�"O|�2ӎ�p�:� ��:w؈��"O��i�m°?Jα�a`�;�����"O�e	�	�&T�vΒ�z� �b"O�r��6*S�����V�)����"O��#�V�}#QC"F����"O|�,N_ި�SB	hB���"O���%��b��H��'ΊW����"OLQ�A�_�y�0Ȑ��?@J���"O�Q��-@Rv�����
<Nx�T"O>m���Òi^Z)�c�	v���F"O永&�X�"�B�	�1M�@<��"O�u˕�ʕv������А)��U�5"OF��L
EX©�[<R��m�"O:�pS�ؑn��"�LմQ�();v"O��R�F[g��cѭ�.i�F"Ox��1�� ,PZ�)��)c��� �"O�T�Ît�C@� �D52"Ob��� Üv�Q�e
�N���W"O���`��=<�P�g�W�VuZ50�"O�PZU���E>>袴/-jHarD"O���!��A`�U�68d6L�"O���bO�z{谧��u�L}�F"O�-�3䄆e���T�h�,�kf"O�l#�n���Xx�K'td�kw"O�k�Е4y��AD:x\|	`"O��P�F��� c֊TE��Zr"O���c���]�F
�c��yr�"Oh��a:���ӱ%��-����e"O��[U�"/.ڜ��#�w�P�K3"O9�Gl��G�N ��!M�b����"OҐ�d�˛RSD���I6����"O���C��<J�U�Jޣ`�!@"O �F��n��ɉ1\���e"O�A��k��&h|�� -K�\~���"OX<
ݙ#D��+ë
���x�"O�}�bO��]�`3��8��(R�"Ol��K�[��e@n� C��-�V"O�X���F�����H\�i*�"O��B�'e�Tف�+�D��%"O�	�d��^'�	�W�Qm�FB�"O�
^5d�����o�ne�B"O���p��}�&cbi����#b"O��Ӕ�:8n�(�&M��@چ"O����ûaU��K�JEit"O|X�횸*��%�V�B�`�p"OȘ�d�Ȅ1�4A�c#*pAt���"O2��S����a��؍J\d1r�"O����o���y�1�Ҟ,L0y�"O�0*�j�0N��:&P�R<�܉"O� �`[�~]�YɖL�VΙ��"O� h�X��yJ�������7"OX@.��1l8���I.��}��"OR�1����Es�HH�5�P�� "O<IQ��##�8�`A���^��s"Ov̘0(�?w��1�؁��4�A"O|�irŒ�=#7蕻3�I�@"O(4�b$�i��DI$��~��Q3�"OD� nZ�-�p�Z"%�F;�D{�"O@� �$��b�S"&q&"O���ù#�
@j�"
g����'�i3�&}z���)��M@�	P�',� `����&�P�nC(���'��� �ӌ�*���O9q(=��'4'&�$q2��T�!8���'��4��ސa�H���6�TT��')��+ҫ�VZ�����50YP
�'ŸAR�*[�wfԡB�ߴ�����y"*ʬ ���ׁոA��yb���yҬO�L���ka�L�O.̣r��"�yr
	_D��o�'?����bB��y�+:;�rH9�E�7a��Ж�X;�y��z{���X�`'0܂A�L��y2�\"��0�"��R�~��`)�#�y҉���\�R	�9X3�BU�Ҥ�y�M̕L���N۪P�����N@=�y��
`�EB	�F�����ų�y�"�;���Ң�,���ā6�y�
��d�x"��'r�(N��y҅��\����ḇ�J��&�P��y��]�{��0���g�8�em �yri�d�abF��x��0+�D�/�y"�T�h�xh��	m�R�� '�y�ʅB��D�����]呒�y�*C�=�j 9��9#��Hpm�=�yb-��(Fb��@��66�=
D���yR)�%�#��«y��%)���y�#G�q�2z�kǗ?�tT#C��1�y��^�:SP\
�I�9q@ԫ�ʃ�y�I�* tX��O*_�L���V;�y��ޕXB~�ꦎ�_�I�6&R�y�`ǣWR>�� � ��X�K#�ybʞ��Bi�Qj߂}ц��yR׸c�"���]H�ӧ:�y"��.�Djw�H�J�Dx3д��y�J��i1�AڭD\^�a����%�S�OϪ�9u�ߺo�2����
<Y410�'�|�d� !K�8J�1�� �'Y�����iD P��d[�H�
�'���IHU����*�lK�#��	�'y�9��K��0E�,�d����h��	�'��axv�\�bx�R5$T�	�m��'��������]�}4�b�'�d��e���pX	F�@��'~t"�AE����Pύ90f�����xR��@�b	��uG���¢S��p=y�}2�K�M'r5��س9��X@�C��y"g@^� ��e�.t~H����Ol"~��+^::K�}I�dMH�M����iH<������ѡ�9)?�d	��-��ɚlQ��|�`D��hU���1AF�y�#WcX�,GybB;Dp|�𲮊�X�n��`�������<��yR��i.hC���|P��VB_��y��^�s�<0!�R�yPH�I�cX��'�az �\��B҅J�z�&����'�az
� &�Y2m�7|jH��P�D� wO L��é��Pt����%�uL�����=����8�I�p'��2��^�w-�-ze�& n���U3��'~�\��R(+
ک�w	�	P��u˔�|��)擞
��Z�H'��ɡ&�=G�.C䉺K"����0XWP��(�?b����!��'t�a����a�V�s�Ă/Z���'��|Sc�I7'lΔ5�U�/�p�JA�k�<��4J��P� ��x�Q���Bn8��Gz�+{W���7��3�8�G�G�y��P6=;�mk�휧�\xc���	b���O*���iρ���ֈ�Ú���'�����$f?�q�A���s��	��}I�*�d܂2{yK�a8S��Q�ȓ.R�ԍK�8�J�P+R� l>��ȓ/K߈GK����R_�E��E5D�����({V�+$Å�����0D�t{wf��@�B�cÅ�jÚ�`��#D�D+��� @��F@ �g�~̻��5D��z�c\;y�l���"x#�D���&D�$�ʏ�,<�A��-���rC�M�<���%�I�"*p�D�L6_�I
#��8Wl,B�I�yG)�q�ֽI�D�B6��9{LB�	*�M��I<'N`�GI�A8B��q*Ԝ"qj����03��v�,��p?��H4j��xc�n+��hr�g�<��"Z�6p9�t���U����	`�<��M�͔4�0fǍU��te��<����$�Ot-
I~
�'���O ��Qt�I��(9�'D8�*tfD+M�p@3�?<d��b�P�ЧO�D��O�T��+Z�vv��[����Z�pY���'�Q�L�.��q,쉙���d��XP.F��y�d�R�H	����I��XZ�E��yҎսNżaye�Pu���MJ�yr.L-Et.E"�#V�t	� �����=q�y�L"9R���WŘ�<4��W��yr�S��@B�š�R�k�K���'ў�OK,�*�@2+M��{p �1�\��	ӓ��'$`"fF���Pp`�&?�Pش�y2�)ʧ{q. �e�X)>�외��5\�-�O�7m(}RU>�}ҐiZ����v�Ņ_z��	���I~��UE8�@��+� j�1x���,(��͹$e�Ob��ԧ(���kh_�>�<!ʖ��=�VU�ĭ�-[��B
�'9Dq݈H`��@�	$^� C�R�t��X~�@�k~���I
lxb8Bg��̒�Ȁ�y���-:�bP���ڭX��ȋ�����5C�1���T>�'�� :片�qOJ��t�Ȏw��+H>������85DԼ3����h�*�e�!�$͖I�����Z�1����c��5/�O���O��ɝ��-+VaЊ�޸x���.N2B��c��	�vEƯ\��8�����N�'�ў�?�cqi)S@4-��B+�Y�+!�O`� �'1���J6L���.	m���y2�'��3�k�	%)�1k2Y�hol����?��u7 T&��q�G��NѴLq�ꈐ�y�߹/��8a�9=��T�yR�;8�h�b�D��)9��Vƕ��x�ő�@��mמ"f���k
�!�D��Wy>C���,!h%��E%!��
��PH���0$ ��'�'|JqO���$@�4Ϡ���=o��X$�� �'��#=�}��� v�Ęp�!�9 ��0�X�$$�O�|�d`���R�ԳTؤP���^x�j6C��c�4S����h�-��:�O��d|��� Ф�W$[�C܄�h��=V�$��"OA��֥u�^a�r	��i6ܱ`��';�O|UA *�(&���GطU�>aR7�;4�����[��Y�� et<��f;�d��(O���	�ea�ot0�Kb��X1�a"OZ(�Ц�*q|d��@D 'ԍ��>���&�	���Qca�:~B� s�ǝ&D�1��1D������0݈���
����"-�D;�du��u����$Sx��Ս� 2m��hV���y��);�r�sѥ���(���`	��/�S�Oҍ�T��y��!���.W+�ێ��7�'��y{q��:Z#ZpJ�#*8ɸ��ȓzU��	�,J-5�H�f(�$2�F{"�O/� [t�̊x����F��X~��B�'a��A�o\�*H4��i|�&���x�S��(O~�=Ab^�}|��a��%�H�Ūs�<��(���B���E���Q�C��r�'��y���C�`10���*|���1E�š�ybB�3h�`!�PnD�nd>�Ҷ־^�':���'��yzp���!����d
�tS����'���ʗ]�z���FX�X��5��'VĨ�%�O%L�Ѩ3�V�f���X�'�h��!M;�����ԏ0�v��'&V��U�_�*��a��A"t*l�A�'1ў"~B7��� X�H�s�N?j�I��r�<	�@��a�&��!�=;(L��Qd�<ɀ��*t�| cV�Z�2s�%�e�<�P�Z+8�r����ܔb�^_�<AC��4��QQaJ٥ F8�* �]�<��ʯh��S*�#/�0t��m�W�<q�O�sM����^#6o���F[�<!���5}Ӏ��ǌ�tň!����\�<I��4��\��/ˇXT�"GU�<�S.\8�R�����%�,����P�<	���_��Pc�)E�8�:@@w����x2�حsp�t����_��y�
gp������i��M���y"�[�Ii���$�;eN^ŋDjY��y��\�
��XZA���X4���G��y�)�7G����R
[�W���N���yB�X:]DV��3i]�D�`��H���y�C�B�&1��7�A�#F�y2�¤skԠIr�-+*��A�)>�y�ɋ�g�(��i�R ��d���yD�>m�u�� AX�31���y��" ٙ��H!Z���-�y�-�8�bM�C�Ǌ�2�#���yr�Z�?�����M �,TD:�#H�y���d6�j0�X2��W�y�� Z �8��� );�C�8�y�&�P(Z�+�#0��9D�
�y�#˞׌�k�WĔ9I�@��y�b�.m���Ӱ��4�X�'���y�H�����ʋ�֪%���@��y +m��ɪbʕ+O�4� ��N��yG�>�$ՁI��?R�]a i��y��P ��{f퉗9�N%��c��yR�ʎ70l��t̞/	��`e%'�yRG� Xl���k����)ܒ�y"!��Jjp�pŖ ˬM�� ��y�QML�
6}�=��#��yB`�.$�s�E u�FA�/��y�NZ�f��E�h��衴�?�yrB	E"`#v�S�f^���#Kܥ�y
� <k��9Y�bA7l@	$w�][2"O��q4�A[��X�G-
�`���e"O��(�"،<�\���#��L��"O��j��|���R�
�~��K�"O*��E�@ [��	��ڂ,n�]��"O:���/Ò��e�$�
�c���"O��)	�!�|��4���~S���q"O��Sg%�OYq�Aa6S8�D��"O
M��D�:q��u`��+�y�G"O�I�Ѵa�J�2�l[�&xYJF"O44Zl��}(xd���ևfT0q�IA���jG��>�� ,A	)P�ɛ)����K	vl����8$C��YھM���Q<i�V�c�7�lC�ɛv�J��JS9*���T��&5e`B�I?`��ᘴn�RW��HwbO�&�B�I�w��bZ�4��%��NٖVY6C��'p0iyEaڇ|�B�PT�ل@I�B�	�~�~E�M�x�NBa�=�RC�ɑ=r&���MHr$k�덒*��B��]\rB��*,$X��� ��B�I�_Ң�#d��ps2�I0K�-WlB�I�?d��{�"��YB�)��I}PB�	�WiJ���c�o��۳&@�#�B䉽OR=���ܰeĂŠ��ޕ^�C�Ix����fS��Ƚ{����C�	�\�"g�kN����Y�re��dD2p�&,h6+�3#���s(	�b(!�L�BCx��%��#iʸ�GfUD.!��*D�(��_�-X�
�f�9!�E1_`�Ғ��~�J@�R&W�!��Z�r=(�z"�6��!`�&)i�!�$9*�� vG^5oJ�"0�I�Q�!�D*]춈ʤ���FS�8Z�Û�?�!�d��x7��ǅ�T|]:���_�!�؁cM6�Fi\�9h6�+���n�!��c�����I	�΍��cJ,C�!�$��<%�@�4�Y$���ke�X�}�!�d�fq�l�P*�;jQ���;�!��Ő'����I r���堞�0�!���Ȳ����z�]yu�P�!��JYH	�vX)��4����	t�!��
0h#���M�4�N�J3�W�h�!�
�"( ÆʉW�1�p�kb��ĝ[�p=i��|�x���y����ȁ�̀C������D��yR�8+�P���
 r$`r��؜�yba��g�U��׍]��0Ca苢�y��˿@�z�2��8�ʌ�`藾�y�,P)ij����J�"���T�!�y��z�<t��Z�;�@{�i���y҄�f�DI1�0�����<�yr+ٟx4�q�N�v� 8aE6�y�ԧ|n��w��0�R�_��y�-�+\80�!�0��)X�O7�y�b�GHH��dЪ�p���舐�y2�88uH��QH�p�P����ċ�y�R�\�v �gN�?kz� 8 �y�J�87.�"Cl��e��#��
��yr��w����gѾYk�!b��N/�PygT$uh�q�nQ�@�ı2a`�q�<��ϭ<c��(�N˝>���a�<T�ьh���jEcЭ.���Qa��G�<)�d�o���[��+H��YY�v�<�.� )�����H&M%�\W��j�<� >�Q�m�嚹8����'G��"O��hq6^�^qh&��6�"OB1�1K鐥s7��#W@=�"O�#@C��>dh�BƇ`C:x�F"O"���$D�W�w5J��q"O&��&��;���D�<=6$��`"O����F��@8`U�J#4՛E�'"6ѓUGOʦ!���V�����W��$�FL9D�`�6ʓ�8cD��u��	#[h|2�I+ʓ#��l��S�9aF#|���;bWf�Q��/���&OS�<y�LهFpX0&����T0��WȒq8!� �`�!c��O��}��"�j}�&D�@ܮ�r�!������5�E�%)� �Tp�e�Y�O��mZ�i�"��[/2���� 'Qd�x�h@�;�H���C�D�4��Ў��=���$�6�CQns�S��d�('�;�^I�a��Px"
P�;�89���=KV�@5�B���'*R�:1�U�Z�1����>����|� G��M8��'m $����Co�<A�lYJ`袯K.leh�G�&˘��TA�*�ɂц&3zdF�,Oz�R$�
i���j�hX�X�#�"Or�����4�bg^.))(
�̵@B�s}���R�؃`�p�?�c�2C�"i��Iy���p��b��tQ���T�ZT؄�65��Z%/�5<�Θ+�%F'� (`�+W�X��ɞUd���j�;v36�(6�c�+vM^)<��1���;������q�T/O*3�
�@s�L#K�D-����.b� aA��@N?�*I�t��d�(C~H����,8+��Rhi��c�:(BؚF���*H# 喧�uw���q��O�
\��IˏP���!��nPN���@;%$
��S�4D��+e��v�X��i��t&�a�w�=S"�,"��	�:��Q:��{Q��U�N#p�h�Cɞ$q,�}�7e��?�҈��d¦���	��|�B�.LOF���ٽ:|j�'B�%R�ʒ^OZ̻%$ md�@Ag�#%���U�Ľ[FȀ�� v�1r�/j>śE�P�o6�l`��66k`���1X1OhҖ�4T���RJ2u{��a>�8��Q�i:Π�E��2����2~G�ႂ��Y&�%�a�ȟW�:4�W�'�
=A$��B�:���vc���MPBM�ix�䟫vR�8p7F��k�)y�d܇H�*��̃ui��&M�E�.���"�4EW�lYG-Ǘp{��k�'&��"��P���p��Ȝ�:����d�#�	�1�&o����so�M,��ZR͐���X�vH��<����O.��P�ۋl�� 9&DH5�V�3	ۓ$Č�Y0�������e���>a��AKÜlZj�����Ll����Fɱ�$=(�P����S'���l̓L���� ��l�2c	�;yL�>	ѥ<���OÀRX�eڟ���\�����O�z�&��%�֣ а��Y�,����[�f5���e�B�.]j `���}�"�+���*�F1�r�bx�������J0QO�|���_%���N��A��y��A1��� E\/���c"O��K��V�2����|��h?y�*�u�� ��o�2<V�uE��d��iJw����K���ɀ8̞���N��Iv4�C�؞ ��}R� ��ۑ@�R�@=��,�Af��1p�)
� s��Հl�6]1DV�D#p�4�g?i�YX�23�h�&~��qJv�'Td��d� c�'}��Z�O؞Dܰ�q�-�2��I,w����$�
 �鉊\��Q@�hX',�"�N�e�������l�:f�_��s"3��	S��`2=���2D���*@V뵠��@�$���+��T�"د�)�7Y���Pӈ�#+�)�t�ϟ(�H�ZA�P�Wt��PD@ɀ�0>�#$ƣ O4����Q{0�1L�JdQ�z�80A�4��nJ�Ed��ߴ�ħ(�1O(�(A �%h��2dO#CX&��q�$K$;;�M(1"����'9?�E8��z��1O�=G(�K$���R�֡�ߴV8�q�GH�x���D�")`ʽ���:d�*�����8��5Ң�]�^v䤧OT�KtŌ84���I��iat$�F*t�kL��0��h�ƆJ�T80�=8�!�V����S�_�R�� ˗eЗc��,�>C���+5쌳��ɴ�:ͫ�jY��'Q�,L��!ޓ^?��z��U�q]�m���'���G������ҍ�)�M�D�U�I<��B�'���!�%�\~�%K���c3��P8���5�͕
��lARC$�x�U�<���	�O�``гm�2�f%Q#�"�[.9bN�zrF�
*���{Ȝ�"V�"�B�Pj��
�'��|���T8kɔ���2��=����5\����?p�ê�":��`�@ U;nΞ��O�N�E��m�f.�*pC�f�9e�a��&��}i��RCN����pԸ�pNB�2�&�8�Ũ,�8(G��F�&�ɈA@���O �bL��:���H����/ ܽ�B�?�A�hz`NY�$�*p!�N�`�dh���?��<�R@B�lJ���<\�<�ci�O")D�''>2���S�? �ș!IӾwt�͂��XB��ۦ^���S/�*ɖ�PF_6tk�Ę��_�9�hY�r蟛���8=�d�j�%[�D��D�F�8�ΓcH<�c
����D%�~
zQ���=����)� �S��%4)d�]?9��G�6� ��Im��]�n98��6(WX��Ys�r�����3D��Ͱ��ܰ)�p�C��ݤX�����I� f�-�k׹|�Q�����Z���00��Ot��,W�X��'�62�ˊ�r�H15`�:+딜���$��`���K��R�6M�R��qH��țA;@� �c��`פ_�t���IģTϟ�0Љ�sG�}h��'�^�H�IE�d	���H�7��y�'(�9Po�<A����+r+R���b]��L�C��O��b7D?E�5[�Ⴠ��9��S6I�#��s<��_J�)��@�A�24���"sz�݈��!:Ĭ��^8�G�O�$y�� �D�*�@����������0�,�?�Tl����f~"�'�p�S�A�G\J���"طF�ڝ;� _�15؜ 4%�.(-�q�i]�s� #C��BVZ���bضE�εk�����D��7հu �+�BO����MYlQ�,j͛�s����+zܚM�� 4��Jul��a�&\k%J3�Lx�E�,W�x�(�,B�4W�� �Z��=ͧW%��˒B��~�����I!��'P��>6,�I
�����UQ�U:�N�٥�MK%�ؿDږpX��V�4�`D�u�Q) �D�{�-I�hO?m�`C_'����)i ��ehf�h;BkE�S�<�#`⌣�����0"�D0y�8*�Z!��̼+sf�,?޼K�D�>9����v~��'#H$0��C1��D{' ��/Q���ŀ <>��H�s
`��e����^B��C�x�_h(��͈�h�`r��>�0D����8ʐ됼8FY�7k�W�H�aWC�0b`�����6{��i���Q��͹�	�#D;���AY{o��=!��Ի|v�erfHP�s~U`���~
�h֛-��TCR�]&�Z!h�d�<iw/�{�4ـ�Ǘs����C�<�'j��
|h	�ʛz<Pxg�S�e�h�'�5n�0�c���B�	�3p�!��Ő1+|&�u_�Zw�C�^B�Ĝ� ���~&���C��{P�1g"��J�8	�B�74�|)�a_`�����뛹t*^�p��ؤS�����|}��)��W����&Ϥ`���2d��pr!��G 9��yđ�~�%n
xqOց�H��0<1f��(�P��H�.x�ЩK�AZ<9F,��2�����r��j�2���s�<��?9�h
ps4ȁ��H�-/��Z�WA�'���P�; Ȳ�$>�����`� pѡ�W?B��1E�5D�$A��B1����C��M�9�2ð<�O�Z*ZI�$*}���%K��ŀ��1qM���,�:M�!�ę�l�����@2-d��q锘���O^�Xuc�*7+��qOf�'b��{�t��v�ǛS�z$qp�'Ul���"	b@Z�r�O:e�	�⥊Z2l�pvUi؟�bR���u|З�̕J�l���%�?#�i0�޼0R.���Xw�N���D�L?~̀��"O$�X���k�術�����*�]�����<?�2��S�>E��%�(�Lb�B�.r�60�E*���yBB ^�z(��fjyt�{�ƃ�^&�'���J�DM$��ϸ'����4i�%���G�!
�]��'����E#$_JX����5g�^�J��SX~!R��'�:�J#�X/���[V/O�CY9!�b7����N9�=)b�1��lL�T� 1�N}'\B�I�g6Lpr��îs�����L�0B�$E&ґ*0*ɲ��0
�=Q�B�	}2uis+˩E�h�$��]�B䉒$���'$����JL�B�ɗ ���Q��li1Q��ON�B䉂LX�C1�$��c�푰%��C��:iNq�aOU�E�x�5@��|B�ɢC�	"Ƅ�?�v$�E�4B�Ij���鱣��'�F$X��� A�"C�I�&*����¸&a�R3$�+enB�Ʌ9�ɹA�	#j�UY�
[,B�	+u��4��T���8�r�
HU&C�	�TA��c��4��`�
[C�	� �I�a�71`�(+򀛈9�0B�I�7�|��o�#$m��C�lB�I�q�J����0S�x$�Zd��B�)� ��CQ�̮0����P-GѶ�r�"O,"@�<y �ᡄNKo�y�"O^e�J^f�n�A�T+;6�"O�}���'��E	�ٷkɎ�K�"O|��D� 7��̓�
4 �NB�"ONM�� ��q�쐉�`��L����"O������6p�r��
a�}	�"O怚��G;�6	&ș�V�fh{R"O�p�a��\�f�Q��C�|/~ub@"O<%�&c<{�T��fv��Pa"O��Ф<���`����PH�5"O���䖞3�-!4�5[B��"O"Aٵg�<�Z���ɳI6 a��"On���8~�6PQ���+$/0�;�"OZ��u��r�jT6'C0���"O��z�k�5n8��B� ��e"O�i�U����C���{.�#"O"�@�\ �����Zu�%�"O�9�Kߙw�<���d�?'$Q#�"O6yk��4AW
��1I�On�"O��0�#@?����[�i�T�"O����� I堰8a���%&T�3"O�7DM-�r���j��0?j!�d�/O��<)�jF)zÁG��!�+P��+��g��HB���!�E>'e���˃$�P��@K3�!�� nj�h����]�N��S!�!��U7`W8Y�]6v��yb�Exf!�$*8:\�[�ċ'Y92���=4�!� �.��e�ٹ"�Vm��9z�!��@zx�i�6�A/`��D��,��!��2%0��*��%�(i3�E7�!��-0$��Q P-Gt��ڃk��!��֡�	�g��`!��(��!�DK�!0nY	�PjD��(ػq�!��
/�bM���� |�4t�A�Ӡ	�!��}��� @灴=�BH"�I̓:�!�d��qb��ՄS7 �jP��+T�!�� 'n� \����Gɢ������F�!�$���ip�$"j� �;B��8
�!��O!܅���B
VU��Q!�ȵy��$H���\̼J�LSz!�D�<��k�CQv��ŀ�=x!�dF�H1�(�T�`�"D�T/!�$� �e��(a�M
���Ga!���,��$
2��7b�V�k�̎6�!�䜣 ~��ӂ�<2�0@BaKQe!��;Ll@#B'��1�$|��AȪ�!���$y=��#ק�@�tpk3�=�!�J?v��yL��9�6<��@W�5e!�Ƞ����D��4F�l��<2�!�ѲjWnhF�@=G��A�t���O�!�+.��s@ÇY��:b�*:!��O���\��cƙ*n ���;{�!�DV�U�H���J�/�\�qsKπl�!�D_�6xP�k6{�����V�&�!�D��<"���Ց$��EcNߧm�!�䉌�Z��+�@<mSW�ۨ"q!�Ę6x��;+����o fk!�d�5}��Ά(>L�DS� 4Z!���ODV�V*�% [�%��ŐT!��E�t����2`GZ�ˏ!��P�<�z���	`:(��W͌�h[!�dW����[��/���ѐ�W�^_!�� �a�2L��+Ԕ��EK�;�REy�"O�XXƇϒ?�p��E
�+���B�"O�qr��6lI!�	�*���W"O��	��@�s�ڭs�JR�`�6@R�"O�%b�ϝ/q(�9ؑ��\�X=�"O�,r��_���R"o�"UpQiD"O����`�,����@٥X�!k�"O����f�n��1�V/G�7��m��"OD�YrI��@�^�8��/]�x��"O��� �@ u�,�g��D�<*�"O� P�W�+tPBd��	lBLZ�"Oz���aM|���9�nU�_�x�$"On ��
��E�Bq��O��v��"O�HbwGW,h�P�d-��|�j)R"O4(&���S[4Q7L �o�v�jf"O�`�@k��A`p٪���+$��S�"O�\ �+��@�Hae�9Q�eJ�"O�9���M"<R�Q�h �X�X`�"O��f�kh��H ���^���I�"O.qB��ŜĒ�F��R�.���"O2eR�&�5��cgNاRwX�X�"O*z��܁���"�֦F��h�"O���O*n�<Pj�l��A��!�"O��ߒJFar��Λ'�:�#"O����ɛ1�f��¨э
�y�g"OT��f'[yܺt�b�ą!G\���"OLa����X��hf�`�!�I21�Hi���	�O> +f��l(֔#Џ���iKcØ0�~�朁f9���:d�,I9�@]�S��@�#�3sy,�S�o�
б$���?JV,x������l�	���h�d�ұ�wdL�,q����>B�I�,��\¡DU}	������*�(��O%NPaЇ��|+T�B)�7/��L�ᄕ�~���BA%����k�8k�ă�k<d�ƅ@�F��{��V�oV�*tΌi��9z��J(&\t��1h��6l� 0�n�#ϸ�2bEF�FP9c�q��1r����(�y��!5ڙ1$ʎ�2<��i���'52ѳ��Gf���dd�)Hx � 0��6J\yk���9|����Ф�s���z���6�@��g/ݟ�0=y�&�_7��Շ�;�>(B��5nf���#M�[w���1i����x��ǬZ;�(��'
;�4�$�j�q���R� ��!�)A�~�So�1DB�I�H8���
&a'~ArRh�]_��$��Y.�x��"�ʀ���ȃN4�!��B%g-pi���^Z��Pst����M�,�.�˰���v����c��YA�V|l�K��?��<Y��!
��1��B>vL���Αw�1@��0�(�s���?�C��D�z;��C�֐	���3�D$�OD�`��C��x�{6�/"��%8Ř�^-ǚ��Ð�.�ڰB@$�q�b�	�4 Eh�+�*azB�[+��i�HY����u�%��ʚ'	8h���1�yZwL�����D
"maT,�=Z����J��[uo�1�,�T����"OX3���@��߯y�`����O$��;�r�%K�$q���W�A G����=Q��hB�ODV]K�.�<X��mS���z=��gҀ��Ƭ��5��ŏ%L\K�$(Ѹ��aA�gV�Ty�T�L˂O-�g?�녹w�d RC�l|���Ǡ�D�'�ڱs��M�'`7�<��Y>���K�D�R��8�I#h9�e�)ʸ1I�ȇ�	�F��@�l�!F6�q���e����D]����;ȉE��gl�=b�PY��a��Y�rh'D�p��@"�v�jP�Ҕ%�F���������ԃk�
]�{,a  P�];�)��A�EfAh��	�;�b)@�+L�0>Y5�A�\dJ���H/.����?2����\P�
$LĪI*"�#�)>1����\n\n�j�S4��'��@���@��)M7��@Y��^+�>��tGBH�S)�:��d�_+|nP�&)�J>��%^�c���n�+�.����Ɇt��z�B�iC�l{$�%M�`-rN�%_-�<���̴D&8�'�P�B��n�Np�ܴXI��V�׊�5,3}<���L�67�|��`Ϝ �y�g\#pmL�Ӫͽ����@M�1�?���<��ܳ!̚M��,qB��烘t�Sf��g%�)�^�iC&�y����8*{J����7���+0�󦝣_/�ұ��	;����I>?qw͓p$",1��3OR�;��»k0H��2d$���\���`�!ϔ�p`�����О����6c%�-��ܒ)�ě�+�2*��顁���J�%�IZ��ҤG�h�Z5A�
�<W:���E^(HP`,�v�Փ�Kş(JD��/�%+4X�>�{�? D�A-]\Ox\��G <�S��'�Z��#n��Ȩ��h�$	�veD6E�&p ��*X��y�Pʆ!SFPhCdKb������
�| E�>Qn���I���@	�%SS��[�'�p�O�"$Z���X��,w*<k.JQ[�Õ�?~^(�%T33Bxԛ��T����'E#yWN!#3�'���r�	',��1�i%H��ݱ�O$,Y�.O�J�&U�ů�c�d���B����$��M�,�.��� �O:yP@���N��ԛ!�9$� ba�P
j!:��'ȑy�\�F���~�i�>9N�D�c哵Y-��H`Z�o �@�D=O�����$�7BE�Eɐ`�~���^BP��E��`�t)#�@Z�>ͳ£�^RT`)��3��� �?-0^-��'��iĆz���@�H�� Ŗ4r�ZĘ��C�J�G}R)�
\tyC������©t� �h��5��ᆬشn~�J��B�i'�u[a��O�]�fg��aa$�0<ɖ��;� ��U0`i�Ph�gDs?yF敍c��=+�e2=#�m�&.�ekH�8F�X���cBٴj��WF��o �s�N��*7|봩V�r``C��/uAv�0���Ѽ-It-S"zx�B$G
���mڒG�&�Q"G�/tDx�Pa�Ѷ)��R$pv�]5Y�>u���߿_ļ9�R퓁w�b������p��T���u*2���� =v9Ī� ���Hx����@��dA0@��_V,�s���N���1��D~�(�>E�bްt�H���*��O.ȩ��(a�c��KV���ÅÝ*��)r�ʕR�f����4��o[��R��/�:b�n	s����0<�ԆF�h����%���^�NH�2HA[}�L�C���7
�A�D:�C[7B���B�ɭ{/�D	�4HjfHs��U�݃ŉ�'�x�����4,h,��#���B,�����*���l��3�֠���Ĝ�%*E�п	B4 c�L;�\�!��[�T�әw$� L����s̝�36�y"	�'x����"/���A�0d^rai  9O()��N
+�{F�֕��I�wPdP٠�x�����j�C4`�-���!�Cy�a}��fȦ���� TMzE`LI&h슶䙥�h$"$V��*e��M1T��RF�(2xR��G�W�G���D{B#S�W1@���-����a�s��	$U�
oK/:	��1�=�yBG�4���Oſ1�|�闏Ο�y� ]��P�33-}���1dg>�X7�=�3�;uвu��/;8��хȓ:��L�gN �8р��1��@��/K$��ɳb"V����L<)T�.2P0�m�3�B|bc��mh<ɕV8|�4�bt���;��c��Td������0?9�	�Fa0�o��`�詑uF�y�<��
H�ĩp���;N\i!e�Lܓ'����'D&O<L���0b­a��;NQJ�8�O>D(�R?>�%���ս{�3�ʽ5M*����:�Or̡�a�:���� �Սg^��W�I�I��*�cñW6�OE�����C8:uj�ƅ�M�je�'A.`+P&��
�2FM�-F8���.O�D��7X��N��|��$*A����� 0Ō���Cq�<Ѷ�2*c ��菪;�����o9�Tr���ጠ��g�A0Ṯ!�ԧ4*P�T%�}�da����C7@��!6q�e�F�M�ح��ɍ"fv|;��'9��懖U2�*�fEW�a�����PNA�DKȚ��'i�>}�ceE��8Bm�m����I�$�WᎿ,v�x1O�\�'��|�ѢD8#nT�OQ>U�"e��̔�D��)r��I@"O"D�(��Q�6SuB%E.x�բ�
���	�]���5#T�3�	�{@N	��G/J�pT	ǀS
�B�I�zDD�qԣ��F�a�R?Cz>�'��E9�}���R�썡@E�8=V��׬�M\���G��P�y��o�
�@���43�F`h�S�yB���Rt�e{5��.q�y��B��y�+׏lf�9P���ht�A[Ҡ��y�f�&'��Ggɤk��(�A��y­@�fR�9�!� u�K�
���y2,:��M�g����@l��yb��1�.D2GB>a���yR��&&0�r؅����>�yrD��~P�T)T �#_��鎥�yri !3�bX[5C(@����kڏ�ybn��r�����q�TrN��y2��yzi{(�/wux�8r���y��?lL���R"2@�	�.���y
� Fhr֥�'M\��!�%41l�3"Oļ!�D��-�tq�m޴,x��"O�}ʓ"[�$0��D]8��"O�(b(6��!I��V*����w"OvA	�O�&%ׄ4Yd�7D��Ep�"O�)n��[0�131�����"ON�!���:E�H�*da��{�"O�ds�'�� aF�Pd@�8�̠�"O��Y���wؾ�A�@'w�Nt�"O�#բ 6�x0C��F~�@�"O.��F�%��\{��<[����"O"���_3������M@��"OB���
'X��d!1h�6xOT���"O$��s��R�(y!g@�M=� *F"O|t���L=}��,y��H�}8$�d"O��C#��lD^%+���hK�"O`�ȥ�kؒq{�ƆV�l$�6"O��ґ��3Y��X $�(H��xc"O
p���(w�0�0��<7 	Z���,���O�ax,�W ǧF��I?g�D�0L\�	�|8��Ƞig�C�I�g�.$Ӓ���j��1��q*xC�	;�)��b��%nۘwΘC�Ict*$P���n��d���"�fC�	�n�P��"�J���-)>C�$���*��>?�Ub��;x�2C�I%ӈظ�+����"���72C�������=-a��93M�)q(��HOQ>��%/
*<�������ovZ��"*�Wt�4��#\:
�h�ɨ*�]xU�~:����O��8c��G�Q���a�`��L�aY�m̳Y|���6$L�фX��I4�'w,rA�W�V�g�U�a��* ty{�w��s�.�:��b�w��S/:F|cf]"B�x��0C�:r�^�Oz�� c��r�1Oq�,6h�)3�2�P�,@�Ml���Q�¤b�3 �4c��|��c���1�*N�Z��<!��D�(i .^�p�qOQ?-RE��5$,$�ҍ� >0pɒ�U�XK�{rY?��'�O���3��� �1�dN"�>e��O�3Z���鱟<P�	[x�S� r�OM���V�HA|VY�'����{Ǥ�o� m��k�&��1�Qp���`�O2�A�6O�dJ�� ڼM4lx6YԦ�a��	7�D������?A���#8V0j�m�*�)z�-���M�p$��Fl�IGcE�EN�Aۊ��'JR䋆:�!�Cܾ|��ꂚ|�c�>�Oq�bL��O&,dR�qU"�u�\	cQT��Au�5�Iֺ�?��ٕ;a���)W�`����`�v�<�p'��n7$p��(D)Aܐ��c�t�<�q���M)�a��	�y7��brFI[�<c��,P��$h��(T��B��|�<�e�T�?�Ę��� �"�p"���v�<1!��o�~�2`�S��Zt�EI�<i������7�M�mw
�+�`�<Y��}�4��UJW	 P���wdIr�<I����z����l�![x�#u�Mb�<�,X�q����c!���.�cr?T�0�� �<%����U�9r�)q��6D���f�#'
r3)�c��[El1D��@�G �(�`3F/7F����3D�pc��M�yX[�V�E�3��$o4D���e-�3ԠD��L�R`�1� D��Жo�"=��4c�#�;�b[e!"D� q��4B��H�󥄤Rg~���5D��
N�*:A8��R �5l�E�� 4D�hk�1���� /H�҈���7D�ԋ�^�%&xY�D�Sڍ��e8D�����7<�	a�I\���-qU�7D������P>�]�ժY����r�9D��ɐC�[K����
T�w���f9D�`�$� ��z"mR8>�J@z��� >@ڇg��J�J���[i<���"O�x�FE�\��0d�M�H+�"O�9�G
�� ��Q��ˑ?4Vջ�"Ob �)�zp��〤�� :d"O��b��P���Mz��I[�ԁ�"Odܻ��S���U�ӣL��h�PA"O�l�AR�q�S*c2���"O���qc��*�`�W��%)@�q�"O԰6�ʴ�x���� �Q�"O��"2��X"}Z�J�#�r)�1"O8�;v��by92Z�&�`!���y�/��Eg�aQv	D9�^�aG�-�y��ƑE���V�� ��@ 2�y�%F{�`��B�fa�U�^��,��`���
�*�	���� ϯUXJ��ȓ^��x�
�#����.}��ȓ"P��0D�@~NM�cl�EK���ȓ[��e�F]�6$��bFF!���/&����Ll1�	b� ��x=��84��8E�ڰ0`�A�.�(6���J�} ��sK�a�(E�@��'~>��Z#�L��G�3NP1�'���r�m-$�t���/͍/���
�'�ĭ���!E!�Mi&�3*��C�'�F�%N� �S�K).T�z�'j:�9@`�3Q��l@A��i��}i�'%ܸ�ug�=��:6��L��,��'��M�L	�g��ʥ�!=nʱ��'��؈�m	�_�8i��ě�2�Zh��'I�0�Ķm�r�t�	q:y1�'�B8x�*t�0����?R8��'�~�)� %������3aF}H�'�J�10�<c�����N4-��Ё�'�4���mF(�zup �Y�%n�e��'�rX�bBԬ|�"�j0�F-�Z��
�'��]��K��D�k���!�V��
�'C�TE��d(؃'摧�0a�'$�UG�=Y�]��B����'oB9��*�v)�+�	�9�����'�����O����V�,[�\��'� ˶�Ϳk���2��U."`�h(�'�n}���ȴ�pX)����4D�LA��0s@E$���]����Ï<D�hʰ�"(^��Ê�p���*O��)��ץ�ʝ+��#D����"O�-3�i�`��㯓�H&�Y��"O�@�A(�=,Kj� �m�!Ć	�"O�Y�d,��9�V-��-̥
�hs�"O�q�e��/߄=I�U4SZ�*F"O�m�b|n|��+����5"O�!����'���� � [vH�qw"O&�[W+��8
���F�:sR�I@�"O6�"U#۽Ƃ��s]�<$�DB�"OV��s�P?,��"��A�ld�D�#D�X�� T��p[��z#�+Cm<D�ذc�y?B%�t�Y� �,�F�:D��t+O?.bz��-�3j�A�#8D���b#Rk�� K�k�!�� S�a5D�܉f�݆Z�r�����^(J�ktc>T�T�����@�X�:�BM'k��x�"O�����$H2�;#B���H���"O�� �-�1I[F)X6���<�"*�"O������ 34(h�p�Q�"O(=K�䝵hW�q#��Q�/��\B"O� ެ��Ϛd����݋N�.�$"O$tg'�$/K\� �J\�$� a"O.�!v�Y9)z0H����!���"O��4��o7x�h	�f!�|*�"O���t��Es��+wf�
"O��`A0��Ł���+"<T�s"O��*Ů�&�,�CeJ�I��� "O��JseX�zU�!뀁Л5ʾ���"OH��+ҤO�����/$�h���"O�=�b�K�G�sa��;���)�"OZ!R!h��.���ZR"՗mX���"O�	��GZ��.Ÿ"�& [�"O��;�n$mk�\��H��"O�	I�d�:D"V�B"KH9.�ъ�"O��b�Z�6N&09t�ҪF�d�e"O*5uB�<�*4C�55��mx'"O��J�N�5٤���M��Y�%"Ode1-͘*��K��8�zh"O�5��Cԫ=+d���'[D��V"On�)2�G�5y6)��R�8�"O������F������?vcj��"O؝I �� q۬��B/ߪ%Rֹ�A"O�$��bROU���C�Y2�p�"Ola����N�䑱���:!�,��"O:�R ��u����u
�4o��m�q"O�� BJ�L�|M`��զ?Զ�"O\T��(���T�#p	����H�"O�@F��6Et���"�({r��"Oܔ�����,(��̲A_PDp"O�0h7�F����ID�,�`l�T"O����%��f��ߑB� ��"O���s&ȣ%�Lа��=
�mJ�"O%�#<i�ppׁ]�S�|��B"O��3C�q�@Mc�b\ *�����"O�|A2FL�-⊭*cl����i*�"Oz����*3.i�I��v���"Of��pFY"dL�b5���U�V�f"O�Ȋ�%J�E�d`"�J�b���"O0Q�"ʐ�WHViy�CI
K�P(c3"O�@��b.m��Pk��8q��tY"O�����X_v`AZ�e��M��y�!��͛ � �%Ұ���Sf�D��!�$֌v4ʡ��o 7�6(�F��lv!�d�7������=q���g"NWd!����q�	L2!ɠM���F1`{!��4n=Rm`%���	�����@߲]!��g0���#�_�	
�$F� S!�D��&l`�eBt#�{D#��$A!�D�v&���l��XAzQ�D��~!��H$2t��T&�Eˊ5�r.K�7a!�$[�57 �	���=z��(T,�
0w!򄁇{��u��o�y���1f��k�!�<r��]i�G �R�@A��H E�!�䆔%І Kg�>i��ᵁ��k`!�$��(Ƣb7AP�W��]9ԭ[�^!�Շ_�QǤݹP�`��vl�%!��B^���$�$���t�F��!��E.4�~9�����3�=��I9�!�Bop����Q0Bn��r.M*d�!�(�⣕75�a[��|���'�h�v�<t"2�*�`r
v�*�'����n���ܱZP����H�'����Sf����f���q��'h.��׀
4K60�qt�ق}�t@
��� R�Q��<��3aA&(��IS7"Ox��Pf>*^�����a�"Q�"O4�9�lز����h 5rL�"O�����֦O�A�G�#L�n�aS"O���ReU7*���@�26��-Ä"OT):e�Φc��(�#`�5sX> {�"O&�dn��]���'.k�~q��"O�Ȱ�ӎj'2�+%h�i��8��"O���� �7L��1'���)K"O��i�����\����"Ohhad��.���A ДJ5"O���M"k��C� \�@�f�@�"Oցc&�Bj�"�.D��pf"O�H2�A� ��1p�Κ�J��F�V�<iC ח<�R��s��>~�,=��CEP�<��I Fp��zW�>09���E��O�<I���=��\���S�^�FT`�<�'-ã+�\�H�MLj�xf��_�<A6$�?,�j� "��D�5:��X�<)�ғh�t�b���X�%���H�<Y��&SN�RУdֹ���{�<qTJ12P��Ė4�Lp�6DG^�<Y��P����ꃈW�d �6��R�<�0�3q�F�@�^i��d�c��L�<�D�p���p5��Al�1����K�<A��N1NG$M�A��Q` �c��b�<��J1��<B��9�i`��B�<q��[�
�du
�JI�]yQ�S�OU�<��m)h9�)�@H#vLd$9ҦDR�<yUL��b5�cR \O�A(��r�<ѣ�q[p���MRżu��p�<y�Fܳv��qɤ"��F�KDoZG�<AeIBr�<p�]�t�y�@B�<	Ң�@� ���YN�q'�T�<1� -$�EB���-AwV}��H�i�<1%�1>�|x�ñf6@P��b�<I�H����ѥϒ2Z���My�<�r؈Z;���a�H6t��+@LMt�<A��	;as��"��c��S�̘J�<aiJ���Y��:�^��� r�<14膢6���F�\l��"��j�<��IX��5�����~Cp(�ld�<��C�h-Ii���b� 5\.B�	� hl���L����r�`�=)TB�	�X�r�����7}Ϭ�B6hī��C�I9y�L�%k�{޵�E&k2�C�	�C��u�hQ Yd��3����+,C��/�*��2$$��%�r%�f�`B�	�U��@  �P   /
  T  �  j  �'  �0  �6  
=  eC  �I  �O  EV  �\  �b  i  Po  �u  �{  g�   `� u�	����Zv)C�'ll\�0"Ez+⟈mZB%8牶7Zn�D7sF��aH�-똅�#��n^P�Ĉ.~�� ���DV����	��o&U{��	 ���'o¬�a dW�~����
��V�
�[���F��vp2E!B��a8��4��R�rԁ�&��*U�0��I�u�݋3���m�Z0#n	%ye��IG�Fh QCڿLh���4/�����?����?�� &�-�ᬌ�\��e�)���j��?�'�i�7��<�����C�'�?��>E"U�v-�J�5!�A�=\E��	���?!,O~���<�CĎ�a��'CBk��"�@�3��@�8�I��#h@��DG|2�ieʅ�Ԋ�W�:9`@`@�r.�x@Ǥ>9�'�'U�� !��)a���r��w*D�)�����'���'��'��ٟ̖O��X�;��p���޹G�l�C P-%��h�^�o�1�M#2�i�"Fi���o�!�MKV�i�2Գ]sj���Ɏh���e L-�ў,
��)��<dY�q�I,IV<UoO4>�ֹ�C�����Ȣ�Q-�6-P��q�ݴ�R�O5L��T*[B���Ǎ�j'x5 �j��f	�D��'��� �eH|@��)RN�]�$�{�ː0� �i=�7m�����%P7>_�u�WMV�D�PQ�@hJ�M uP�D^��f�R�4V��f��|S"�`�}S]w@�]�uI��F66�!a�El.M���%*V	��H�*����Զiw�7M�ʦ���5Z~r���H� �(�*�K@�n
x�����=�te�FA9;�T�޴!$`02��Ю J6, G��>L
�Z����E�Q*�aVM�%��P�"�?q�B�'�ҏ$rM&7��O(��V�	�j�!q�%^��\5aH"G����O�ZR�O��Du>�(r�=��X��'���=;$�7���6�Q*f���U��Q�|��&Y�R�rb��3�P@o�<��\ѷ�D��,c���
U[.Yʀ�C�J���0�e�OH�$3?�oI�o��\�S"m�)Z`�W����	��?E�TCX?��x�0��:�D��o����?���'��-�G�%�F����YW"�S����'t�ܠ��iq�Q���0��l��!��#a�k"D�!��(o�J9qN�z
�Jk D��%�����g�S�|�ȑ!1� D�X9�)�0#��,ڱI�7S~��S>D�(:�j�]b5iw�� o�H��`C/D�,�0"�8I���wAǙ}nX�� �O�phC�)�D��d�D�/' `�({q�E��'(�|*�ߍ��1����)y�`[�'���cW4Th���ϑ�?6>��	�'ˎ�iσA#ʨS��;�@�	�',�2q/(s��l(q��.@���'p�����z�*� 2%�2E�(Oҙ�'��:��a,�BVOȖI�83�'cf��lP*+��B�
��|	��'����I��L�!&�%:d��1�'��${ ��p�$��%���0��M��'3Z��"eB�C�`5�ul��.���ϓe�Tݠ5�i^�'aH���jK���p��X!pn��x5�'�"o�6G�2�'�	A#���c�lV�V@yeF��f�Z��E	&��q�dL�!�4%H!EXA�'k ��7�_<J8�DM
�
$맊���]���� H ,*�╝.Ť#?���R��I��p�I�c�`%p�(��nn��Xr��� n��'��S38n���P��Ē�{揍#�t����̟�H�'_Τ�Cj�,\���e�O4�3f�.�'�y7�
1H�(�;��J�y��{E�>�y�c	~dMA���x��������y2��P�&��#�	u'68I1���Py2e�
o!��D!K�'�^-��MNt�<A�ۓ`'������I׶��E_n�<Q�i�2Xx<�
T\V���(�Mc���?��xӂ����̀�?��?�ӿ[�EJ��Hɡ �+.�p9� ::�� ����8�rm#�a�� ;���F �C�hج��#��d�BŚ������ׅ^N��%����(����It�2\�^u�r��6&�A���%�'��ɴ ��D>��O����OF�����~t�<8uD��<�8�&�=D��X�		�PY��ԼY^�wB�<���i>��IFy)4i�pİ����c�,=p!��l�@S�+�1;���'B��'�r������|���ܸa"I����&�L@�%%N�����.��{��9�zȩb�&iwdH�!�[<AU���d�r,�C?��℆��3��	J<�����UB؀����'oIv�h�EP�<	q��Q5�x+�o�p!Th�WJ�I��M�N>�(Оs�ߟ�1fi� ^��u����**�F�s�ǟH�I%iyΜ��ܟ�ͧw���U�H2��]0���P�6�� ¼i��c�a�uǍ�s��'���6��&����2,4*�B�rӼ���@/�2��VO��0<������	m~�ȓwPZ�j��° �&�RU�����?yӓK� :U�ƍ_l�(�a�T�Z0���	 �?9��QrWj�ۑ��氹@����Д'�6x��'��>�ϓi"��k$��M�A��k�a�,�'����8��+ËȽ_�f8J��2)Ӣ����J���&�^P���ɽR����w����MO�k��}����b�1�G�������~�nG-�����*G���}*��Z~�U�?�t�i`x6��Oʒ���iե+ʉQ�j�>B�,���Q}����O����O.��D�	�1��Y.$�ʅ���n�џ<�����Xlh�+ǏI'zc��(��9���?���*�1G�,�?����?��{��,�Y��qkf$:UƂD���C��œƌ�>�?M&��|�<Q4��^b1#�d* 20r�Ovc�5�6P�@�gݲE��b>c�4Xt���)�� ���q@��"$�O��d�O"��O�c>˓�?�"���Zt!@w��*}�iY7�^:�y�J����11�)]*}`��&f�0��$WX���\�M+-O�qP,8G+�-)s/̠���K1�Ȁrꐬɳ"�O����O��H������?y�OPazQ��;ZU"q0'��$�*�p�b�hi�<�6#�5���=,Ot��Eˏ�mϾ�kpj�N��=b  �X�$��*W5"ü�J7.�}X�T�/T�vƎi)�� �!B�Ae���X��d�O���:��X�O� ���/���B�jRh*���'0*��i�j��t��J7`��(M>7�i��_�a�-�8��I�O��0�OC(�D����@�� ��O���c/V���O�擼)wF�P����P��uQE� ��M��M\ 9\���A&U:��i5gX����&h(�1�����`"ݴ
�r� @�^�_A�
aNA!�x��Ɂs���O��E��Z󪉿HKm3�%[�kD�M'�8�	[���a���@�44��.V�]p��f9�Oh�	�J�5)D�>�6��Ҧ͑5ھ����'gFA���	s�1��Y�>�(�;u�����s�&D�@i1��[���)f�Ķ`S:Z�'!D��2����	�0��j��E�`���;D��*3(���r$��z(����7D���e���x����B�X�g��x�;D�����@Ÿ���D�mT�โ�O^T��)�'h�L 1�%�LH�d�����'>b1�E�D�NV����bʺ`��1i�'x�
Q���B'z��W�,C¸�@�'��4��T�OaLm�ǀ��:�Ƹ
�'� �Ō�]��[�B[�h�	�'�`�"��"1ƍ�$)�>�L	R)O:����'��`S�� _T�t��N�1�h��'2���j	��l����=)�FpP�'4rD�T�*�PV#����'���cvGV�L�p ��L^+}l�)�'?R!�P)�,� �T>��\�
�A=(��gp�K��O�n��P��q�j��9�f|3#�		|ت�+S]�(1�ȓ=��yK�ސ$&h�L�3*��}��Ub�����^�L��	ϯAj�q��'� 5�w�\9���±?04���W�:�s��*T1���I��PE{�*
��p���?u�|���@���M��"Ov�ѥ�ȞC���P�Ղk���"O��p#["�����G+fj���"O�������Z°��e.2�<�i"O�đc��^\q��)<���a"O2�	cN�X3"����$r.�r!�'��z���&�F��t`�GR���2������ȓضȳ�dڅnHb)��KX+`����Qh��qE��5���&i, �X�ȓl�h�*BL�3$f��Y���Ipa�ȓD 
�;�JD�Iް���.#�\��e*���枃���"F'\|�&l�'��Q�SCX��ȨeS��I`�K�6�\t��S�? F�Xsiܯ:�,���F�HbZy��"O��IU�M!̩����-�
E"Or�`rLE�����R�D#	T�9�"O౐�.�,v�����M�ji�'"����'�E���[^�\@��l�X��'�����!���u��`��-�'B�jE��r �1��U��h��'���V��0�)PF��s�'�YP��_�V�Ɛ!���4���'�D�A�dN�s�� ��������b��i6���%`�8wp��7��!�������n��=8����!�$�VM0A�v͚)pLe�LY��!�d�%lk��r%�N�iT��k��!���:uj�B2x�)��U6$�!�ۉaT|�
��g�<U�#,�7Uq�*��O?Qq���B�ajUX%�I9���T�<�,F?9�hTC?L����R�<�@̧F�d�%�ҕu�<bgBJ�<y$��()|̂v�W�T���Jz�<����	#n�x3&)��VVLz��A�<���_
!#�[q�6d�j:��ɅO����+��]��)rx0l���Ķ!���$-X����E=�X-$��5�!��f�n�a�֣ln���.־:�!�%'n��B�Gq]H�Q@�)j!�?�|,ĩU1cJ���A^�WL�}���~��
'J�Q`��OVx(*�k�y���U�m���V�E*� c7���y�	6egLp��Jt�n
g�ӑ�yr���¤k�ֶj���S.�8�y��.8�$��Ӌ1�p!B���y­�i=vhB$@����)mXK�ў�!�3��lE�� �iZiP7��#7����l���A�$:b�$(Yʸ��F�J��bY�t'$�!��?v�^�ȓ-[Z�r��}o
M�aù)
f�ȓ9R���JӷS�fu��
g d��a&83�e�%�����ZێD�I���"<E���:]9(h(� W.M�^�s�+a"!�D˦��d� o�"0�\�x��9p!�D�E����҉Y 1��uC�� }!򄂌Y�V�;�i��y����l#;_!�d��S���\)4���DPZ!��-k�̕�� |�rf(\ d��	�'���$+�p�B@�����-B?o�!�$���YX!ѓ�-�j���	�'M6Uz&�E`hb�3�iUQ�� 
	�'
��
T��&����A�S- ��p��'F* k��?��	���B��"�`���B�f��"Z4�n�)�c�ai�y�ȓ{��H���:y`!c]�M�ȓ��5SF��S�x� `J�3քe��hb�U��A#	w�ha�-P9G�؇ȓ �U�,F
x����R��0�����Q��qf��s�z�R�Sf=ZG{ң�+����@x��Ⱦ����юD%\���#"O�ȁ�-��F`���� �j�P��$"Ob)��m��4B�X�# ^�"3BD�E"O�=�ЋzȌ�"4�D'p�"O:عf��N؄�Y"�%��Y�"O� ;�  ,UX���ρ�N�L�yV�'���;���w� �2��:r�R�;��U�E�V9�ȓW���+���%g��8�*OS�h��S�? �t�A(���څB�r���A"O���&f�=�P�KD,قaR��Z�"O� ���J�+2�\�B�D�l�S"O�-�$�>4Ez�*��=����X��+�.�O��rb��87�!"R�H�+���á"O
��E�Uo�u�#f�'qj�"O��pk� R���V��b%l	��"OT�@UG�W��ɹ��W�)���"O��g��=W(x �ȍ���i`�'6���',r�X#�^�!i���s�U= Px�'��:S&\�n���oJ~e)C�'��u��܃&�@z�/� r��i��'�$ s �@�R���U!b�"���'��}��G��14���%��07��Q�'&����W����*Â.�������]6G�Q?�rE ��r@����<�<,�!	"D�`ô�-RHy�T+�;G�
tZO!D�8s�A�a|Pp�d��ع��>D� vF�U�<��J�@k� ��>D� (�)A�&xLs3�	
%���T�>D���s�	6�~P���@�j�X�"�O"m�D�)�'7���B���:FdDW��|��'5���+ �f�)g�.KzHdc	�'*蘀�  !�zhVn�7G����'�p!`@%O�a1N��u�B�C��(��'QdH�f�-0$��F��B��l�
�'+F%��+�',�p��єI�v�H*O`M��'*0Y�'����,|�V���<s|��'=������&8x���ɍ�0����'E>թ�h�>�Y����.6�C�'���t`��
� E����ȣ�'�,U�Ӎ�duF�[��H(~*4�������dJЍ�F�����9UA��rT�d��EH���	B�ĉ��%^�k;�M�ȓ&����!�8 � 	� =X���*S�:�@	4�9��8|
���mz�4"�'%��鳶d8�b-D�ܹ�E�Qb���D<@�6�Rtm(�^���F���2n��(��iX0.��[@���yZY��Ȣ�K�.G��Y�IJ�Y�VC�I�=�b�a""�//���
�=�2C� 1�\��(��u��L�6L=C�	ni���L�%q��SDț8�C�	4>iT��fK�'2&h�O"����
�I�"~R�mQ�* ��B��-�d��.^��yrlR'Rt�1�ˀ�Z�2ͪƤ���y��Q$1L
��p�B�B%���L�yr^�WCL�	cd�48�v�1����y	�m�=���+@�̢%ڍ�y�E��FX(��R��y}� �`H�4��2��|bI��x���(z8x����'�ybM�]B�����q~,��7Ǘ��y�UT���PFbRmlꖅ7�y��J]���HB��Z�#6��y⇄�R(ĩC3��5��ek�^��>��*�x?�Ŋܺx$tB�j?>M:���P�<i#�
Va�L�E��[츀abL�<�$Ϝy
$�����{�z����`�<є��94��f�ق>6&�"�^�<��$@�A��+7N��|	�av��n�<Is����X�g��'HD̑baWn�'F,aJ���[Y� Q���^�<��{�+ �!��M'TB:L��gT�R�.=a�	,E�!��J<V�]��Ͽ��p��(��Py
� � �N_�#1$Qb�kF7v�Y �"Oؐ触J&}E;$�U_��P$"O��2�T:%h��0l�Y�M8��'\�X�����(c���q呇��b�Ŗ0n��@�ȓMf>q9G��GrR$
�YS��ȓ>�q�'<���/�,{  0�ȓ/s.�h!E
	T �#I$@v�t��U�i��"G!3���u�ß:�p�ȓ2�������v��"��؞s�H}�'m$\����<�wI�k�x52�dG	'�C�ɏ5���4j��A%�X��ɴh�tC�ɕ9��Q�p*;7�,i�bI�o�hC�ɳS6~��B��#�x�JCD��/�JC�IBm�Y��#�5M3�i��T��,��$�f+����{��ɈTo�2�H�鈰y!�$�T��!�WꁟM��%���=yd!��T3E_|������+D،"��\#V !�䘺E/�� ņt��Y���L�*�!��z[h��7 ��T�!�Fi{~=jcf?@YP��#u�ўhxf�%�P��c A�vH��!CL5��m��lhƀ{���*x�>�s�&@����)s��x���a��]�s�D1T,��cF���G�bg]�F@S~І�+zDj<0�$�"��`Q�X�ȓ ���RÓ�})�l��$�T9���V��"<E���ܡ0���q&���Z6<=H��Q��!��6(,~)i��/ �x�G��;y!���$�a'C�
f���&�k�!��f/R$Qw֕HR^���+cv!��T�T�P�I�C7����%a��3]�@)��5�Lp����B����_���Q��D)/�N�FT4�'v�uRGc�&��pXc:*�P��Ą�t������(
�d$>{`MC�L�b��f�K�Ye:A
��;�I`D�1s�����8#��Ĉ('r}��m�&π=��Lѯ��O]q�'���V�(Ze�"-�r2��23��ay�	u���"PG	�*�X�IG36bl�g-0�O��'� ����*F�ѱ��R4��,O��@�2OH��0�3}��ƹb#bk`+��y�����y2Ǜ,2����AZ�aV��S�O2�Z=!�0�;�F�'{�Nȝ'+��|v��h kڥs��)�8mHГ�@�M�L\��@�~��ΓJ��Iٟ��䧫�䖷sJr�B�_�~Ix4�Q�U�w�!�dծG
���`� �uR(�kF�Y/�ў����iA�M��pր���VJ�nB`m6��O����'7�2(����O����O^�$к��e�*%��	�<Rx]ْ��G����.�H�[	�(wʺ���I�n00�Ɓ��W�V@СHhUXPkr��ڟTc��+�����!)FxR�ͰR���5)0q@����d�7jS��'Sr��h>� ���� �+lN���'�!���BB9j'a�C=�A �?���+��|�����U�1��*�#I%R�q�'�����@�@W)9��D�O����Od�;�?�����f�nגe0Qh�@H�@&M+*��Qp�.]/ ��(��S��	Ó^���y��"e��@
�U��l�T�J�W1 L`-G=���2���{���A�O��P&�8lҹ��F[Y Ř��O��d=��z�O��㡠	�f��� 
n����"O � b���c�ѓ�Ȗ}�db1^��C�4�?�.OL0�nB�T�'��	�-m����q��],�QE��-���J V��'tC6W!r��ˀ{]�ק��%3�F����52A�hE��O���GR3c�Lؔ��{�SS�d�"�02�H��UPR�#>1Q*Vş��J�'b4���Kj�����M�{R��'[a~��^��\��)ݏ~ޜ@W��>��Z��b�(ܞ&.�ܠ2���,
X%	�d�<9%��&�?i��?�.�z�	���OD�$�<kk��5��6}hP��Uǘ�$T���)g��Ԣ�Ĉ2K8NAA��[bdz�O)1����DOW��}�F⊢"���V>O����S�|Kb�B ��o�n�Aש�A�Ok��렩��[�
y�3閿
uX���'�<���?9�O�O�)� ~���a�u�4�yB�/r4�7"O�����N(�Z��4)T�&�I��ȟv��b�N.�
+�$�v�P����[%V٠���O���w+Y�E�d���O��D�OR�i�O�蒱�V���s�
� u(����
�){���(տ7�2�{Qe��fj�'H�O�Q�HɉE�ly��_�E�0��5fR;�f��)чv.mZ5�O|�����'e0� ���Vؼp����8-�^���O�u��'hr�I�<��ǔ�d�@,��=$�1�+�T�<��ɻ-�؈$�%u��hAmYԟ@ ��4���D�<&�vU�I0!�A%N�ܹ��I	#`�5A�-�j=�1��?��PT��O���a>̀��Y2lQ�"��w���R�De��� H��i�m$��ٰ<��^o}����9��tp6(W�J1����.��Y_�
Î T�ay��]��?!�m�FnD�S�ԗv�&�q�c��?�����'��>���*�r�a:]��x����z�<��eٸf��4�"C4F��q�My"�uӢ�d�<��FY����ӟ4�'غh��Q/P
6�p��9���>@"���ڟ\��.�RLzǄ�0c*�-`c��$XV�c���%�T��d]���Ҩ6"z�	&tǶ-{1��[4��C�B��J_w @ q���7�pu���J�B`���� 	��'@1�r���	�y��d�j
pi��_����I�L����O�f�v���#TV���d�\yr��)4����ɐ�9j�䁂��D�O`���O��?��'�� �$Ll�x����&�2��hO"4���0AnA!��7Z�j��d \��'#��ұ�t�Ӕz���ɦA��>���摟 ��'��I���<Ѱ���Ϛ��q�S�|�Yp(�w�p@ �Op�OP0cR�>!Ԙ���?>D �#ALI�zt(DPRC�%լ�O���h��d:����p�ۢu�mq�ǉ$eê��c�>�r�>�+r��R}�dgQ�dې,޾s�7�
�?�@��I����8��?qp�ߴ	��!�K��NR�I�MH�P� A4}�&}������	�M�vj\�������6��Y��cPSy�Gٞ��	��ȟt�!� ���x�a�=0<��$Fd?u��g�T>片w?�����x!Aظ��`��{i��'*��-�I?z��ʉ���Oa��	+� Vw���M@�R�U��q�$��'i�S��'<�ȣ�'+x�	��q�����ژR6���"�������G+�H���/zh���.B!�$�7&1�)�<p9!��PV�v�'��'�(�g~P>7�����1Z�CO ���%.��?��	[�]����S�*Zr��0ꄊ�����!�䈍RXU9R�c���EA�2:�!�G&`������M��J���*+�!�ʅ2�f�Y�K��`�r�=�!�$��ܬS�!�W�C�D�/!�d��֬%����q߸Xh'N�"5$!�۶h1V�yцh��P���>#!�䛕^�Y�e�_ 3���`�-ҏo8!�Dɹ62�B�ˆ;C���C�!�Ć�X�zd��gĮuW$���L�A�!�d��I�2�ChĵV�I��)�!�dß;"�P��K� h�%#�B$n�!�H'a&��SfP�?��]�f!�� ��O.,�Q��F�d�M#yo��#Dl���i1 ��20�(Q���͟5d:M��MD��c������'�!�����$�������ʭqJK#� 9"!�S������9l&�%��ʁZT@J0�4상�P�7(�(���4|qN|��hL�%��&�(Ӗ��x�^�K�a��j��eB�4D���'�N=pg|1Ҳ��	����4D� �m:N��ۗL&K�IJuA0D�̈¢���
C"ٕ���`��.D� ��;�t)a��Vz�3�:D��Qr`�z�4��"��Ĉ��8D��:�BX�J��N�!}*��G�8D��(E�Uw^ 
pjޫ4HX���6D���BᘞQ?ƌ0�F׀@���e+4D�Hk�!
�A���b��i%��i3D�`(`W#m��s���T18�S,>D��AT�s�t �D 	!2pC�.D��B�̀�- p�a3��W'Y�L�!�� �ԂsG�4TR�|��ۀS=D��"OT�6�]M���1�Z�q$$qa�"OF<���ӃVq�ݒ��6.j��"Oȑq��=����,#?>�A�"O���#��(8�ıZ�����\z�"O΀�4��+l�X��OŜ�nȰS"O���ff�!*"(V	o��p�"O�ӒOUD�~��`�,Τͩ3"O�5�d���R�@��+���"O<er���
�J1PҀ�C���"O����Ψ	�y����~��g"O^�+��Q<y�����G�<;d"O��#��{��QQ�"08����"O~�"�nC������u+�Ȁ�"O��h�*��A�^�k櫆�>��I�"O���w��;��#'
J�Ij�a;U"OV �wJZ�[�*=a��S�<_�AJ�"ODM�Q��,��J
4Ȝ�"O�M�&	(t���!�J��B�"O:ez�A	�&}��B��C�Su"O�=;a�޷}z�y��L�>�aC"O�M��dȠh�j���^�se:���"O�D��oϠw��� �,��r"O�<AG�T�*c"����ؓ
�f�g"OF���Ff"d�a`.�	S~ʵ[b"O���#J�xO%q�
�yhx��d"O��5ܜ�x�B�C+xh�0"OT ��莎`�,a��i.���"O�S�K�,C6L����O�m`�,sE"OJq)�@�>B!Ι
���-tm�ݹ@"O6T�#�N�Jڲ��RL	yv"O���J�?� �$F�%<<���"OR 	Q+�B���E�>\�z�"O~�DQ�i��,���K	8R�Q�"O.�9��ko�x �@]��!S"OF�0S#߲x���{���:鰅��"O&����T1ZŢ�YFŗ"�P�Z�"O I�A�=4���e�^��a�"O-���c�ʔҲf˥cI�u"O�-��h��4���&��}4���"O�5 ��δ89t�K�o�R���A"O�	 �#.�r�smɇ1>��&*O�}�T�ܻoL��Ri9n��S�'3�%�c���$l"�Ӻ4[�D��'�tt*T��+I�B4�0`�B7D�|�S+R���Ŝ��$RG�5D��ó�B�@�V D�%dVt[ע2D��Z�ɶ>e��B����*Ъć%D�����ʊɤ����=P-�=�Ɗ=D�({e��"0�OZ�@I�ݫg�8D����
�!R�X�J׉
n���$�3D�4rCB$+uИ��LU;/��$Pl2D� K���0�iA)�,>�����1D�2�V;�*-cQd�
�<�)1f0D��c���=j~e�Bw}l��蟞�yr��_:z�{ �M]4<8ê���yR��2�٠u��B��p@�-���y���%�Ɖֵ2�p���6�yB�'^�d	�fI�1Lj�X�M�y�凵#sV�#�hA#+KFѨGh���y�m݈UvV��J[V2�`�M��y� QL�l۲�Дz�v��"	���y�I� j��5�%�J`h�)�-V��y�ɟu���P'N�U�̐���]��y
� j$y4��r�(�i�T% a"OaI�o�5gT�7�8t#Ҽ�D"O�:���_����0	E�>��2"OdpZB�:���c�(סD�@"O$�٧k
���a� "�m{s"O�U���C�=� �B��ۗ����"OT �ԍSE�F1�P�{0ؒ�"O�;�
C����RՀ"
��)�"Oh��ц́=!Zy��@���
AA3"O�D�q�
s�u��/�(g�X0y6"O��Is���D.A�a����"O�	8u^�]A;�,NW�> `"ON��Ɇ�F���V,�6���(�"O(yQ�-@�dY(4RǫB�0����"O0�Y#�P�,T����Z��ޤ�H�<1��҆rے0���3<�1��,N|�<�$��� ��C�č
e����NC�<Y4�џq��5+2���/��S��Vj�<�4� ��0/�?dg�a�"��d�<���)��K��g��Д+`�<�jU3J�b<1��ɱ8渹��C[�<�����.��=)Ea�8ke%���Q_�<ypc��Z-$�"��ĞI��icŇ�Z�<��͈[ڂ "jЛ7]� �m@[�<I'��	�xG�H�t��$@��GT�<�p�]Xs�U�ǡ>I��}�V��v�<��T1��)�d�:;�9ks	�I�<QQ`օ.y�0�� V�j��7ͅJ�<��$�>	��c�lG�,��2P�l�<��3'�T` �@E7�����,�]�<��/4?0�1CW ۄM.�b
�\�<���_1X�j��[�&A��� Gs�<��ӫ!��'K�r���r�n�<��B�9U�$iW��k�d3��i�<wAQ{	��BL�������b�<Y��_5E��pAR�^��##�\�<iC-�D�<+B��-$�!L
W�<��kF�Fx�`��b�0�<�˰�Yh�<I���?�M $f��$J#�a�<�/��qx6�[�#��v���9uO�_�<�4�Zs_v�Y�(W�Dg��'
P]�<�sHQ���v�x��_�<sL]<��%�3F�č��a]�<�4t��vɛ;Di"�;�ADW�<	Q�K7Ͳ�e�40��2S.�x�<ic �kj2,
RH�� #"��3�L�<���'S�^�iA��* 〉�D"N�<!�N�r��h	){�pA�Q�AG�<D�ҳ	�֘z"C�;/�x�ƌZ@�<Y#�:O4hA��݆O�u����<Q�!�)@D>��5S��B���
S�<ѳn��_�@E{p%_9r��-�Hg�<�M�� % a6aɩ2XT�Y��~�<�ǁ�=g� s%�p�f���}�<�v��1�M�6dR�8����&	|�<���C�z��Y���>Ⱦ�Y�z�<��O2!�0p �D�0*��|�A�L�<�2	Э7cb��Q+�0L	8�0�h�G�<#�A�^N�9fd��HC�bOJ�<�ւ�2i��
Q��G(���Ԩ�H�<dm�3n	��'��RnJxX� �B�<��%#̠��uCԝ6��/aeFB��5/�]A#"��d�<C�(6f�^C�*8$"X�f�Q
s����,X�6C�)� (l	�Uqʦ�K�%_�1	�A"O�塢���9n��1��(��K�"O�Ȋ�g�7I�̡�×N��pڄ"Ov0*�ˏ1|���7��F�����"O� BK)5Lt�J�]�y"OV�2ĉ�]-u	��*'N`�%"Ol)CeE��D+1�'4=.�j"O|ha ��_�V�3]��ۢ�Њ?!�dϭ%e�0�*��:��aܬ}!�$=Pڊ�3iD7!ܰ*`�W�k�!�$�%��	�F��I�ިx�dD&o!�dPhݰɸ�#� =�Ȅ��$!�D��hq�K��y���e�!�$1,���*S���t���¦�B3h�!�;kr����X(^��k��U��!���
W^��[`·�`\�2r"��!�DC���X��G�Y�P�`�`�!��/u4EY߈Omn��S�7ZC�	��,l��*�����5m�Au`B�7��l��U<EZ���d�YbB�	�N-�����:c��HÂK[7)`B��Q���1��	:�ȓW)�c>NB䉝�޹h�d�7}�p��R��^��C�	<p�:�)�(�@�j +Ցlu�B�ɻ0|��g�ѭ,	(�!�aN:k�
C�ɏd���0�Єe���9qB�A��B�	3^�
��F�Y�{�{�L���B�I8{�� t�W'h�����A Al~B�5}�T��ɝJ2�J� ��-,`B�	.g'�1��cJ�j1�TK4�?V\nB�	f�v�1��ވK����SeA��TB�I9q�8�e�!h�lp��oDn<B�8�Y�E�G-�h,��i�5�B�I�r�U��m��e�u�O��C��?WѴ���=0���h���;Yn^C�#;��b/�?8�Q�Q�^�I|C�ɡ@�����4fUЁ�rVC�	>:��0;�j��G�"����;�C�I�VnjT��%ΏQ�P�+q,L �C䉹 ��I�Y�)�$�ۓA��d��B�ɂO͐xk��s
�Q;�*Jk�B�ɧ�Ψ�So�:"�`�� ��B䉿�r���=:��́we5�B�Ia�j� ����t���H!+�
��B�ɀq��Ȑ�'�'ʜ���FS�B�)Nl<sE����@%j�X��B�ɮ,�8LzsF�O�\�)E/��B�I8(�")���:u�.!a�0&|B�I;3w~�  Ȑ�=0�کiKzB�	)���2��4(%ܸ��G�B\tB�I%Y��R���V/�U81��kcB�I:8�H8c��/�����˂�mc�B�ɫ]�L�9U�F�8Ĵȡ�
�Gq�B�)|��WǊ��B4�0�V")��B䉅$�p1rK�����d��/&JB�	X�l��iW� 
�J�	�B�IEJ�=�U��'FL�� �$�"$EV�u�B(S��I�2����0���\N�ZQoB�v�D82�B�/4d!� �8LRp'�]?R�ʔސ1D!򤘂M�bL�� U�]h0;@��>`�!�/[oDH�b�<O~9��a�=�!�D�_�X �q�]M�bA!��`�!��J$kr
���	�&�r�&�G��!�$�E�
�	�cѢq�$D����c�!�� PL*GY�(h����ɖnu��`6"O�!���&�h��R�XU���"Ot�f-��~=�4��.Tm+X�@�"Oh�aTB
J�����8$��4"O�p�˫hh�`� �֯)-�i�"O�ZUAw�ڼYS�,(|�"�"O4[��QqsD��؂>w� �"O8h6G�?d��(���mj�i��"O:�{�AP2NHbL���F0fPBHrs"O�(�S�J���a�� '��+�"O<�3���?c��,#��"Nih���"O����dɺ<�8�H�LZ�=�%"OZ��AU�N�ll�HJ�zH0��"O�!�R$B!B:� �3�����E"O�̰2�A�w��X 
W �d�+%"O�P�G��Y9�i�2�Z}"O�с�/�?��3�n�q*��B�"O6�X�kZ�n3�Y�����z&����"O4`[wD<C�D}��m�&K�y�1"O ��։�.{���gG��t%8"O�M�ckN�9Xv)��%D'6e�M��"Or�[�O߻NÒ��5EV�3ü ��"O� ��IU4nQ)���X7��u"Ot���_rU�yBd�^�&�(�p"O�(#�U 63�$���	,x.�o.D��@�fN�#�r���y��*v	:D� !�c, l��%,�2C�Ь�f5D����M�cCt9ç'u��*�>D��e杉
��!��ݨ4�R�!D�D`���C[�`�7�O^ʵ뤇2D������o�tx�lDo���x&D��sS.�?@
9կOe)�dE/D�4��i�s3ʐ����=���4�+D����B� ��D�ƻ~[i"+D����j�D{�ȟ7}�$k��*D����R�/,�R�(ޓK����H)D��ɷ��7|f�Ia���[+D�$)T�5Ri�u�ņ��}�f5� -3D�����"w�(�`0�G� �����A?D��j3����,��*�#)��Dr#�=D��9"�4k�<�Y��IY�p�A:D�$��߽-��0[O�%R_l��6D������P�Z�1r��#{4�w(8D�̒�(K�WK� D�ڡa��9ħ%D��@ �G;�՘�
Y'ь! ($D��J悃l2Phu(��|�R��%�-D�p)ǅ��`1��a�L��4�RPA)D�0�$F|��NӀ8t`:D�(D�pf�,k�tT�Ф!z 0�D�(D�@q� %*a�I�q�&��0���:D��3� ��?������^�I2�P+e=D��q@%�H�\��G܈Qä���:D���ݜ:-����^=�����$�y�$�3�r� An�n����Be
��y�c�'lu
�;�E��p�N`�RMӘ�y��^�T��uP�A�'h����u+�y2c�=�� (��_/uL�Z����y�L4`LI��ř-ZdrdO��y���3��`���:�bm�Wg�o�<�1+�>z��RrI4,�^����J�<���e�L��LY,h�K1BN}�<yBeec��� Kh�ň��X$�y�� 5�CHO�D�<h��c��y��РRtp��@�>{r��2i]=�y
� 5XGB$v�4�:@�O�OF�=&"O8
eL�.:�������p���!"O 8+e
�WDҝ­�!�J�ʲ"OΥ� ���#R<躓���4�
�3"OPm{���t%B��囹C����"O� �$�ڤ:;�5�.�J@V"O�52Pj��@Xj�'P!�D܀V"O@(q�f���0�ݠ8���g"On(8���)>�X8	2얙l�"��"Of�Q��$⚱x0#�p��P�"O��9�h	<Khx*�a�&G� �k�"O2!��;|�(�0�ֻF��ɰ"O��z�F�6.�����2��lk�"O��Ǝ	 m�|XT���A���V"OB���Ha����L]Cq���"OL(�Ȟ�U`��"邔g�(h%"O\z�@45!֕��#:�j�Q�"O`�@��1�yC���O3̱�"O��	,I=��Rs��0'�A"O�,"SoO�sC�\���*Ƅ��"Ol��CE\8��=*ѩd�D�z�E2D��k�9^b^:@�
6,
y��`>D�h�'N�;i��M�7 �<yR�A�?D��aɌ@*��6�I�S\"� 2
8D��@q��'>3tP!U�Q�`!����L�<���\�V�DYJ�b̰<F�:A��@�<�����L����0j,��q�Y�<���_�E��!��w&���@��M�<!"Z�Bf��af�0
V	xEI�q�<��E !;uJ� �垉���iǬ�r�<�QR�5̸Ro�ǆ\	�-�O�<ץ�'JB�*F7Np-�tHN�<�kE�%��YPpꏰ@�T���G�<a���#���5��	<��P-H{�<Q�)Q: �i�f���Б��g�R�<���5�
�8'�Z^K ��3�VH�<Q��N�\��� b-��%>��3�G�<y�G���-IG�P�#�hdS���i�<�IW8Ҥl۲�UIɈu#Ai�<���
X���PoN�mcx �n�<I�e0 �{�*��j�42�LE�<�S�V���ԢcA. � %"fƗ_�<� ���J�D`[A�8� ZӁ�D�<)��D�w�pɣ��]
d�!��@�<� ����Z��s�ę2u�a�<��S�S�H�12�Y�D/V"b�E�<Y�mܚ~�<���H�Tcv�+2)^�<�p��egR�C�I��� ��\�<�G��'|��T��<H}�ɻ���o�<���H�b\���'�Y kd�+U�f�<�FjT	~�h%���>#`5����~�<)�o�3z6j"�B��S�b�p`B�z�<	"烀5�X���Q�L���'��u�<��%ī(��ѡǷQ��):7�Vp�<�25r���Ve³g<8�K�<9gG�f��`��(��>	��E&Gp�<	����͊b��kD��Y�
�Q�<9 �<A}�qh�a�d��qGH�<�f��,yr�0�f�Uy���n�<� $�'�����ϼ{@��"�g�<)����x��gR�4"�4�K�<�1(�~�htjB�"�:!����J�<��F��5��
�x s��TH�<���^�S�q��1`�ebMH�<� C�K��m?�1��C�z�|��"O��xuG�1B���7H�#r��ؖ"O���ŏ�X`8 2�':���8"O��+�.QށF-R�X�p8�"O�p�@��->=��Ð�gV�t��"Oha$lT3��iY1�K�B@���"O�x2�V��������u�"Oh$�f�Y��4h
��]�&����"O,X��X4h��]�EB݄}�ʨ�c"O�Q	�`ۨm�x1��Q/-��x "ON�2AL��q��D��'P�y
"�`q"O�5i�F�/a���Y"xޔ��"O� wi
�(���;��7kor���"O�4���_-ae�M%�\ 8��"O�m���	�e� ��\���"O�H���]�����Vp�b1"Of9�CG�{���y�ܲzO�1�6"O@e�0���Y��Y�fg[��r,��"Onݸ�Jֳ�b0�D�,t�`�b"O�L��iS	Wx��㡤�!L����"Op���� beV��k��64r"O������v�=���R)����U"OB0z��<71��a�(;���7"O�E�À{;���0O��v����P"O����SN��]��L&�$<¥"O�����2\7P�p̈́-P3��S�"Ov���FW&~ߤ��C�#Ӕ��v"OZ�j�'�T���¤ǒ/7~-�"Oj��D�6窐�qğ\ūv"O�m�G*ԿR%���v =��iU"Oj��:~�n�2a ԯ^V��"O�]��
�;7�����S�-I�iۤ"O�P�lU�!I�4x�"C�̠��"O����8.�C�@H��ZUs�"O=K4iM�	�zG.�&���P�"Oxa��̓���s��k�r�q"O*�x'�`)v�v�!Zܲ���"O���j��q���5�A��H��"O��ՄK�[Р�������P"O�K@���ұcŁ�`�L�hc"O05��Ax2H13�R��0m@�"OJءqc�(�m���$��ӡ"O@�Ռ�
J��ad�/���Q�"O҉A*¦A���(��A��E��"O,�A��r(}ؐ�׋� �;�"O�91�߹4!4yK�b�*:Y�=��"O�q3Δ"�ʑ`f�����;r"O�=RSIΕRB#�CR��Lir"Od��l�Y�3�hU�]Ĵ�+t"O,�i���Uw�s`�Ȓ/�l�"O�M�6���S�L��󋅪|��	0"O�M�F)z!�M̓D�:�qT!�2d�!��ν.�(����ڟ2��I+4A϶]�!�ܶ2y�Ǐ�iZ9S�B�;�!�d?c��	�q��9:�6 ����&�!�˞)�d� ��G�4r(-`E{+!�D@�G��(��	�L����]�!���C�$L�a,öbM�(�a�BT�!�)��`B��O��M!0�̥`!�DY�k�"تǎ�r��)Xj�F�!�D��:&�:E��5�r'�>�qO����
@r��1��9r��S�|�hݲ1����i�7�"8x ����y��	̩�	�2px��L;�y"�g��1��Z2#���;��R5�y
� �bS�jXĐ�#�׹�(@!"O��)�@�9?"!ZB�ӭ!�l�!"O���Db8
���ѫ��ͤ�"OP��w�F�VX4��C�O�!Tj�8�"O,:��<$����		_^�0�"O�\;�J["`�>]�6
vJ�}:v"O�$B��-:� 	��O�Y�@�ys"ORUPH9Z,�"��"8�0"O(���Z�A�!��8Q�j��"OX��G��83��1/}6��`"O|�swƜ�>��	���!_ԍy�"Oj�qMG >�	�q-Ө}X����"OR��P��@*���
I�YF"O��ڦ��	2<2��ߚS,�2F"O��p�_v�V]�OA�N�v��"O��"UA�(g�1�����aL��Y�"OB�J�jN[�j�x��SQ�i�G"O)�t�(�l��/ڥ>L�Ыc"Oʌxଋ�t�4���.V�&L�"O*TS��țs�P���M�N8Ep"O�U��/ҡDX����!�4�RK.D�D�"H3o�݉c�^�0�\�$�9D���c΍*O񒬐��Bpp*�N,D��(�
Ų�xё��<U�,l��*0D� ��P3{�2��G�G)x�0D���ƇU�G���6`ō\���C�N,D�D�s�/2v��U��2:5�E�%D�H��bY�#n���&P>h�1��b#D�`q�űp����K�!s�(#D�tB�BC(&�5�3ę�}G~�`� D���d�����3|�d�P$=D�٠ڵO� �Ã��c*2�5.D�����,+��%;d%ϟj�QC,D�8sdă�){@�$O�8J��cS$=D�`��%S�Ej���3�X��h*;D��Qd�xY;�`I}���/#D�X��ߎ;ͨѤ�J�iߢ�"S�?D������&��˄�2JԵ���)D�X0e�C�2F�0�8-E^���N5D���afߨAP|x B�4k�dujF	(D�@0@�V(E혠�V�V/=����!%T�d�WȞ,β]aj�;<攱C"O��XdAӸf���;ↂ��T��e"O��
�=�Mib�ؙ<��A U"O�Ը.�		YVeȻeQn�z�"O�1���	P�6|9r�{=� �'"OH����2e�&����.%��W"O-�6%]���D�Y$B<�Y@$��X�<9�D[���ׯ�#?~q �n�V�<ɦ�A�ΐ �iC�_>�pd�w�<�t�/8�da�"&JD�>��Ƭ�s�<�sC�>SVa��ț^גI����U�<���>]>�ӑ��azT�UD�N�<9�NAu�BIy�.ӕD�0�d�K�<�hɂVx&p� ��K��+��O�<iR Uyd�С
� �f��P�L�<��ъ�D�1 �<�R=���F�<�v����ɗ�ߍiv��w �@�<��AO�sh|��� w�p\�ƦYb�<qV�`M�d� ���>S"ng�<)Vfʁ0p!C�D�Gq��2�l^�<!���:LG�xeGA�o;ڼ��ƎX�<�R������u���r������kM����KӚ �Ti`���;H��=��S�? jX�e�f��H�`�Fr�K�"O:�J'�z�-*e�L5s0<��"Or�˖ ��vT`�9 ��:$:4(:�"O�z1e�(cȰ8�� �*?��"O.Y��F�Z�\��һ%v���"O�u#�"]$rxd0	N�U<(��"O�	�dmM.~4��:\hT�r"O�hB��D5��	 F�|
Z���'���r@L�`L꼐�F�Oa��'����L�\��D#L�l��	�'�p:D�[���j�*��1)���	�'a`i�c͍�Ed@$;�e��~ۜ���'Q��ٶn� j�@�-�z�ܸ�'̰(��FA�k�8D�䊈�s�i��'L�0�f��g�J(p�'��:����'����W��J��+�@ 0z�4�
�'�, ����X^�9�P�č#lq9
�'�h�b�
�D��((㉜"�t��'��mr�C�y�6U�f��=0y ��'BΉ��@+ux6�*&뇯�6IK�'�F�ekS9?wĭ��H[�aSl���'�Tm!s�W�Y'vmPF�>U�M!�'Dq)��2Y�\�%�H�LLd���'ٴ��W�S��0��+�71/��Q�'�X(��f �r�#W�˒(�V��'�Z���.I P>�(dX=!�ЕB
�'�p���/	�d.6���ӟc���	�'�b��U��"���/ܾ#��t9	�'VDrǂ��6���Y��sȘ�r�'�P�	"��|)4ِ$�=��]�'�� ����1*�t��c ������'��ĎݖM�lĪ'L$u2��q�'BrĈ�-A)hfy�#���3�'�X�Q�+K��C�J_�j��'Ȣ����HS2I�陒R�Е��'z���}d&�R��	b�0 ��'���7`ՠeǼ��g�9*�ظ��'��p �C�k�*���Q5 $B�'�2Ũ� F�=�(��elCk��Y	�'<�-ɦ~�Phu�M�z�~ur�'�b�@��) x�<�3�ǎgF���'�`��M���q��_��a��'�R���瑜\Q���)M�dm�D�'�4��|�t�XB�����.O�!�B.Q�F�a�+ߏ]C�uY��Tm!�$W���(`�F��3�.�RC	�!��ӻ>����W G�A���	B�bt!��M�@�㠀B9֬I�N,a!�$�Vef���D��M�d+n��B�ɚ�H,��@#�2����G�i�`B�I�GX���Q^
K@�ƻd:^B�ImV�`t4r��E#
(B䉢L�>��r�Y�JBB�B���)ݰB�ɏ'��I�H�v�ĉ��LW&��B䉩k���ˆn�%�1��픪QF�B�X�&,
х��so�Z�R?�B�	�k �� ΐ>��у��T)aN�C�N�jq% 1q�v :�'��P�C�I�b$���S�r�R���"~H�C�	_�%��,Y>ej�� 4鉮	���)ړ�v��w-S�����G��޽��k3`(�ᇀj�r�q���� L�ȓ^���l� B4�Q�D�U��lvXC���,h�T�c��LɆ�S�? 84(��Wv�l`�#��1�I�"ORQ��.�w>����T�"Op��Q�b���8�^s�6ls�"O��R�/ŧ-˒��/X;D�6���"O���*�nh�h"�G�{`���"OTT#1�YT��,
� L��"O&m" �i�)����_�
؊�"Ob�2�C�X� '�;D9T��"On5Z1��#M^���MFnJ�!�"Odm�e�O 7����4��3&1�"O�9���r)TC���<c���#&"O����f�;,,"�D+?v��!4"OLu���֯>�8Q �T*����"O����H�K�D�7_��js��`�<���N=O�x4eT�B��Q�TG`�<	�bYC�����	��%'�b2�X�<��Ɏ�g�j0 G�Y�#5�8q5� T��x��U$Xb�  a�do�ᢂ�(D���DXU�i�èՠab��+(D�,�uf�
o��@�ҽ(��es�
(D�h�2/�T_0�ui�9Cy�M�q�9D�0�#斲��Q�MJX\1�D�"D�x�'x��i�A��3,�(��"D���s�p��P���TE�\�!�5D���'ϊ$�
�$�k1��8q�4D�䒁�u���HE��mhZ<�C�6D���7��$��Z$h	9n?�Y"s�9D�ZgL��T�� �-����}���5D��zc���1lZ0�dA47�ba2D�4BѬ�%INJ�I�e]�q�L���1D�Hb�j�(*e�d%�"g,a1D���!j�&*dD��j�T.��pF0D���c���%E>��1!����E�dB/D���Iɢ1��F�	�<}"�D�!D���T+��e����Eۗ_�ͺ D�|p%١M�JpY�3�N���#9D����C�5<-is��Ԉ�Ä2D�0�W[ 9#�9����c0D�x�e�#~�!�	��W$�� $#D� ���?�^��FŔ��br�<D��V�&Oʥ`�lP���<D�����W	��B`�nY)rG;D�`Bp�M+JN��§Ĝ�L��)Ua:D�x��)��43�5�c�� h 9��(+D�	�㑺�v�Qun_%1�&XCGk4D��CR<�1��>����1D��7M��_���v��7���k��<D��r��ݯ<cL��!ZbI�3�;D�����_�U=<����Ҕ'�|<�f>D���c`مY$�r����-Jhb�k'D��{��
cZL	rcLZ�#�PK�&D��Ư,�LU����(B��!k��*D��@oT'6`�������w�%ᓠ'D���@ߏ.@��4Km�f��&D�L�u��7p%@]âI��D7�Ҥ�.D��r�ND3w=6p�L<g���Va,D��N-C�2X�A2N��EK��)D��@���/���%�9[�\���3D�\��C���p`��ilVx�0�6D����ʬv4z�A�$�(8	8��6D��S7"�/8߾�K�ϲT�`��Um4D���2aX�@I��/�U�$lj�.3D��� q/ �8�
��AI��i�+3D��5
�"##>��@�
=��U�6�>D�� ��X���GL�{g�P4�TxI"OhABC!ʬ4�0+6I�%�X�9E"O�����sR,I���Q�S��\�"O�X���NJ�ԡ�H܂]�P��"O���hӹ'ٜ��&^��P�R"O�([�J��hY�ާ2�HRC"O�13�ݑ$w�ܺ�%O�cz���"O�l���Рis<Tcu��1.���"O�,js�Blr��c��
[ifd��"O�-Y��#'("�b�E[��N�a"O�q�� �7ufp�$��>dQUi&"O�$��c�l�r�Ň�J+�ɸ"OʰJP���0r�Z�$��D"O^8(h8(�H-�d
y����"O�s�N�L���0L�oF��Ф"OX85'%����*F�h��"O�{�'A�T�a)� d���"O�y�Q)[3;dIS��-xr�`�"O�E��DK��2m��I�I\�в"OD��*E)<���B�$�]7�!�"O�T�SD u��)Kp���A4x�#�"O���f��A�!
Y��u"O����c��+��(H6˃A�6���"OD�Q 
�.A�b��%c��P�"O
1y$F؅TY֘栆a���%"O�P����J*�Q�5>�8���"O��#f\튣'��"�D<�NC�<�옆3����G�$
��)eNW�<Q�,��5�t �"H�h	%�R�<�&�]�)Ef����w�6���@V�<��-�s���¤��L���r���O�<�Q�;"��0����=��$��R�<�����YF��E/	_9�13��d�<��␁�.E�i�	�2��4AY�<�ߋ{���`0�c�a�cNK�<����
���+u��Jt�}��'�B�<��CO)SU�y�'?�襹���@�<y2��>��hd��<H!\����}�<���]�]j�iJ���[�:���HR�<�BR�8�
t���n[L����U�<�!�?p�QXDCx�ХQ�<9R@M�v=r	r��#IrT�DKMJ�<�d�:%a�1 sH�:��-����D�<��lH$nejl���-�j S���}�<q�Gӓ]��A��eߊw;�+��OR�<y�ş{�x�Ǡσ@����Ys�<Y�Ø,��XS@�� t`�-�$
{�<108��TJ�ۤc'F�ÒM�u�<9&ƅ��x�$gZ�a]� �Bu�<�a�d��'T�"�����u�<�qi��G���S�Y�9�<x���Y�<qv�L%d��;"���P)�f�S�<Y6�D p[0�Z�s_� 5)�C�<�Ħ#3�n]�֫C�[��0�΋~�<)$jՅkRdr3��� ����2`�A�<!qI ��R�����(c����i�<y� �S� �X��*,��1�o�a�<�n���=�0�$jbh)�Pa�<��[;U��YY1 l��MIE�<��[7u������:<��A	6��F�<�æ4JS*MK1Hĳ�lԸ��IC�<a�/�Z�
P�S@�V�4�H�JQA�<A'D�
`��h{�i0Wy�&g�z�<�Z�C ����a�)C�YX L_�<� <șԂM&@����!�	�E���3"O�ͩ��+w/脒2��V�pYC"OtU0��rg2h4�^*�eX4"O�-hQ��u�l���ՐY�-�@"O��#b��j�^�B�-Пn���A�"OT8#��s��ZM��n���`"O�����7����+��lv:TC"O6Pb� ��F�jأ K�`,�R "OȤ{��h �(�$Ɉc'�0��"O�y℄�3Vb�����<���F"O�uX�-X?<�e:D��4����"O�v�϶;��,���]&�<�RG"Opi��fYNR��;��ҥ%�\t20"O�,	�cD�Pr
C�g�J�ف"O���&�-{�j�\6u�h��"O�(�S��!(�J��)�t� 6"O�0�E
@����C;�R,q�"O�\I�Ė}��8��X�"��f"OP�!S��{�X�����dS2"O�j�l�Fn �"���[o���s"O���Ű�$-�e U��Ad�u�"One�b�Rc�b}	 �ܖ*R|��T"O��#$��2�50ÅG� +Zݳ�"O��xT��$s�T��@$�6-h\ȵ"O(Q��j3�+��^
��d"O�h���^!��A6�<�F���"O�����84�PbT\T��4�"OD�ri*mc��i���p�
"O�X�ΛsR��p,�&Lf�}�Q"O�X/ݷlӊL�a)I+l�`)�"OR()��P<Hi~a���;�
Lҳ"O,���K�+��I�DZ�>ɒ���"ONPR��"	�
�h@l���B���"O(��c#�;Q#�XQ2��~�v�`�"O��a��$
�B��� ?�A�"O��$Oa���SiN� $ڡ�4"O$�"%i�����F�?�-�#"O���G!R4j�!��4�T���"OB� 2�F1�811��IC�"OK�����H!*������Ȩ�y�L��7&F=3 ��4-�Փ`Iډ�yb�$)U����G�	��#����y�(JBI&��-��jn�2�̈��y"!�)�di�I2s�5���yrIȨƜ���F

&j�p���yR �L�������"}�(e���yb ��+���/��FD `� ��y"g�{�X����1*#����y�䌀X��a+sF5`����!�y"`ԶH����ك,8� 2� �y⪈�m<D�r�GG�?B2�+�%Ϋ�yb�B8g�Z�;Сǘ:��!m@��yB�ƐZ\8TЃ��4V.�p$��yb�?{�4Q��F�0��ѹ����y"iV�	&��Uo�9t�LH�#bC<�yR�4lO.��c���mߊ��h��y"K,�|�PiލRJ�,�	���yb�A
[���� _L�(�2���y�GW��d!���.~�Hg��y�KUb��L�B�ԏH���Ԡ�yB�X��P=���KX�pc$n"�yŭ}f��c�CV�8�b�'�yRŊ%���7&W<q��x��jZ��yR��&�(��W�dz��CL�4�y
� pQ!P(�Y�$%Z�l�"O*�zF@S�"��炚?9w��!"O蝛�� x�HdPV!	/��� D"O���)H��
$"���@l�رu"O �z�� f����({]��@"O��A�T���⠓�0O��b6"O���Ç�z����W�R�10*G"O��r���s@�R��u���"O�y�#�V	o�XIX�E�2=����G"O0��C!�ws�p��V'l�c2"O�)i3i��!kȂ¡�q��LP"OFWJG��ڸ�+�) ʊ��"O:@ O�5Wh���H�V��i��"O��ӀK�p�0�ԻqAZU"O���`�7�°��ؚ.�F(9�"OFY��,X ���e�-��À"Oh�pӠ�Dm�aب���IR"O����B6W>���%�u�vP;%"O II�$G4f8<	Z��S.aܤ;e"OJM���ބ<���wĆlX�s�"O��(F�U�=�0a��c�-R_4�#g"O�`�l
�u:Y[�(�")>�� �"O���E��2� �AW�O���"Ov`��l�!m��=��!^J����"OH%c��ґE5�9B��P1?�.�xT"O�`�@Ԛ"(��Z��6j��5h"O�	�Vd�)#W��9"�ӑJ��y�"O�сv�DCҌ�U.�<�E�5"OZ�آ��D��­�Cx36"OZ�X��G97�d��6͑'�9Z5"O<Y���;es&E��	�(�ZA��"O�ؕ���M���ËR�5���%D��w�.@D5@O�pu�i9��!D���"鄈G𩻶A��:�p���3D�,j �N=X�J���<IL�d�dl.D���GR&��\��7km>�V�0D�,��-O"f��d
�4k� �E-D��Q!� �uw������X�cF,D�Hѕ�o�R��������n+D���G������bUH{%�6(_��yҧO47�� B�"G�w���⠃ؖ�y҅�z�:����9XN��a�=�y2��)���p*ƬG���#��[��yr��>�D}�oJE�h);��R��y�%U)F=����N�F:������y"G�U�&�Z��̑=�
��Bٖ�y���D@�ѣ22���bl_�y��QA3|�r���-�n��G
9�y�ȞH����*,���9E�Ǐ�y�ڡg ��
�Ň�(d��C�yb�Ku�m`�� z	Qt�S��yb��q� �Ȟ���L�Cb���y���n�4`eN���5�_��y�選w��{th�}!�,�5@Ʒ�y�g��&�����#L��$����y��p���c��)B	<��dž�y��z���c	�9�2����5�y2�ۨI���au�*��Ha��yBbȫj�P�"Ą�8���Hq��y2 �����f �>GV � ���y�B�09����G;#�ؤYS˒��y�lVL�⸳���!*X����@��y�ˇ= 1eh����.�%�d�ʛ�y�_��j�c����!�BA�y
� �L颮�<���;��ÜN���c"O|i���j���s#2S�pt��"O�����+�J4slƦQ{�a�E"O~�ZՄb^�mS#�&_L �b�"OL�n؏2�t�0�A�A<��b#��ҟ���d2m���)I�2�ܘ�S�@�86-�`�aqO�dB�9+V ��$��ZV �i�Ν�[���Op&�زؽ*b�I�f�Ôi��]���%	��c�Z���آV焪P��m�'-���!��X-�]y4*ɵhT��Fz�m���?���Q՛&�'\�e�<у�@��`B�ܣ����q9������I8�	<&�����8-���!���>����dKǦ�`�4�MS#
�\��T��
<"Ւx�E]?�	�X�F�'+�i>=����!A�� �&IE�eKbo�>��1 �M |s�УW&���� j^�/q�J��w���ð��A�[#L(H�6B�⦭��fH2���j�Os��������H�k��������˕�n�)��Ħꛆb��?q�e���'�?7�� q���W)�#m̱�����J�$�O<��5�S�S&g�Pp�#����� �hxv�<q�i���ig��]�-(5�`�V�����F;�LʓyTFX�c�i2ayb!$TD�&�ج��ӈ���H#0��y�b�nڴZ�+�D���Z�I7�/��H�	O5U�E`���<i�X1���ԋn��T(��f��D��h��c/��ZP��Z8�ze��%�v)LM��J���t������8�ɬk���<q����Ĉ~����f��-��ʴ@F�%�$$��bV�� �:Y��_�!h�		6)n��6R��$�p�O��	�7�9��f�&g�� p!,(��d�/$��M��ԟ��I⟐�Re��x���`r�D0/ud�[��U��zW�ـ:ԑ۔�Ǽ>k�xXvm�;D�p�AB�I�eS:p�g�*Z����W���@�6�I�@�B��r�L�5N��tO��">!D��Hn��F��$��gĬY�,\Y����K�i��[��IJy���*7
��T�N'6m���t�!�D��B�b�b�.C>Ah*0P�3��D��5ܴ���o�Bmn�$>X�d�#;=����J��<�6B �!�	ޟ$&�*\e�f�4`?qx�G^�7b�i��	�ډ��-T� � ���+� �HO�H
�%�\����e��xd.XP���|
 O�h�Zš6��GX hdnx�' �8���?���T�i���(�պ�(X;]$Y����/�?)��O����0�B51��%#P�Һ9J�A2�"�O=l�M#ڴ���2H���!� m����l?ц+ cԛ��'0RX>iSvGG؟�����鉂�l�={W�qerh�Ƙ {<T�5�ݻVI�G�ʌ�9@q�?��Oa���j<��-܇It9:!F�w-f�{a�i|lQ��7WV.,Bb(�{ZNe1�dT���k�ѻ,�!���B�Q�� �/X��E\3�?���3�6�'�?7M�.1�̨#Lɍv��wNǍ18���OF��$a�\-bm�+t��Իq�I�v��g��'�M{�����I܊[��-�3n�|S�)%�Y�Guĵ&�Ѕ��9� p   �