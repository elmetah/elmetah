MPQ    "^    h�  h                                                                                 �}K=���Z1��0��uOǅ�q����"��U��R�%'3PP�:\#��5�������B�1�Pl�5����x����2k���P�����-����H,�P�~���t9�E�U���N����U8�`�0s���ɱ��_b2e������	<���h��J����ꦂ*gi�џ��KԪVl�] ���%ј��ڄ���H��J�V�R�4$ ��l=�w�q</s�% ���� �-�m��}������5��mŗ��)��x3}(%��u�.Z'�ƨ��?mv��n~������Y�O4����OvS9���?D�|$��М*�?cE-�T�z�+_�\������K�7E��ėB� ��U��Fh��du����Qű�:����Zˆ�1�Gh8ZX�<�*(�'���^UX����TtTG�)�\�.�ɒ��T&7��j�ј����uߢ��g����P�-�o@��'<���4��b���ˣ�"�v�{>2iaVh������OA����,��X�n�n�
j2��V	mz�n�*�b��Ԟ4\M���k��E�S���� {�D�an{+Y�B�{�J�N���
�Fa9�o�j�܏j��qv��,Ti����o����g"ME�+爕:�O�vQd�%G�XCŋ{^m�̒�~X��y��[~:9�1�T�S���&ay/���峯!J�g��=IC�tܓ�X,�SG~����:��Ϳ�x�w�NvF�����#S(4ϵ�d/�j����	3� "`��	�&+��y�Γ���0/�	S���_�?���!��\0���D?�}a���5���k��h��&�Z/�η��B]�+F_ƍ���^u_�ODE
����c��&:��*�D�ْ��U�)_���8�����.�{��
����HU�����_�o��b�@��8U��\����lw�e��xZ.$t���[���q5k�N=�ߒ����j5+���r7v�L��K��szd�����T��s�-{�ԥ���G��l�d)��y��v�Σ��,ۙ=�S�P^ΞLE�o��nL��c�~k�
�#�HqiBv��quKM�CǓD��Ƃ8<����ѧš���}9��#��rnB��Y��]V'c{��Q�����T�(j�v$̽K���q�.Bi�\=��^֏P��YIint�+狟M&C���!*���d���ݴ=�U�MM�Y�pJ��\���5>}�S��[�>�x�� ~#��Z�k���IH��A���cxs�6l��| !����w�KY�V6�6�h%/�W���][l-� 2Ϙ��"�_�^�u�.>X+���cS�Y�y�ؙF��>�C�%�!���>�;��<
��h�?�H��KAO��1�K��J�}@�x./���w����߮x���c6X.��%X|��;��Z���'��4����qm�����r�B毹m����t�o��{'�1-	�M��t�c6J�ve�(��X� .���� 9�@P�%a=�v1s��u����?n�7`-��o��f���XH�]\�z2�HzG�n����	��C�t�ȕ� Fߒ
�=�ֵ4s�W��y�?�)E^�-��y�T��M�C&`��\�(3�xN}�+ɰ�EHó����R�A&��~����f����v!LZ_%��mȷ�.�Q����:/���Q滾��/m=P���ú�%�0Q8YSL4��ͣ
o����y�C��e*n�L*N�YhT�a�Pν� D�$��{�����!�3eP�K��Z�����EEU�c��ƛ(��������\"�{�vyY��1Q*�s��F�R����1�A�#1�B�HiMC��ᵵx>�cg�E�����=���߹��2�ϖn��gu�J;��-s��$�&U=����"�TSF��1���)�� K���e���%I�	�v��B��_<9�A��Ա��P	1?�hF��3��~�0Ӹ
/B�F-�������NKmh�_���<Q���=+�"�	�,$�#o���:�β�g��Sg�i��7>�7��8�(�l�(�u�����s可��}��Q]�̒����#��U��э�������[�{&ZٜO����|���O��O�W��QH���]6�i� ����]�rM�MW�^{g6�`��O�^z)��=�2[��/�]�,Dp�Ҟl�Up�[`�p*�,ҫ�|ß��;mb�����l/�)��Y���P \Q��ؙ��ǛP%���_/?�픒T����}Dfq�m�'�Ł]5:f�Hh6ID�&g�1�m�ډ�7o���~�f�:�g�i�c�l�s�6����4A�߰�>͟�Z���&u39\��j��=����U���s����c�B� ��k}݋�dir�nad����V��*J�AS�b�TvD���y�:9�b�w,�w/��շ��MW��|�B@%�~e�-��K�l �	fh�����W:��s�\c���Ab89[M9�.�k���'t����o��(Qg���8l`r�O���IP%�ܓǡ��5�V"�4>f#N��[��\6d��
��r��;����~��Z3��)�u4��U������G�[�)ԅ�@I8u�'�+��S���)��P��K��.�ݓ1���3m^#����g���yJu�Y��s�E��p��^��f*��@\gY	n+�iI��P��>��H�]�����w�r�����X\��w��#�+��mFO���@�|����^����T��3I��e��	�6r]���҉�?�oZ�l���Ś�lh�蒬�׶G5+�`�6��O�[C�w݃ވ���k���v�p��*�E�4�X�ֵT��g�PiF�?���x�(D�'��J6:wyƉC/n>϶�F�J�D����v<�,U�\�D���'��z⸶eH�e�]:������BP 0;3�,���J~�y7��q˳�����fM ^"-Q�؟樂$���ח���E��4������x�]��)�[+�Rß��J�=c-�[d�q������������sLԩQt	nI��ik�q>{����E�)�T�$�_bQ�al)���_jp�~�_0gB���52mr�2�9*u�Ff7��l3�X�kr�Q�yi������rKV�)�!!��~C�����W��?�����W�x9	=����H.�7��ݕ�����;�/�b>,���z}er؞CX@�����V�I�Jq}#h����j���M��Ī�I<�只w:8�/.���j��W�V i'T�mocZ�+��6���\) ��.���/Fv]}�ꅐL�����L�Z�/�Z�Z�nD2�4�O��dB�tO��J��ZJ�|��]�����S E�}��u�^_�J������-�՝�Yx��;�;	�Ut�Ih�sZd��ӣ�����RG��a�c����Z�>�%��'p��%�t#T��f���=���)�͕�ļ7�ϊ���:�;uZ���BON�9�R--d@��<m���H��ԁR<��\rv���2�caQn���x���ϙ�A,G�F�I��E����tRmu`���bf��O��M
��k�nQ�?���h�`@v�C��m�a�ْYZd({_��N6W
:09����7�%�Qq������o�����E�����:H��vl��%®}C�2�{M��ݶ���yU��'}[9+9�=v1jWxSj��&�p�=�g��L�|lg��(I^���R>X��G��ۥ{c��,@��j�2ҁN�;�����[2�Sc����oU�ei��;��3{�X{��	��2+}	�	B�f��|�;��?Q	:!3���~�e0r���}����0���	���#��&���I1!��+�#,�`?*�Y4G���$�@������2�~�Zq��͓�P��__���c���́寲�L��U�
.�Դ)o(���i��򯲭����E.�\1eA��xUNt!<`��L���o���ۺ粮���j�
y��m7�����
����dv���_��"o�-����;�GOW��J}�/���߸���^��j=*!'PYO�L�]�p�!����۳��ӆ��$B��q �����N{���&<��͸�{� ���)�}4��~��r)L�t��]�C{�ip�
��c0(e�$'�B��̃q��i1ģ���^�)Z'YIdc�3P�����j*��L�m���9{�O"lU��*��/�J;/x��9u5�zSy}��H�D��N yf��Xgk<x7Ic+�Aq��cS�g6�>6�6�!���mZ-w�Y����%�^h 2/W�z�����-��}��۶"Ucg^�J��+d]�c�c���'ؔ���LbyC���!�j�;���E����<�CE��\�kO�1؜���@_@�|>/�������:(M�v8�6sj���7W��;�%(�����9M���(C��
0��k�	]��NӢdO4ѿD�oS��'f�	�$�m��>;"ȫNebЭ�S6���bҠF��=-����Q�2e:u.� ��섒�x�@nс��`���3�ž�Oz͈(�C�GR�}�?p���t���9���>=#�/oW� ��%��Dӕ�t�T��돹MG��`��\A�"�3�a�Fr#���ÎXȖNs�R> ���SY�>�!�S�ML�v�țt)��=��h�/�/?���n���R�m����_�����%hŀ8T{n4�5��0����y(�C���;n	�*�M�Yc��ge;�l�;��$�ɱ�V����e��y0ZN��6ĢE�S�cryt�c>���w�H��A{_*`Y�!�Q��s\w>F�k�8	'1�8��~���ihY��\��x��gj�ŕW�=����<2���n����;��`s�$���k����N�}�#SE~1Ő�)K�7�3���ʫ	�+
��K�_�=A��Y�,`kP��?5���v ��b��R-
ꬬFHm9�L��YKW�ɭ�{�7���LF�+��	��w�h�#J&��u�-�Q*��N}N�ҧ7������ԕ(�wGcwu_��TЏ
�T�C����e�Gy��M>#�bB�;j����#09]=DᖔU��B��O�SRk��̹�IW�1����߄䂫 ��]XMP������g�KM�����y�;����5�j�]��p�߶l��K���Y"����W%�9ٷb�#�����/*���+�k.\���t�����d%I����? �����£}��H��� 5y5ՀHc�D�S������މ?+��>�~'%m:4�i��i��.?^��П4��n�_LD���I��u.��$�j�����w�Uz�s�f[���.q� ןqؽ����i�a�a��y��41V�,崽ANZY߯O�P�y5��ỈR;/wj���R'�MRk��U�aB��f~�w4-Wp�K�&@�D[�o��RjG���+ctڋA�Ԑ9���[(�.l���"ol����oz8>Q��~�l2`M&wO��@�c��%~�[���I}fRV=Y���F#)k�[�)	����֛��9j;N|����7A 3��!���^����r<�U~TG��)�l��*�8P��'X̅|���P<��@�q.���^x���3���h���b�A��{r0���ː��]�-w�.�1�'�e���g�e��u9d��˳�[P@��d/]������wbw�ʘlS�"��v�����[f6m�Ҁ���|�5���r��	\����@���D�
r��`�ͧY?M�'J\��:_l��m����C5�D�1rO!dʢ2��ޣ:a��m�Q@��+�,Eb�:X��jT���������v����bVNJ�Ey����H�q���eQ�D�,�����g�*��}o'�p�zԖ����e^-ЃĄ_��v��S06H�,r���{yR*}qF�\��Bpf��M"�y�Q��� |N��UX���+I��I`��N�/0�]я	��5�R~�0�e�F=��[?E*��F��{���d�@$bs��Q��I�Fk�ܑ>�y�����)�O���{�4a�F�Z��p֔h_k8`�p��5-yI׍J�*0�fRnfA�3�k��^�ͭ��x<�n��K��)��7!��lC|w�j.ҋ���e5��kW�9$�̒�H	�7��Y����i�lG5�=�>G���:M�"C�=����1�Q:���t##��!6Q��S�_|v�)��Yt����w�� /�FN�ϐ��� D/q� |m
މ�����S�xګWfDp(ō���^���}^��嶌䪊�<��u���ՋC�I�.�oڂ����n-O,�d[�>�up�|�������,�QEc9�p��_BY��u���H���-���z���vH�U�h�md+M_�^�-��w��Ɠ�<L����$Z���� ��'ˁ����*[�Tj���c��\�Ģ���T�79�S�Gn��UZ!uխ1���t�M-�˅@�M<z'����7���͜^�7�v2�2���aL���qɮ�VQ�'�,�- �$	��6��,��mpQD8+Hb!�"�j"mM�x�k�4O�z'p����������a�W"Yե�{:Nq��
�M79�� iQ���q�nO"M�So6��͝�yE�L��>��:��v��%=�C{�h{����Q��tr��/�[�r�9}p1�y�SEb�&׳���QR������=grm7IyǞ܉�LX���G�X;�#0��n�M}��/)N�PF��n�6�,S���"�S�`�Ė�36�����	��*+X|��D�<����䇖?}#!N���{0M����v}����+�k�drY���\&������n����+�F�����Tk�����=�ƀ���s��ֺIݒ2�}�K3_]H�����*z�q���Χ����U L���)�o������G���1�����a�e�I�xP�vt|{?������D��ە\��8�hjk"��xH7,8��W�B�.d����:: �]��-���{2G���ڊ��J	��l;���T �AE=�gPT�L�ӻ+��<W"�t����R���sB�N�q�,�x�	Ҩ���<<y�����է;�qJ�:}/��١�r��Ӯ��G]L�%{q5_�E=���(`�$� ��9Cq�4i�K��l�^L����I_���������Y�	���H�f!�(��&�U�]��ǩJ������54�,STJI����j� t�&��k���I~�9A�Y�c.Cw6�4�E�!�B��G�w��>Y�}�h�T:W�i���2-����N��"��^1��$�+?+]c��<ů1T؏p�ԧ��Cic!+|d4[.;qms�$�ʞ�q�>ԑ��VOOXQ1���@Ռ@v�/�׍DdX{F�����1�6������2p�;�靸~���^"�FXe�i���Q,�������%M����Ѻ4_o�w�'!��	 W���?�`*l[e��R�N����W�[�%�Zҽ��,��m0�u��Ԉ�+G���#�d1�ќ	R�ۖ������zh&g�>�0G�/���~Z�
$t�Uz��+���&=����*�W;�ꪍ,�_�o�#Q�/���ʥ�M�
w`p-\�����Q
�a;ޡ;��i�Y��jiR�ލ���.�ǐ���1��LP���v�z���!����/����]����m35��:���0�%zH8O�,4SP���c+�.!y�����>}nG!�*Rm5Y^ ����U��)K�V*$�@�1GT�,6��W��e��!�Z	 іQ$�EK��cML���/�+�U����s{��Ym�Qg|s7��F���i�1������Ӈ�L�i����׈�x��gJ�]�0#�=��{�o�q2S��n�k4s;hmcst�\�����<����S��1��w)���K���ۍ��[l�	� �����_��A��lԧ:�P��{?pם-C�(����
�7�FcOs��D����K�-_�����2e���+f.�	Ŧ��B#%���s���I���7�%�����e(�����u�\Q��U��e����h�wv��*�##��"����Ԕ~{\���"yْ�����KΎ����\�WN�����9/ф_� m.G��M�J����g���`�,��"���}_������_0] �p�Kl]Σ�Ѣ����"0�2���t�b&������/��2��b�Ɇh�\G���O�{���%�@�Ō?{���jV�9�}:�\�#j��;�5p��H^2�DD�ͳ��f���ʉ�>_����~b�:ϒei}���P%���	��˻47P
�:zK�Wʟ���"u)7���j<�c��]�U�#fsf?��مv��� Ҏ�3��]�i�2�aZ���`�VVX���SAI��
I����y8��/!��-j�w����xoMM�ﰥ0B�d~�^-��K� p�p��),r�M���)'c/eA�f�9��[#�.V���8:����Yy�o5��Q�p�.�`(V�O�#-��N[%y���WCj8��VX�u*�#F�[-`������L;�(
�;	X�����3���\����%���y�Gg	)
��6,�8+��'Y�D��b�����9���b.�$݉���^��3�쳕5��]��/͹�{���q�i��a�m�iI�����1g���}�6�F��6������]8�J���w���S�$����"������m|.����|>��������)@���w3r������?vJ6���9����l^c�H���,D�5au�,{HO|�Ѣ�$�޾�Ӎa�5�,t�f=2E���X�^;TUS����M�8K���Ի�5ώ���Jlq�y����J�,����D~+ �c�����y��5�x&'Cpz�kH�� Me�҃�c��41��01}�,tF��0ym��q�����"f�jQ"M�uQ���[{��~@��������~ � X���*]�Z��`�R9k뎀�O=Y�3[%3�
"�����f�y=sµ�Q��I��k|g~>�_ �5�#)��x��s�Haa���[p�ʳ_�)�
�5(�<���J*�~fm\M���3��%k�ͯP���o-�Ʉ�K�&)𥳐!y��CW��'r��&���'��a�-W:�!9?���V�H�:=74�ɕTR������s���>b���p��(|�C�Z��P`E�Lsƴ  �#��<Л�`1P:	��d9���d�۵�w��/�Y�T��M�t g�S]m�x�������q��f��_�a����Ak��}��A��Q�?�|����ِ��PJ8�$@�ƪM�� &����O����鐶�|��k�a���g�VE���ky_���0�z�c-���U�󱧩U�IXh܇6d��������.R�Hf��ۘ��F�Z)I��w�'&0ߏ$k�EbIT�JЬS��҇_����7�M��	��pL�uP�}����˯q}-cS�@��$<���CE:�R��Hڣr�vN�Z2:��aGڿ���D���,=���C����	���mkb��[Ob�����M �!k�ݣ�Ⱥ$����,-��u۴a���YPS{�-N�H�
S�v9{�+�{�+��8�q�����X�ZPooqd>�8��E��b�I4:���v�`�%�}CV�{�D��숽�o�C���[�ڭ94��1`��S �&�-�s����R�2 0g-`jI�0�MX��G/1ϥ�?��Y���	��Nǅ��wG��)S�}����)�[�;��S�3������	x�+3c���������-ԇ��?��!i�,�t��0(%�ʭ}2���&�E��%z��&���?���ӷ�+���6�O˜`$;t��5�Q���N�W��X�͚��F��_�Q!i��Eۻ��L�����U���ʾ&o�Cx�U�(��̪˞����ew�xK�	t��>�>��»p�����p�s(!jZ=����7���m��*�dl)��z�Ϙł-L$e�vDG�>�����e�܅�Q�q?�J��=`�PO�WLV�D���əW����^�����WBG�.q���^���H��{<������ߧvV����}*G-4�Or�����]��x{L!���Q�*([�[$݁ѓH��q�:Ii'���^����z�IZմ�<,ٟ~9�i���6�#' \�݅K�U���j~vJ�T��}5��S/7��vI�I�� oL�k��k���I�ՋAg�@c	��6E���g!Ɛ-�#Uiw@S�Y	g�Q4h���WJ�M�.,�-�
ϩ,�"��?^LG0�9+oc���J�؊T��	PC$26!F"��Ą;L���L�9��9���� O
�M1�}Ļ�@Q��/@w���
)v����z����:6�B�喠;_9;R���S����s��<��٫������1���`�ڢ�(-ѵD�o	�)'���	���c�P��b>L�e���I��?��2�?��������ud<����}�H0/�B�ѷ1��V�鸞��Jz䝩9m?G������/ft���q��C��=Y"��%� W�W��HS��z�4��׵�
w����M}�s`w�\�{B˩w�|$ᡶ@�Dp��ā�Rt�ŁŔf��חTX�L��L�D�Q⻷Q5"�M�	I9/�܂��3�ﰦm��a�y&�k�/%�N�8J+�4��c�;���I)@y�����n�Y�*�YYS��j�����q�r$�����gy���Qe��
\��Z�h�l�E�:�c(? ��}b���+��}m{%{��Y؁Q�5�s�WFH�n��1�@��4*�s˥i����R��x�g�����=�AE��*g2�!n�QJ�y;Ca6sO�<���R�� ��3_bSwN�1�Ȇ)B�K�.\���-�	��Y�ST"_m8�A���"5�P��8?��=��Yz����A�v
`�!F~QU���fw�Kͽ(�0#��-�Ӽ�<+!d�	��w�i�# F���鲇�D	)z��7o�`@��j!(m�E٣�u�ʆ��v����b� �;��=�[�Z#S�ׅq�E��rڔ���������D���q;�ɪ~� 'K���W�>�ym#�T�
���8 HzK�̟M��"��gG�ƺ�q�����u�����l��1C]�#p�Y[l���یZ��'��iD�IK��s�b�����u/���e�ɡ�7\��*;��L��%~���U?�T������T,Z}�����a��v��5�HY�]D��N��� ��5r���da~�c:jX�ixn�����f9����4�α��⟒� ���u${�m��j�m�dU��usA8����d�� ͝1�z\���i�#ua��S�;\LV���AAD�Z�ebB���yS�c������w��Ո�[MH����Bq4�~��-M��K�����������H*n�*c�obA�:9}��[��".��P�Ӂa�v���o��5Q�l���`�O6om���%t�ǲ��'!VsI=���#�@�[h���-/���̃�M;�S��w�-��3�?C�9��~��5��pG"��)%@鼱M�8'�'�q�������a��|t�.8'���9��3d:��� �X褊>�����:��R�<[Tޤ˴�]cE����gj~;\�������h�r��^�]����}�w�(��h�l PӜ���FKm�-�왼|��F�V�&�����4���D���r.����C�?�g����{��ll�F��#E}�g�
5���'��O��X��xH�ٰN���	�����E�v�X�R(T��)Á�G�Sƙl�����J�ؾ{J��y�f'@���j���s�D���>��b�-j��s	:'���zJ`f���)eT,@�zbϻo�!%10,�*,�:|�{��y���q<c��v�f�Oi"�r�Q�ؽﶚ�9K��(^!,T�a�Ї[H��e�b]�E��l�R� ꎛB!=Ԟ.[�$��EK��q(ذ��xs}�{Q�Q�I��kW�>,f��NV)�1�55��a�2��P��p� �_�:X��B�5#�K�C�C*��f�j�\�X3x��k#Ĕ�J�����Z�${�K���)
�=!��,C2J:b�X���b�	�����W��9Z��̈��H��v7o�-���q���"�`�`>}�q��4�~ZC	���D�G��[w�#�kW����.��Ye�������wK��/_���!��B6 �����m@3q���ч	?��!)�zp�Ń���D1�0�}����w茚{�����٫����(9�����嶪�������O� іo��|�4�<@��PE���f}`_������~~$�#W��0�M��&EUE�ch���d�~��$'�k���%}�򉛞3��Z��|['��T�JT$�`�(T`�Ї�ݿHgx�����(7�����5Ƌ^�u�8v�������-��|@�c�<0������m�T�ý!��!�v�h2՜�aB@��'�:���ә��,�䗨ڞ������b��mf�
��b�2�����M{�Xk~ ������sD�������0�7aڳ�Yˈ*{�M�N�t
���9v{��֕ƏV��q����5�[o�;���\E�P-��Q:y�Iv��p%3�tC1�{�&�݇�f�j��J[jb�9O[�1��S���&Mn��[��ſ��'Bg�r�I�{i��mX�m$Gj)��L�� ��cKDN�����?E��vS���XO��VC��Lі3�V�$�	��+�;����7ǡ�����LA@?�Ă!� U���0{0�x}��!)<��:�T%o&�Jպ]����+20��1�ՠJ1g��}D�=��P�j��):��0�1�h�Y�A�t_{�$7E�`�e�g��vlb���UV/���s�o9�G�N��C�����[�yVX�Pe�xFn9t2Z^�G���}m�:�W�K�î�xj������7�lv��b~�Eh�d�y&������ m-�暥q2G`w�Pl�ր�bR �LJ�ۅ�W=�I�PJ��L��6�����r=�jEc�v�E�4v�B�_�q�d��;���2{�<o��s[������Ԯ}%���.�rZ	0��W(]BY{'-���+��N�(V5$8i�snq�i��Ћ��a^�n+T(IU��؝�9E��'�u����������� �?U��k��UcJl��(�5*3�S
D������ j�����km�I�ڥA⊛c䒆6X�-�{&�!��M�~��w�+�Y$W��D�h���W�U��ɱ�-�DJ��"�.r^g"�xx+�&c?_p����؅X��]��C� !a��*N;'�j�����n��4R��mDkO�+1)PM�6^�@,HO/{V�z�QqZƧKT���J6�ޞ��_�m�;��I����A��@YYif�@��y��r���|�5�Ѱt�od��'��T	6j�ފ��	�yLe3���DǏ�[���")�t����Ⱆ�&�u���՗�������r���y.��8��s��I��z��̩4�IGcp�pֻ�JP�t�b��y�r�~ϲ=�j�� #�W�2ܪ�7��!��F�凧�@��MR�`	��\R�r�dէ��-,�1:��,���gR�U����j
��R���g�@LF}&�,I�w{�t�1/Pr˂=��
��m)������æB^%9C�8E�}4	?+��(x�d�y������n��x*��YT�,�xK�<鑌X�$sà��(���,�Re����JZ�u��D+EA�xcR��"�a��oȃW{�-Y9cWQ	$~s�P�F�w	��1���Ϗ> �.jbi�[)���)x�x\g����fm=��J�%�2ɶ�n��a�;u�s�rBՒo
��j-���S2�1�)��K`��Q��ڑ�	�
<��G_(xbA�(+ԝOePuf?�=��G�I�ȸ���K
��F�s����A��Kn&���m�(=��]�+ܹB	��#�#���&�D�"2��?`��7*�v+Xɬuf�(HX�j}u0X���y�`*�tlK.�͸��k/@#�v�����~��4r������8وՆ�]2������޹��W��4�t�o���U�� #��I�M!����%5g��S�֌���J��1Þ���$J]USp���l���G���ܦ������
���pb\����/;GW�E�zɼ<E\=�����Ǉ�n%�Ν��?1���@���o�a}0�x��yӱ�5���HT��D����	$-��P[�����{'r~��:>is�z�޿_*�"4-me��5
���5�Buߡ�nWj�P��[UxֱsQv�O�z�CN ����\�Ӯ�i�4�aP*3� V�++�ȇA?�e������mzyn�A% P��'Gw-�#|�MCZ
�fN�B,$�~��I-�ohKg ���<�_V�C����%Zc��A��9��"[���.�,��n� ��co��Q�ʎ�$.=`��Oq��4��%o�������V��� ,p#�[�[�,%��lD�����
�;of ��Ĺ3dlҺ��/8���F܏f��G�6)@��,�08�9'ϜQ�M����%���O�7�!.S�M�����3Y���9��SbE����a���-l�_*,"+��md��L�����g�:����;y�<�u�E$�4�]n>]��e?wsͥ�Ʉ4 A���m)�w���5m��o��L6|���J���A���k���z��݀rɿ�����?,���X�!�1��lTJ�����ע��5����"��O2=`�c�<���эW#��9�����E3w�X�f1TZU�<��n�#��ٻ��v�� J�(,y�E����Ϣ�7��4�Dtԋ����R��@��n��'��Yzuh��8ne�[�U�ﻪ�f�0'G6,*O��6=�y���q���_@�f9U�"�7Q� �ڌ��ub�C�*��[�<Hч�X�� T]�P���R��,����=O��[�D5��8�L��ӆ�Q�s8�Q�VI�?fk2ݧ>g�x�k<�)�ҍǐ��N�Fa�u���9|pg��_l2�A�	5]wמ��*aIGf��'׵�3S�k^ ����������2KB�i)%�,!o��CT���\��/RW�k�9u���E�H��7�$���e��p��},�Ž>��m�fޟCD���I5�B����#T�ard)�VL������X�UHm��[�w���/;��C�� �60@m�)��"��d,������ ���;�pgg2��}/Aސp{�����m���4e�F'F�ڻ�� @�Vg��ZO=d��E��Ƣ@|�*��a���}E4,Ľa�_SD���<��Ν�둻Y�'ƴU�6�h��d<��ӏ�y�#�@�>���X��n{.Z_���{'�ny����{ЏT��^�b'3��}�X����/7J��x��Ʀ��uF���"��%�x-��@�z<�����<���d�>~5���^v�32p�Oa=�.��9�����8��,3�5���1Y3��*(ma�gI�bR�v���CM��kYF��+kZ|�X�CQ���^a���YF*.{�mN"�
�H�9qb+�1\!�<�q�i���ʀ(o�2�n;�E�T�ON:4��vبo%��IC{9)��"���e�\�@��[%
e9j��1V��S�ww&�{;���ɯ�ntg��<I�K��ǀXs�G�A���!���c�^tT	�N�O��mX��SO�е��^�Q!ħn�3gL�P	n{�+锄��:�Ҽj��_���	?=��!�K��j�0��sk�}hve��N�u����&*)��5W`���+mṱ̍ԠEp?��$�'��k���P��k���K�<�_n��߫��{�w��KGQ�'�8^
U�����Ho��	���^�y�a��T-.�1.e�nxAt����4B��_�����&{)���-j<)♐Y7=7!�x��`5Kdb���Y[���-�ɨ�lS�G�l ��֛�;����'u���s�=���PE��L��\	����|��KS�Qt6�o�B}q�0:�	�:���M	p<�;F�N���n���} U���rK��Є]��{Y�����݅(Q�$�����?�q*�i�b���0^���MIP���b����B�z�P��
c�n�ݻ�`U��� MpJ'�N�-b%5���S�p�4��yu e���!"'k(o�I���A]S�c�j�6��(�a9!��J���%w�$Y?g��X�hl}�W�3q�dW!-����_��"A�(^�6���+�TCczH�ŀk؀|�Ը/�C�/r!|�A���;��1���o�a�/A����O�Œ1D!eıR�@̟/�U~���ld��M`�b?6ߚ���Üy;Ȏ睉S�����We�%�0�Q��&�M�g���2�Ё�ѫ�;o�>'R9	Q�՜Y``��c�l�eή��?��շҌ��Drr��å۽��Ru�Ab��}��Zf�����x�Ly��N8��+z9��/�PG�@��+�2�e�t	,�T]�߹W=��µ�WWL.Ū� @�;7�������{*�M�%`�\��b�ǜ��V��������:�R�:>�����[��.��L�u������X����/����%��m�|U�˼��ᯠ%�W08@[4d����T��uy�k�]ubn�)�*#�BYOy���%��"��-\$�붠�~���_��(ve�Eq�Z:�^��)E��.cބ��OzW��o��x�#�	{K9$YT5Q�2s�.�F���K%1�ȳ�ꑶ��(�i���H5�x�Sg�:��F)=�_�߀�2� �n'4���j;��Ls�!�-���/��!S��811��)� �K;�A�\P�,S	�?��	�k_��!A	����{PP��?!G��������@
֗'F���u-�eKC>X�f���#弸/}+�/	Η|��#����a����t��:t0h�7���Fp:���](#�OP�u����U�v�q�/��I!��3S��Fe�#�g�����:���I�O�������8+�?�b�V�����W_�v�ZV�д� �q�7M������	g�����������k�<�y-e�V6E]�ep�S�ln���j��UL��n��츦%��b�u��=�/��� ˇ����\��*��4y��ل%������?�9��s�Ί1}��8������A15A+�HO�DUI���|������+92�V
�~^):�CLin���y{�%�,}@4�+%�����F����Quc�#r�jm�k�7��U��s��߫�"�� ��D�����i�e7a�~^���V	�}Q&A:�����<�y����Y����wV� վ-�M>?}��ҞB�3N~��-CZkKBN`�0p���!��>j�:թc`��A݃9s�9[�q�.���	q��q�j�.of>Q�y䟮�`���O�e����%j��h�ii�V����� #���[���c�h��W�9;2;:�^��#ۯ3?�$\��� z��"���+G���)[\���8�(|'
I��9��,��l����W.nN��O����I3��Õ԰��N���@�����7���!����0��V��1�g ��T�Кf�������oم]	����m[w��Bʄwr;���b���RR�TmMmi��l|O?��2��\���C��bD�0��rd
U��_�?����+�L�l�mO��J4�ݮ�526��VO�������\�ґ֫�w2�ɻEΗ�X~�VTf!���'��ͩ�b��o�R�N�yJ=��y�DA����]�����D��C����Sa^c7��i}u'T֞z��N��eJ�`�0����2W��0"ܽ,��p���ey�F�q2xғ:*�ftz�"�{Q�x��l97���X�^������ш"�N�]�{��"��Rj����<=�߈[��.��s9����|��9s�w�Q�!I
��k��>��R�J�)�����	��a��n�F pB,�_W����B5����*��f���R��3.]�k�\�̀����i��ǂK���)@�c!�8C�>�G���e3�-��r��Wk��9���~�$Hu��7�ҕ%�}]ͯظ���>������	���Cri�!n�=;�ƒ#���^l�щ2�o��r���ׅ���%wdk/�=5�Ӥ�3 �κ{��mv���p��9ڗzx��~�yB�K�mM�}ʦ ��
�P�R�(_����F��E_���[�˂�7@��>,O��=G1��H�|nK��Q����E�g�\��_��Բa1D���ֻ�N4�b��U{݂h͕�d�r�Jΰ�>CT��˨Gq��EoZ�O��'7S������7TV3;�=�����0�ݕ���7���3�_���Iu�Ck��g]�`�D-4�T@���<�P��tv$���<��^���:v�l2"�a8l��ݞG�B�u�S�,�������lO����Im\U���ebJ�֮�Mq��k4��fl���}L$=�����)a��Y��]{��N]
$܄9li׌B<����qSV����äo"J"�	:�E����+:��cv�|�%)$�C�Ty{tK�ݽe!�`&#�[��F9���1�C<S�i>&è��D���un�C��g^��I���u�?XN�-G�yå�a�|낿�Z��oN�c����YS��f�����LC�,�3"�H�	��C+ć=�0�úm�+��(���y?���!�����I0��s�v�}���1}������&EIհp^�d2�+�ض�g��@�S�q��l1E�
u��P��֦F֒�>��7C_�-0�@p����]�,���s�sU��xͻ=�o����Ǐ�y���[a�/wζeH<�x<�lt���ޙ�b_�0���p��$y�j��ș���7�!�C���{"�d�z����I7>-̎�g��G�q���vֶ�G�X�!�����;=1P@��Lg_��U왨� �`rO�,j����yB�q��oex��l��h�&<e�Ҹ)}�'+��;}�E;�rЬ���i)]8�;{ݤ;�1��"��(L~$�e8�y,*qEg�i��`�_��^8��ag`IK\R�M�'��T�]VP�*0���,L��VyU����{d�J���H��5 N�S��e�o�W�i� `��|d�k���I�D2A�;�c�b�6ξw�f!�:#�4=wq=�YZ�쌋�hG �W�1���a-��Ϻ�"�Uc^�8�UQ+��c�Q��4��{����BCU^�!��� ��;ݐ"l�I�
�w�*PM�#�O;�1_��,g<@�o�/�t�����g�]�g��P6�v��_���;�y�$�*��2P���M����K�n�o�~(�����k^�Ѧ4hou�'rA	l_��U��3,ﬗei��:0Pp��G�0_8�ۘ0�Y��u5���˃J�Y ��P4��j���S�zI-����z���*�SG1M��-�]t����/j��q�=*\�;-W�IN�y���˙t��쳛	붖�MN�`�K�\����U�͟��'�(����u��RE�~���6 ͙������@L<�/��v �\�)��ߔ/�����о@��m���[�=�%o�X8;#?4���lnU���y�4d�8rdn3��*�+�YJ���.�@��`���"�$��v��&>����re��m�<Z�b����E7��c��j��( ���~�0~�;{��Yo�Q�`�s�,6F���?,�1���E퇤�i�B�îlx`��g6�Ŝ�=�
�ۥ�2?j�nBյW�U;���s ���ȼ���^��D[QS��a1L%)wK˜�6��2i	��t�dѐ_�W�A$�	ԓ�P+��?\��}������R�U
���F���~T�aK~.������z}+R�	1��ڑ#��F�����X��5�c��f7��|a���k��(����Vuf���ٙ,�р9��>dD
ͮ�7�!��#y��BEטz�����*m����~X��+�z�b�񱭹��HW����Rd�Sh�K�G �9��AMW����:gX��L�� ��[��T����h4]�&;p� ul�?۽Ay�%+�!�Ӟ`�Zb�Z�����/���-���X\3�?ػ�-��!�%P=��?�۴��a%Υ��}&9ś�	��'��5��HJ�/D�����Q����P�1�~N�::;i�ii��0r����G�|4#
�q	�C��PC<u�~�Yj(Na�R6�Un	�s����ŖO5� �����I�"i�aF�Ճ�VD
��uA5<��vn!����y�!6_ψ�e�w�!��Y��M9Dl�wnB�c~�U-�d�K�Ѓk �^��9:����c@3A!�$9�,�[ov.BM���	6��Ţ9o!U�Q	�,�O�`�UWO�'�jْ%e`(���$:FVġ�}#p��[y|��G�нP̔�d;��6����3�mH�e���~���GS�z)vQ�"rI8��n'E/��i����B�r�iR.��uT��Va3ωƕoo�If��R�׮��R5�U9(���U��.���Ȏ�g{
�܆�ܔ2`4�����ƍ]�G��ԕw)���?��V�\�ݨ��-p�ϧm�l��^|�������wsR�<��j��k�r�t�?�o��ՙ�g;NlJ����7��5�>��9O�m��3��*��M ϫ��<�R�Ei��Xy�T���ò���W�ݱ��J�ގ�ˆJ�_Wy�c(Q���hɱ�pDj�G���>�����M9�dg�'���z{���/e�� � Z>�I�0��,��ꛬ�*y�q�2N�4�f��)"��XQ��X�Ǹ�j+s�yDR��o��b�ٙ�6�^]��m�}I�R%�~���E=E0�[��w��ή��Yɒ"ls���Q��I�Vmk�ґ>�8���w�)�t��F��ķ<a\M����p�_�.��w��5�"�T��*�V�f�T����3	��k��,��A�|�J�5�K���)[P�!e��C����Ғԟ�o���W&�9�����HPV�7 )���xj{�3eb��>����\��C�C�ʥ����8�l�*#�Sc�xW�L��|�Pܪ��V�ǁw\f&/��-P�X�9�B ����`+m#!����g��RSw��X��Z�&$��}e,[������$E�������0�<��󐷎Ɩ�:��(���BrO�JD���|�����
��SmuEjì�W�_	�����1���tg�����dU��h�/@d�K=��˱Y�ϩ4$˃VD��/�Z�O!�K0'�W��{�h����Tѝ��{�����q���7 K̊�*��Txu<�g�d��˛�D-ϱT@���<A���/P��M݁4_��~�fv:*2��Va32�8$^��]�nPw,)g6�ko���e-�3�cmW��\mb����M�(Gk򵣡�����x��ژ�a6�a+�IY<͹{� mN�9�
���9g���H���:q3\��l��o]�ͤXpE�Ƶ�O�:�8�vq�%��8C»�{����X�2�[�e��q[��,9��M1L;S�{&������������]9gk�I z��ªX)D�G�'���w>^�����kN3���c�}�>S�JQ�)O��G=S�]	�3�=��i	d��+��f�k�����k�]�V?��p!�A��`��0�T��R}��:��Ǘ+3>ꅡ�&`��+���?�'+�\U��z�;N���8%'[��kf�9n�����f�9�8�2e4_$�JU����KԌ��2I���r�U't�ͶR�oJU��V����u��
�	\%e�Jx7�ptC�}�x��.�T��c�܄��_)jrxg���;7�+7��Wі/�dX+����(τ�$-��L�b%Gq�B���n�ѡ;��䔣�*��6�Z=̒0P;�L¿�����Æ��۸W��Ȇ剭B��Uq�(����ǰc����<�>��>�bQ��}����er�.��#]���{�;�l���ZA(G�A$IGp�49^q`�i�ʋ:��^s�G��0IF�)稝�j���x�p����nHI���lU�5*�֛�J��c6n5�S�*勪���x� [����Ƈk��eI��ASDtcuzv6	��L6l!�ؿ��bw,v�Yu�>���h"�W6Pe���-����N�"�"^�s\���+�Xc�z�Ŷ���v$#�n�~C�>!������;����ʥA��%R�~,O�X�1z#mħ��@�3�/,���K��b賧\���ش�6sA��TyZz;> ��z�������خ�f�����M�Lnۢ[@ѡ�0ou�'��m	�1��Ok `�$*�e^T�5x�*���z�Ž�dd�s�z�	u�ƣ�Ʃ�����#��B���Ud�����zo*�%qRGtA*��ɬᛩ�t���
ɽ�/�[=�d��W�w�4.=��ڕ��vz���"�M�,�`��Q\cU�˕
ө�����ðc���R����{^L׃���#�L��VȽ="�=�N�q���� /aG��n<��[�m��y���7�W�a%
�86
4�B�'Az��Ly
����nnz=*Y��YE_F���m�T��7f$w<�x�@�S�C�^<Fe�!H�	�Z�K\����E��^c�J�����2{5z��\�{� �Y��Qz�[s~JKF4���,�1��?Ϡ�Ç_qi
~�>HPx;sPgq�C�7�I=����6d�2��>n]��j�;�p�s;�K�c�A��I�DaSc�n1g��)�?�K���1��bt�	�	˧��_Y��A?���_LPd�?��LH�(����
LͽF�n���&Ҋ�K�>X�������n�+{_	L��r�##l�׻P��Y_�0�/�r�7[)�| լ�J(�X��|�u���: �,A��o~�C�)����0S#?��ݝ�ub�E�n�e.�8Ʉ��IX��4�ε���u��/�W�,e4��l�� ��}��( M������g��:�sn��3�a��/��̺]&��p��ul$�&�x9�-�����yg��(b-_ڑ�M/L���v��k^\�� ؖ��8�M%�|���s�?B���qo����(}���j�[�b5w�@HE�-D�:�ő*�!�[�0E~�:�:֮�id�y��5��5!�b��4�ɰ�?�~8����>u�W���j����m�QU�Rns�[« +H�6� ���s݋�pi/(a�����+DV����jA0����,��[�y�}L�>��t4�w�˻���M4i��w;>B]��~"B(-9�K�!Q�����0� �4*��c��A<!n9i�l[J�z.}��?���\� ��oܺVQ$§�u`o%O"ܷ�=%`��^��*pVߩl���#KlN[TOV���и�����;���Q��h�3�G���� ����:y�wB*G�)��ü�8r�'�,��5���+��� �h�.��'������H3
���
NǨD���C@��-�m�p��p��6Pސ,��ɥ��Dg�/OH�o�ٔ���}[���ө]?�m���gw�C����Zq��Xv�����.m�����%|��{�mɒ���T �b������r��_���D?=n��lق�il�r�Ы�S�
5h��lOC6w��3�E����ӫsS���E9�Xtb�TԘ�m`���.�X�+�%���HJs+Ay��K��I��Q��8<D�A��������p���_q!'
I�z6sǶ"��e@�1���[�>��0fA,;Le�g��y��q(V��]�f�$�"T��Q��o�"X�%����&b|��f�GIE��x]�1����R�����7=��[ad�1Jx�<���7b(si�Q1rJI �k���>�c�<��)�uǡը��a)�3�<�p���_Ϳ9�e�5a�ׯ.h*�Cf��HJ�3�>0kurͶ�:�w"hܐ�cKs/�)vɪ!�Q>C�9�Nv��-cd��՟(�W�q�9�YR�t�rH+-�7[�G�[��s����1�Ll�>����>�oŋC��>�W��3��ǔ�#�6ò���d{��a��k�&W���D�w��!/K��kΥ���4 f^��3�m�]a��lǇu�.�L����o^�����6} ҍ�������F���"ѷ��k���ћ=�'9��f�ON������^|�����]�a�E?u�RyW_dO���D����iD��6[��c�U��h��(dME=���ʱt����ca�^��:�Z0�k���'�{��6S2��e�TL(���T��4�f.��T�7[�������Nu���?Q����x-j�@�}<�%��Έ��E��9�Y!�vuU2A'�a.H���Է�U����,,�Ҙ�FJ�������umR�hZ-�b��o�5cMg߮k�w����+Vs$��,���aF��Y��A{\Q�NӅt
Zc�9b�m�Bo��B�:qN�
80��[.o����?�CE����`��:e�v)��%3RC�B"{�����V�$�Q�[V�9��x1���Sg��&9cg�z�J������g���Id��k��X!�GVJ���@Sr���o�%O�NNo#��avXI�S Ώ��9�B{?ĸ&3���8e�	�eY+z�����κ�]���G��"�?n�r!��F�ۓ�0o2#�n}9X���.����@`E&{��զ��$I+����!�6�0�'�E���������IM��˒�K3�-ρ_`E�+�̷�S���'��,#U�uͱ��o�)��:g ��q$�v����jD!?e~��x2�t���3���I��&�d۷�{����jP���Zm7NV��y'ѱ\�d��p�\��Ͽ�_-S1�]��G�t�<�����N ������q��=g@AP6V>L@ ��L�މ �Vl��i� {uBNq�T�%�5�kz#��s<[�o��e����"8}�v���rF��1�J].��{��
����XI#(B}a$�H���evq{��i����=^�����xIAV}�ʱ�%d%���K�/��jP��f�݌�UU͍L�1�WJXb+�~Ў5�MSv�����e�P�� V�i�2I�kYx�I /�A�l�cP�f6D���I!��h��ww��zY�WN�R�h�ůWq���5�-�h$�p&+"r�d^����Z+a�:c+���Q�Z�q�����ZC��!�@���;���=��@K� Γ��=�O�R�1�T]�"��@�r/g���+f]f������9t60����})T��;ymz�Z�A���O�h�BE�y���@�e�������͢�w�ќt�oг�'���	�#	�ʠ;�Me��e��I�0��Yҽ�N�����u�N0�ϓ|uk�����t�
��u0�>��ɽ{�0�g�5�0z
x9� �MG�q��\��\*tz�J�审�j��=`�ص�,W]�@���1��g�C�Q=�,�M�`�`�y\�۳�P\��)�,�Ë[Ֆ��UR{��������>d��ӗ�L2��Ș$�x�}){���9�/�#��)���vLm�݋\$Ò��%�Uq81q4u����3Á�[�y�/Y����n�R�*���Y@2���%7�(<V��l�$�Z�S֓��������eܿ}#g�ZkTq���E-��co�w� ���0�uS?4� {|�"Y���Q�sY��Fo��uM�1����K:�%�i%t���`x\Wg��'�҈�=���ߑBs2���nxw�Mo;��sv����Y���_��MQS`1���)m��K�(#=K]����	�����_�xAZE	ԉ�P�M�?�l��x̈��N�
�F<��tť��K�n&�7�m�)��n>+�P�	g���#GE?��������+��A(T7��x��a��(�C� �Yu�����Ϗ�!I�`[B��ͤF���y#z��x�p��Rzܓ�S��t[���u;��7�'Y]�߆�Wp( 6d�ۥd�Aj� �Ւ�5��M�B����gUH���'�6�܊��
�b�-�]�yNpԺ�l8A�3QM�H#�����TRV�֥�bȃ����/�d!�1S��(e\)n�q�'�s %�����G?����,����eP}*B�Eӝ�n5��H@&Df��Fk�E�]��SR��r~�ع:q�i_�S��R�Ky�}N4'��\-I���S���Yu��4<�j��8��bIUd�Zs��;�;��kr
 ��-Uދ�U�iJ�wa<<���oJV�hm"�A++�,��m@)y���>��O#�w��ՏM/����B#�~=��-�ټKӻ��S��7?�/:��K�Yc�sAWs_9�7�[%�.������.���{�o�@IQ?����`JO]ǜ��^�%[���y��;�V�Ѽ<#&I[�E��4��гP�J�I;k`l�����3�\�������v����(G��)��^��8M�d'�݅�p���P�(���#��.�t �k���n 3E�H��Lը?�S�QU�M��B�K���}���6��d3*ɾ�Ug1l�L\!x_�(�#XM�� �]�У��EXwߪ�ʵ�)���cH��� �m̧��Xv|`�8�6k0ɭ}�����=ڜ��*r5������?����D��ٝml@���jÏ׎9m5��Q�O��O�7�`�.�C��N���tzE��BXo�nTw�D�(�ơ�o,����� ��s�Jcy���ώ[k�"yPD`�4�����O�4�K�Z�'e��z�Z�=)�e�Y���<ѻ�.3(�0[=,��ߛ"��y,jq��˧�f%�"��Q�X"�}���`��(�G4��[����$�l�I]����3��R����"��=;1[<��l���>��)�Ds$Z�QLJ�I{�$k�H<>Se���2�)�����F:/CaD�"��PpӭI_qd��=|5
M>�
��*M�f��ûT3��ukJ1l�Ql�r����*�K.�^)�b�![ACy���=B����S���tW�^�9��
��;H$�7��p��n�K��B�Z>���R�dJg�C0�ǥ�6�.#ߴ"��#@9��&�B"\�����/��F ٽ'w�\/�0���/�� AV;,'�mG�y����!���d�!���IN��2��}����򓠌a5��Y���2��2a��F3���Ԃ�i`�٪RO��1x@��2�c|wj���ܼ��u=E��u�M�k_�=V������I��}m�wڦ���UL��h��md�^�{<���w��*�(�9Ժ�Zd�Z�.��t�'H���" ��,~T����N*�o1Y	���d7�	w�dI-���u2�e�����-!}@�J�<������s��gv�*�}�4q�v��r2�ٽa)^��s�W��@�,^�!Eʗ���i�mMh���b>�u�'�(M�"k��0���@n�1N�`��#daaJrY2��{7�-N�
�V�9]>�ם�����qi�P�?�|W+o�O{���nE�
��: R:vD�{%���Cx�^{%rvݎb��Q�_쬊N[�9ֶ+1B��SB��&t�H�"^�m�T�~g���I6nb��=�X�$G�⌥S�mDI��}�
@0Nid/�Y� 3�S;q"�_D��=��$�3S�#SE#	ZI�+U 	��3�>�?��C�k�?)'�!���V�c0J0�WB}�8p������`��>U&�A��!}a���+YŮ�8�1����U&���׍!�y��p���WT�o��(Y+_�) ˾_��Cь����&��$iU]�ͬ��o V�������­�
��0me��x-�Lt�����y�d(7���Vے����j�G͙|E[7��M�t<�̩7dN��7�6����-�Q�Xk�G'���ϊ��ۅ�;?��`�۬��=JP1�`Lx�r�H�������ѥ�����[��B�:�qؠ&�g��&�K���;<��������y��&}�9V��r���L��]���{nH���-�W](=_�$�i����rq��Ri	���,�^��G2t9I<M�^w��;���c�f��ER����'��U���j�J�g���W5��-SQdt� H;��� Q������kf�I;��AI�Vc+
�6X]��!�ֿEE w�GcY��E����h���W��)��-�-�AQ���"-,^�I����+<L�cf-���0�lL�$��C���!覚��);n;�����	�=�4��OllN1���ĝd@s/��K���GX<t�su�N��6K��x=j/�;;��������ቬ�6� I���������Xt��xԢ<�ZїD�o+��'>B3	�5�E����-he:���+�#a��x����9�x�S�)�M
?Du�E��UԄj0V�F�Y³�8gf����pD!z��@��DG*�d�a7��/�t�2���ߥU�=��e��VW�[������t�� ��,�Z�g��M��`�@\�����;ݡ����f��&��RuP�� D1�Q��`ȹ�+NL����s+�����Ĥ>��M/ z��+�����m�F΋7� �ͤs%@�a8,;t4���F0����y �U��(�n�J�*��eY;%�?x��ٛ�$m~�.�6�ɬ���ve�}�~��Z&}�E1E��>cJ���;��h�p�����{7H*Y���Qp��s4�%F�����1�X<�VQ��c�i@��4ۛx�dg���m4K=����@�2pg�n�x�ȓ�;e�:s��ՙ��軼��Uw!S�j51�ql)��4K��Nx��ژW|	{S�un _ϖHAu���MP�W�?XK�N@�{�c�U
�F �k������sK/�(��P��tټ$�+�F�	��9hl�#"���MR��)���&�[��Z7�
����/�(�N�;)3u7�!��ܛ��!��g��m��-��|0#�lz��A�k�L��
�5s��n��������K�+����\	���W�d��W����N��� j�w�pYM(���/�gi�5�}���Q_r�WR���H��B��]\S�p���l��[��cR���<�/�U�C�bc� ����/<d��&�Cb\�p��L�lǮ��%!�G��y?��&������j@}��2� ���N+5��H;��D�>���u�`���G5���W~��':�iZ�)A��-��)c4�e��7;A���M�!��u�]���jY���(iU�Essc�e�v�U΅ ������z�Yieja��]� V�G�iA&�߇��(EOy����]��*2�wB�G�*4�M*"�-$�BӲw~X0e-/D�K�u����f���*j����)cL0IAr��9_�O[ E�.���u���8��Q�oR�QZ\���`%%lO��խ;�%VR���H�Ul�V��e}#³[�[f�π�Ю��̥<�;&�h��u3�©� ��6c����Ï-��G�X�)�"���98(�g'�9B�T$������l��~�.�}!��A6�[*�3��Ǖ@k;�:�}���0e&�|��?M^�n�y ���&ɹe�g����3M<Wm��G�3_��[N]u�q����w:2��p����:�Nq~ӾF�>x�m�+��Ϋ�|�H)��h7��2�����B���r�tˡ�?���=ٸ�Xl�;E�E���ɧC5�LB�	:�O�&�
��{ڍ���)����E:Z�Xj�T����}����R�N���s��:��J�"�y��Fb?��I��=ڬD�*�`���?���QمU�='�;tz��жXu�e6)��������Î0p�,�Z��;�y*ccq"
���f`O�"�^�Q�8q���!��+���Jz����p����8�m�]�g{��bRV#x�=�s=���[�4����Sau���O�s�:�QgB I��bky�9>�+E�r��)����Wvc��a_��2Z#p�Å_CB#�H65Y��e%;*�tf*_>M�3��kk���i��m�W�F�DK��)�!��CT��$��c�������U�WWk$9��+�j�pH�:�7џ���E�iQn�D*��{�>S���%)�Ck�d��@s�)[��}�#�[���	���t7c���'�\Vٸ*)wm-�/�4�x����| ng:�m�2j����+��ڃ��qW�e�*��YA}6}ې�, �������Mѭ�<�!�V�G���]����O�3�e�M!�|�S��^����/E;���H��_L��M�
� ]���R���N�PU��h��d���6�u��s���B\�C^����Zf�h��9b'�$3߬���TB�%Щhп�������Tx7����d�-k�u��f�����Ls}-���@��+<Rz��`�k�%o�� ����v�2w��a$DP�It�.Wk���O,�	"��_Z�Xh���mHY .�b����B;�M]��k�っR��a��i|n�,5��ʿa|�BY�1�{NI~�
�jT9X����)���q�7��0��Ws�o���ut�E�\{��`:�Jv_�%��CS��{`<�)L8�L��G�[�0�9��f1��Sq�&��>�v	�U���QgJ��IQ���a��X�:�G̚����h�X�%��ŝ�N�y�ԲW��Sv4	��n��8W��na.3��nE\	�L+0������h��׌�n��?�!&����0%N�b}o9/��P�<���=	&�(՜�Е�+��i�Ӈ�,�����X����N���K�֒C�
�0�#1_5���w���I�>�E�_�U�،ͧQbo[2&°�����l��˛�X��e�.
x(%tT����a��$�T��m�����jC_��wP79�/Ŕ���d��^��5�5��-���SA�G������"J��D�v�n+����r=��JP,xLӠe�����`�LL����\����B���q���Rs���ԯ�<Q����@k�\�"�M}(9���r�s��g�]$�{I������(8a�$Z�X�eSq��@i���ˣL^$&��rI7И繂<��3��Rg�&� t�� h����UÝe���J�GȆ�d�5�S,1��[�D�gT La���yk�s�IV��A�zc�76����f�!�2��2�w]�YƗ%�x��h��WW�j:�ks-�:z�&7;"�$w^	�R���+�c���Ň6�g��@�CAY@!-�'�;I��XF�v4���ʗ���O'��1����@N?d/�1э�S�ާm+�	�a6f'���
g�;�K���9��@��7�g��
3�[������-���ђ43o�r#'��	�gɜ�k��0��e�T]�&IB��3Z}����E���/E
`u��ڈ����u�<76�tʆɳr���tb���z@�@�8G�2����B��"tp������6:=��
��W���e��7R����J��(뢇tM�'`�'9\tHU��_�9١�3�A3*�a�ER�S�� �Ҥ״}y�	�"L(�S�NRȷ_�5��./r<j��ӆ��jXm�J��-��%۞�8'�4+{�Xy��Pzy{�����Mnc�**�Y68����-���%�.7R$�%n�	*��O�/|�e�[}ف�Z��ǖ)��E#S�c%cE�v!,��)k�>�U{��Y�EQ�Z�sd�F��,���1���ϱ���Di[�V���x̍ug"P�  =�ZZ�G_2+Q�n���C��;@��s�m��4ב�ơ���S���1�}T)c�K�j���3�r	v(����%_��A�)�� P��)?H�>���¨ܷ�l�
}.F;���j�c�/Kj/_�mȾ�
�l���+>\�	����ܢ#�$x���Q�ġ��!����30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�%ڜ4�z^��2�Z�n�;:�|͚�<���͟E9F�_6���(�(F��Z$����8#lfuP��Դ�I��O����Ŭ[:v�,�82�B'�l�(�,YB��F�2�%xd4��o����C�ƶ=wS�%һL>[q
�\�������� �1}?M6�h0&�	 Ic[:������  Ll|�A5E�Rv�/�h��]��
���Y�������le5H>�Q�핥�'��Li��?��?�.';.���Hs�o����=L#����ިa0׊���[�1죪Q�)�0����m���獖l]v�%���6騌 .�~
�J~ :��J�?ą�@vW1}[I���Y�G���w�qT2n���_Hw�V��Ԥ�M�z��ް؛��eB���b]�=�o�f*�.�_��e�b�Lo��n�|uwAB��R�k*�H�3��<�ێ ��X=۔�,�͠����
Z� 9Qi`N*P�&�nI+AEԌ.I������bWӔ�iW�(�G�5;����&E�C9"DDtl��s&ۧM��(]'FxPF�Q��їCj��ȵ�f��.T��b)��^/U/P4rEu���K�4A.RI�1�I�I�������Z"����*x����پ��]����[ʸ�1�%WͶ�T���62I2<?�ᖜ�M����V��|��%Quc��^�7��`8�,�oʭe�h��"���������^)�JCX�p� ���울���Y�%���O\0�����x����e�Ɓ|��Ӄ�M[�Je�?�t,�E����fӅ!�kJU��WZ) V){_�p�����Twz��$% ��/��lc%f��.3_>|�daL����1��9������ul�Y^t�{��a�����'�G�9r�h~�Dx�G�,�<���;��Cޫx����H���� %{���<C=I֘�͗e��W$$����.D;� ��EJ�w��8+־z��o[�Wp�Ʀ���w�Q�:��k�"�H^q�z@��R�p�
JV+�_��B~��Ǘ�/̓:i�X��R�x��boE��tj�yf���EЪ�.+k�|�ء'�!�3PsW��<*{e�G|�aO. g	uB@�<W_ա���)0�{N* !�d͜�ʌ��Ui爖v1��bן�� ��]�yQ������T�U�N�}�'�F�&D�/a\�l���#8G��4�_}�����<��r]���/a��4�cK�,�}�"5�	����YS�<�5.�6H��nu\���`��V��� 	MriN���v]YZ�����-�:ٖ�	,{	�����Ǐ�p���_�$5d��Ph���5��*�^�X��{�QY'��
�Q-��FJ;�+��νi�ق�Z����\��U���<Jg��S�-\%:��6SN�Q���hGӗ��g��{U�_ �(� �qc?2����S(I�=#6�Q�����I_��q�ζ3��C���4��K�L�����3�y(�^�/��X;����V�K�����E�x�\�L%�Kf+D�X�@�}߳��*V�I������+�%�K�����9��<I���w���r�")�|��Z �c l�)�-���C�1�#jQ�t����ـ��~��k�_�ϖM�!��}�Offm��w���П�J��Ρ*!cQ���S����f
�DKZ��x�TT�T�T�"�a]�O�"�r8|��_�\ĥUm��0�έ����-|�:�Rt��dt6*����z�t  R	l�_��^�Y�gH�%�7��N`��i, �h�k��t X��Vg]RYl�{����S�gA+5���t�kD��#�{��a�ak/~G�A]���Yu�Z�}�,kג�!����峪	��\e_�^��(z��ɡt���z*m*��,�yK��ې6���(��vM�G�-��K.`��<c�7��������HǶ+��-���Pͧ������a��c3.�V�/	��2��G��á=!� �`D�-��jcU���x��(��n�~�M�%46����V�v�BՀ�ړ{TT��I����B��7��6Av]k�H*/^g�虐A*�1V�Z�51����ex{��Y`]��A� ��o���d�"WU�������nˌ�H]?��".E/N��.ze�7�:��D����V6O������`S�D��ez��7�~�<�!���Ȥ!py|J�}h�DQ��|6q�u,^��������������V������b��7�� �-#�[�����gR��s��x��z�.��2p��j=�����&ŹN�Ղ���TqC���׎�g��R��3�.�Lw(��/�U��n��|�� ��$RpV�}��d��!�Ҭ����Vu��I�o���Z��|0u�yV�:Ç�(��QA]>�+�yd���gW]
y]��ȩKc��2�<S��T�3Y8��;!o�7&U` �q�S
T��ͥ,�Hd'��-OV�n}�`�v���A���BQ�O��i����-����h�̐>��~�n,��ĺ[���K�����k`u���5��#1=���Y�)��6��3Т�p�uG����'n����[��BJ&�񊳒V�2O��p��jاn�\�SLU��2%���}�7�i����D@�P������q�Tg{�ɮ���1��?jZsax�Dd�"��Ǖ���Z���g��f��0o���~"�}�����4��`ӗ9�|͒Q�_I�ol�@t��V��� fRiIa�i
mΪ|'0!�*��K�aJ5�ڼ�7�TI8��D�2�њۼ{#�~�$����b��T���#��0���ч�##�(è� u���4�����!�>��0�,�U6D�\��![������k.V����·R`��0���נ��X�%�������h�tM;��q�B����%i���>)�m�h�����P;rG���N��.f�v[R U0r�>vބ� 
)�M�u��&�As�د
��6�gP>r�n#��AP��?o�i���ɴ9l]V��M� ��[��`�e�%
�~8W�l�i�
�*�p���[E�M����$�e�9�*2Ӟ7�_?6�.�?�(���J�Z�W�%����L�6�m(kl?OG%D:�Ƒ�{^�̣,u�ڑwjL����Zy�l�j�n�;�����*�ĵ^9�f��ijDv�e��ca�eL��6۸* ���� ]���]���"x��lE�������C�Э �W�%?���Z���~SZ��;���:9��X�
e:������Yn(��AZi}�����l�	�������4����&�� a��q��8j}�9� BL�#����Y�R�F���%`����o�&��m��ۃ�S�%�� �|[v��\$������W� |�?rяh�%`	�Am[?�@�-nV�EZ�law�5ʉ�v�
h{�y�롤���Y>�U�D�ݣ�$�5�3�v
Q�8YJ���]�9���' �PԀ�6s
}kp�=�ڊ�7?au�堇s�
��v��e��W����;fv�So��-b�-`�.��7�G�:m�4�OѪ�*Xv���[.�V�U���l��<ĥq��f� 7gHtF�ԉ����)!���NЪS���bbF�3~*�Еz����bA
o�On]�wF�i��4�*K�
$<�sk۳�O�j�����wkjo|�U��ֽh��Q����U�L�2)��A�?��K��C�f?��LQ<�p�#�mW�)��+���,�y��$��.� ���-8�׾�]3�+2�z9�},�<<"ID���F(e8J�]���{ �)[�����sP�ux�[�{_��PuX�����G�Q`&z��6G��T&��
�C�>��?���<�T���5U1��p�H{���z��}��$�~�S]Ȱ<F��NϹH���b'q�:\
VRY�R�Y����F�R+��X@h w�D���Ar�
��&�I^C��Mu�*۔m�f��۠YozŐ��2Н����~mX�@znmu9i2&ň?H�g>�m�G�J�����vN�_Yz����h<[T��u�C�G�3�Lz2��8�xT�!�	o╠XTk*���ԕ�S��65_�J���!�/efŌ��K;r��{�C��*̮��|����i}��y��߅��2J������5M������?C��ق�-�:����+�7�br�&C�-���X�@���@T�
+R���m0�b,bR4�ǡct6��kQ������֯wzִp&��)@�K��J�%'��L7a�=N$-ya��fw�]G�#�^Η�'[�B���t�c;�d���Jƈ���(뤝G��p�����cf\t�5F��N3�t�q#=5�g~�Lip�[���1�h��a����Ք��q��=����&��&����kߘQF�ʝ��/Z����	�{��$��$E�U�����5iY�I������A$J��ɑj��&�c�cV~���#��I_6��@�|�"B{�����ڙ�~MLAc 3c�h������1=jyO@��W�-PTI�:�m�㵖���C����'���%<7jA���ԣ�2�D��6���j�bNw���v�r�� @I�2Y���P�D1�,�A3���q����Z옄�Ԯѹ�OZ|�Y�-}�E+�aq�1����s+�!����GZ�Y����	q+|aX�ge�3�8�4�����/m����UGB{@���#��3��&��+����D�u5pQ�NT�@���e��GҊ\1K�.��1�{b̋��0�/&C߅nާ7���RCh�������$����K]��%vX5C�sW���x9�'Sx��-�d�� &���
�Ć�ueP!N�Q���	�3�q������ĺ���9���ƎN��31��`��c��W�p� Ih[G��?^ ��`p���P�u���Fgu�6�M��:D���1�������u��:
�G�X�F�B�O����l-S R�g#�f�}���\�0�}T�O�c7T�@�P|j���/)bZ�5\�� ���*����ܶC]D�)G`nA�a�ʕXz�#�ۻ��[�������#ȀOc��C8�{�^�̘��O�U�f���j�r�I���o5�g�m+�mjj�D�K:_ݕ�q�Tè�DT��@�緑��8�N<j+��ϛ]|q7����%aA���u���]��M	D.\H+�W��V'R���G��iC?�VN55��T߉��"��n��C'ch���?Sk�_�l���J�"��0�	oO��xo�^A�Fk}�B�-P��G|�|�٠E�4��{#�x
1���J
�eiN:��V����Wc҃#��)�6H�{n��RY/�Ĝ��i8"�V���52X���xg�������coŒ��Gak9f`lI�u�JR���0�R�O��yx��6��kO%�b�ǽ�|y�E��j�0t�xZqe���
�UQi����+�����E�� 
���}*���/���{�F7���{���^�~,j�/M�21���$���q|���p�����ĺ�^f,t�]��]��C^���������O��H��>kG��.[5Jn�V�ri�ԯ����k7�����P����kN��xd�3	X���%8I��DO�:��rC���(�)�r�.�ѹ�}:/�����5n�r���~~��Ӈ�e�u�:g�ʟQLL����pm��A���א��J׌���O\��� a7�"�u�����91�&�����AVO��4a~���MF�3^6۲�ַ;Έ<���f64�G`� ����WH�v��Σe;ŔE�o������L��=@E�V%J�H�om H�I9`AѢ��σ�d�#wBڈ������b����v	p;�@��'ʹ�08S������0�����{�A�e�ak{�����H��r����O�� m�PV�w(���?�#{e�<���z�O�54���Vz��;��h+���S�
�QC��ƑW(�'B��AM�Nk}�4��G(�X���q�BE��v�
�/��)}Z}���B�&�OWlN��eW����9p�
��oR+��T��hd��N���3W���\��0�F�聧�1��%�"��d���	�W����ˎپ�����19��vbʋ=˂���;��E������]�(���ˮg^�'�38�Ӑ<@]*���R�m�&�}�8�=>��a	��Xr�hKS����Mu�|�$Ŷ[|߿.�@�LSr�X����넱�+#H?̇Nz�c|̿���U�oj�1Pٙ��Zmg��1̴qn�F^���=
�&����AÙ��Vޔ�*k��B��s���t�xN&�I b8�)hW�0�io!|�s`��J����Z�$�.M��ݎ�ꗀ����z��+a�q�Z2ڜ�S�0�M��	�X7V���=r'������tp#?܉�ք���q4���Up�b'��,_y���B1��/�'\-49X�b���oE��&i�$d�����<F7,��{�R\݈�!�z�?�؎To"s�h�s�E�M�r�@���@�B�jq�`��J-Q�p������;�N{�Fp'�zd���Y�B�3�#�
;�8��zR]���-����*����B�լ���?Tl��\@̜6r*�����JϔR��� �� ���i"p*RX{���A�lE.,�ׁT���WU�i�>�I@;�oA��?�C�ZcDF��'w��)����'Hq�P����t.%C,t�ȷV��T.T�n�^1�dPvh!uC�F���A0�M�sۋ�DV���)�s���M�q�x���(����q��[�M6l�%�Or�����a�ItǪ�c�y����������`j�l�|ue��^Oo��������kb��v"eU��D(.����^k��Cڦ�p~�����n�?IY��]0q��7�:�������ƃ���F��eCJ'Fv�vߴ��&�K����JW\�W��V���_sm���x�w�g�$�1�1�l�+Ӎ5�@_ �d��W ���^9m����8l�<��7��=Z��cv��i�'V�)94��~�N��L,���+��y������WثE��ϟ g�o�-1u��F���e�m�$�����.F	� %�aE�*����:-�z
��[<s��}��J���c�q$M����H`R�z�a��"|�̣�+��ԄP����Y��̕�1��7Xt���:��bq�mԶ^Py��Tf�E�O�.Vp$��׺��NA� �cs�Ӛ�-k{'��|��A.B����@I|_�ٶ��:h)��w{e� #d������QU+�_�xKa��1��8�t�P�yS:�����ÜgUN�y�'���&��/����n��]�%GY��!�-���W<�z)]>2a/#�4�r	�n����1	x�(�[J<������0NW��趖%j�"�	��N�۸?�Z:6��������<�{�4��V�"ǑK��䕑��Z�m�h�|�5Z=����� ���e>�6���؞���Ja��+m[:�+@����я�̎��ŗdQ�C�J�8z�ժ�\�+��8}Ф�J������\����� ���(E$�q%��2�������IMR�6R�����'�_�gYq�ұ�5��CH1;¶.K�+�L�A�ط����5d/��`X}�O�
/HK��y��Ԣ�E��\_��%��f-��X�2�}a�����I�ҭ�4W>���%ygp꠳u�N�������Āۛe�d�D�����kcv]�_�-�6��8��JQEJj�Ug)�Bx,�����k�Q�Þ�	}�؟f�qǗH�٩�P�c�GH�*�%Y�C T��e�fL��K��x��×V��d��a��*��R�8~���\�'�j�[v�ί�u���T���R6	�fF�x9�]�n�6�rRL�_��^cBg
�j�9����+� �,�Y �mf�tbZ���8g�cl�ٹX����uA�V���&t4�#Ɵ�����o�Σ�?/ e:A|��
]��$���-���؍�/ft�,������`M�(���#t��o��|�mmlY�,`[����n6��T(J MJ�!���$M�9�+�Dc~{��cb���������wb�ϫׁP*ł+�瞄J��>a30���qڲ���Ϩ����`!�C`�����jeE��+iO���4nV��M�F6>ޗ�\��o�K{�f���ꃆ��9�G6��r�f�H�jYgۜ���^f1؋:��}�뙟է�X���]V����O���q�� �"Dn�����N6�]�]v�"0�C/�|.��u7���F�*�6 �O���\-}�b��D��e��7���<�BR���`�&u�;@���DD����z��7�����굳� �2ZK�V�����b?��OF,�/m��F���0`�)Z,��s-���������p�/�=SOI� ��{���d��v@�G����i��R�93
t�� ��1���'��l��>1� ���R��N���$dRłDQ���O�أU��5�����2k�0���y��:
KE�j#Q��V>���2�6��g�^�y�9�2hK��4ʴ�=S�`�T��`z�뽄a�BX7 r�`b�z���S����%9�n�#d��-��n��``�B�o����Q����娵�"s-���xX��-�T�W0� �>���*X�̷�@kR�@�f��րq�Ef��=�k��EB�.ƚ��nPi�Yվ�ݑs	���K�{��_|i�d.�/��
@�r&_G�j�n��)"�.{�- ����N���CU�/|��
�􅭨�<o�y�&��m%��0IU�����'k��&6wf/6���g����<G�����験6�;<D�]�"�/��K4�>�D���N	�}��˗s<^�(qKΠ�� %�q�g��:n	aNc�y�(�uZ�ۣ�0w��/���Ewo{��V�Ƃ�����u�&�
��uhA�%5���v�񽐊���9���
�_����Y;>J���+��]���A��p�B�S���G���]@JÅ�E�6\W���1��a�Z����L8�bC:��H(�l�q�)�2&���UI�R�6�Ѐo�����_ �q�(��4C�S}�&��K:�'LfN%�H���k8EDl�/,�uX��z�K�u��_������\�.�%�.�f�jXc5r}�>��\?�I`����s���%�}���e�����.�,�H���K8��Ըn0�Čd�c��b3B�-w���uk9��Q��%��OXٲn8��NWN����S�
}-U�f!�����9dX�㫷
!*6�����RAf�
�KL�px1�N�Ɖ����EaO`�T�8�h���ė#v�˼��0�2�r危�R�	���蓈��m����<R{��_A�^Ӣ?gz#
��V \`9d,2����ZWt����<g��l�T����E��A@�{+�t��k6��U��[���>/p]�A��"�z1k'���o@��t�#e3Ο�˳��3��Kx�Б�(,�ɓ��&�Ġ�Pm��.,�3���}6�@(r��M�w̺_�!�ʂ���c��I�Ӹ��U0]�ha���bk��Pxs��L��=�G�3��%�������3�-��5-�!L��`6]�=E�j�I�ܛ����3n�usM�X6�.�H��t2�!m{i��;^:��K\��'�6��]o�H\��gK�Ð��	1HLL�gL[6#�(P�x��]��t
,�!�صV1�"����}���~E+]ql�"�W�/ r.l�Z7-z�����*O���̓�����DaB�el�7Л<\/�?A�Ȗ=X�6��HD�U�n�	֧��Yw�Z�8��Uʑ!V(L�UP�bx/��D��9$���փ�ث����5��*%z�l'����p9l�=����&���iGY��@�kc~�"q��i�RR�@3�b�~Y��Z���&�`�w��C eһR"�a�o��d���u��PM��HT�{T���@��K0g2y�J:z�����Q3>����.�%`gI7my��?���*K�M�$TS��?T;H�{�-��G�U7��~`Ҏ'�!S:��؇>��X�dI�-��Dn�?�`Ч���?�+Q�;�U����J�-�?�|�~3Q��w���r���ͺ/��m��'M�k�����5��rUZ���YvgB��*�ե��t��"〹g����W�u#�na���q!��ƚ&d��D�12Alݻ�a��ˌn��QS>큀d���Z�����i���?@F�kj��������;],��{���RKZ��{���k"ɘ�����_�Z�gf$�f���o_M��"i�`���k4����	��|3��Q Io���to���� X2�I��
�r%|�E�!^��E����p֌�a7
g�Ij���	2�f9���#�75$#��֠������������0q"T�y��#��%�t��ue?<4z :��5P>^R_0?uU(��!�����Wk ~U�F�0�)?@ϽJ��vM��x�X�)�4i������B��;���N�~���Wj�U�)m��hx������r�O�� ��� ��v�e�U��>(�I����!�x�_�����E����>$q#�/�P�K�o?��h��9^vڋ>�T>���&2�R��e�]�������X*�=�S�j��[���8�e��*���7�F6��L?���~c��oJ1Wq�R��w�^��Ln��m��?���D��������^+���tL��>�ޞVr���2�3i�����^����rOj6���>�0��X���]�\���Y ЋD��b��0�x!��E����%��6���B� n%1������I��Z�I�;ߡ�Q8	���(������ϧ� �(]�bZ�࿉Y�l�E1�q���|�&$� Ьr`��#��8	c�k��B����nmY��F �M%��z�	�os�������M>�Sb.
���[��U\�){�i�ߟ� :��?��Dh���	w2�[q����c�����lS�h5��Pve~uh-�P��da��&TY��N�� ��5����躤d>K߿��(��6�'�Բ�ss��"=�A�$����a'�P�y���:������&��-䍭��v�?��ˏ��_ x.`ip���C:_1Á:(Ĝ�7vNR`[ �b��C��ވ��ʭq��o�2��H�U��-�{��1��G�\����9vb����f�*�]p�m���=b���o{z�nO��wx���i�*�~Ϗ
��<�[t�%�u�� ��Rw�5|O��ɚ��Z�QֵT������)��sRt�;ut��B�?��	Q5Hu��#�N���q+˾�,�fޑq��=��D�I�R8�J��O��+d�����}�
�<;���0F��Q8���]���ʭ�)�#����'sB�(��f���9�=��`T�y��`�뒒���rꎤ-_2CH��hM��߆+��e��1~LLp��K�3�z�ϝ�U8����~D��]:�F��Z�̈��z�ԥыІ�
H5ӓ����FE�b+��Xr�ww#���DAd6�z;���y5̤��m���\�~���ł>�275D���@�0�,�2*�m��B2�9�?��e>�ƍG���6\��(Z�_K��ݫ�	Tk��u�n�G�1L�a�љ^�j��!�r���TQ������1<Ũ68��1u��!0if7����r�h_���"�O~��h����	,�`s�m6Ue*ҩ����E��'�M�M���a�qKr���_r-ﭶ�0�R���b$hFC���s���2ǧa�s��o_�̕#0E��b��Ǔ��th������������o�����$�@����>%J�)��T��a�&&N7+�-�fL�]�w�o��U�<�	@�[�g���/�cGT�d:�������(G(��plʾ�t�c�����#� �dt}'y=g=t~1Gpz���ː���=a@�mʇ���c`=��=sI9>��s�ɘ�{	�Okd/L2��-��{O�@$zl.E�X��@�����T���>��x��LD
Ɗ#yM��qrR�ז3�&z��y��2��;�A����{ �kRcS���dC��ZZ��{�)���|>��k����0�D�y	_:�G���oQ�[>�U���s�D�g�>�y��"JUKִ��$�S���T'�M+�)뎥^�}�71�`��V��1S;:�ب�٥��dz��-hAn*�v`��z��p��,��Q1io���2�Pő-}���%��?����:���:��ƙ�N�)��̨�k(n�qY05v�CV���aY��Y�G�VN΢v��ڹH	)��X��D�n�������E`�&�i��h2""����N��}(nδcS��Ҁ�E���,Ȫܝi��a��"�@g٣�,��r� �����H#Ȑ۷��Z�&���A"
�Q1o��j��Z��g'�@fz.�o$I�2v"��a��Ѝ4~Ӫ�F|@��2��o��t�1��@ �4�I�2
���|�8�!����q��^%��c�7k:�I��N�W9'��Ԛ���#�O($D�:�᣺�}�rG�6
�02w3�Z��#�|-��s�u�J4�u�|W>���0 �9U	Xe�!�E��){k������,�ʡ��~Yξ����X1�j�u���)��ï;�|��61_c`�XF��vn�)�c�h٭��A�{rZ�����ۉOv���U��B>it�sa�� �D�����x�F�7���6>eP5#��Pp"�o�D��)n9?I7�?�K4M�����0Jebmf��v<�߿����*�Yp�tk��@ ��Ae�e��u*Et7F#�6s`�?����
򰟈W��ys�����L/�*m���?�6D�c͑�@�iR���Vڤ�7LY*_��<ޟI��R��t��#��l^L���3v�j��?Z� ���XZ��p޸�vd��&i �,d���� axBzE���fͷl��`� /�%�[��U��j�sZ�;r��Җڒ/�%�}�����ҧ��(~-�Z\Tٿ�<�l� J����N)���@�(������d�v8j�ā�53B_P��`�Yz�
F!R$%�j$��o�!��{�\RY�#I�:jk(M5���z����ӑ�{C~�y]@�F�)�R������ڍ&��o�
�6��6��lF�+wb�X���w)����.�A�]��K�c�8��?w[��3@m2��b�є����2}3��w�����۸�Fm�K2��?��_>.:�G1��<�%��g
_��OYC���LT1�u>G&��L��љ����h!GYQ�߄T�7L�P�����Ů��������!vw{f=���EQrjN���A��U�Ѯ.�8�BQ�U�?�s��+�թnߙ�\D��,"MK�-1bշz~�.VQxG-u�.�v����Web�s�CN��Z�����ۧ'. ��Ǜ���0K�Nb�Z�4�t��"�g����W�z7Q���[��@!\≄J�3��*_au�<N}?�-��n��wf̉�����[e��v�c�N�d}����(c�?G.�p2�cd�c�g��&����tj�=���~7C�p@!��Q�p��KaFG4�MV���|=8�C,��tG8�dgD�ɰ��A;/����s�{U�$@�fE'�E)v(O�/i�����w�1�C�R��$�1#�	ǁ��΀��v~�x�ߛ��01u6R���dPB���˖��R�~��4cxː���X��ة��yǌ�Ϝ�P̓.�3��[~#�pi�Iϟ؟/����cj����L�F2!��*�<��Sj=!�wFo�v{,�%�� ��X2�q���D�NB�7��o%�C0ү��%d�1��,�YO������n1'E0/����+�CG�pY6̛��+�։�߉:3�a4�ʧ�8���X%Y���C�8@�i#���31��ZFL�8�D$x��ON�rW@oCqeZ�� �1��O�d� {�\;Co�ҧ���o��D�V�h��O�����Ne*K����{_�9W���i�k��9EyZxRv��f�W�y�`ٙ���1�e��~N�4��Y���'��c�<�O������NR>3�� `+n��	��- I�G�� YxR�ةg�\��u- ���	���n͆�F:�뙩��.���M�up�Q:�ozG%��F4�O�+O��=�{	g�K1d� �Lf�\V�}�v�Ou�#T"��ȝ��B+')ڹ��RB\X	�g�����fM\�{ �ՌH)���n��1�B�1z��SP�VZ�o�Лi����D�wRN���D������U) ���F�!��^��5#Č��n�  �j;F�K�j��33��񑯼Q���]ַ	;x8#��j������|�nt xĝVR�8���n偼H�	�[H��4�G��R��Ŀ�"i��oV�y15u~�Ws|;���ֻ/ac�MM�D�lk��l�C�3,���06)�Ob$x��E�	k��V��"��UD|�DEL���)�x}���/,.
عiƼj��{���R�E�
�ۡ�r������Q�щ��;�7����ޡ3�!�,��M����$��7q���sW��$l亦Mz,�y��	׾�_~��.���3���+���>.I��Q��J�J�U�b��f�1k:�\�㬶������Mʣ��HX�JR%��a䥟����5k��I4�ǵr��4��(G:�n��X��ܘr�̬;�~��|MZ�Y�:
c�TM�LD-�3�F��G��a����ee��x
����ar"�֮��!�9��Q&�7O����]O��Ja�@Ǧ��3�"e�G;�N><ɋ�	|M�JZ� �f�޵H��G�Q�J;�H����4�f7�L��N�2V��H�m�6n�0�9�עE����N�:�Keu�"5���d�ݐ�p~	�e�wf���S��U��x�������[d�A6Ԁd���/9��a��?ʡX�
�Ƞ"m@��V�|T��j�Ɇ4�c"D� ���ף玤'tV�$;��h� ��i�-`Q�i��w�(��\�a,����}T�
4r�{,���bB�]k���L
)��,�}�kxBVE~OzN*�%W�%��|8 
1�RoU�_sɻ��md�N��J�LW�k	\B?/��M����1]�n��Vd�rE	m'��i;7�}��$E��FK1���v%"�0�Ԃ��� 3Ƒ���A����]ЋP��k6%*����(�m�]�N�������[&���[�=�\�D�	@��r|��S�dJ�yª�
�A���I����@��rl�����.���#�p̪jc��ٿ�0(Ę�&�P9x���UZ0�T[�q�"�^{��=Mkv&0���a�!���WY\k������s���t�k&�`�Т8���W�����o!��ts��:��F�Ũ>W�'�MS(���2��������ރq6tu�?!���FM��F�[y�L�a'��w�ɔx���?���9n���	4�kU�AO'w�b,_C�y��ȸ^YG[���4\����!����ޥ��$��>���p�dF�g�Ӟ�PR�����܂U؎�|s�xּ֠k�,Y�c�T�ý��M�`�p-��U���~��2�q��i
���LzGp�ٜMMBs'�#�rz��A�z�t� ;Ն�s��B3�L����TϹ6�ȃ�Y�ҽo�9��_������e� ��zi��*���=AJ��.�s������!WX�_i|a����;�ճ�+j�C��D��
��6��,m$9G'2�P�� ��+C"����i��hT��N��^�^�P��iuƤ���csAs�U����j@�;y����72��M�T'�x�nJ�����54���[ҽY�%\����g�;�@IS�f�w�r�>��'��3����O:u�r�^��� 	��Q�������#�"�qȫ'լ���O^.vC�L4p���u�{�b��Y���@��0YM���5���N�����FD�8D�R(�J
Y ��N�*L��N.��FoDJ��W�~�V+M_V���{��Rw�E$J���l�델eU_�-dRmر�=��ѩ9�.���el�@csK� �ݦ��ƽ��'Y.�9�pm~��V�͎�>���{�������Ot� �$������a�'9�ev�#$��	�.	�� HY�EO�̲��.p��z���[?]��C|���a���^������PH��*z%��׳��/U�+���ԧ�v��\�<�
��WN��Xwd,���b4�z��g�y�`fb�>E�.�R��X�Lf��b!ߐ�� ~f&����[Y�2C����M���1�Ս��+�C���-�\�Li��Eg�b@vjC/���0x �N�'�}k馘������0�Bb ��/7It�C6y�t�ֽ�ݐ�[����~4:��F@7��Z�J���pS4a��NSa-#���w)�މq��Υ|{[�7�ڌNcc��d�d�r���(9|gG���p��=y$c�*��C�r�͔tE�=�~�;mp�,@�g>���aܚ7ʣ��-=E��C;U�i]d:�_:j�k��/�u�I+�{�h�$���E=����7�W#i�zT�׫Y�Me��J$,�_��tiz�ql=~� �߱���G�6�M�JH�B	&��l����~��c�l���$�����6yݐ˥#�Pb�O��q�#��qm��$������:�j�����}#2w`i@̝�[˂jӓ�w�4-v��I�TS NQ�2'��2D<K�͠(����YVw�����
9ч� �m�Y%Qk��݌/��1$0���/#>�j��G���Y����.+J~ͪ��3��,4�:����nҘ��Fy��@���@u3�H���Z�c�~D:q���jNb��@��Tep�����1Y����{�u����=k��S���5�>�,%�h�'��R����{��$RK �
�d�:棢���"��m9���xh�����3������v������$�e^y�Nf�3�����������yR���UϜ�l�Nrx;3��`�����>�4I��Λ��� �af�.���r`�u�I�T���TB͜1�:���?Ҙn@����uF�:jcG{ӖFJ�O�&��z]�g�^:[���\t��}�$OK8�T��t����X�)���ꗸ�\�B�}�l�x�������y��)g QnOji���\zn)l,N��Ŋ�@���v��%L����U�]�Uj	j!ݸ���3��59Jˢ������j��K�Z���Ƣb0��c*�Ι���U8��j�`��)�_|��!����]5�Ny�DD�޿�	�}H����6�R�V4���iу7VZ$�5�(�+3����;��Q�c�@��Z2k�l"��"��v0�O�:<x=���$�k�5J�;L���x|3E�]���vzxӾ��E��
U��i\d��$���7�E�\
^�H���a>Ԡggd�t�7��䴟G��j�,��M+AZ���$u��qu%�������߫�<<0,�:cѕ�¾��睉xW�������� H>�m@˧LJ��+�`Ԉ�|��<kP\���'�Rx~��#�c"�����X� %18����s�������b�f��<r^��ђ�:(���D�n(
rG�G�" ~'Iz�R���{�:`c��j,tL��ɷ1�B�>�w"��"��{Э�H.ʣdaHC�"7	��4��9��y&mj}x���A�O՘a��ަ�"�3ם�#-�;���<_O,�_���`[ ���}�H�F�g��;~gH�H�M��c�L���y��V~�Hb?�m��=��Ĵ994â�����q\'���o{�x�����ﳛ�po���ȹ3=��	SL��̉4���Јl����A�$|�z�v� ��]���ݡn����-m�_VV߀�����\�[��țvԨ�79��S6��.	VszZ;�%�hd��W�ð�:Q���Z(w������}���Ly��W��
��B����Oc�
���B��}�?'B�O�7�N@=W�����:
���oki5���>8OdQf�`��W���\�ͩ? 7���13���{�ed�L	����?�6դ���z��^1r�Lv����f��u�xQS\�ž�����[E�a���]{#n���:�^Đ�H]#"�;����&3Xz���=���*G	�A�rҢ�SZ����f�.���ȶ��T��>�@�t�r�{��Q���h#���� F���b���9��.�ec��P+����Z��̪,q^Q&�=��&��A�-�z��� ��kr���3sq�zt���&��2��8�i�Wx1��6!;s���#a���H�=k�M)�X�5{�� Y���便q�o-ڕ���3��M�<�Q2�Ϣщ'x��_���m	�?,��@<�s:4 SU	̼'Mā,���y�/θ+
ގ �:4�.���a�������~��'��!�ņF��W��R���ڰ
�)i�Mùs�꠬���ڵ�UG��i:�#�`��-Jش���ŵ�R��U�迁��-z��2��B�Yv#��I�qa�z���v�ۆ��Ə�'n�w;B��է�ҊT�O�����UĽ�hW�V�o�+Xf���� ��]i[��*�y՜)&�A`H�.�z��!���,Wn��iR㬮��A;T%=�A�WC�R"Du� AA�B�a�0`'�$�P�6�C��Ȑ�MT�c$f�^���P���u�J9���(A	:��l����+R���un�c���*Axl(j�����(��h[hR���%r����]��t�Im5(�|���H��E�S���4r(�%��u>�^HƷ�6��'�%�7�#7�"��K�����2�^d�<C���p��7������[Y��߫�	0��5�0㷼�*���C�ܰ˸�Cm�hJ����O��V�d3�1J�WLWt�V&��_,V���x�w$ +VÊc�l���λ_���d蠌�P����B99��7�Ot8lhury������<�6�'oU�9mz�~%\c*����"|N~��s�����]w���� ����Ɗs�Z��e�\$�zS����.�q� ��Ee6�i���z)�[U����+�ZH��z��
�ǝ��H9]z{�)��R�7o+���������}��n|$�0zX�6�sq�b����/�y-�f8<�E���.O���z��"43�y�s���!n{��|�� .;�k�o�@���_0��w�`)K��{�� �=R��#`�7s�Ud ���i� ����c|=y,�b����õ$2U�2�u��'t�&_��/��Gw��V׀G6��Z,ޓ�<M6!]�\P/�n�4e�m�g�����u	�yʴ�<g�Qć��tF��抖�ݽ�/��	H��NL�{�1��Z�Gq�yhp�ԅ���k{�ਏ����<�~ڭ�?�q�J��h��5SȪ��y�Y���s9#�ߵ�j���s��iJZ&`+�Nm�d�B�����K��#����.��eSJ����V\ ����㜤|ŃZ�"�����!�(^)�q^{�2D��=�I�;�6��ؔY�Vb_�u�qݣ���||C�4��O��K��8L�~_���z�'�08/�X��
��*qK<������>��\x��%���f��Xl}�rK��I����-Ag���W%��{��������W�������sV�]aP�T�US�ct�8<!-�KJ��6��k�Q>2�n���{Ӛ�B>&2��m���}�Bf���ǰ����jA3����B*<���� �u� fE_K�C;x��i����ݘ�axj����8W��9n�@A�������#�;7��{*R�@�?�q���v$̍o*|Rd��_J��^���g�kL�A���U��	,�� ��8�t�wL�,��g�L�l�D��Q����A	��	t�Bj_������ď>Μ��/��AX9��c�0J��n�g&����(j��E��W������(5xɼ�o��Uu�meFt,y�r����6��m({XM��Q���R&$(�$�c�e���2�>K~�q���>�d��P�m	�$�b�"���Y3�v��mH�(�^�a[Ԟ�!���`ߖf��j�ܤe��Cw�n�SMc:6�S��֩="����{���d".�?�Ȅ��6|S� �H%G/g4 ���,$1q)����"�uՠ`۔!I�]��<�]bא*%�'�"�=�|�t�G���'(}]:�M"���/	�.���7vn�����/U�O0X@������Dj��e�7[��<�+���Q�?Rt�d��+D��<������q���{�9�����V��T�^��b�������?z�6ְb,`����3W#�����ad�p�M:=L(J�9Ŵ�{0��I$��
d�k���B��R�R�3(/�G�;�C-������R����� �e4R����wd�7^8��YjL�q���O�[-C�+�n0��yQ2:c�z���Q\��>B���s�/�g�z0yXPk�j��K�J�MDSB��To�cs~
�֩Rn7yA�`ۖ#*ϞS�+����!�g='d¾�-J��nr�R`٨օ!��th�QyK1���0��YU-�,�m٤��-��A�6N��p���q����kp�+���5�$��3�b�Y����Pk����]̭+ϒ���jM��~pn�V��.��9&M�l�M��2j�7��e�E��n �S�_��-��C�m���i.gu��M@����?�̺7�O���$����RT��
�Z�~�b�"R�hy�����Z-�go�cf�VXoJU9�z[l"�A#�9݃4ƪ�����|���z�)o簒t�*��B�� 	�I\O�
ȗ�|� !5a�5���<I����7��qI3$؎���!<��36#��$�V6�)�,�g��4�~�w0z�AѢ�#�P���bu�φ4#�����>G�0H�6UQh�ט�!6���5��kɸ)�I��������ޠ�ŒXy����q����;�j �����jנ��ܾ@�)�~�h!2����|r���	VU�It�v�#�Us�>������3�H���a�h��4G󨣋���B��>���#XΗP��Wo(�ŘqM9�A����+|w��Y�����e��u�ل8�'�t���*1#���][�;�Ӊ	Meݱ*�JH7��6��?]&��NF���;W_��hz�GU=Lw$�mC�?ʏD�"��Eб�u'����D�L�Yi�����j�I�s��K�4 oΝ~^��J�{mgj_���C��h𦠵���̸%�+�B ��3��ù�h�x���E5/D����\�� wq�%Z�J���p� ZL��;�E��t�wTJ��	[��2�K(Ɨ�Z���2YNl��7J��@g�O�W�c1y�ۺ���<U8��r�4��B�fZ����Y�d!Fi#%�d8*��\p��)NO�fh��qQ��ź�*Y��ۆ-Hʍ�Pp?�ʠ������e�O��Yb"�
g�s�kS�T���5a�B����`Y�&'�sӁ�!h��@��nh�3ӑ�`��A5Tn���=���@&0;���c2�Q��\����nٕ�S
����& S�5K�i�?�`L@���������u��i���헥�Z�~ι�1"�p�牕5R�Z��4g�ٙfe�JoM�}���8"���\�z4I6����-|�t��k�o�Ent;`/��� $#�I߭�
��|%f!�� 8��1��؋�7�c�I�U؎�i�0����\#�$����ڻ��'�=9�a5�0�d�E\�#\Ĩ@<Hu��4FI�G�A>*ʆ0���U�����yQ!������k�b��������	H�ΩV���X�y���,�P��r;Ș��
�FJ6*ףv��!�#)��^hD����dr��
�Lӓ��v���Un�>ta����Q�����DV�?ED��B��q��ɜ>pua#{��P;�^oR�����9*Mk��i �����2de-����~ܘj͗��׉*4����_�K�'Ӭ�+e`N�*pw-7ы�6^�i?`L{�J5��U�W=j�Dص�*��L���m��?��Dxo�ܔ%��N�����ׅL�Hl�p����6l���h�$\W�Q�6^wz��zj�N�b�����c�ދ�*������%" ;�~���k(?x�E�ugʍ͂=�J� ��%��ݒ��Y��Z;ݏ�͝ݒZ�u�E򞂺��1�()�lZg,.�U�li5��K�����F�f�٬>��ot|8�ր���qB�+����Ye�@Fl�$%[�6�t�o?q �FZ�v�S�_���)�[��\bg������ �� ?�!�h�}(	C�@[�8�k�^�C��l~�5Hh�v1�{hy!���:�6�[Y|.P�B$,�}	�5K������^3G��w��P�'޽g���%s?tOi"=o̠p��u\�asj�E"�4�:����c�7�ɽ*�]�H�y�v���ח�r髶�.,�b�5�:+����6��hm�v���[�!a�ӅK��2�:�Jqw4��~:HZ�^���G�}�j���ШBK����b���R}*����r�h��bAkoǗ�neBw�.e�5d*b��� <B���V�h[u�[%)w�Gy|�����&]�Q"(.O���J*�)�Е�
�7M�A>�?`cQ�F���s�#����+R,��ݕÜ�����8����+�ͽ���o}*2<��#�8Ff{\8H_]R����u6)�	{��b�s�wʹ���Nq^֏o��Ň�`dݟ�	��>��y�UC}��Y����ҟ��1�>1��pvQڹ��zY�W졵}���,~�ɋ]�zF����5��_�������
h�А����F�w7+��X�Ľw�0�uHA0u_�Q�y�9��Ő��}�m8a��(哠W<�N��2���O���|�n���Pm�ћ2dm?F@�>t`G7�9����t;_ِ_"r��B,T���u���G,ypL��w��=�6�f!M����Ti��@Z��yh�t��H�tA�!|��fO���UUr��u���� ���g�M
[�[z��9�G���Z:�b(��ő�M��faߺս��[����/-�@!�|~�u"ubp��C_���`�r�~�����{��f��0.�bPg��_�t�������'���dy��sѴ�O��k�@g�K��o�J��ϼ���a��HN��*-S ��0�wY�����]���[� Nڼ�c�p�d���HS��M�(ii�G�jep����Cc�/#�s���L�xtI|
=�+0~��=p�U)��kL��av��]��/u/=>�I	7t�>���^j{��EIʛn�/�C�y�}{��$�5�EmK�/0��2iK�s$�7�����$H���O>㶤.��׬~�����6$�6��z1�B95�˜����~K��c����1L�CH�/�&y���HNP��8��ܡ���7��5�%H�� j���y�2��pS9��8�j�nw̭	v�;�+�2 ~|�2W���@K�D������z������%g�Mw��eYѷILUKYU��E�_yL1T�6s�_��暠�G��Y<����g�+z�t�%K{3ֺ4���$˞��sn�²@@���37q� ׋����Dj����N���@�?�e����6�1��^��b{ �I8r�m��߃���e���\��h�r��E|��R��T�mKP3����:����l9�1h_9˔x����{�UI��o���Ʌ�7)e�$ N����B�^���c�Փ�O�Թ���ʜ�G$N���3�J�`1ϷÉ'�n��I&Sԛ/� m��^7�����u3����X�4ݚ����:� ��o+��b�@r�uv1�:H��G���Fz��O��YЪȟU�g�UGj8��u\���}4�O{-�T�9��N�����)�G��kF\�[?�4#��O�,�öFc�)�=�nM~��#zNqHY�,\IͶ�롛�������=8�6f�ډ�J<X��"XU��"K����1:e���\�T��,�E(���D:yʹ��V���]r��b�~$~�c���::�$����L�9g�zCĔ�"�hX����|���ٙ��;pwaٝ;"起���9��&~���)��O���aHJ��W�3�!ǲ+!;�<���X���g hJ+�k
H�.�X��;���y��)eL%�
*ZV/ȧH3E�m�HM�肼9j�¢�g�c��텨ڒ���I٫��֜���pE�Ѣ/�n	��i�S�m ��S%-���H��"©A�,���#ɖ`m�R�!��Q��_�i���lm�}V0J������b`�G�2�{��j��2�V��;R�_h�j%��H�T�2Q͌����((��4�h���=}Q�Q"|���+����B�z}����
����V�}J��B��O�N1m�W�9k�C��
�h_o��D�"���Od"t�QU8W�vn\	�5�����U<1���,Id�Ζ	ti�P=P�ջ;�\[&S�1/�vll�W ��������Gs�Bv���dB��L�u���<��Fq]t�Wf7��dJ�&��V��`=�4v�+�	N�r#5�St6��|x�\��hR���׉�@�!�r�8ׄK�{s#R�I���P��pt��.�_����P�8�aryZw��{�q���^bso=��&�\ ��T4��_�ޞ�.kև��	W�s�^�t���&;y���J8`�pW͸���!l�s�c��T=��O"����M�h��ܚ���!�hX��+q�A��Q���MU�����{�
��'�k��9Oھ�a?���젱/�$��4�$�U�'^�,&��yGʎ����oq�1��4�����������K"�R�A�~9�FA�D�Ŵ�R�!���j�IÎ��^ss03�=e_�W���2ԉ��b�4q�`��0-���f=B�`�X}j萟���z.��c%�B��#EXK���z\5�G����8��~'߰B�CA�%bT6�k�f�Z�����v��g�Ӕ\2E�J�� \i�i�*\��4AQC�.���"�=�fWߩCi�\�SVh;%G9�2 �C�,�DP"|�q�+۳����|'R�P�A\����C�o�����VjT�����#^;u�P���u�h-�ר�A:�+���t�U� ���&}��^H^�(��;cx�'-�e��<��;�u[����%c�t��;7�I�ۿ��'1��K,��#����%�i�6>fuo٣^�-���=�Ѹi6������A"���;���^�$QCdnpHK����V����Y����' �0 b����Ӽ'1ÅZ|�ƍd��_m�Yv�J�gj��:-Ѱ���'	���YJa,�W���V��_=����=
an}w��#$��\�;Yhl�I���_ʐ�dY��@�=��97G�� �>l9b;j���f�m��d#'��9���~�\"44�w-Ȁ���
�hC���6�u���G� �`�������i��W�e|�$0Ԑ�o��.P� o�"EV�t�z��7��zTYl[����p'����j����Ǯ ]Hj�	z�wg�^�N����+Χ<��ǧ����#g�̟����xX���Cb{��� �ryݺfI��E�d�.�&���W�����*�s�F�O�{�lp|h�.��~.S@_��׈H��)<�{�T� -M�(ǌ� U��������P�����tjuy]���G_��&��U�T&A�'E�S&P�:/�9n�x�=�N"G��d�뻺���<�_]�f/�^S4������p�.	B
�e�h<8��B�����E��yx�K�]��!	�HpN��q�pZĻ��Z���(��T{� ��Ǜ�O�OU�0\��[Yh���5�C���+��Ds�$?��ݚ��S������}�J�bm+�"��*���捏�������|yJ�ԯ_N_\�@�B+m�ݹ��tR�&>��y�����(ϱ@q�-2��פ߻�Iה6V�	��fՕ_)�Xqn;��?�C��f�@[�K���L y��"�q���k/ưZX����EmKMoA���g���$\��-%PE�f7L�X=J&}�����I���~z�7��%CNH�sJ�c_�Hж���f��PO���d�������c%���x-�����2���Q�Jy��p�����q��5�۵О���}�a�f��x�!<��s7��k���*-�X��H��Xhf��Kf�sx����`M����airg��6�8�i���sı�a�%/nιp<����=�R <�p5����vQ� ˫R�_��^�g���C���y ��,�fL�wOt���T�g�N�l�����V�_��A��\ŝ�t~��Pڧ�Ji��t��9�/�ԜA��b�׶�W�����k��G��y�`���o��_2�j1�(�Pɭ�i�OŠ��gm�S!,���j��6�LH(LY}M�� �� W�؂u��c�h�-A������Bh��EK�u�P�ӂu0z�(����G�3:Qܻ=I�Ry�r�����!&�`P�Ʃ�A{jo���uv��4��n �M��j6Y���bHީ���${��U�؃P�ĄC�`6�%�w<�H��Sg��G�Ϳ1bރ�Y���O�����F] ?��א���puJ"�I_��Z���_˘c]�P�":��/���.�Da7��_�P�g�j�O��&2�lK�D;߶e�#�7l+<�Մ���Ȱ�oG҉�=Dݴ鈭���i����4T���7�$��V���/a�b�[����9�8���~���Q���G��O��p������r�p� �=�A���I��E��᪌�~M}���|�o�s��R,-�3�/[�ؙ��1x��D�zGM�]� �Z`R�1����ud��^$�*F��bhW���o���e�|[�0���y�o:�n��(tQM��>SL�!���5�gcB�y��� �K�I��>\�SS
�T����\��GR����7*�
`�5:H�S����!r����"d3H�-�tSn#m�`��C�����Q�eغ/A��	�+-V������XNz���9��M�,��&A�`^́��k!�z��5��x�M��`>YP�И��Y�/�b����q(��/�ׅ|-n;$�ϋ ��L&�׳x2[P���D�v�ngd�SXN1��?!����ðvi&U�%a%@���De��+�Ε�M���f�ȩ�K��*�Z���PB2"��P�co�CX�Z��jg@��f��o[�"�܉"C����n4Wj�ӣ�]|Y��k̉o���t	M���� r{II�O
yj9|�0�!&��FO��m��f��7$*#I�峎P�(�����U#��$����z�ѻ���K�#/�0K�ѓ�#'q����u?{�4����U�'>�7*0��UB�*��J!g.��!�k:��������ϗF����,jJX������h���A;����[��+�ױ���(a)GmLh��O�c#rS#���ȉ:��v�ʦU<��>���,G	�٣]�|
��$ 䒚��Ìs&.>�k#�H�PI�3o�e�BG=9x����BVݪ��lh�e;����ј�-���*BM]���|��-���Ezen|�*>g�7_uI6���?nт�\��IV�W�|?R4����LHm4~e?ۻ@DF�P�jC)�"���O�ڝ�`Lr��񾹪��Ƚz�@��4���_k�^E4��L�*jP!��qw��n��Y�)�����>�� ��4��T��ye'x�qE��`���͐Q��� Hi�%K������Z�w?;+�6ͫD;�(7���B��i���J(�j�Z�@e���lww��:h�g�E�@d�tcݬ/���6�8#�ʁ�u�BX�մym�Y�y�Fz��%)z���o��(�T�r����S<ge�,#�[�b\0��U�	��p? ���?~]�h�3�	� [ˉ\�9 ��Mplm��5V��v���ho����l�Dr�YJ�L�О����P5Y���.p>%<e�6A���E��y.',���${szU���=�}?~�ZC��a聠��4�Bu���z��AT��Ԯk�6�GH�vtw���鹖�.��&��P�:y8��m��6�v(�u[:�&����x�i�ș|q�/Ì�IH(�u���ԕߪ������f��6�<�^�b�F폫-�ꑗ��nn����AB�:�h��
�����}2slB�6�O�- N��W~<��+)�
��(o��9�Y;��cd
�9hW��\�n�xs����1������d��j	\��8ս�=����1�5�vTP�?�ɂ�}oqT5u?�/��*�����c�#T4�������J��.�]\�N���L!&̧�j�=������	﵏r�\S\8����*��wz�P����<�����@���r����lx�c�I#:�̹�l�Վ���M�GS��P�
�I�\Z_��cj�q��^J��=�S�&��\����p��ކ�k�X[��D<sj	�t��&#~���
8H�$W�t1��16!��s�v��<���7{����pM��]�� ���ǥ�%��	�q����|-��s�M=\��@������w'qNK�xy�ڦ�?�q�����w4ٕCU⭾'F�,g�y/o��)kW����~4kb���l��ͳ��[��:���n;�f ?F)�ӭ�RR�'�ӟ��1����Ts[B��%�E�?r�rۉ�������`��d-����N��g�z�@��x����zց�Km2B=V#-:&���zD10�/����Z���#�`�B��fTTN��N��hֹ�^ ��O�ȔDJ��2�� ��Mi�X�*D�-��OA9�u.���ɢ��%"W��i˳�;��;�����C��KD8
��Y�Wۛ0Isj5':�XP�Z@��TC�bȩ&�>��Tws��^#y�P�%u����A"Pݪ�z]�=,+����F1��.C�#&x�Gl�M� �.�#��[V�h<F%K&��f���I�`��I'�����_���{���хuWɵ^�E����Ѡ05��ӣ��"��C��𓬮l^�y�CL
�p0z"����qO�Y��«cA0"f�i���w�B?�u�)�G^��A��J�2�hb��Չ��̅���JIAW�7(V��_%��͡I�wn��$�}�#��l�g���_�+�d�ձ�\�%�R9z��6�l!��RL����p�Uo�L��'��9�6�~�p����%J��d��
�P��loG�]���~�� �Y��������և7e��$�9�W�C.8ϼ W-�E>5��b�D�z<��[�(��U��.
��3��Rǖ�xHR��z�t��Fhތ~�q+�[Զ�;�sl��r\̇��GX���:bc�r���y��f1qE�4
.��&�p���f���s˟��m{�G|��.t����@�%o_ɹɈ0�)$��{A �l��Ќ�L]U�ݖj����!q����\yE���/d,�G�U ���'-��&8?6/xL԰`8f⏻XG��h��@��1�<�R]�̬/��q4~q�������	*���M;�< �*�^�������3a����	�_6N����wZ�I|�r��䱰X�>�{�[ڨ�ǃ��7.�   N   Ĵ���	��Z��wI�+ʜ�cd�<��k٥���qe�H�4͔6Z"<ɑ�i�6�3{�\2V��<d���fJ>@,o�$�M3P�i����d��f���{�9ݖ<Z"��5�����@�MC7����O�5��4_@�,F�@�x�cB�c���'��l�������.O8kq��8 �"/O�!�k޿q��	QǊ o"��>�P�޴4.��O,�Ӧb���u%MHy�A�{<:1aO�)1[�A�΀�H��(]��'�n�	B+�C�'K���=�XUs���X%�h u�c��'���ቨr_�'|P
�g�=-T�8�F�.��Dڝ'�!Dx�_�'k<|ku�ʣ,6��À��+;��@a�5f(�"<���>�1���"�D g.m� i�d�i��Ѡ�O�8�{2`S�`z
��1EDx��9�M��0�2^|"<�G&��\ᔰU䄎׸-�iγ
m�I�>a�L=�2�`�F;� ����*}�H��ӭ-XU�'U�]Dx2�JA�`��9�e�QJg�%�=�.!�?<"<��O���`��3+�����_�* �)��@�O �L<Y1N��=LdY����`�e�ÉMd?�%+=�B���<�1��UVU���'HD�8#��ʟt�O������*1�n�q���y��5jb�
ED^'�U
D*��d?h@$,Pi����$��xr�x�ݠp_�Xh 6'V�h˃�&����$���u� ��G"�E�P�-�W����u厭-��P��̜��y� @� d  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   
    �     �(  g1  �7  �=  CD  �J  �P  	W  _]  �c  �i  (p  lv  �|  ��   `� u�	����Zv)C�'ll\�0�Ez+�'N�Dl�^T�9O��Q�'��(�bE�f��
լ�( h�n��%�~�#�)�t�6��7�5b�ͱ�~�e�E��?i�Ǉ�?�K����D�Ιx5 Zce� ۲l�.q���`֨S����� .:��թ���uB� ��t�'�:�+U��ڰЩ�̀��հ�.ءD�0�Ă�O��v��$|�#�ѦX�D�<��ܟ���ӟ�J$��E����Ɵ6bx�4��՟��I�M�1��0����O�柆�d�OX1af+�;�,�+!*�06N�O�Ġ<y��?���|���'@�͙p�rP�U��*l�lJ��ԋAE!�_55"��f J�82�	��oε^��	�<I>��'+��^a�$�Id����DC�	=B�14B1�?Q��?���?A���?i���'I�,��"�|���v-��;����[(��ep��=oړ�M���K!��"vӰoZ�M��B�YHE��X`Iy�	ε2��!q�II>��V�ǜ ��˕�~��g$��j~)b �XVؠ�[ܦŋڴH���O{�)م#�҉(�!V�<��i3V�)�V�A$��kL	cUV4�b��q�84K2�T,<�8V���)`7�Ħ-Rݴ\�Du��<F��8❢B�>j!B7if8ċ��ގ_&��B~�*�l����zo�9��+��P3:���
2ĝ�~<4ys�����-#˞)qg)���yb4`u�rnژ�M��i͇&�5:��_�|7Hy�'�;�@}��k[�!
(�A�hG�a/�!0�i\PC3��1L*Ѐ�����'��O8��C��C5��Q���]���I�A�O������(d���M�Ο�HJѡd�
��O�^Кy�4�'�I��D����p���$u�ĸ���Q&�+�1�jU�UE�.z,%S`�V�3f��	=��Ƞ`�#�P5�2�B����%"��.��ZH���	��O,O|q��'����8G�T�O�� :#

/3J�����OL���O�㟢|�'|>������'5���D�Q�����T)jL���H�"�q	�&~�j���h��eV�)G�D3�nM�Vo(hᐅ���/��8�f"O��0KP�Z�B]0��3L]JP�@"O~��e�O*� IR��/T�y�w"O
9s�Z�8����r�Дb9�""OHa([z٢%�T�;��2@"O4��ǁ\�C�X	�\�k�'����`:�S�O����O�3�����y[T�1	�!�גNhXBSF+�ř"�
 p�!�d��H�	Dޞ��L�Rh�p�!��Q�l�P�R��-I�z(���J�b�!�$��j�P���.V?J5�򀅆�!�	y�L a�!A�65���1$��I8{���D6W�<���Gv�~X�D� �!�dF�J}P�A`��"E����@M9�!��=YQ��	2���?)ڱ`w�Մ�!�$*�Vt��F*F�~���郇�!�D�'X�J��'J��r�(��}l�y҃�u�7�1?�Ǆ�ߞ0�� i>I�`m�ϟ�'2�'_b���86I��
x�$ܚ#�O� ��+�Xk�5�p�qlv4�b�'1�}���J�T4ڰ��D-��)�\��e��oJpzgN�	�0<��j�ԟZڴX��'V�-#E��C�D�p�
?^�&@XP�P��s�S�O8|1��U�9���PQBܭh(
���}��D\�N��-{%I�q�195/��?�H>�5O��:��|Γ�y�,ǋH�@��]��AD���y���Q�Ӌ\~�0���.�yBΛ9L�ڥ��kͿuJ8ȉ��-�y��������Ǐo����D�3�yB@[/�%�,�`:Eaԩ���yB� %2A���H�^d�y���u)�f�'�B�'�<� �O��3�'�b�'���##��� �>H�>��NU�/��[q�?���#���#���h!]>���i��'�~���/�L� ����Y�r���k�.܆��'-ޥ��Ejg���m��)������h�L�󮏲8e<�P�$�6�`�:��?s�6�ey2�ՙ�?�����?	�#�%h�XZ� �c�h�,�sϓ8^�O$�#]�6 y�L�T&hy��]�${�4f�V�|�O���Q��
�D�i<������}?.9��Q�O[��]�`��ˉt>���,	2���h�#�1=��C�	)�����ܸR�����L����#����n}P�sg�@�}Y�Իr����z����e��U����P?)
�b6D�L�`�! �LH83�����};Ѐ/�DNĦy'�̉������O�h�ߞ-���k7�N�sZ�]5��O��ā�
s��d�O��
��H�3�¹c~�cv��M� �L�R�ˎ����F�50��+��'��!�H�\�0��U�5T6�)f ��@����xy!F�aaxr� ��?A���dЛV�I�AD� a*���qb�s��'?"�'���!�ٕ�pЊ���<9��EK���8�l���ӆp��1�Co��?A)OFl�B
N��Q�IҟԗO2�-��'| <���<aHe-�j[j!�F�'��۞m��h�Wc�M0ʄpwW̦�'��i�&D�Pa��BB�fe��:儍&8�I1���v�G���ǯ���H��l�#(	7` ��gkx0�����ra��O���/ڧ�?9��@�|"��b�
�� �+�y�%U&r�xk�i�76�A`p� ���O6�E�Tj��`� (x��9Jl\�a@N�����'���3�����	��x�'�<%(TI�:R`��E�0j���Z��@F��:<��d��L#�p����Ds��� 3ցY:H
 �fy ���l����s�'M��I��!��Ϙ'�|�:G ��0_��a��M�d�r$R����������'�ў�����~^���f</#�q��AM�<��\8Oͤ�@g�uId�i��My��?��|:����D�zijؙ+4�T�%���V��Ĉ�ƦM�Iӟ���Ny����?|��ٹ�I�$HoL�@��C�ę������� 	4B����ڝ1�6@����w(4�J)Lx�*㏎�j���G;(�n��dN�j��)[w��gH�AR�b���,0��'E��^�'ћV�M>Q�,�2�b^�P�|�"Ox8B6O��`�)R�̃-�DT1��|�CsӶ���<I��Ø��O���ӍU'#�@��蝗a�l�������O����O�4���!g�Ҝ{6aT�ki���FJ��m�=]�4�efK�x�L��d�>R0Q��fզ:�@���O�L��B%��Pn1;�&�c�'.9 ���?��OT�,Ш�U"�P.I���ԓ|��'����	���� G�C��1�	�e����5��0�jS"	�N0X��6�?!(O0��qG�On��&ʧ�?��[�:*�P1�T|�>h�@���?��3��(��&l���!W�	]��)؃T�<[4�"Cd��3"F���ər~TtK�ɕ@�r�C�I�Ok�A(����v$z�L��Lp��O��H��'����<�7Ddת�'��� �P(#��b�<ᧉ��.l��(ʀJ�Pի�C�S�'9D�}�7��/>f��:1��9��b��M���?I�f&`�Iao��?���?����y�:���˳.��n��](`�G�r��V'�@7�٧2j�@r��D�1V����)?�(�0 ��|���+w��u�uo�10e�pr��9�3�	�^�ꀸDcXm�X�Q�ev��$"?�f�Zڟ��	؟x�?��/��s����c�'����r/�2�y�N�xw$�E���FU�1�V���j�����'e�ɺH��y8w	��G��`�!�1
q)���M���?1����8��K���T��J�M���zSIU�6@��Q�G�2��`J�)��sϓx ���b��P�e3w'=Y��LB5䚄mK� #b�-�M�T�'ؒ�	��^�J�ԓS(ȢC�@� �!� �?��i^O��O��� ֍;�����K38*,Q�W�<�g�v3�賆Aٓ{vđ:&l@R�	,�M+���'[p���O7$ t��[=L����PͲ	�'�T���3h�� �c��zM���'*���7�X����a����'�T	���hD P��䋸G���	�'�`�+ �"s��MI�[�o�$(��'���Ț���H�Nõj�\#��dǾC^Q?sg��>⒔za��=+t�:�m8D�p@�̟d�d�7��Wl�3ä D��h���F�J)���Y�,t��n3D�H����;���w.��N�2� 2D��[Ԇ���a�ǥ@�!j����
;D�����;N�G$�*p�����O��F�)�'��a��쐆`\䚧Nj�=[�n2D���@>�ma�L^>�(P2��.D��@�]�A�@%�c\�����,D��#wh��Q�^h�B�1T/T�� �>D�$�mR�p�����&WJa�o!D��*���-<�|�w'�o��<m� B8�X�+�!CbQ��@-b��Z�d:D�� �����P�����_�+�<!rp"O�D��?�n`�'N.W��K�"O<}·�ܫ{I�- �%�:j�thf"OĔRc�E!ĴXd��>�|�S%�'S�]��'���!`�](<��JՠJ�X�
�'s4�6��9�t,b�5D��$	�'�IYv!	o��C4 9�,�y�'o~5:��G|��!�d��-��`�'J�jAӗE�����G�2z����'v&�ң/Z>6�H"[5&������dM"6@Q?�bi� 8�k�̶/_\�X�0D�$�OڝW���vF�':�41��!D�4��!�P�ݡץj��1�f>D��` ˘�� AA#�,<��C<D�`٥�ՙ<��)������xh�"8D�t�ү�F<f<�` ����'��O�D�3�)�BYiQTJ��k���$0��Y�'��l�U�>��ђ�m\-q�Y`�'�������]͖���͘V��D��'���@�ȧk=b���I�H�L ��'�� �WEX7�
��F�;Of|�	�'#�e�w�XL��e�$��q)O���'�'�vj�-�)D`qs6�Ƣ0~ؐ��'��l��GT�j�n���*ߠ{l�\b�'�,��smV�ekFB
��s��P
�'IhGoG�h�����,�>`ntc�'�6p�v�\(|��NWT���(�&��QԂ|Ӈ/ �^IT��DȄ�"f�مȓ��5x�˛0ޮ��0͞1VF����{� `�	�YzA��F�*2����t�*��ܱ|G�t�vm�PO�!��#y��ǧ��:� ��O�$�"��ȓI�6���F�jVn�9PԘO;P�G{�����!x1H�,�x�P���3`,�,��"O\�qw)��}[��C�╊`"O�)��[��#�(B�^��`�"O�:�@eX�i"�EF0�0D�"O�����r�����6G_j9�"Of�#"��2�A���iW�D���'�̵Ҍ����h�%S�H��Pۢ�[?�0���Բ6a׷6���e�����ȓfΒq"1��q̉�%
�SN����IzR!svN� +k���B�8�L��0;   �U.I� [1Wz�ȓ-�$p hX)��(+C�(JO�`�'Z�����ɋ%���04;�+�W�M��$GxU
�խ,WfHI���(.%�ȓ�(ԩ#	D�C2<epC�K����_֔�k0KV*V:�$�5����ȓp�P�bY�n�p��g�ɕj�����	*�	Ss�(�!��W&ށ���t_�C�I�E�̭�f� ���X#��D�ZC�*8�D[a��Ki�hУY
�4C�	�
����D��×K>B䉐y�b�0

�@Un|���#2^C�I�G�Jy�FW
0A�����O��D�=�Z,�~�#��[�j�;��`JPڤ�S]�<���&�zXPo�Pa�3P�Y�<qS�ɣ&���R&G�<6$���jV�<�f��l�V�3��M:\^�Q���\O�<a���H��1HE����6��N�<a����!xW	�2���Z�j\ǟ$���"�S�O6h�!lN��d�,Ϸ{�6��E"O5J2�H n�b��*�y(\�"O� X�[7��(D�cjЀ.a�}��"Ot���e���x ���.JU
٠"Of�$&�^���"�ǖ)_>v�؇"OP�h�~��i�[8�̓qW��#��+�Ov�22��+�V0k���14�u�"O���Ƃ
mF�`@�,���q"O�X�1EF�M�qc�%�m)	�e"O"<���R���:���}7�Q �"OB��E��5q�nP�HU("P t�'�ܭ��'�!����b��Z�Hc��6D�(�m�?8�`��%O>!o��Abg9D��aOH-�c�@��$��4D����D�%���H�͍7?���AӠ>D��Q�4���"+0�\��>D����Ϙ�-y��� ��Ytq��!ړ{N D����ig���7�T��|�!F�.�y���+��P�T�����D3�ym��5.4�2��&��G�U��y2ID�H(c3*N��G���y��6,r�ؐ���Hޠ����7�y�$V�.�;7�BFԨ���H��?���A����X� $h�Yȍ��A��	�Bi�&�3D�h�6#6.,��Jk�\���3D��z`(!% �B���:o� 8QN7D��`R�Tq܎$h4�Q�*���.:D�K�BȤEd҅bb�ɮW�*�(.�!��[3uѕ��)�V�#*Թ@S創TX����S0u�μ��M�	�&Q����"@!��IB�98PLR�M�r��d�"BC!�$͸p�s@�S6ԞpB��u%!�$�'��<�"�R1T�̅�q
�'/!�D�A����EڝcԦy�GcSc"�}�����~�ޮ]��I�H��dRQ��7�y2���=0��Q�r��4����y"i��'��T�à��X�4�q��y�Ή/w����O��L��eA�n�<�y".�n쐨K�׎L}℩�d��yB$XNȒ�Z�I�I+�Ւ�j��hO8����SLi�v���a.u��k�T��C�I
&*|�7���f���#4�LC�Ip~���7Fү�$���[�KDC�	�	�ڌ㰏	*]�mA+��#K�C��5~> �F�E�  ׄ�2!9$B�I�*�ec��Ǜ[Z�r���a!�����y�"~R�I �V0��P���8��ԃ0l�(�y�CCN���#�Ї1�u�w����y"S�z��`3��.-%���w@E9�y��Q(X� ��d��|�q���y�e�y���%'8�"�؆�ڛ�y��\`�$(����2�N���%��dU�qk�|����_�
�Q�JR7tNa�e`���y�bZ�&z���11�LQB	:�y"��Nk��y&�Ex����˵�y���"���!�kݔ�#��N��yb^�)gFh�qgޭg�h� &Q���>y�ɎM?�&gʅ'��!�Fϫ�������d�<A���8�H�k��\�(a}3b��]�<1G��)�<X;�g�p�m�WRV�<�R�/ؖɀC�#tY$C�FS�<�mɏu��E�aN��2�\)(C��s�<�r���W�$����r8�T1Dj�s�'1V�ی�)P�{k��>��Г�e� ���'�~Mh���o�����C׶8J�!�'�4tQ��ud�9���J2�h�*��� X��fo<Q�`�AE-�@�*�"O��K��8>��	+lPk6TӒ"O��v���A6�E���5`a"����'�������SŨ6���Q�s�T�����"k����P�k�р4`/,���Z���B	ۧQt����E�z�<t��F��1����EPl�3�?@+|H���dy��
��Zq\��c�B:b$X�ȓ�����خ{l���I��tb0�'DL��j�&y����fLk��-3�Ņ�H�V�0"�T�l�HcPIP4=Nr!�ȓ��aA.���x���(n�D�ȓ ޲g��'X�<�z"儤,�lP�����fE	<-�tH@u�8S9����ɇ,�r��+N���Kr�ģZi���cZ'Z^4C��+|BD ��I�G�6�h� �'f�B�ɚB�@)��g�EC�S�A�S�B�ɤf�A[��ߞ0�!�I	>�B�I�E�����90��(I�J�)g*:B�	�z ⳅX]�j�I��F?p��=�7E�Ots��^{|�D�@�{7�X��'�����&����]�rE��'�2���1[0ε!6�ڏ�>��	�'�=�dLN7V  A���!�����'2����vD�F�F�g���'�<b�B��q�dQu)��_�����)֚�Ex���8A�Bݺy41�P�4#�dB��7\V�H"�Ċ�
e-@tLT/K�BB�I�Cc�-+�L\�W8C�̒�W% C�Izt :��Q�B\py"�O�o��B�I8#���a��0:�(�`f�_(LC㉔:�TbaGH�H@�r�K�K~0D�ɡ��$ץ��$֠ n�?	J�ׅ9���Ʃ��rn��b�Pgy2�'��'��]`懃:dLJ�*��/�~�4�8����>G<����q~x�A�	3h �\��j��b��\1��V���2�l����Y0��bRC���O�<Pf�'B�]�k�b\Á�2vO�n�c���J��dk�
O���{�D�#)��]
!�Ov��'8��:A�^�>Y%�ā�Y?\�J/O�����Od�$�<�+�D��O��{���Uh�@F#:؈��	�OlABM�m ���)�f��)�,��� $$�5���0ĄY�*l�j-*D!`��pl�E��O-�蟌 jfH:e�,�T^�g�Z��c2O˄��?������4��Dz&�� 0*b�B6!�Ny�tL"D��:��>k��T�%@Ι"m2Q�p� �}E�?ݩ�Ǜm��Ⱥ�@��*���O��ܕ'ςH���vӬ���O��Ļ<�'/��Q��Lӏ`ڐR%��
I�H�A�Ծ�?�3��2c���?U������6(���&�+�����JY `��Od1!���J�v@!��?#<����1ޘ�����d�BT�I[~R�ѣ�?A��?���5��$C� ]�9i�KG�"�4�"Oh�iq꛸Jʖ�� @˶ra��  �'X@"=ͧ�?�*O"� ���O1�$�tn��'�p��H���09c�OZ�D�O��BѺ���?��O�P��b^��0U��F>b1��.�T�K�W�}�����'ؒ2 �ZJ�r���i��&� �I�h��(N�r�/C	8����'/H�z�!�F4���MZ[�=JuDS	K*1��?���S(��i�B�/��p����>����ȓJj�L��N�	{�(R��; Dx	�'��7m�Or˓�E�������O��?I˦9��'[6���9dk�4W�T�dN-y���O��D׫~�4h���/ �jaX����S�:&�W �h���\�H��t�IR`����4,�T�M�p�tLA�IK�8��i�kf��#E+�O�%�1�'��Y�l��%$̑ �d|[�J�2��IP�����ǒ��9� %�Z�P�c5�O�l�'SR��g��t�����H��.O��*ZЦA��🄗Ou��@�'��	�6m��y�慴 tdK�
݃b.��-��
Q�K�P��1S��O�F̧ � kAc�f�f�{�)�(#ۀl͓>[oҡt��;q+E��h��A)p����-D�[�3OȐ�'�Ҕ�����S�? t4�R����xg˕F�.�0�"O�U$i���%�֖~/���	!�ȟ&Z�h)��Q2�m�N����O�˓R�V�
��?Y���?�-O��_�e��J�eB�y��cS��)0�8���O�X8�iC+&
FB1�?#<A�FB����dQ�Dwd�v��d����t"��2�AB�\����O���A�
sP �$� �ԙ�� �O���5ړ�y� 	R
�s"���l0`�O��Pyb�#���Y!퟈L�V�z"��۟�i��4���D�<I�NG]N�J�d�(?X�u�.ɪ��P4sQ~e�I֟�����$�	�|*cJ�>�	C ʼ ofl�EÅ'I�Z�bt���$0X3@K��<��4Jp�S�W�<o� �b�M�0�����&O���0��)��<р��ӟa��Z�ξ4���	�|t �a��ԟ D{��U�I��� ?��Ek���!�zB��!si��@4%�8�iwB�"X=��CÛ��'"�ɛMKX����$l>=@�'M�*+�����!��$
�
�O���B�O���OP|9� T�f�t�	�9!���i>�8�`Φv�؀���!4�H��i&�1H�h�7�� C_��*G�ˁ��i\�V����ӎ�>�Nlr�e�X2����j�O��D5��A� ۶�@�O�3v�=F
��0?���L/{�41���Ξ=O¨a�sx�T�/O��+�IS=H�h��BFv�����O
�$�Ov�?�'1
�CD�R�|,��D	����1Ó�hO2%bV�6L!:`Ν�t��B�$n�.O� ����+�:��4�϶:WR5���V���DJ?���v�T>�ɹd)�Y)g�S�5�)��� Qaf�t~�	 }���!���ħ/�bI˶� H*�!���	!�4��B�)}L���F��'ݚ�y&L߹Knq#�� �DM�S���	���	0~���'�X�9�aA'��G�0!� �!Xd�	�w��'D��2��	�2,D�P���2S���@B���t�����5B�-�=�N��Oz$nZ@��$@��;@l��#f�NӺ�%8���O�`G�D��^F!����"0P� ��_�)�I�S�pӧ�9O��@A���Hb�̫FHh�n�=�Pi%���"δ�'M���OR���	� a��E�M�%N�8T�[&e��J�^?A��Da~ʟ�D4L��$F*��	�#�)%�8Cf��(@���I[؟$��.\QP<��/��C��C�.=D��J��@(p̩��	X$#���h{�b��.�$�v��O������*V!;�
11*�wn1�F��>�O>y��T? ��P6G}�ȁP���Rp0��v�4D�����)_i65�O�v}"��T�/D�:H_�zG M�s�C;���Fm.D��(���a=��I�`��r�7D���O�m�T<s@,Ҏ2������5D��z�;@�+��QQ}|!��b2D���d,�%	S%TG0�p�.D���㟛5����2B��)<�IĦ1D������/j�A)�D�:,J��e�"D���5��B����C��8Q���?D�@X��ET����"y����H<D��IFl��#S��@'n�2l��ꆠ$T����̜(>��A��/-�����$x>|�"�F�1v�་� 
 H��� �B-\t�L���3?,<D�<3�i� �C��dl��B�4N����>��$*���)%W��B��"���@��N�,��̒T�[0&� ����įw�@�Pc�,_y�U�Ҍ�t�f����*;�c��(����艵B՘]!�'�f�����J�I<<Px�	�C�*�4���?A3������1K�,oi�i�G��~�bC�'�ʥ{�眪=�,��'��J�@ћ5Ҥ\"&�*=B)F���[�Qք�UJR���%�ē?����	���F���i�y1e���&`I����?q�6�Z�a=$�X(�lX�&��h+�E���C�8OdiDybe1V��!P�!\
*b蜚4`���M��Oz��ā� �x��h��.DV�Ѷhρz�!�ď�hEh���J�[&�šC�T�!���,�����5��i��NX�w!�d4i�䲱*R�Ε���udĄ�}�<���_2&��DjSV�U�8��L��Ec�(Uƪ剐�sH�����d�+�lQP
X��r���S�? 
Yb�
�����M	�k�"X;P"O��F�TP�����υ �Biy"O��S��6 �0K�kПo�9�t"O��C�J7Ux��a@+�+8��"O�] �	Y�IQ�m�%e�UW$ɓ"O����"P�i,x ��Ë(bـ��"O�t�%�h�TX3�g�$^���"O 5p�k��d�l�2�K�t\�0�"O�x��V*K�D��ӯ8C�iC�"O��I5k��&,�<%
��>8��"Od�ʁ�1��A�_�6�P#�"O�JD���K\�����$K6��"O��t��f�(|2׃F;q�&p��"OI��'��:�C�:��!"Op�R��S�E[,�+��� �E�$"O�����`�<��v��	7"O��PY�����Џρ ~�iS"O&)p�
�[tt� ��ZG���g"ODkQ�A#\!bC�J*����4"O�J��C+(��!&`�h�"OF�#%�*��(� ԀW>��f"O6�kP�C�%�5`��wAX}�"O�0C��S�t��� z%Ȼ�"O�p��ƞ;f���2�A�M��2'"O~ {3�Ƶ#LT�0lAy+p� "O"�!�D�2�Tz�銃l�-�d"O����MJ�%�^h��Y:6����"O6q��� �|�4I��QP"O~	�3N��&����^u�Y�"O�y(sƀ=P<�7�A�Ǡ (�"O����%���Q���&ǎ��"Orp�4@7��BWZ�Z5xB"Oڈ�QA�5&Ĉ@w��aiU"O(�4�Q�3�D��,�6E��qhC"Ol��&e��.����G�Ÿ@lru#�"Od�QF���{�Cb(�KAЄCE"O��2�D24�p0>B�A �"O��s��N�w�%�F�B,B'���"O"�����L�a�`�R#���"Ontڒ-©h��p )%����6"OР��Z?J�����	�!I���"O����N������	&&B��0�"O|�Ǧ,?$�A�a��[��Ӕ"O����j�
�,�;�+��lM`�"O4����]e*�(�Lݮr-`t� "O��� 
�x%Ҕ�+�tIK�"O�m�D��"U���h4�;�J���"O<p�$E�D��  "iL5~��(�"O`��Q+; �\�ϟD,�K�"O`q�ca(m>��g�6� 2�"Ovp�+B$+�4P���Ԛ�LP�U"Ox�����M�Z��EG�r���F"O�HC�K�P���*� oub<��"O"��-��	D�4Q2I.y��a�U"OD��V	ղ{�.�� �!ZD�x1"O��(��тlHj �E8@�雳"O�R��*\*$I	!�̅DZ\�9D"O�thu͐)���A����p�\�'"O��I����(�¤sd���H���"O"�H�L[0>��4�	.}����u"O4L:[�����܄Z�j�s�"Or8���j���I�.@��(Ht"O�<Rmڽ+��D��6'c4p��"O��ۦ݉W�}�ԧ0]xM�"O� ܊`nʽ8� ����Xp"O�� Kӊ�@eJ���.w�T�A"O%�����$�c!��&�͐a"O2)ik�$��ԳB�g�*��"O��R��56 t�k�aЬg��\�"O���'�4�d��p΁)m6m��"O�iG���i�m���	s�"O��j��Ŗ��}a�Έ�#U<�q""O�l�A��H�D{�+�\D�Йf"O쁰a���qӾ`H�*ܹ`?j��"O��i�E�)x.�b��1s(����"O��C؂q�I��J�2H�E�"O����fԩ7���z!/޶Z<��"O��`DT.º�;w��dcp���"O���$�K�!~T	Ū��zL8�3�"O��Q�l\9A}�-[ChR'U՚Y[�"Of9��e��U�J��Bb�ad�Ih�"O��cO�� r�9
CgZ�z�>�B""On��$�B�	Ͼ�i��4[�����"O.��	�(Oq>�cD�פ<�B���"Or��a�E���!I2�ʥ�l��"O�1��*^�a����D����F"OdM@���'z�fPz�-e����"O��K�䋙�hm���Q%/����s"O��@4iC'�����Í����"OR�hR�-�^���?|N Y14"O���4F��0&Z!i� HF�t"O�q�v���rJ��q���-�QX�"OZ *�I��麁+q@\�\���V"O:d颅þH] 8C��d��h"O�}��7P�Y���6$�:�"OP@zgE�sfT<CVj��r�"O@�	�"XL(�M�E�]�n.i�"O"�Q��L�Z@*���4�a��"Ol��ˀ'F�u벇Tf�j���"O�����-%ax���cJ�ryB��"O�Es���3�N���@�,:
�a�"O���/ߤ�d���M�.a�
`��'"���T	A	����s|E��'u���M�U��֮ƙYXJ���'Ү�r��oR�P�uB͖��K�'�@���E�I��e��$��'b(���-�ɳ�Z�/�A��'�qp	�3Y����v�!����'���Ʌ�M��� �&����
�'kTI ���`���A�>t�tTI�'8V��Gi^���٘ե�5m:��'uZHXSF�	"M��f�Ҏ_?�h��'㎨;�
�$<�AJ���_�d4!�'?1���'���:%J�9Q�ȁ	�'�BT�h��nnX�Y�Mm���')ji�0jsܝ�+:H5ځ �'�֝�D�y����ȥv�4��'�UK���l��Q	�X8rB��
�'zT�"�O`B���i�.n5X%�
�'�ڽ�QK�8��B� U=`1�)�'���p�Ûx�4P��a�$TA��'��P7��]�Ƶِ*
+[�P��
���&�і��@�+�.�`�9D�`��T�2������T[�"Ms�%D��' �@�H2��<*�1sD�0D���E � 7��C��ް��t"D���Bɨ"9�aI�(�$R|�#�O D���욽$�24�DMZ���?D�� x �M��<'Ba�TA�;(��B"O�p�+�$� ��*��Q�"O�z�'WQ;~���R�l��ؕ"O��
`�@	���a��ұG��y��"Oj�XC � m�Z)��E�D�1�2"O [�A8B�r@DcS"i��%S"O�1ffF	Hr��E��H��XG"O��ס,(�8���+�ܝc"O�;C�G�:�y�Ɨ:0A�]��"Oh	�O�+h��,�ue]2/H�*B"OL���"Q.s$�Q#�#E f+L�"O�b��i���p��Y/4`a "ORQ�_�$�
�'�!+��@�`"O�}8��B�_2�%�g��[���3�"O@cv�-|�x�`/�ZaT��C"O܄������RI�ŀ�aX��J�"O�=��F�"7Y��`7oC;es����"O�m� ���(<Tx $�g(�k�"O��W�C�T�D�M��F-�4C�"Ov���!`m��B��%
��U�"O�7�,A�v�q4����"On�����6Cryנ�O�x1�3"O�e{��/M�t�i'��`i����"O(�z5�5��3�ϛ�t>��w"OZ�pܘ8�ԀW�f_�d�"O$��Y.�ph�S�~�̰�"O�d;�J�-+��I1EiKX��$�U"O�PґȂ�,Ҕ%�զ�5F|�#B"O�.4�8��!� b�D����!���'_��*��m���y�o�3w!�dȝ҄����a�f�7� v�!�d� �L�KS�(v��TY!��!�$^?7���D =/�����:'!򄗉5[A	9+�dI�nW_ !�]!��e�'J�e��-:eAG!�Dt|�QpoS�)� ��-D�O-!��%�q3e!��W��]�Q�L�!��8v�pX �ԓ~6��2�ʼR�!��F�X�ꌴ>z�I��b���!�$Nxe�10�g��f\��PAm3C�ɆyC����<��sF��
w��B�P����TMݰ��0���]	��B�I7%��`�f]:��H�X�1�pB�	��"l����Q���2kl:B�-<�j�)�KIp_�%p����#�>B�$
!��$�c�18�iX/�:B�	���[��۵f ԙp� �&HB䉮��'g�;f�n�X���'l	�C�I-z���ql<C�lxy�	�7��B�ɞPT`�!��8�n�` �j�C䉨=��G)-=�B��U"I�\�TB�ɓ+�B0�-��:�ق�lH�i B�I�Y��T���%s�Dy�13�C�ə^��`s��ݦ(��� cQ�L��C�I�K���s��:n����
�rdnB��9ft�xP��]4D���R=�6B�I9q��[�c��I� ̙��Pg^B�#����)R�Wԑ��<�B�	�R2jŕ�?���v��c��C�ɛ:���U��;[�|�Ӳ�r��C�	�ozZ0�HI�'P0:�dɎ;�C�V.�0�ˑ
~�m�GImt�C�I�7�e�-B�����#����y�ER&o��J"����牂K�J �3c .�PePTm�6 R�C�)� 0��kɒhW��I��ȒP�j�"Olm��H�q�rR(Ѳ2G Ȳ"O���j����ؔ�>A��K�<Y�C�E�.h��MY#_ˬ��h�^�<�a�#�l���i�	i,�q�Y�<�`"�z6ݠ�lQ�%'���&d�Q�<`$��z! ��'Eyvy"!HE�<�]����;x	�]Ҡ�ߎ!4B0�ȓ+tpx�@�� g���lJ�.��0�ȓ �8�C� ���j!��)X�W9ā�ȓ!0<J��L l�V�.Y����k#D�p�!%��@�ВcnN\��[fh"D�*7N*lH�dk��=9�	.D�DRvi�PCh�!�f�i����!�*D��{�O�^�"M˷L�H��<��*D���/�q�J��b��p�(D�@3��RX���� fD;��qb�(+D�8�FT%-�L�i#��!����aL)D��C�߹[tj�a�#\3X����'�*D�(�Mۓ�֬����++��[�,&D��Q�U�(������hI��!D��RHJ�T�yĢ[����%D����A�	K�A�7. �a��]p��6D������r��e�7�֝T D�L 4�D@���@�i�����m8D���拎H��d�rnG) H��)0�&D����eR �U( 4C����+$D�D�%�>'�|�� �[�8U;�g,D�0��L 1[��;@�m"R����&D��!U���m*.h[S��X�<��$D����_��\�[p&��� �."D�!:?(}k5�=E�v�
�:D��;�/:%,�pF���a�-9D�$1��H�^sFD�w�OX��"a;D�#g�B�M�=�P-Օt^l�	d�3D��Θ��2|ya�d��U�>D���Pb�>� ���U3��m���7D�0�3'؁v+����*�W�J�
�+D��ۢƃ8KB\���^	_R����!(D��fl�]�2��%Ȱ<E�U�"�:D����/����%"�$����&D����i˕5�Hy�%��e�@ٳ�o$D���VmC��ɨ�A��%�(�F$D��9��7vw ��a+/*/�e�/6D��`F�S�颂�݌f����U�2D�,J�S�O��(;��,C���S�+D�\+�X�&D�ik��ѱ��5`p%D� �d͕)ZL�[2н��"D��"�l�.��Y��*qԠ��u-"D�H�6��>�P��,mxA"D����I4\ڂx��Q�V���!D�X2��W�A�X�k )�jt(AA�!T������¨���Z�;,���"O")�b��hj9▪D�=T"O <�Qp���I���`���AQ"O��J�l!.����0��]�~1��"O��I6�G(߮�Ҵ�՚w��1)u"O�0K�M�!e�nLQ"h�,KP�"OK�6:�"11���p�r���!�yBM��oYZ�K��(d<@�"� �y"!�����c㙹a���J�G"�y��ёNF ��ҦL�t;���1�y	��'���hë30�0A�LO��yR�Q2��b�/�5z���Ŝ�y
� ���q퐑W:6���&��ܠ0&"Od�0�.ɚ�(y�c#$ֲ횠"Ot�: ^VN���i��;�"O����J
�2��)�ʌ�g�~a`�"OQ
C�DBdTx'�آJ�$y�Q"O"L0�+�)O\[�*��"�B��"O�%�T�ΙE�n�rv/^(%<09��"OD9{ �֩C�"Ȓe"���"O�x�`C�g~��)�VB���"O�8�ƙ;c<�
D���E��Uq"OF�� ��x@���W�H�J�"OX�h�J7PTn�ҧ��	[�8�%"O�,���ק%�
 �1 �Xs7"O��C�A�%y;�8벇�1e��d�0"O��7E�6�h5hζm�
Q�"O%���̞[<��D D�$9��BY4�ɂj@.O���8D��l��D�A�䏣 Z�@Y6*O6pH4�R/$���Xw��O�\jd"O~�
C�0G洠��e�)Qx�c�"O$�S����$5�A���@��� "O�[f�kx��D"�@쨋0"O��[�LƩ$�:D�Q��|t (0"O�m�%�F	�*�P4�1Yڭiq"O�
WjX�T�jq��Ȥi��:�"O����G� q�˦(��Iy�� �"Oj��s�ţ|�x��v˿g�9� "O�E�A�K ee�xh�AH���5"OBQ�P�H	A�����+�N�PT"O:m�F�Ͷqob��v	�ou>P��"O�HH2��6�N		'i�l�T��"O^��%HGʙ(v�к_Z�!�"O0-�C�E#ihః.]e�� Xq"OL�YÏ�\z�,a�FR�?=T�b"O��pG�е��[c/$mn�f"O�TC7`°[84�^	
:K�"O~�83�1Ʋ�2��Ӵ�L��"O�+6'�9��Sď�>wL����"O�����M�^�B��W; d�z�"O������ r�Z���#'�D` "O�]{cb�g�v1K�#�	YmD�Pp"O��i��UO�5J�`�b<4�i!"O�|�1���bI��d��\*~irp"O(��G�Z4���������"O�`x�O�=�
x�'K�s�i+q"O>��LWXTc���K
��d"O�z'�O�j�~�9��Ѹ4}�1C"O�uy2��X�V�����"����"O�k���r�81s(�+Rj�A	�"O���Cͅw�4�h�ET�fh��"O�i!�@A1J� � PxH��"O~� ���`|��H��4=D�,zD"O���BNڮq�e�1�1:[�sB"O���DL�{�:�ѵ��- %�1q"O��B�J��%��H�N�v�ֵ�E"OΔC�d��\����E���T)�"O(�:ԥF�D��5KوeO^�� "O��{R�׋.����G�T��Q�S"O����ݼ)/��戤U�Du`"O��Y��Q(Z�h%y�Eȩ$d)�	�'G�5b�(M�I"�գ�8�'K�t�1���eb�	��퉧���
�'Y�8`c#��w#.رW�\��P9a
�'d�<���i��)0�/�3TVq���� zD�7��R� ���U�4��p�B"O8X��nXI��L�#j�!<�B'"O�j�I�H&.ȋ�땣Y�U "O�	v���$z��S`X�re�\z�"O$�KW�Z�#�N���L'(Y�<��"O�!�G�D�h�x<9��c�.8�"O$�`��?}�d҅�.K��T*�"O@��Ee�P@��	kX�l���"OT���	48rH��#��W�F��"O\��@ŗ�z��#�A��"��5��"O��`� �>�FR�)�/T�"O�YC�iP8$ R��4F:8x�"On@X ǆ5jK��;�薆+D|�*�"O�u��&J(7��Y��M�CZ��"O��"SMH0k��(r�(FR� �w"O6H�!C�K��c�.�3rWd,��"O���Pa�,e�F��o/��L`�"O�xkA�p��p��/дC�6��"O���fU�8nH�)aL���D��"OX�v� ��ڄ8� ��M�j��#"O�Ec'I�35��*C�A ���3�"Ox���A��/t�Ay��VV�:Ȫ"O�IK�Nc��я	��|H�"Op�c����N �]AEA�m>�5�s"O
��q�ā$�|���A�/;�P"O�q��P�z"�uڔ`;4D���"O�1�Z�>��ѐ��$n$���"O��؄�Q�8}���vbP�9�|��"O��kW\q,�{U!D��9�"O�q�Ċ�!:���Ta�_�v<�Q"O���#�T�crZ�u�h�k0"Oȑ��C)}5�P2f�����غ�"On���gͮ9��$)�C'#��b�"OR%
QM�;u�d;�b�)����4"O��[ N�;4^!f�+��X�"O���^
n%�t���� m|���"O�i��#�?Q�0)��^�'Z�tˤ"O�$j�o���l�0W�ر"O@فI���A��ur ]�a"O\{��D�W�P���X!CyV�"O�U��Ί[���(�1K����"O`E� F��^~� C���Q�"O��@�'.��crl��,q:�"O�y3G	��hr.���i#����r"Of�z�AG�&���N���h��"Orc�F?fв��Δ!�f�a�"O� �7!X�?d � ��:��p"OR�a��� `-rg�]�C��U��"O^�+�eݠL�fh�ե��=Z���"O�@0嘐&���ڤ%�<NEV%�"Or�{P�<^�A*U�C�'P��"O4ܡ�h�����P֤D�Q�ȉ�"O�L���ݢ`�<�ūٍ���[t"O�e����~�����꛵�F�۷"Oz]1��޲[
�� "ɍ�~(��"O���h��]R�*�HG�-�ؙ�"O8y��-��fGf�v�_�n�q@"O���Ǉ5}^���]kZx��"O��Vb�=k��#�'���yg"O�#���(�"y�f�V3i�ܨ	&"O\���O+1k~��7IX�@�ĥy"O�P�5bC�G�4�P���q�&�B"O�|�I� ��4� M͒g�h�"O|T�p�Yc謨Ӥ��y/��"O� �}��O�)~x��dN .~�	%"O�)���U�6.�YbQǨa(���A"O,����_-;P�hro�l�x�k$�Z�:�~ճ!���A�t�/<OTxzf �6��A	��S������"O����LH.
xc��ʒ����d"O��y%��^�f%c4H�I�Xy�"O*$r��K+TTq��dN\4�a"O�y�̰g��,)��C"6��"O| �
�>i�tucS�h��`"O��qw�ۼ<��TXT-1a���1"O±	���_Aĩ������D"O*q��!�R�S�e�4U�2�i$"ODTw�J({h�h��
�9�����"O�Iw	O�yl�ը�
��E Z�V"O��1�L�
����&Dr���"ON�x�(�=[ǄQj̝�6wn�A"O�)��^�k_@ ��*Ӕ%g��"Or�)N;�N<��K(HZ]��"O���ǉ�r��	 ��wq�%�"O�eK"��,-�jgK��3�8�"O�d R�=`�<��U�^ . �4�',~UXVbB1{+��t�O�n>)��'��bfFH
M���C3v¦Y��'�"I)�0�ȼ9c�H)[�z���'^�p!��)z�P�3h��RQB�'��4s�*��kk&y�bң}q:��'�d��U��"~�i���@9u� ��'4�p)�䉣	*�	p���qu�YR�'!�0J�雵Y����d��d��x�'����oBR�0�A7gZ7J����'��1
EN��n�����>�<ĳ�'�� a�ƒ>q~*=h�%#RZ���'�D��U�Vj&�@� �J�K�'�p}ɰ G�(∑� �M7����
�'�b�`�^�q�^u�U��WP�)�'���%�e���"��S�����'�阒.*Yc�����w�����'-P}��ǙD&l(�B*�6FRRT��'�=8���&�#A)F�/�`@�'��A;��͗'1�T��]6-��,��'vB�z���UNPA�G�-H�ժ�'��5Ə
ls�(JpG�5I HS�'T0HW#ڼ�����Y>�Ę8�'��h��M�hpL� �n�"�'.n�q��gtA���4	dd���'�(� �l�.%yl˕�כ����'I pS0�]�>k��
�^�Pܺ�K�'/�BC��1}t�Cc�]�6�xk�'ì���,��w��Q҂�1lj3�'@)��1r�|���˄4]�F���'� �A�nF�V��;R慺[�zI@�'C��kQ�ϳ���I��#�'��BP��8kT)Bt-̻p����'
��9W��/
XM���n�̴��'����2lR3^B�`ƃԟ9�ɱ�',����eP�8�pucN�1��
�'b (A֮!m����əR��{
�'DNI����ڠ;�gO�����'J�02�BlJ�QAI��v��'�\�
fKL�3ŒDq�N4af4��'�ԉZ�-��(�`ѡ�P��&ѐ�'n�!�f�gO^d�A
Q �,E�	�'@){e)Ow�"������(t��'^�P��ϨY2��L�vzp���� �Q#&��bS0�R��[�Ԕ٥"O`��͔>�� �#L�����"O�M[Ď0N�n����@��qh�"O.����B�_j�#NK5_���u"OLjD��8G�:=a�MԈtN��t"O����s,��e�ÔnV�I��"O�qKR�	8Wu<*#�Z~����5"Ovx)
�y�@��4i�+]��<�"Oĕ��!h%���[W� `�"O���V�4�ԇp��"S"OR%#N�1i�	zjrA[�"Ob �u��#k����H�>f.\�E"O�e�#�f�R�!fǝ�	G���c"Oh1���hy>���y����"O�AS2���rG4��dL�y,Q��"O��;7H�m�^���@.g��`�"O���B���Y��5i#1�fMSD"O^�(3�W�&,��+��̫?�|hcC"O\ءU�4^�\ HRI�D]3"O��J�*}Hd]��G�8XD"O�M�F�H<*������1���`�"Ox��NՈB�����8Ү1r"OA���
�,C�ɱkZx`�S"O����g��S#�#�ڌ�"O�����+W¦Б�ݸ'�<�h�"O�y�D�1�$QrAd���e"Ol�bV(�Q�\��!��U(�"O@�I'�6PBa��ŲQ�i�f"O��kU�Q�C(4,�#@�?Q
�"O�d�5�[�:
4�FŢ!7ȝ��"OtC�o_u���х�W)^#ĕ�"O� ��#L'.���Y��p�
��"Ov��' �;���iw��<�,�r�"O�ЂdN��Cغ ��m���	�"O0�Ҫ��vHa��Gֈ=}�ّ�"Ofdȥ�P�dV����g�1:Sz4�"O|��`�\l���G.Oh%Ѧ"OrL�w ܳqL̍�3��.j�,��"O�t��)\��0�I�Zڨ��%"O����8�P���źS���"B"OD8�B�	]���d�O�H���"OL�{�Nk��)��IJ�|hBQ[7"O��vc����%'�(Y��"O~1���*OC��Vd�}r��)q"OVq�5�΁l�P�a⡄�S&dK�"O�b$��x3	�����#URh�e"O�R��9l6���+W�2F4]Zd"Oj�p�mɛC���BEZ��%����y�$p5 [�JR�ċզ�$�yrC�v�l��0��@�`m�W���y2L]��mPD畋6�H!�6�y�nG�N�����Ð1�0H��,��yR�N�9%X���"y�a���\5�yr�T,�>}��/$�R�%'�yB�ú���A��	f�:թʛ�y�eճT�Ay�B���b�D��y��Q�[E�D1��
y���d����yR^�҅��5���*�εy��M���]X��h�@�9>��Ú�m�(C�I Y���&��"C]8h�gg")xC�	/}"�N\:R@��W�RպB��;���q��b��"���e��B�IƦY�d�� 	�4����C-.�ݡ�)%D�xP�+z �8�@�l.�PWE D�� �d�ѠA3yG��qǮ�3\��Y�"O�܉�'Lݜ@��Q�>=<��t"O�j��(N<��Q`��=#�mA�"Od�)��@0�>Đf��v�c"O*�!6�]�Z��[ŭ�<t2�Sc"OX4��/hrv�"猟> ~��#"OZ�A�fO]!$���-C���p"Op�a�bOv1"��X���X��J��ym�1&M��Z���<]=@�o��y��8v;� [u�PY��iԭY9�y��1�8U���ڝC���3J��y��%$x� ���_n�0��KK�y"��~X\U��AUx�t�����y  k�j��P��wy�����	#�y�
��4�@A�߯9[�0` ��y2L�_ѐ��"$��b#\��$&Ԩ�y
�F�.���eA#���e��y�n2zX)��)^*�����y��\�XϮ	pU�ӄ�ih��S#�yb@�.G<)�`I)!�$�4���y�G��a1�aP�@�F�����h��y�e�/ADoʄ>� �C`�Č�yB�R�1W��R)�3�8�Ѥb��yR�-c�d�2�(�����.�y��Q�L��Q1�@�0L^�S����yr"X/x�L��IJT�I�#d/�yB�T��$(�oܾEK:�S⎒�y����n/;�X��&���y� Շ0:4	M�h^�Z��� �y�l��)�$��TB�ZK.L�@�:�y2B��z��$�	;T.�`{wKȱ�ykG�Bϲ)c�MЈ�&c	�y�b��d��I��3m�X�Z�"V�y��&���3�5j$�93�̈��y���[�J�c��]� C:}4����'H����D�0�%;�Q�pk�$��'�j��$AΔ )��@,[cQ���'�|��`�v�M����׬q�	�'�HD:��	4D�V:�D��%
�'?���PΛB�ᚖ��8i�<�	�'�*���@&?���a�FI�Br��'ɢi#���:T�%ٲ�D�Bv8�x�'���⣩��F����`�51l�ʓR�PѺQiK&Ld� 1���?���ȓU��2t	�EB �li(�����܀3撁3.���H	}~U��/��ؔ�O���`�˗H����ȓYbJD�1%>q=����K�=���)d2$�#`�*fd`q��G�
��P�ȓp޹�t�ײ>��LHAiJ&�I�ȓDMbpX�gV*i�� b��Ʌ�R�Z���6;�N���.�kX
X�ȓGR,���)��D��I��9��I��f�E�gcֈL�Z���`^�|�N�ȓ{��В���W���W�͆v�H���~�|yI�.V,�Z8`�LLj)4X��'����3�K<�s����-�@�ȓT5��s�![0��܋����(���ȓ0���s���)2`*��v��܆�H���C53�:�v&Џ\��4�ȓ9v��{��H'q��sJϷ]Y���ȓn���Q%�
�v6, ����ո��ȓR/��B��X����(������5Z85�V���z��������4Qx-��S�? �D��F\�a��Q(r��t.n��"O �'Z2���(��P ]=����"O�3�DW�j���kɞ�*OB#�"OdH��tEzI2	ʖ_0$9P"O���,W��e3�M�uMx$��FN�<�7h�W��h7�� 
7�J�<�	��~�$Q����&J�ð��G�<�v�Y�O�<���i�O����P.Iy�<���]+L@�EA6�L"�v\{S&�o�<�aNQ>+�h����e�b$��Yg�<�� �B]��ZQ)�,�^�*���f�<���G�%�q�O��īFk�K�<�J3M�����*Q�p�� �F�<��O�{::!��FR%#5�0W��g�<��Jٸf���d�[$h{hxU��e�<1�o��Q��{�g��i�䁋�@�F�<A���deȅ!fZGp�CÅ
�<��E��@���j� ��u��|:��{�<!B�վJS��Zr��1;�\�`�f_�<���D	;F���*<<�<`P��r�<A��WcX��:Ӎ�#!3� H�n�<��M+FV���o�!?w���ᅝt�<��K�,;&m1�K��	ː� �(�G�<)'D��R��	$�A
`����Gm�<Ѡ�[� �{��ʍ4�^�:q���<�тʡ^D�UCA���5=&�Ҕj��<���X,�8�R=1���x��Vt�<A�G�o��(���K��<����T�<R�T1}�Lu��;Y�(�+GEQ�<���J%6k:��EG8&02��P�<�&��8�^�����.0|2<���L�<�fi'J�%(4�--u�4�S	�K�<�ҧMb�l�cCl|���	%��q�<Q$'�������o0
���d^k�<�UbڜI�F�Њ��	��ȃ��1D�����"8��Q��F�1���.D�,����*qh$����>V4��6�+D�@ a��~��IQej��.����s�)D�P+0B�Út!4�)���uE)D��9@d��kW��j5ˤ����%D�dr4GF�0�b���E��a�b#D�lSucZ�/x����k�A\����%D��B���B��$��f��Uf��+%D�*c%�.o�NpP���V�fa�C�$D���FmSn~}P���6{�h����"D�ܫS��:%�X���R�9Q�q�%-D�L5��
����
j��e��f+D��yGܴ4v'�*pC�ѲaE)D�,U��
s6F��j�=Oa�y�g9D�L�&e�+8Da ����JI� `�8D�H:�JF��C`��fD&�y��:D�������<�U) f�:DYB�(8D����� V��K��ТX �8;�7D��G��	u�ʹ#��L��`�c�8D���b�S?v���AJ�hа�1I7D�\ZA��%�f����p���+�?D�l��'�Y�8����& ��h�w#D��r��}��0zwG�:�x�n#D��8JW��q���3�R��"D���+�o��P��.}b���,D�� �
&(gXt��/
(��%�ve(D��2��re�x�Ώ5bK���>�yB��1?��y�7.V/BE��B���!�y��1Y������D?eRtyओ��y
� ����E$+����4D���"O��b�G:�|y�	W'G@�D:P"O
a�t�XXDB��ŽVxl��"O���+�? ��#ꊡgM����"OB�����_�����ȈL/��H"Of���
k�:phǇ6-����"Of�i�Ȋ�R�������O�D*�"O�\I���1!0��B�)����$"O���n^�#��I2i۬�{"O*݃WFO9>�����k�6i_�l��"OPdP���FY0lT�X�v�.ّ7"OB%�b��cT�(�d�Ƹ��"O2�@�EP��7�}��`�E"O�4ITo�q�^�j�Y�a�����"OFAn��}����@_=zX�x�"O��r��)KiD��$o\���\�"O�B�/_=2D�JB�_, A!A"OhUQ�*P�$apY����u- �"O^MB�&D�c+�)��)h��0"ONU�pfަT8~��f����Lj�"O�5Jl�
B�H*��N@N�QW"O�l��ח�Μk�Hў���"O*i� �85g��g�ڳ>%�"O�I3�
]
���2k�p|,�"O8��E�[4K�D0��L�{����"O��X�g��Ptsfi�$k�<m��"Ob8�@kP���Je�]"X��i�"OVĻ�T�B�����:!��"OPA�zz�p��1.d-�"O��p�KI�=$�Ƌ���K�"O>m�%ΐ�S^��aɮ
(Ļ�"O6|�7O�g�&u1�S"�i(�"O1ۆĄ,l�����++���"O��b/� c�5����+2�N�Q2"OL]���>���x�J��?x���"Oh�q �=8�+�'��,q�ٱ1"O��
S(�)�L��F�����[E"ONM��l�(�^Y��&�vZ�#e"OV��NP=�*hXa� \�"O���smV��v��fț�1�"Ol�+<��y{�J]j�D��"OU(7�f�)��ѹ�DpV"O�Ma�-˄N\��fB;0�� �d"O�x�&��,��9�g
�����"O>@Y���N��Aֆ�2�≛d"O���A��0�y��G��>a�"O �R��[�/�h<�M��m	P�{4"O�9��_�9�L�A�	�q|i�"Ol	�Ql���<H���U`�Y�"OD��Յ�.�n�Sbf��e�ذ�"Ov�k b���l�c�ܓu�le��"O�)�P�� ����c�A��my�"O:܉0�� ��HC�J�#bʬ�2"O��Y�C3"�dP������i�"OP\s�P�&���(1!ݞK�P��"O�C4C�V��(�r��+�bls�*Od9!U+M�+o�i�E�:?�S�'�d�yD�X'Omz���j�5ŸP� "O� �C����&�!@
���Ջ�"O4}�uA�P;BD8㨍""�h��`"O  C�_�x;(�c���y,�)3B"Ob�RsE��Jl]KI]�j"v�"O�AJg��=O���p	Y��5"O �l�C�b�D�@"Re<1p"O� ���H
3p�a���D�-al}�"O�m��	�JX|IU,Z�M/�$�1"O�L�k��Lq2=+��Ww+�i�"O�m����>}Z��W���>�xy�"O����\-d+d�A��$�p#�"OZ���
ۇ�8�#�Y/��z�"O�H7I��q��E�^�x��"Od�j`��7������.|%��"O�T �N�B���"�I�=����"O~�q���߲E���nF�[�"ON(��*@�&��]�F,Ƃo\,a�"Oح��� W�İR�E�BU8�C�"O�0s���SnJ|�I�M��})D"O4�G&��o�I9�H�'L���b"O�<I�]�P�@�ف���pY*@"O\<�b�06�
�
��A�r�Q�"Op$j ��5s�u���m�1��"Ov���#�(>1�islY%!����2"O* ��V�/��)�Tj�'j���)�"O(UQ����l��@�G�C�(�b]!�"O>�#R�ޘ5�u��E�V{�k�"O�ժ��w�l��B�5g^us"O��@w�ċ4¢��@��'yq`i:�"O����Y-f��R�˜�WW�5
�"O����囓0�z幱��c��)c"O�5�B�p)�d&`�~�jE��k!�d�!��-��k7ܐ�"�I�!��ȁ}��cv"-�����'3�!�D�-�!"Ǐ[##�ޠr�GV�'Y!��ąx���$�ʼ&��\�r&�#2!��z�\U:��"^ވ�)�"
u!�$˞b5E��+>*b�he�8>!�_*j*��Z�l�(��Qt!��u�R�J�L�5&���+�;D+!��Y� a�e����<&0�kӈ2�!���Ak��":�V%��!��?t<�4�	.�.Ȩp	�-!���WWzA�"�ې:U�d	$��i1!��_�Ku�i��(D�8�n��O!�$B�i�I:�,o;��Wo�G!�Kh�j���p3b�I��+!򤛩|0��$,�-j�tt9�P�
!��[<	���b�%��|b��E�۬	�!�Y�0��:s��g`�yۇ�g6!��Z�>��M�#�J6M����T�)+H!�D�2<�	+J�&��Z���&?!�> �n�����*��14�Q�!L!��4���!A#�ZHy2҅u!�D��qOH41fU��8��%��|!�D���v���n͐$��`ǉ�Y%!�D�� �6Q ���>�W�"8!�
�%�f(�H�m� �(dh�)(�!�C�A�L�H��ᖩ��N�!�D�?g��� P8z��1�7n��^�!�ę�Y$�����&��ܓ�џz!�$�? 5jX9�������Ӕ�>5�!�d^5U(>T	��I4��d��<!�$WA-�p����Z���8C!��ƑlP�R��J$n���p�S-!�!��6��0�� �iW�����#G!�d�(a��="�j!L1��{"�O�!�^�eb|�� �ְ'l��!��To!��4F�> c�푃"�����V��!�d7;��x[3烿$�>����\��!�� ���ZJ�\��RNX�HG !��"O�hKbN�w�LD���AGB�)`"O�t�`薡c&�����D�)H�"Ot)1��L�.�d���h�;�����*O�� GE�;n�xz�[�P��!	�'��|xW�Y8o� ��ڥMM���'�Q�c˜��F�C�<EX@��'����v)�:r�9�+�@eP	�'d�my�o~�ĉ��;��IY�'UV��T��9h����3��5@	X�'/R���Ǜ�5C0lЂ	w��D���'{<T:Ձ���5է���E�is�1Ira
h`�`���h�X��!
�l�U��JI�a��
;^q����w�!�!��OO0$�!mT������4eZF )���UvK҆����k7%`�F�a�E7�\c�P� �ޮN�����)j��ڴ��!�I��M3 �i��s��(�A���a#T��W/�;���4�O���%�O�eɴ����f/�bGTt�P�O"�O��lڭ��O�2�̧a�֜:��{n����7DpY�(��E�M��9F�m2���d4J�Jg
�lڱ! >It6�xu��dUxd+��P9G�ԁ�U�';|������"�K�m&����C�2;K�@	�������"�����I��e�&Iį���V0Dt� D�
f
�d��j�-~��!�\���OړOP�D�O��A�"i��&W1s,����G�d��I�4F�Obf��<x�*Q��ʶF�����CP�M�����|�����$�-�3�g��`y�'�պ_RUE�%~�����OrVB>-L�0"�J(��je���:xK����5�fd(!.V:f�KCU�'��a�7.
BN�&�fU�éU�a�8ⅭG7%I<�i���ZZuA��l����=��F�@l�����A��o�R�!�Вs�K��xr�')�T>-�R,�95�! C�ŹK�QХ�ޢ��xbiG$)^.A����F��������~�pӜ�lKyr��	m7m�O��į~j�`	'k�6y��ĝ}8��@�&0��v�'q��' �p�^ R����D��I6�kR���|�BC��?���T�g?D m�v�'�f�b�ʗ>�B�w���@�E�v������d=�8z�+Ɂ� 5ZAe�r:��QU�Ā91b�'c��6��+qfꔐg��f֊�z� ����IM���h��׮#�ْ�L��h�b�v���p>qB�i��6�w��x�'M�5�n�9P�G�_˚��~bA��e6��O��S��x�ϝV�\ݹ���3�4�q��=Sk� L؆{�����G"1`d:�!��OU���1pأa�IN:���JqH!n�Af� "�C�&ڌ���E+~O�`���σ�F�Q��~�1 /��jA�4�Y�1���E*�QoZ�U-����O~ԕ����i�*��d`�����Ò��4��J�O��8���<y�}�
ǣrִ���M�u�~��	��(O��lПd�I�M������P�k�NE�t �Sx��@�n�
��'֤s"n�<-8�'1r�'��J��
Ta�|�u�E�Ro(���"@��]���K�d_���c�*���4���$X�l<�T�1��=Yb��+.SUP�����U��d�8B�2u;�S?��ٴk&�
�-�<у����3wJŅ�g2X)�'l��S��?���x��'�X�L��AF���<-��4
+�	R���'-�̰�!�Y -���0J�+5�����/s�l$oZB�i>���L�I�ɺ�j   �   ]   Ĵ���	��Z�t�ʔ*ʜ�cd�<��k٥���qe�H�4͔6Z <���i4�6�<�TԇK��,���I�q,�m"�M��i�F��D�J���PEK�=������0��1Ï���M�A�d�2�O̨ٴ4e`U�5��nzneP'�R(f9�'���1�.���q-O��qo��k�<(Oh�:���*soұ �dV�O�r�2)��P��-O��I�b�[%�?�ɤ3eR`�W�MW�|t(fNM/��`��e��'��u)����4~ �KW?2A�1P�@8RJ/u�u;k�E?�eeD�P�?}"J��l�~	�M~��
S�qĢ�x�-[��n1����<�@�5�sv"<9c�Xb\uA��B%N־t��J�~�T�%ቕ*C�I�lS��Hi~�Cd�!K���'-: Gxr��xܓ~��IՄ�4�!����FG�\o8V�h��� �Q"q�Z�	H���$�,\�28ya$7�	����a���1���;P�:0���H�Œt�<�H5�����zqO�l!�,�v��)���[�"Ԑ�x�	4/�����y5	+�PB�K�Ϙ'hP�Ex�
�u��%}y�9����	�pH  �?�*�I�5��hE�xb`��l[7(2[��Q󴅈�^p@�(�OP4�-O|�雡4�1��q� m��~�MK�j�*���wv*8 %g�@y�2\>�� 4}�i��|��J<�
/�����Դ4�2���"�0TH@"��s�	 7T�"-�^���/y��DM�]_�����b��B��1kp��  �OV��?1��?���ܠ�JaJ_�*����u�P{� (����?�(O��np��IƟ������a t[�HS���X�����$�g}��'0R�|ʟ��2d+[�p���)>ԑ�U-({A��3$� 
I�i>��7�'"�D$��X�#ف:E�T	T#�^�9���Wşt��؟t�	��b>�'7-�4�($� !��"�p���V?��E�!��O&�������?��^���I�O*��K��LD ��*E'���	��@����e�'�R�q�#�Qܧ
NDR7�Z�D� �s�g����$�O�$�O����O��D�|
!$Q�!p�)���U#2L��hS�n��������'������'7=歷��F��k5�墎�\��͉�e�O��1��ɏ \մ7�}�@)C���X�s���    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   

  �  t      ](  �0  7  _=  �C  �I  <P  �V  �\  #c  ei  �o  �u  -|  �   `� u�	����Zv)C�'ll\�0"Ez+⟈m�R~��8˔�DBA��a��/60yfN�%w��U��&��*ADu�mJ�+Vi6�;n�$QA��<�Dћ��n�r�rgȓ��V�J�����l t�T�-�O
+~u�7�S=3�̬�#��L�s����<�D�{G�4ӧ�4��r�BL5i*��DÚT�z �	��:�dIM�0�R�Kݴ�|L����?��?���T��?�~!��ˑG�Z���?�ȭE<��\�X�I�+F� �O��D��$��A{��
2�� *!��ln��d�h�����Oh��B/[' �	׾MD���?zhȞ|lE�Ƶ��5�QjP+�!�7ns�JvB̔T���C�x��I�<H>��'YREq��Q�d䏰�Tu8R��w���qAP6�?9���?���?���?�����v�KhR�kC$��m֯.�^%2�� ��v�h��!oZ��MK���&NnӮo��M��W�����Q��`)#�1�L��#�	^>u����\Oh݉Ƅ_�j)�a��>~M ��(LV�����m@ܴ{��O���������X��\M����5,���� ��n�1�90L�!?�S��LYr�̛)%���۴o�$f��t�_�e�t�#d&F9h���r��R�<(�7�¶Zg��o!�M�Աif���E�3.P���Δ$Ё��oȿj� i`�%�@��
Q��3��٫FM�� ��k��,n���Mc�E�����F반Q�+S5*��q�ë�EM������(�ؔ0P�i� �%�!GL4����P���';�O޹�`�Q Rn���tŃ�x�N���-�O���	۟����M͟Dѫ�
D0.����̰v}rQ�6�'��������������R�@20�Tl�p�*��������|9Hd��蒥)�����5W�hX�B�N�W���)BAXܟ|CS
�)Y>�A6�øt��l��2O�@�B�'2���#�h~d8���9#�1�?����?����)��.���'$�*g� �s �<Z�R��O����gט(����'@1]|��'�'N�OX͸f��Լ��LW� �yQkě$n\ɓ(�V�<��FQ�f��\��(�o���e�[x�<iA.�5?5@��Q�s����a��O�<�&�(��B�@�'؈`�KPS�<�� �$4�R���7�>��'*�X�<��e�TԈR�J��`�F�Vҟ���b7�S�O�R(X�&�[����GJ)T���"O�4��I�>
���f� p��x"e"OR�����Q��@3���	R&"OD �gď)`��у%��P����u"O��S��&6B�CTTM�P`"OL���-�=l�t�r�̸1=�(T��(��4�O��zqj�$A�q�����e"�"O����j�$= L�9n2Ջ�"OZ��P�Z�h*�1���7?V\�(�"OĸjP��7����� e+Nh�<y6����,C�o�r1�T)�"�Jx�[2����M��O��D� �^��� %NJ�u�f�2S�'%���|�Iɟ�x�nZ�N�[s�ft{���O�a�`��Z�Jt;7G8�cA�''�m+�0 ��\y�hR5�BH��08` !  ^�j��w�ӿ�0<��؟H	�4Q���'d�̱Q�A>lZ����DN23.�P����Y�S�Op�\s�`4i�
U�Փ�YC���2���Q��Z��X��:���6�?AI>����6�T��|Γ�yfN�Fh����(I����4T��y�H\�}�*5���߹=z5jǊN��yB�6P�,�*���4�p�9vɄ��y��B��x�@�ԅ8��hUҕ�yb�.	��G�Uy"dhJsn��y��xc�HS�pbd0��I^5.ٛ�|2%��m[���'��'B�	
�P����M��)&g���)��͎ xX��44,��cg�����f����XR�	d"С���
G7J���O��5OZ��5��� �HdWŖ
���wA����Pk�6)��ٓ���|��6nM�!S.O>�hV�'G1���'d�	@2{�,�x��o�ذ�А<��	�ly�O*�k6{�@��E�߁/p@
�Q��ٴ}��ƒ|�O�DQ��P@���W.�x��@?2m�1
�e�;j�0�IU�L�F�
[C�Ҥ����k�,� �C�ɟl/e�T���$
�.��`��8�s(8�x�TAQ�vT-�E�%^b�q�0L�}��$�r����`�:k�t��b��O�� @�&D�d ��"T �h�3ǆ:w@�!A�#�$YŦ�'�����2��h��s�H�
�� �S��Q�H(�I}y��'���'�z��a"45� �r��?(Cn�n:� �E��j��T��4��EM) ź�D�'`�l;"��
%�����P7-���4\��j��H��0� �]axҁ�?�?������Z���9�ɛ!�`$��FϚK�'���'hR� ��%*�ʹ�FA�5CA���
��V�b�촣��h+��� �ͼ�?�+O$L
"e��$?E�O)���=��,��#ԥU��4�G!�=6�2�')��˶JA(i{�\+&4��n:§'��Y(�$˘��"������'P��K��փ!Cf�:��\�?l"}�0i�.X#�5*t
į9B�x�s.K}~"��?����h���䗽a�=�F��8$!0��]�C�	�v�]�3j�;C�n1�g%^)A�V�?Q���.i:0p�6��x�JY�&��lǟ��'	
q�6�O��'��Q�p �OI�@ڌ�cCD�Jaj�F3��y���&=���O�xb@p���y��i]U�M�`Xą��;��|acm�A��ߴ(�P�ATH�g�n&l��6��%r�l�bb��`>h��D~�����?A���hOBL�$�S2F�+���cF���)D�@���]�����Ӝ�`]�Pͦ<���i>y��y�a�+
Ӗ����ƦB�`Œ$���u��=h My�^�D�O���<�|BL�]q����^���T�KRҹ��!M�y>t�2��9D/���ĉ�z�Ɒ��G���D�	u_|���ϓ;����c���N�T���I� vh�᧤ϔ]ƌ��$K<J���g��O���*ړ�O(7��1��P#���,E�L� D"O&��F������L�|�VX�I����u�6�'��I�B��K~Js��2M&����L�2ND���R�h�'r�'��LYJ���wf��7��d�������7
Y
?�ŻuB��W5�T�=O�Y��S���=�bnļj�$n�Z�rͱ������	T4���N%Z��'N�	�t�^���ƛ"D�]��3��O��эs���q� &�X��t�� t}�"��O�܉�C�'k�P�2Eg�;SH ����' 剟Y�%�	C�S]���'8 q
�ۇP3z�� gP��A �'A2��5���O�'�����٦#|��(4��Cޛq���Y��n~��!�����Ϣl^�`�)ҧ��p"�ȗ- $,L�P�ѣ}
B��'GNX����?)��)v��㡌�O�R�(@��l&��È8D��r֩� ��W�ٺ@��%�gh7�%W�>��G�ޭ,�f�� %FQ�g��ۦ��������)h(��1������Iߟ��I�c'�ϜU�Nhz��*,��M3a��9E�lXP��	=�?AP���$�
$�|�<�F<r �@����a��#��9]pT*Ć���?���ϫ	L\!�|�<q�._�����J�h��:�h�ڟ8�'�!����?����ǘP~��CN�V����	P�1�B�'%��p@�oL�����3��A�'�T#=ͧ�?�)O���ъ��!�`sv��
(sL�iR�ݶ+���cP��OJ��O�������O���"�D#��!d��w�daT#�>J���R�i�1)�A��w�	�%K�;tӌ���@L��p�aA�n�r4o�) a{�훠S,=���ȸgإ�E�͆ �q���?ُ��?v/r��cK٥|JR�Ir�Ė:��͆�p�i%R�+葒�!E�&�li�4�?����^���4a΍4���VO3��H����yB��]��ъ�F��2�N��مȓn�d��V���hh�h6�*K��х�3}�̣$/1R�(d  "��Fa�ȓL�J���@ug.m�� n�Ʌ�PC�u#�ƞ)cQN`{�E��[�9D{�����r���)�ĴC�\�g.�u1�"O���h� �RIc��Q�B����d"O�����ſw3ޱY�B������'�Vmے�կ~~B����s���1�'�B���&YXR��!ޗ��
�'���
�%��ah�.C;}��9��_��Ex������LS&�ֹE��dc���.�RC�m�I�� �Z��HЁ[�0C�ɛa&v�Pw�ćC,Ҭ��k��k��B��[�0�)#���j5�Ј=n�B�I�m29��AAb���C�uI�B�I���d.ŋ&�*��n_�C���k�d���	�$j~�^b;�����C�bB�)� FlZ���):�Qjg��2�2�"O> A�V�8��6fC��h���"O��$��:z �%B�$��q;w"O��C ��5
�x�E�$`������'b;�'?�)�Q�5v^�q���GOnͫ�'�@9�S���X �ݹ�e����-��'a�2R-"!m}� !^8t����
�'�\�[ā_-?�P냷�VAC�'5�\��
۳1�Z����&Pr�'㰐����qK�0���d�SQ?��qT�/�v}b�A�J�JԢ��&D�̉ѣ�Y�����k36U*��+0D���E�?.����.G�����-D�����%[d4��닆o����-D��@S��TFh	� ��6����'a0D���b,A	N�>��֪�i�Mp%l�O�i3�)�;�Qd"ќW� +�L�#�����'0z	��T-p��=µk�:!�n](�'��R�ډrl��8� W �	�'V4E:ȋV�D��Ч-�Z���'A�\�2ß͜�ae�W�x�65��'<����JI?N0��qb��w�р.O� :��'E�Hڃ��4A�j�����in L��'Q(t{��1bz��#�ΣX���'�1f���)I�vV'R���	�'��a� �$�9�Ḿ6^L��'{�HA�n��Bi�W��6j|9��I�����\(⁼{PuC��ڔ"�vԆȓ&��0K⨀�^ٜ�	f�C�o��T��jbN�Bc�(D.8�  ڊ`��مȓ8�Tq��.-Y>�
v���	t ��ȓ>�*����Rj��:�I�)bH�ȓ�QXe%�S��8j�DNv%&�G{2 _����@(H�AϯR��kS�@,nM���@"O��"֠ފv���aU��rCr���"O�x;AL>lD�h۲�X+�
�"O ��HR)YSh�DFS�,��qB"O�`c6�؅D�p���+[Jƍz"O��(�
P+K��("� 	d,p��'S�HI����;|��J�e��S�%�(2�ȓ-���q(�<Qe��[i�1@8t�ȓF/�` O��R���ǍX�7�Q�ȓ8�~080lڿİu:RfG�f����u�[0l�2^��ae.�G3D��:k���T�	<�  �#Ʉ^o|��'٢�5G���0�F+i�$�4��)8�N�ȓT����bA�;ak�-�$�=����3J��m���������11`��ȓ/���0%�$L�x* �H5`p��ȓjȘ����Z9~ $�a�X<?�΄����@0��Fw��Ǿu�~𚳡��|B��h�TT�``�'C{!.�z�� D�PY�
��D���[[�(U�#D�HkC��.W������6O�:�w�4D�s��S5���5�K9	cd��0D�\�!��1Ͱtcvʎ@�i��� �|蚵F�Dm�~fX�dǗW�@pȓN[/�y�B- f<���gV�@涀Ȓ@���y�BY!G�>A�%Q)M���3Q���y�'��;s41c��.��\B`��y�Ȉ�|���o]�s����T�yb�G�0w�9�-��]hU�G�P#�?�hEL����¸9�E�#d��LK�AV�{����6D��2��6���j4m��$4D�� ���� %�����+6j40	�"O��J��X+��,�0��gh�IS�"O�I��F�Y�F����Mt�-�D"Ov	f���вG'�Qn�Ш�[�(q�$!�O�����0� ���B�wz��P"O�!���ґo���'P7
~J�0"O�!#�,��`6D%*l�"Ď��u"OT���o��AԱ@SD�w����"OZi���?�*8Z�a�t,��v�'��<Z�'؞t"�v�Аe@�5q����'3p��T�Y������.�LM��'fJ5k�m�V*�]�s�p��EK�'�*��Fe�F��l8F���r��$ �' ��z�Q�X�ce�ޫAkĈ(�'S���M׬lR�-�8w,����d+JzQ?�X�
�>)�ݡ�F�>�U0�� D�@s7@��l��ʇ�(}o���* D�l)��=q�`#ՎU� AxAE�+D�Hb6'NH[�m1��؍j�����*D��k��G)v�@i�#�(��P�t�(D��zw� ET��!��VZX�tQҬ�O���)�'
�@���|X8%�!.�8���''`lA��"1��w"��6|�x��'���!	�՚,��+���p�'9�pbbj.�®1(�h��'� )�Q���R���J�Q�'�������<P �a���W��0!*O��Cp�'n\%̆='��h�@�8�p���'��!�
A6y��� �Ց.�l ��'1(:Ŀ��S,@�p�Y"H��y�㏓���M�&4as6&­�yRǆ�}�� �� Δ`@wg�%��>���Z?q3 �����H7V|�iæ�c�<A�N&!J���^�*��T��Ny�<��H ��83����g�a�U�x�<��`���\��"P;a{d��u�<��g�4���ݴC�J��f�r�<ٳW�f�Aӡ��Zy����kC�'��:����
=2V�2���V`�e)݋\!�D�k�N4`
]쥹pn�4[�!�䕤d&(���-(_p���G���!�$��1C����/��T^<1�A�K!��[d�� e��!s�58Ո]�-�!�,�EP��JlH�Q �0vk���O?Y�f%���CAHXom+M�`�<"V��B��M ���`�<�u��Tw����^q��u��N�V�<�dȃ�y�l���,T��X,�u��H�<AP��,�t�����=�H�b�F�<���;��FC�hu4�ACCy��ǲ�p>���Zd��!���4�s'�e�<cQvo��q!c��f[��@�,_�<��Ԉj~��P�b�="l�����AE�<ai��@�T�hR�ĶT���2�HW�<��')P<Q .�6-�F���o�kx�x0�����5Ő�*�5�OW��}b D�L�b	���
!�S7W�vi�`?D��*f��_:nt(r�V;d9�G�>D����@�w�ų��40�~e�C�7D��A4�J�?O؁���U�=�8 ��5D�����($��eSV��!g�l:!
4ړ/�^�G�4ƀ�,OA�N�D(yH�8�yb
[�	0G-yR��8'���yb�I�[�`��I�5xl��6��y
� ¨��*%���®�X|~�{"O�HU�YB�<l"Í�lx�j#"Omy�D4:F<F�T�f��J��'�������SY#���]%6v�X��1k��%��o�$a�q�;�f`Q��Z/G*I��_5t��H�<.�<��*�*=�� ���A���"/�B����(zm��ȓv|�5ѧ�68�qeF 4^�-��sD���5FF��(�6@���0�'K�Ly
ap�ӎ{�}�L����.X8�3���b\4�b�Ύ�|���N�p%R��ʃE�R@�螬7<�܆ȓ]�sg$W
/��m(�l�%Rd2���
<x���1M*� ��cZ$0�!����O�b���8`��H*x'����JR6�
C�ɔB���#+�=S�)P�E�"B䉧V\�xaP&�f���B�n	�<�B�I,w�©I� ��@��;�a��rF�B䉴m*��s@ţgz���F�.C䉆'Ex��dD�Iv)�s>\��=�S�n�O=��Ȳ
L?��V�
�3���c�'��{C�Ǌ>�Νk�W�/ںܓ�'n^��A�	&�q���K!)а�	�'�� Ц�^�m�r��hESp����'Q��*�=������M���'��Py���<#���p�ŕYd6l��h�5Dx���	_t\Ȃ�G@��<)բԟ^Y\B��[Gr�C��R?s�,-�/ߵw!�B�I�D�(�%צU%ș0�)
�;o�B䉴E�P��� .,��9%L�\BC�	�giN�!g��%�YX�l��^�C㉋i�B�ʁ��Ir�q��oL� �ĝ�I+����#	���&K��I�B��4�@P80Ț�B-�c�ɟ����O���O��!�"'4�g&�O����i>q�2,Y����Q�Nz�8af�)�&>���ƍ���H���Z���)�?Xn�bcbXB:��yd@�%�����O(�!���bx�glC1�43�	�$b��0?��BD�&u&l�u�j�0��FNEx�`0)O��� 91��T[�n�א%��Q�`+�l���X��Ay�Z>���� IS`��,�ĭ��*-kT)A��0�n��y��U�2��+v��,r�S�O�2"Ìҳ&�0�8�AD�WQ�x�'���"��tP㗛 ��?�p�K�'3 Լ���g~:xQ%k�`*B�O:��5?%?y�'�r�b&9�(��@�S|8�a�'2FDЀ�6u(.�a� �R�b���dXs�O�q�5Ma���+J*Wjʈ
��'���4N�)ڴ�?Q��?(O�IS�p�l�!�Ҕ]r�t�r`�L�U���O��H��G�>h�ax��Oq��=1�G�x�����LD���A�O�Vɱ��0^<��b�.�j���O�Y�P�˭:{X�{���Z̨�@ᔟ����O��$�On���'!����'H\�0�F��T��y��Q���ʷj��]�e�"!P�X����	�HO�i�O�
6(��UΛ�[�BA�(�1"-���
ɠ䛦�'B�'�)擇+��A$K�\8DigH1hh	�A��E���
Fꦉ(�.�8��u�Ζm�����ټZ�P�r
�>H�@�8�d��9�Hu�ϓK�@��	�=ƀP�`M	TJ��b� �;O��������?���I\� ��s�=|����2_�C�I�:���BV@��aXY���o���'��I?Mb%p��D%R�C㒌�����t���o��!�I���I�\fd�"��.�m�tܣ��|��'Q�G���7(�[� mp�h�J�'!*���ܖk�Fźq�^�:��?Pi"ڑ�F���%NV�%#�">�7*M�h�IW�'u@|ꡩ��L✽�&GϨtY��'�a~��4C�Ȍ2`���0# 9j�� ��>�Q��0��?,� 1S�Gެ\�ި�&��<!�̌�y����'P�I`���'Q����c�����8���15�[�A��B�(�"+Bw6�8�'�O?�i �M&)�b]����x�n�3
a�$�q��T���H
���4D�4同>,���b�Ri��
�Ʉ�y�B)�?�������$��� �{���I��KňZDb�iP"O������,�rQj�g��g,hy[�퉸�ȟp݊��ΡD����hK���� �Ov�C��X����?���?�,O���8S`p:�B��C4�3"�H�wA����O��'�N$3=B$x#�?#<� O��/�h���䙌)k��aq`ؘ>� ���7 vm�Q��%'��O�u��\�g���h|0�V��,����OJ��:ړ�y�D2G�Z���+B�q'v�"���yb̟�S��Eˑ��lm�=
O��?���i>��	pyFO�"��mC�O�" �j�kӷ>^���'�2�'�bQ�b>�CM��]��EB N��%�pP��%p��Ag�7´R�炜��<��OF� ���ñ��=��hE�!A�\d�G/��H�����<)T�G͟��pJ H��j��n� �'&ZßE{b��7:��d�¨�8>1<���I�
B�	�Y��!i+<�����`���"S��'x�>[x���f�$c>�+�śj;�%8uJ�'&�:��OPФ��Ot�d�O��R�/�z@�9�nK���4�,8"%@B�#�-BE)�#K�F�q��p���t�	�U���qO|�S&�4?v^� ��,�
Ѓ�h�'t�D���?ъ�T[�JIzI�5�ʙ�7�µ��$9�O�u`r)�!�t����O}R�a �'���`G���
7Wa��A�K�",$0�'�R�'�R��8?	ǌŖ\D��ۥhN�Ux�r�C�~��F{�*��!�T�Q� NYE˓�6��'|�v�x��ģs�T%'"@k�z#=T� �'פ�I�T�lӧ�9O��W%�(���d�6a��6;3��lR�{Q
�O��'>U�r�_-\�ƨ!Q�\�,q�%\�*��:G��=��<�w�A<�t� V��8fײ h4�P�b8�O��O�ۥ�>��[?5�F�5Qz$qA��H��C�O|�Y�>��
J�O:��RF��=8"@(�@�ղB��%���'c��{L��#M��H�=}��h�4����	M�~\)��P�V�v��t]��aE#})%�'��*2HL3B!Z�<�H"��Q�S��[�
.�S��'��,P�Otq��m�,�t9� ܾ)�!���${�2�q�X��'�|�D����:����tE�$oY�a�K��?�C���`�L3?��y2�נ�~��]2vR�`���_�/G\ԋ�����?I�.�O��`�K�\Y��gG8=UjE�"O�]3��Z(8�0��� ��6iXL�v�i*��|r�~�'~�s�"��A�&@��"o��
d����V��$�,F{���QR"j+w�4��R�S�aOly��"O��1A @�A-2�#v��;�ܠ�"O>�zC�����B79g!�"O����>0ߊ���d��iG��"O�Q���}`�=:��	+:�Q�"O8i�!"ζv�U��
�i	��Q�"O �a�䵩w��)�P5�"B���yB$G�`򕇘5W~���1�D%�yb@�P�� ��
�QGҀؒj�y2g	,Ӿ��g=_�VHJ�!��y"�����S�I�(KF��6G]��yr�Uh��4DD�+�&�f��y�fS�|�ڱK�"��#0��i�����'L�]s���Z��G��+WVD�;���0I�� 
E.Ⱥl丩���3@��Q�A[-$��k�%B�M��N�O}le�A,ìX�h	�a��)|�l�Z�FT3�
�*�)�_���2ƍ��ܐ��؆H�Q������bF�
\�HE'\�4�9��MT.5W� [K>amU-,`���C+9(��KB�<Q�\�/�(<��H�2.��1OI|�<ɵ23D<�"��R/6}Bt	�E�^�<����$�r�@1��6+��b��\�<1���1iHmX��[�D��T�YR�<i����.�2w�+V�h����s�<����8'�>̂.�#y����ao�<���޵c�Qe��M�l*� VS�<A���.�ƬI��0X=��qE�X�<�t��Z�X	e�N�?�`���XU�<��LIq� �JÄ��mq�/�T��L��8�Eʋ�SNzQ��a�9/Z8a�ȓ0�6Q�Mܤ6�D��+2Q�=��S�? ��	� �񉄧�-[�ya�"O|�2���"��]S�6/[��q"O ��Vg]+<y�tRq
:���"O�����;	�r!�R).�6	�"O֌���W�Od��)�3ژ4�T"OZ������@C�%
�'�@X�v"O"��r	�$;�nX�N�%�����"OXԥhD�&��$�H(��"O�5 ���T�rC�+��d1�"O��
���("�a���b�P�0"O� �5Ƌ>m{>麂���,�"O��	s�\~Z���Ň�+; F��"OB!Ja��
up� 2�J�Xm4H��"O�`�dN�,P�En%XkZ�"OB�;G��e6��9.[%qw�iX�"O���t�6X�����-ݸX���@"O�<x�Q-���0J��W�r�Q"O���#I��S�� ��Ì��\+Q"O�)�m�/h����({ߨ���"OLh���|7JP�`� ��"O�賔m��GQ�� �K.�,�6"O���ѠM&pa\���*Q��:�P�"O��E���E��D�7�[��T��"O؉H )�+��Z��[�4�
yy�"O��� KG�48�����c�>���"Ozt/ץ �P ���;4����"O�P2�G�W�&��/WX��-�"O \cEHJ����6��x���aW"O�D��*�	3.ā/��"O<rtl��\��!g��Tˮ\�"OT����|2�%؃���ZA*""O�!B�������B���� H�"O"���J�rf8� da��M�\U��"O����$��
FG'~�Y�g"O(IբO���R�_C���"O���cLB`El��T䇀	Uj�`3"O�5c�5����֘h���s"O~A�� �#���.ʛ]O�tS"Ozl����sҠ��f�(FN8T"O�ܨ�# �+�*��KF�45<�g"O����c��bdt�ȧO-�%�"O����R5���+%�A���My�"O&$��/��XQ������&"OA���ړ@���� g��!�q"O�ԛ���9��#hֿz�����"OJ`�D1VB��BgΌYЪ��"Oh\�6&�:�$SV�@7n�D{w"O|�I�'lU~���.`�4#"O\LRaEX�["9��Ć&U_��b"O�HW�s2�;t#%r*`��"O����֞;�6�@4�P�0e��!�"O�CP�ɀDK�(xd�ӉB���K#"O0����>3,l<��IĥJf���"OF0�&�ʝS�2uP�)T<�`�7"O��z6#�=��a��f <��UR�"Oؘ
���?rФ pgF��d��"O�}낉EU1��1UH'��H¥"Oڑb��B�d���-I�nqɵ"Oh-ё�Y��9��J2� �"O�,X�k�A��x ���t��Y�"O��7(��W��-Q!�J�9�:A�"O�aߧGK:���u�b�p�"Ot=`�Ǒ'Q�P<�!hM*�Թ�"O�@0WbLN|�R�銺DzVh1"O� �+��*+HT�s(O�o�D|"On|@�ņ	�Vh�&

�F9"O�4�3Ɵ�v��D��.��3��[$"O`�rAd�*�z��I�	o�x{�"O,�Yf.-�f�2��-g:�Xf"O�����ҡ|`�Rc'���p0"O
d��C6(��G �B�q"O�`I�(�3^+ā`��X5u�ꘓ�"O��Q�)��=
�n�H��C"O>d�C$Qٚ  R��+B`]�r"O����9~���]#J:��`�"O������43Z���"\3hh�"O�y���M=i%�	:d�ө:V��r"ON�8�DM2T���U���,�"O��0@J��b9ubdQ��#6"OP�y2b�bZ���A!�*Jjј�"Ov��T�h��t�M�U)$���jĖ�yB�� f����(9c!��H�h ��y�-�?����hV2Z��3��:�yb.��IaQ0/��"&t�qꅘ�yb�R;���I�L�/쵐��Ӷ�yr'�>\)D��5mI�f�hA��3�yҠ��`!�
�яul DT��y��S�a�~� W�6X:�TnC�y��L�E��90�L�s
��s�6�yb�@3h���!�&���ȕk�5�yR�#b��	��~�X�um�*�yD]���22��A�䜩D�P��yR�-O�v%Z���	*l�j�o��y�I �+�q�M� Xݜ�1�d��y��<Cx�\ؔˍ)8�N���C�y��<in��Ú2#����+�yb���vB���'*Q&3F@�5	��y��
	hy��/Z�:B��%��6�y�	�2��RC�=*��3���y��O��eH�)g	��.I926x����|c���	�Bϛ�ɇ�pH8�gi��RO����]�b'�`��\}���]$e8��&�5M����ȓ,�z!�Fa�4'�@T�J�XEz0�ȓL�r�ۖ�W��`,c"�^���ȓ]I�2��
&qG�Ia�R ԅ�'90m�"�L�t���N"���ȓe��X��͖4^Ǿ�U��*C�t��6!N$Y�NG�=q05�`��H��܇���q{�Ƙ:;�$�å�4�^���.~�x���RL�(�.���9D�0Xa	IIw�y��L�`1C�$D�,5 ��ED��!�S,h�4���"D�be)nd�|X�R&<\��?D�X #o��;��X�`ݖ	����o"D���"�R�e�X4�'#�aǸ��ӆ!D� �eþT�b�%����#�3D�HA)?mQV ��E7���B�2D��zƥ1��Hk*C30��l�P�+D�����
'P�������(N?�P!�*D��"Ԃ�H^:�#!���֨���:D��Ð$<�r8т"�"�X���D=D�H��
���pr`�P�5�|� �l<D�lȒ��%o �}�E�Z����:�7D�p��L�>9������}t�Q �'4D�ȻP�G^ak`?���ӥ-D���v-C�\ɖ��Q�#lp�SV�8D��j��7�x�kL�G�$D�� �z��O�"TQ1ۇK̄Y+�"O�1� �tG���1��*��1ر"O�]3S �y�`���x���"Oa��$�:9�T�,Y�X@"O�U*����J����唉]��"O�y�����i�D]�B���ʂ"Op�:���:W\3�Dֶ�bhq"O�l.`.\�)O�!��p�D"ODE� I
�+-l� HʐfH+5"O�AasGA.e��z���4�x�"O����iֻn\$���Č�=�c"O�|��P�����.ʊ1���"O�a�&j��8Y|� 5V�~��@"O(���VT\� ��)Rm8@"OB��R�Y�w>آ��K<r"�0q"OLQ�����
�[DF�s|��sb"O<q
�k��H�� �ΚSi�4a�"O��цhӵg��=z�+σ)i��j"OF�X0��8��@l� AQ�؉g"O.MᷥU4���!e�FF��	�"O��YT��_�vH��
@cx��"O\�w��	f��5"D�)��"OHк��p�F���ȏcM�!��"OJ�1$`=LefKS����9�r"O���oK�z8��	^; ��"O�p��h�5rN����H�R"O�����	����C��T�~\��"O^�3�I0K�̥#���u��$C�"O��č_ɔ�B��ٰ/��1��"O�H��#�L�X�ɾ@�0��"O����G�%���C�uʠ�9$"O���TSZ�	
�832"ORT���'IV~��c�)N��D"O��x��P���̀�d�����"O:ݫǎ�'9S:�'J�.7�NA�"O���� ���
Y-M�X�+W"O4�7��s�R�Y�(c�)c"O$����+yE�;W��	�Li�"O�	�0�)`��#'��9�tի"O�E�� ͯD�Ys`�������&"OJh`@�"'��訧���6���"OvPP$d���`���`?+���"O �a�+{&TȒ������"OT���Ɩ"q}3���Y	�(��"OXź%� ���s�N;Vd� "O��� �<GP)kE�PPըiy"OB��⛜tcxm���0g��JR"O��`r鉗/��ՋZ�J`�� "O���c�?n9�zp\l����"O�hB7g�6&��{'�ճ �
�W"O����舃`(��@H� $�NՃ�"O���6�X:�,d�$��'��I�C"O���2�H���)��+2ݔ)�"O0p����`���b�Hu�B"O���%C�p�������n�4i	�"O���Zk����`(>?J`z�"O���Ӊ��u���U��%.�H�h����@d�4�B��nԔd�q��"��'�v�jŁ�>RT�����@X*�H�'�b�I�/RJ�r�ʄ�ހ
t��'�"�����/��
d�Q,z:^	8�'�pB�O�$[�ŀWBT�q���'�"P�!�����[�?��	h�'�Z�QD��6A��!�Qbذ<0�'q��ࢫX�#T�b!��K&�	��� �5I���.i�l�%���"��V"O���2�ɋ4qZp	d�χ|dj���"OV�����8;�2&�5~>����"OM��J�H��
/..^�a"O�A��F�Ik���@ߺU(x3"OQh"'Q
*����G��	�朊�"O$Y�LS$*G�4�G�G�\�,��"O\1���$4��ڲ	�G)F9h"O�T�%��6?RJŪ��>ZT�U"O�|ӑ��387�C���B���$"On@V�P�1�,��MQ��(�FJ�<��X����f�M<�2K�)I�<9b�&~ǔTk�C@0`�>�ȅ��}�<��]�v~�9I���1D���D�<I���<��u��O�i6�����_J�<ѵ�N1����L�J�ș��Hr�<��E�c=�����v��hЧ��O�<YS뎘oAZm
��ECfA�d�@I�<!tg^;m��m��Z$db�FO�<M�;���IH�Xp��FJ�<Q3+�7F.��C�U�������@�<���ވ:`����W��F�<CL�\n�0��q�
P��\�<	�b�'|h�H����>͒1!f]O�<A����x�d�o"P|��
I�<��_�9;�D���zL2�� ��G�<a��еBe�������)#R�@�<!�FώB�@D"R��4/�Z��U�<�7B#b�=IRϔ.u/D�&#^T�<��%F�D*��E����	��H�<�'�@�|0ITf7Ji�U�;T�T;�GA]�
��e�No�����5D��be�D5�N`����"n#�x�3D�����'�x4�P�t�B�A�2D�(�����8���U�����c�<\j!�d� �\�EŎ΁�d��D[!�d
𲁋���/�L�T�dV!�D�&|i�f�Ox�H�Ԉ�!�d�d�r2@#w�LHB�#!��<&��a�*�9H���
�B$�!�$��7(�H%Ƅ� ��}�'d���!��%gJ���G����d�$x5!�d� ���G�
�lz�P�a�"O��@ߘx᠐%
W�Z���q"OF�1R�
	(d���IA[��-#�"O.���F��ACǯ�S\<-"O:1�-	
!'*DQE�S��)2�"Of0�2�S�}�h�*q�D"&�$��"O\ K�f�z��q�!e�nA��"O$�  �B
���X�LΤ�+�"O�uYv�� T.�`�.�&WP��"O���B()D�]�3ۈ)�䊲�!��,����2�L���1�V�w3!�Ğ�A"L�yb�Z:}��z
�/!�dZ-9������c�z=��c�"OZ)�7-No�XE9�o��+����"O��)��Y����`'I>�����"Ob����>e�h��U(x6�
�"Oh��BR�eӎ�0��W�x��.�!��� �2����f]�l� ��P�!�Q�|�Hբ�jíY*Ua Sw�!��`ĸ��u��@k��#�C6�!��]�L�:T*AU�Kg�&�L��!�D=� Ȳf(P2[�d���%N!�� ,���-H�����ZcW<Ͳ�"O
<#p��&y�:1 �+:�a�"O,����4?�x���ڥ9DĈ0�"O$"2P�4�40�UG3r�X�cG"O\��t̉�k�ʜr��ѴN���k�"O�tQ$�O���y��ѣR^���"O�A�7%�!�I��L�1x��V"Ob�b�n�t0�%�޾g�r��"OR�{҅���S��C>蠁�"O�V�d�"y�	ʺi	�(;�J�<���Y������7(t� u�HP�<�$Ɂ�G�^�aO1o$��0ABo�<)$G�*TJ��ߊi �0��Vd�<�#��@`�=��Ц�(�MMZ�<�4(ׯF�J�S�ˉ$���r�g��<i5�[�_�����ʤ���<��ٜ����<x��cQ�~�<Y�ڢvt��S��[��ċ��C�<ٶ$�?-� x��K �>4НS��GC�<��ޅ���a��:��aK���u�<)ѪE�(E����6&1����^s�<9�M�{D�ш��~T8�E�U�<rÈ:x`�9�ǞWu��c�%]X�<�o�8�<�Y��-6�0��m�<��C�$
��ivK����� (T���2恧~MbAFM��bu���*D�����(aT�Y���J�\����,D����O�-4����e�+���y�f�r�E��ʣ;�L�CA#�yb 2/����Sd6��R- ��yRą*�$q�ƯZ/9:u��@��yrCE�&��x0�kY�4,X��p���y��*V�TCJ�`���@FZ��y���aG
��1'�.6`������y��b4iW-C�8?���UF�y��8RJ�a"�fz�@�mR��yB�V�,G�xW�#lu��$���y�K�$@�i�P)I	ke0;į_��y.΁ �0L�&!Sn3�`I7��y�кD�^�����=.�ǬS(�y� �:�|�$��#쉡F*�y"ǁ7X)l�3��	�!C|�"FON��yRWI��\bQ�/]h�3,N��y��H�s���@��M�b� ����yB���nm20���R��|�q�m��y��Ύ(0�E/E
wZ��J��<�y�E��Iؐm)����p���x���	�y�C�
+�bmC� �pt�ȣB��y� Μ.X"�۴��g~�8B�ʒ�y"K��\I�2�A�4�>M�%���y�.�%6�pT3F��'�V%P�C�y���v�"�ҰK���5yA���y"��7~��H�$��	���F��yR�[�6b86��t��0YP��.�y"�;B�L<ӄ���䦉��J��y�c���Ba3��S��@x�3���y�ǁ�U �ؚ@���@iyb� #�y"� U$���!�.Ҵ���_��yB$F+
�q �"9ԅYBJ���y2�
4]^R�  #�l��cBeN��y�&W��� I�v� ���M�y����bԘ�ʚi��,h��Ϡ�y��.,PM1SW��b2�S��y����!H�t����+�֝�����y
� ��ñ�S03M�5c��Ʈ�@T9�"O�0@#�+A*]A�M�#�t��"OH�/ .P�Ѓ�@���ڢ"O���E�M�c��q�4���#�"O0DbWj� /�Ra�"�����W"ODX�ֆU�A� ѩ��+5�8Q"O�-�o�5.�S�*�?�L�s�"O�bg��^��B�(B�xT�v"OP#lȁ-�Vm���Ʊp;��S"O>���;h�����%1۲�z�"O�ܳt�\�'Z��3���(�r�%"O��I�BW�v��� �՚V�\D�"O��0ӈO��r�r�DA'�C"O�ih��ݨ#l���f�#&�q"O���F�F2�rZ�D�x>���"Ot��s�ǣI���FD߽ Lҥ"Obt�䢗�?Ҏ��ej�z|d�A"OR2Oړ k�["	�xJ�8"O8� S�Ɓ<�:�n�#��)D"OF��c��JL�'� �!b�w"O&az���z&m[���*R��С"Ot�Q-��m������e&&8�V"O�y*Abǂr�xH� F�u%�8�"O8�d㝧���(�S�\�"�c�"O`v��d�D�U��t�|��"Oi��	�~0D�R`	��p��"O����a���U�Ո���H!�D/o�2��AIZ�!	��+��p1!�D@"_H��d���<�e�+� g!�D����%�"���lġ#l!�D%R_����A��g#��*���m5!�D��$�X�*g��Y-"8R%��.'�!��8`Nx�!�� x��2L4K�!�䉺c��h3Q�6+��Y�rmK�&�!��ن&!Z����U	A�L�����'=!�L&hP|[��àQ�ఁ`��z0!�d�G���Q�NC�nU�pb׫k!�$�<�x��蛃�@}(fh��.!�$��C�*��MH(4��3���	|!�[�T������D�a�����M�??_!�4ܴ](�K�4]���[�#��;[!�$�>
z	{�X2.�dY��on!�dPo�ʃ*�̾Y��-�jk!��Nwb�i��L	 5�`S/�f!�^�2��pR�L�_/�<9 	;O�!�ā6 Wؕ[�kZF|�O��!��ە�.��V�/9�\�(b�@�!�A#!�>�:`G�A�"�8��Ō3�!��
}����n΂O&���Bǟn!��D�G4l-���C e�iѳK�@}!�d�kT]�]
A�Z��0`��w�!�$����k���i�dqł(D�!��Px̱r����9��	�!��-7�`��e�2�J�3����!�X6ɨ�?m�i� B-2�!��φ%H�����5����� Q�!��Qn��-JԢ�S���g'P1p�!�$�qJ͠p��]���	�e
!�!���(���b#L :�*4���%}!�S��ճCl�V�C���G�!�V@��a!F !����dW#�qOH�p����q�� �
!20�`b�|2c�v��P,�8FIPC؉�y�n�'![�$�DC
"��8�-��y�-@+aV�3elI/"���0�y
� n��*�/H��mc�%P6Q�� �b"O~�iF�׻`'����T�>|L첶"O�`I���.>| ��!���\�Nq�"O��h1��D���A�JO�h���"O,$Ȳ����W�)8X��D"O^5Q���J�AMܫg�)
�"O4���'H�4 "�Ī3�z<I�"O�A���C� 50�hp�6X��"O�D�w���V�T`�
�l#�Ѓ�"OPػVJ�?b��c����R�"O49�#a͝>y*�z�	��3�ܙHG"OP|"4씦~a�ֈ� @"O20d�րl���(�a��A����"O�M�'�	=ͤ��e̝Yy��b"O���Df�[�,YQuN���Dq�"O^,Q��E��Z���&Z���"O@����y
��`�"OTP�ƣ�#���$�B�r�����"O�%c���rT^�*"�H�0R��t"O�D�7*���لCCI-t�"O�����(Jb��@$|�4��"O��ӡ^���#կ	\w�e[�"O��7Х/m�9�w�ӊ1���8�"O!��@Yv�^XjG�A�D�bH�"O��k��.qe�Q���:ua���`"O��1�R�ap�Ñ!B�.J63�"O�lj�H:N��x�FF7��@P�"O�:���U��	�A�O�(�>T��"O�'�Bf�5)�oܧ2w�IA"O~y#1%��r���� O�(@]��W"O��J���)�����NI(I�S"O�XS��=��p��7F��"OjY0�
���� Kwkb�д+7"O��	C��@����dL�5_<�9Q"O�8cB C�x�6U�J�q:�G"O�´EH*����i�	�^��"O$u(��=�x ��= _:u��"O����B�;���j> 8�"O 9j Gч{��<$h$FMa�e"O���C�a�N� ��L*se����"ON�����;ah�!��H�^be��"O�����bC��ʀ�-���7"O���ʱ_�䁛�B����4"O����%1�����A$c%�g"O��AgB_W�fQ�V�z���a�"O�i��
T��b�eݍ.8�9"O����	��R�CW	m,�"OD9k#��+�BIS2b@�x�
�"O��8��"-�9B3 G�3�ƹ*�"O<Z��S�>,��O��<�tx�"O�tS����`J���&o�`�"O0��e+=�t �m��!�x���"OI��*���q�F�%����"O°)W��A{|���D��\�7"OUS@��9Xw���ΑV�~�Y�"O�=�P�����MJ��Z�xQ""O�HʅC�8�jR쓼t��p""O�k�Av��XANNEȮ��"O",�'*N5ev<��,���\�G"O:y����:��U�G��i���1�"O,�P��Z�p��ݫ�#��2��Q"O�1!�f��_	��EI�:a�<(�"O�q�D^�C�����Е"O����Ɵ6}1H�#%�ܯsA���"O� 2�3��	�V���M."xq�"OB8f*OX�����>��A"OZ]S&&� wb]0gς6:�e�"O�hs��@�h}Zd/ǌ$����"Ohi;G*H!k�>�'�8R"��3�"O��)RH�1��Ȅ �9�0��"OT\��-)I:��ӧh�;��Q�%"O8�v�	pe�Cr�R�S�j�B"OΤ�P�کg@�cԥϥI����"OҠQoQ���h��6��̚�"O.]Aqf	I*���QAȐN�:d+�"OH��J8w�b��Ə]�L)�"O
������x�'nQ��X�%"O�4Rt��J�� �@F[��#�"O�� c��HC����ٰ��"O��b ƵX^\�Ja�<)���"O�)�b��2�m1B����G"O���B�L=^�R�Q��S���m�"O�u;���~�8lÃ��8��yBd"O�4I���1�n8����kNve��"O����%مa!܄�K�
6L̛�"OƤ��HŎG�B �R7�Q[s*O�jS��5�2s�@����A�'�cc�߭>pF��A�[�z����'��{1�ūrb���5��oA�x�'&�*5#��$����d����'��I	U�	�$`b5�O#I��) �'�.mk�"l�fQ����:B��3
�'���K��E b#���s,Y�4p�XK	�''�Zt(h�@y�+�!u�[�'��=��(�SJ�S�S�g�4h��'e|�Ct�/n��)�� \�Q��'��$�w$  >t����n�Ѹ�'!� 
_�G�B��2V6}�'g =QEdY	6
x8�e\�.4H
�'.�	{���=�@-x�H�%v,�K	�'6�L���7:��Paf杖u��'�������l�j��a�xͪ�'���$&����\�AF�-bqb�'�.8q@��.Lg���M�7&�F4��'��J5 ���{!�"�$�A�'�8Y#ǝu��$kR�8�,Z
�'h�Eٷ`�}s�M
e�0Ӷ��	�'�\Y��/T�B ʡ��vF(���'�Z��%��֭ ���n�� �'RX�22�ԉTh}	1k�`j��'����Z�>�4K��	^5z�b�'Vz����!Ax���ǯ\�^�z*�'5<����J�c���a	Mdwzȓ�'O�5ۅ��/g���"��\3�'��x�ӭ��Dx"E�1n���'�$8�1�	?�F�1��5��'�T������3�)1!�<��'^��;E�P4Q�=c��0x�X��'kظ(�ZW`ʜքE�+�tp�O¢=E�T+$b�L�rD�ӐdM�H�g�T��yR[��� ��Rk���u�ȓpڙ����t{���-�9MxA�ȓw�fPi���7>�j����ӵX"z���+S<0��U�Y�*xҲf��,��5`V�I�A��yF8����ܭOwpȅȓ.~�C��/%�Ԙֆ1z�����wb}�hڨw����+Z��ȓ*����`��@�i`�Q�$SL��S�? X�B%�(-��4A2#��P�"O6�٦.�+�d����Q��Q"O�	�dlZ����Oz*���"O��x4�P'A�2������P@"O^(��FSM�t��2��h��lS�"O뇃 .V����͉E��t�"O�P��j"6�>]qEL��}�"��V"O\ixc���^���
H�2D"O�X03B��بƮrjJ���"O�5Z���� �.�sEh0+�p
�"O^Db#�EM�.��"�гi&H@3�"O�EuB�=b���r&�K"X|��"O�R�^�I�}qQ�	V�l��"O�e8W��'!��U8����""Oz��U���:f$9i"��V���
"OJ�i���,�č��͖)��i��"Oh�`��' �@	av�Y�*l��A�"O.QY@��L��s�+A:���"OdP`�X��l�1�c±#(���"O�90��.gP����7O��0"O�1�H�0�Q�t��>�" �"O
��q��)T8�����+3��'"O>�%[�&���V�H��E8�"O���cș5�R�H4g�r�dx��"O�l���h��u3�FRzp�"O�� �B�M+�A�ReߏHY:X�"O�%:��͕f\b���dx� ��"O�52�J;x9�3!��-jX$"O>�KH_�`:�ա2�D�b< d5"O�}h�+�yd��*���,YȰq�"O� �ٕY[,���֔aM�\��"Otp��l�j�����G(����'D�TH��ؙw��9
��]�p��9��)D��H�υl�����o� �I�'D��{E��::��D�n��9����� D�����u���!g�V|���rd?D��)wmG!�tC%��n��pH�c?D��`f ��s{�؉�D9A�g�;D���WJ�H�<�uE�.m�(xPF/D�<�TC�gB�0�#�"W��R7� D��7�B�(����kI�%^�C�
2D�0��Ϛ�r
P��ň� �S�1D�j��՟ul�U��-΢<� ��G�#D���UG�>��z���}���q�f D� ��-I��%"P�5C9��Z�=D����E% hc�)��S�Z���&D�T �D�i�ZՀ��W[��IKA'%D�����Ua08���R�*��<�Qn.D��xË�;o���C@x��j+D��"�*�u�J<�1o�s C+D� 1�m�T��It��$��l9��6D��j%��8�@�؈E�lip"3D���" �@=�"��@���2D�[�J�-̮)�qh�!j)��*2�/D�T��ܲ���߁e%2��&�-D��;�ø* r��qk^|��*D���fc��B~N��&O޽ ��H7#&D�4�ԂA��f^�I��$�r D���udP(�'	��X��t���<D�8�dՔ4��1(���4C��C J9D��1��9@�P�ӰaX�Z�:76D�𓰈��#�b�*h�"MхN4D� ��,?<��� u�aR1>D�ԁp/Q��
��a�>$q�C�)� �*5��i<����Y#2Y*=J�"Oz�1���6�|y����3QVZic�"O�}�O�+Q��p4�RHs��"O�$	T�Y�阄��'�,Th4�"OxQ'��/tNt�򧖐S�nTɁ"O8��F$"qo���fF<L{��D"O�)uN�a*�;C��<wpv�0�"O��ҧ�={o�e+d�>R�^];�"O�G�SW~t�RF��Kрɡq"O8 �$�N3�)����F�)3"O~��Z�O���11d��Q�F���"O�`�@Dʙ�
��#N�v� "O���,�^iQ�lվif&�"O*ݛu�J46���r��-M��)�"OJ)p�t�MY�S��x�����y�E̎d��+ .όB�d�*נ�yoB�,a�q�$O+�(�ZW&�y�̊DG�	G��~�*ٓ�e�>�y��O :X�@��@�|�H���yr��&��z�'\�&7��S��F:�yr`�x�h5� ̐O�@�3�_2�ybO�F��M�c�	���F��y"��I+�USa� tL8a�lJ �yҎ��EL����Ѫf�@�tMC �yR���>p1p�ބ\���g�5�yR��U��H��%��^D���1�Z�y"�D�=�=��"�&+� <c�N�0�y��}�F)�(ΓX.b����yRo�1��82d-X$���q/��y��[�!��8���$�W��~�C��8Y��, �]*�3��v�C�I�cw���VgD="��'����C�I�T �5��@�&vu�7
��!�dB�	~ٞ@;�a�.�JI8���5	`B�I8�z���ђ1�F9°��(B�I2Zw 0Y���-L�1��*7B�	$tAk�6������j��C䉜���paL�'h�q�-E� ��C�	�#.����j� 6ŝ�f�nB䉭8lp���]�t!V)�'�i`FB䉔�`�"�±h@>	���;R��C�	]~��JDώ�/�6��`��S~�C䉾�tU3��mx"%�N�F��C䉧c	�� �H-b���#�Cͫ(I�C�	>U����F�����lʻ~��C�I�s�HJqA�w�ܼ!r�\-�8B�I�dO�)Pfӎ39�C�l�5#�B��0=%�Щ2ᔲ�D����	�"O ��8B���*��[�R����"O���f�t�ʽ�$΀;>�(�u"ORYhq�����2�
��"��X��"O��h%n_�V�,�◯�0u�^�h�"O*	[���	����&O�	Z\)�"O��ےkI4l��x3�Mʄ&ٲ��2"O�}#r��W�𘁡
��E�8耳"O���V�H�K�<�X�3�Rp"O���B�#"����F-�t�iE"O�0S��*5�
H� �Ӷ	oh@ѡ"O&]�mC�I���k��߰tO؜��"O��9�L�I��m`Q��&?���"O���f! 4+�f�H��ڸ���ó"O.�A"�T.�m�Ffr�l�+Q"Ov���.+08��D�#I��С"O�92nH��I 6���M���1"O� lD9�n-Rc*�3z|�D"O��9��>&~��)I�[Nt�B"ODd�e�W�f]D�����3OX�I�"O�@T� {�Y��k2_*J��'"O��au��b��� ��l�r�"O�]����'����K�6��x��"OJuP��1r�b��Cb!g>���"OzP�Ư� }3(:6k�u6Qh`"O����Ke����Ծ6l��"O�Xc1�ɟv��h�G�7���'"O8p�A*�`�x�'K�7�6y(R"O�U���$R�~���ɑpt�#�"O	�GE�~nPp�Ҩ]e����"O}���[��6�(wh�8cxdk�"OhA�գ9NUf!�#�V���|��"O<��C7l%3�'�|�0)�G"Ox���Dޥ5/�s�)��X��"Ot`SE+�Eg���i,?��zP"O��3��/f
|R�AE�|�t5Sg"O�| a�ΑJ�p`���"�(�14"OB�K�Oݳ7.ؓC��Z�B�)�"O4�C0(h�N(���#f�D��`"O�l(�"��6pi���oʈ���"O2���K	\��4�A�F)@�^ ��"O&�Q�C�8c0�T�0���jt"O���6$(�|���2fIv\+7"O|���ѹ+jԔYp���$~�p�"O�]i�"��g�m�f�&*l��"O`��SE@D�{V&��o&iX&"Ol�G�P��8\��&�0��K�b$D��K��Y%��ӳ�WJ/JJe D����GM�q��0⥄��GQx��K?D��ڕEE�'�8ҕ�(�t�)6A=D�`y�GQ \�Hʀi���X�Q�g8D��8�Ȳ�|�홌~�&����5D��I���&>a�e!6��h$�?D���aI'.hx�s��$�*���!D�D���ސGG�Up���2���A��3D� ��L��[�6iWG�:^�r��?D��1�GF�O��i�g$�oĪT��#D���M��tf�m,�8�D�>D�4a��K�3��`;�ٶ�J����;D�����4<���r-��@�"K��9D�P`�/S:Pu�uC�AōP�
F�$D�paH�&�ft9a問D��Ѫ��#D���c�&P�Xڒ�ԜI�6�@/D����/+fM�58�%S�MJ��cO(D�4�A��b��Ѐ���S&)D�� ��1QyHhda�1Q�����&D�T����W��ǯŧ+���W$D��p��P�u~H�z�!����(APj<D�t1��^Y|h\iץPQ ����o8D��`�_�yĉ�aiۍP���%�1D�� -�~C��;�'�7� ��*D�(�g+�*���A����J�*D��e��.< �$��q/� ��&D�"�NF�/�LXc�j�=+�f0B��(D�l����\�8���� (�YO'D����y�5K��>%��(
�j7D�P3���ZF��hB�
J�(P�	6D�PA�*]3q��dH�^L�ೳ�4D��;���"�P)0�?H�D��8D�lpT��/!ī�ׅJ����6D�4	T��
��U@�&�:=�n`��l5D�� �` b�KF�=�f���x�U��"O��3�	���4�C��	b�BU
t"O�x�"7e�tN�o�B0"O��#���d".j�����f"OJ�3���7<Wf��oR��t"OV�j��)x@`X��A���L@�"O���OɌERF����D6Hْ1�4"O�|��Bٴvl�����/�pq�W"O��h�&�5g�zx�n�;*��M�Q"O�A�̑�|ZBip�l�>���V"O* �b̯3�vq�T��,Q��S"O6�����6+<�� R��l=pDۂ"O�e
��<�~����O�H.4��"O�42(H<,.�k��#Ct��#"Odr��[U��	U��N^��B�"O�ɣ���K��\B-�&�b���"O�)�&$��}��i �&Z%p����A"Op`S�!^�Q���Eh��� D8�"O��K��G�$LC�&ה}����w"O�QCɟ)�$�[eZ�~��P�"O\1xI�<� �j��B�vp"$"O��a�-���L��%M;|�C@"Ol���#�?�`R%N�E��Թ�"OH�їoQ�k_�)P�%�a���{B"ODY�u�E�
�&�*�΂:,ई��*OH�r0����|)�&ٹx��K.D� X3 ؐF�iK j�7Wۮ��a�'D��P5)ש
��Y���Y�q4$8�'D��tꛋt�̉��؝340���/D�h�aF�3D��00���N�<��D,D��0�F�Q������`�*e8��>D�̹�{�T�i3�۽>��(�Wk8D�`�`É�W�KV_�v����)D�T��iZ�L��Ȱ���� #G%D��� �	E��r�WS��'@#D��93`?r8*�;��T')Q�0�?D�(Y�O�4|'v,��됴-j����)8D���cچ&�ؑi$�Й@�~���i9D�xbJP� 8CV��	J��$	7D�ȃ�E�<��0K�
) a5D�j�a�N�x"0�̠B��(D�r�
�#�~�h�+�-cc��K� D�p�ٸe
B�[%`.|�`���+ D���@�P�
2RQ��j�i�(t"qJ(D�\:PjT.=�֡��eH����#D�(�Dą���!�t��):`/D�d�1ƒ=��T2�����(�ק,D�Tj��O�& �*C����X�(D��3j�&�Ɯa7h99�f%D� 0�e� s�&�Q+R�?~�AB1�#D�����U�2��QF�,I�tXɀ�6D�xr�I/ �rd��!¿"���E?D���	\�k����3N��R#��t�;D�����:V�6��g��	~�c6D������{��AҢ�
;%�����'D��9�B�63[h���N�@���5K#D���V�ȃ �>L�GDM?��YY¢?D�l!wjʮ"��l�n
�f0��b=D�X�%nO.�@� ��{C&\��!&D�����]�*d.�Se��4%+@��1D�,!QA�V�����3��)D�@{����
z!���N"	86<D���P�=Q8I(����6�°��h8D�\Q1�����2"LΝ	2�9D�� �,�$�2%� Z�ԒS��h�q"O��a+!2�fDI����'"O>�92��9n[>u Pa�0��|e"O�E�"ŗw�E��S�B��P�"O��B(��`��܈�#}�"�ʗ���p��sɛ�'J�_?���e�"CŚ��@���`��7�+[Tv)R���?�w�<$+F��*r�ڹ��
bo*@3\���l\$%�N59aΥ\&D���Q��HOֵ�e(q�|�S�V4:r������|� N��QBB(��at��ǗN�'�pT ���?9@��D�i� �
���!��}��.*Cm[���O��"~j�4c��p��a���t[A�����ˉ�d.��O��6m���oZ0j���3Ѡ��\f@����A�H֞���S��X��iQ��']B�O��`y��'�·i�H9$�̢U!� �5! ���x+ѫ�u��[G�XA�h��,"ɺ�H�O@�S�?Ѯ17�
��$˵����td^�ﶈl1p�؈�@'+�f�k"�+nr�s����ޙ���Q dTFr�D�4�1��iy�8����?I�i��s�$e��I�/5����Ũ��pȻd�ON��,�Of��rY�.H(Px�I�)Hҍ���O6�O��lZ��H���]���x�0�Vp�$8�'
@#L5���?A$,^�_��p@���?���?������hӄ�I��S�6�n�E�/D����F�3_��r̚�nԜP'��_���4��@�)�/y�q cAU����`�ĝ`�8yD�:x��C_-��'"�����ޅs�2h��ސQi��9��C�\��II�\��Of�&���	Ο��'�<�R*Y==���'\�uے�؍�$=�'&�.��A�{�Ɉ��8<�
�b�qӠXo�r�	g�X��+���O�0��5jH�$����3nb�H&$	ß��	���	`�� �I��$����Q���E�#�ݺ�e�iF��K�ˠu��U
�rX:�uB�&#���	�k4a�2]�A�\������Av�U����-f�d̹�o=��yPg]�(˰#�}�oʲ�?��4J�(P�@�V{�\c��ȪI�$���O���*�d7��R8N��]zcaIf�~�aǙ*�qO�tK�)�IYŪ �6I��,� ���y�]����M����?���M0D��i���'��;�4��� (O�̥:a�2A�X�n[�'p%@(�fD�v' f�q�B��8D�̧%ޠ��4O/��(�4É���Dz�K
?���4H�	H��S��֎5���Ӹ&Y��ھ_�8�3,V?J�#=Abl\ܟl�I��M�����T~1��@��a��ǟ9#�6�)Vj�O�"~�	��̢CnQ�>�(W�W2$8`�'�7�\���lڊDt�(��L�[Qn�rdE�*B�����jZ�ʒjW���	r��K�]�R�'�Fń5�U�ө�I D`��Tn�X@�iz�R5Kʑ4y�)Cė���|��'�5֧�J��5a"FS�G�n���h-�M�Co9*����א)��u8�B5��>�X�cm@)Ë�k��i��-�&uF�7-�� >��'����"|n0��%`Pl�Yl�	[�Iق��P��jX�D��*�>8o���*R/��Ps�:ʓNT�V�'r�x7��[;�$���C�D[�D���љ>�J=$���퉟t�jp   �   \   Ĵ���	��Z[vI
)ʜ�cd�<��i*<ac�ʄ��i�)m�@x�a�P�mڙX"��xP�MPy�p$eb����4\ ���b��p��IhPY㒩D[���1�N��z\���SV��+<�ɋS���{��i��,1Q�\�n���۰�Թ�0��O���A����M�]��P�#6B��A\�0q���%y1��̅g̐��]Jʰ�P�T��;��|9�B"ΓN:I�A��؉ɀ�Y`����nM"v���O�@��f"z��'j�Ea�DN��~BF�:��\S$�5���#�΄ �~�"ș�y����Q�<�Bf�,|F��P!$�<�L�BPD��<9`6�&r#<���N8b!Yf��oP�AbJP=5 ���W቗>
�	.� �1!	�6�x٢�� �'�nEx2GR�=� :���Z�prHͬMj�oڿA������I�5 ��P��`�x9��KrCr��0K:�	�\D�l�e���Kצ�>jslY� 	�?(��bl�<Ib)<�FI��) HΟzEV�y��*;��L@6*Ԯ�x٥�	/Db�d eh6��#TJ�A�	�Ř'�Fxr�V�ɲ~6M)L�r��r3勺o�
��`m����x�M��\y��R�=�-� N�y%�����O*Q�ṟ��pN�$}�b>JTe�'e�0�`]��*|h\��@�P8g�4`{��Iq		��wEp�S8�:m
�зϑ�4�n�������s5#ݏq��'�04%�݉��'�H9�6�����'ڼ)���S?�!�dދ	 �  ���"O���t)!I<(	�@P�N�N�Xa"OH1B�ks�r���-$THpH��"O�X("͇�%��$�Ɓ]tބ� "O���$B�D��O#�>���"O�B�O�;���9ǌ�<]�Lk�"O�<(Ѩ��\Sl��6�L�7y���`"ONH!E�]����Y�끹���!"O���M�
-��
Y�md����"Ocf	%X$�ʦJ�6l<P��"Or�;%�ݔR�y��n�	�`"O�GEC�.��V(H4SV$<I�"Oԍ��(��ialT
QS�q�t"O�5`C��0�< k̙P���C"O|QX����z|����O��9w"O�Ԣp�L�G���KƤ!K�4�"OZM �'�{1`��6#�l�j"O�m)DO�к ɍ�dc�Q:c"O�YҒ�E    1  u  �    Y!  �'  -+   Ĵ���	����Zv�Ll\�0R�PΓ����I5&�H����O�����a�B䉢]dx�󠩑9b��)ؠO7)�>��F8�:ݳ�i����sboѥR{84�+�0q�N��!M==�N�Jtg���X	B<�,�(ƧNR�jАeL�O��t"#O��hh�d��)S�l���I*(�|IhG�KF�0P�O�A�l���H�)�0�q�[:e�gʉ5,,rP����%U8����'�2�'lR�b��I#'�0�P��$!����@�S2�x��7�B9;��[ lu��2�)R=#��3�&#δ@ �~F&e��`��<q����M[�������E`���(Oj)��L>�N��BQ�*�X:bU�8#e*�Ob���O�㟌�'9S�P�ȅ���	�jJ4�ȓBK�hʣ���rx�`�)�%P�mZ��HO���O�ʓ~a�� ���m�0A�Q:��iZu�k�`���?A���?�"���d�OP��b6b8@��ֳ����ʣ6x�;%���j5)���)v�|��
˓>T^i��`�@�S��	r���`V�
�0�Rr,]8{d94�'�a"��B5�����,���r��:�ժ��i!���&�禙 ��5�1�����Z��/D�thug��2t�#S�EK��0�>�a�i<"Q�|�v�G���	�O��S�.���͊*a�օ�e�<��6����O���Yν�CE��%n��ԟ��8Q ��#��y��c̜ct�LH��	�^P��ye
E `ִmy�!�D���̵"9�D�R�G$��Ѣ�*�hO:e1s�'cB��ҊU��<��CF�7�����<R���|��� wщk5h��`�S�P��Y4I3�O�l�'���r`̶n<ցyAV�k ��O��a;O����O&�' ��r���?�$M�L��Z3bӿ;�2�8p��!"��h]�db�T>c���p�**�yj��\��T�SJ�O�ñ�)�J����}ܼ�f�HD���je��	��S�O��y�s�H'�L#lF쎉��"O��jS�4Ӹ��Us�*��b�	��ȟ�* Ǟx����&��6�p ��"`��h�Ó
:*a}�o�o�jH�F�2ւ�y�D���yW]@t��&Q[�":�yr�̽N.���L�,ov�j�L���yRô!�����0xdе3�!S�<i�'$R�$x�5��l�( �N�n�<����!��%9S���c�*�/i	JC�ɵ2�Y�o�0��%q�	^7+��B�ɗx�8制�/Vu��F���#uvB�*��j��Ł~�ʕ�h�'q.B�Ɋ�^� l�*¢iYWɇ�DB�	eI �
"��T��I����@¦B�I���U�)	+^m��pT��#a>�C�*L��͢�H�>Kn�ٱA�D6��C�ɹ>��T(EJl�3}/�C��1\�FM�@/C�g8�)V�V�j$@C�I�!o�\�`S:^�X虃/5k�bB�I�EM��q�߅z@X���G�?'�C�ɽu,�)[3חnU$t�"�/M	fB��AP4��+��9�ܫ&.�)�,B�m6�]��H�\.N�+$�l� B�	uT`��Z�2�uS3��ZS�B�<�����`�Rb���Gb��
�'�6�8$/U�$���s��:>2u��'�NL
u��fS���Ҩ\1HӲ��	�'���@7o�9�\�8"i�3���1�' \$Q��<;�1��K�&�^��	�'
������(3��D��ǟ[sE��'w���H�N�0�1�̃R�"=1�'�<�#+5kv�۠oݺI�9��'�*I�t+/H��x �M6��H2�'nz1E�Θ�L��c �W8�c	�'ɮ��MW�l1T.ߐY*����'�P�����d,�͂g��.Wf4��	�'ά��Sǚ=C9X	��J]>W=6�r	�'㈘���P�x���	W�,� 
�'�t�cLM�p`Y��մS�tĲ��� b�J��ƾ-��k'���v�BH��"O���i��4�2dաQ�@�
a"O~��pD��%��tӡI�%
$!��"Oby�sς?���9F��#҈�"O�iҁ��0z5� �O�`:�i�"Op���Z��)����+*"�P9�"O�us�[F����p\��IJ�"OJdq���*/i&}SBL/���W"OnD*��	9<�5�v#E�C""��0"O*��pK\��䰳�
T$h�0"O���j��r"��CWc�� PF"O��ca�[�YK6ҥH�}�x��"O2]�S���M�nU0O�~}$ `"Ou;G�L"w���{���VN���"Oj���Ԣb����q�V��"Oh@�5d�m������B�6�8�A"O��i�/�HR�4�� �&�݈�"OZ0P��K���qyv�R�@���+V"O<��`E$Y�u��Jxi�"O�t�s��X[��Y�&��� ��"O�P����'(��U��K���8�"OBQj��/\��pԄ193YH�"O�Q������W�6�te۵"O��G�5��`*g��3�ؕC�"O"�R`��">R�٧��_���"O�|1fƥxƲh���K�.��܉$"O�CRN���L�D`�3L��aW"Oj����L�d�����]8;���a"O�pP�\�a�r���O��!���&"OT�6��$v�0�(!mѬBb("O����*�:����[�����"Od��#��4Q���7b�} ��"O�M���s�����g��e+"O�A7�C�@�%�qI��z�%�"O��p�e��2��JC�R����"O
�Ta M��٥�ٽC��4b�"O���t��z������_�Be���"OPx���^ 5���%@ւ-]���"O�ɢA������H��=A48i�"O����M(0��$CP��Yr`�w"OZ��g���V��H8Liڵ�"O� ��	,p5X���E�t �9 �"O�0�c���ܘv��'9a���"O�` 	�� w���5J�:q
�"O�8��#�5�T��C�u�bH�"O���agɈa����.
I�f�;R"Ot)����^t�<�lބaL)��"O�M�b��[�bUꡪ	f4h�"Oh�)�7!�6�*�L. A1�"O���@KΞ�Pm�f!P�z�DX�"O�D�M��C7,��p�Nꄘ�b"Oh�K�@V 9���;3*��~(`�"Ox��7�B�K��@�/�dcn�$"Oδ!R�PP<AB��v:�1"O(��M�H�:��c�]-^>��u"O�1S�I#t���u�τ	K���`"O�̹�ڀ쐝���1 ��x+"O������{��}��n�_�<�rE"O�����"O?���eM���0Z�"Oh����A�҈e a��K�|H"O�â.ȁY�,`�P�&MZ�j6"O
�BiƮ\d�!��I�W�\���"O@��� ǰ(F-��Ҹ�j<3�"OzB/C�d�dZ�6J�"O� q����}���Ud�=n�P"Of@��Å�U`"i.gdb�C�"OҘҁ�K9&@��soD�dZ�z"O
 �UNW(a�B���YT&��"O���v�P�,P��1"��� ���&"Oj!a4"v���$�ڒ�0aa�"O^x�J������a�B5X��A�"OD�3���{���c��[�8� ��"O��BE�Ԍg&H	�V��g��Y q"O��(�%�:Me�C4oU]�^�w"OX15������-�k�蘳"O*�SDd�ZH�����Є��g"O
i�CN�R�ؐ�bB�l�~a��"O�ؚP+U�m��A��h���s"O��`mU�4��9@6�* 10� �"O�a@w"SP}�u��k��#L۲"O��q ��4mQP���Q �m"O���c�ϬLoΥ� [�sj��"O�E���֫>���h��Ø�B�Ҧ"O�	zs��!6�PS&ٟD1t��v"O�i�����%U�z)`t��"O��y�g�}�:�u%��y .��c"O�}k�IU�H8�x�≽�"�"O�af��!Zȁ�O��{�(A�"Ot@�E�ҿ9�B- Q�.��z�"O8�BЌ	B0:H�"�=(�l��"OB5�����H#�(q�"O��pJ���`�l\a�d��yBD��>�R'�׮)H�����y��U+1lr�3c��Y4}*�K��y*��a� � ��nI�%��y��^%X�aC�ń&�NT������yb��=O�]T&Q�%�|��@i���y"�Hf��s�]�,�l:3@�5�y2��	2r��I�,/!5�Y��J�(�yB�_�P��R�l�&V��+�E�y�n��L�*}ZV↸`�H�z�k[�y�@�-N

���!3h	�#H�y�
�p�V�C 	<0��Ń��yB��&wy�<�e�q��yDm�&�yҋ�9+3|�����7K�y���&�yV�/" 2u��n��r�Ȩ�y�c0D��!��)R���p�� �y�A�a�`u��OX�0(.�(�@L��y�+��Z;��qB����B+��yB��d�nܓ�鏢oҼ �I�.�yb	Y*�C� �bH�M�r����yr'Z&jK�#T��ض*BH ��ȓ9�8pq� �7��)����\����3��X�HT�q��y��&֥�ȓrц�+�k�6!�&�Q2(5M�E�ʓsl��Ks[0��J���hV<C�Ia�8HK��ȯ�	��k�j�C��fZ��Ћ��P��1A0.�< �C�I�]�`ȵBɨ-I,l2���00�C�	� �RlE!^x��"��&��C�I"] �R!�I<S���ɀF�X�bB�7J� �D�����	4�>X�B�> q���"�Ӏ]�� ���:DB�ɗ&B~ykf�'}���@/^�O�C�ɘU�j��wL�.?�,@��zXć�dҲl��C8ˮ]��R;U����9\��4Ô�k�9:��6>�=�ȓ�h�J�)ҞG�!R�a,Y�8��S�? �I[aI | �  �
�����"Oҵ2�1�0x3�^/.��z@"O&����I�3P�y��H �q�P"O4�j�m�+DI~,+PL�*4?^-zD"O�a1���c�y��, ���c�"Ol���P�X���s`,�1X�P��"O*	w+A��j�Ag!�FOV�;�"OZ)�E�{����bၰN� ��q"Oⴢ��Gfz���JFiP���"O�X�v`�+$x^�����4)WN�U"Ojy���sG�i��جtL�m�"O��B�ʫ3�1Jp�z���U"O�L�p�#���bD,�:��X#"O��R@B�q�<Q��� ��T@"O�ar0�N�*�y���u�ؐ�S"O`Ļa��>t�,��/ )F*f%	""O�@�`��Y��{�nC�](x�X'"OP����'SVX#���\F�$�"Od!(�c068��׈�B��Z�"O"5���W"!����Ө	rB�\�"O�� &��Cr*T���̂ܬ]�V"O<���K�<�~�;� 1#�� �"Oz�+T�s�<��U9��|�"O��`�c�/]��ʑN�3�`��"O���mP�K��ͺu�O!��,0�"OryT�\�4`2Ӡ��,��y�"OP���-
��<�"�"m"B�J!"O4x�C&�Z�d�k" �	�e�"O:�Y��-2l`�u�W�E�*�"O����n� �И��F��"�.4��"O����#ԙW�Dx)УT�~��$@�"OP� ���o��VFy��A���%/:h�$|X� �SŇ���I��
/�:}���%D�L�	G�>�Ф��gѷT�!"�)D���1�!�����ΒVz��)��1D�,�� W�B�+�ט� ��.D�3c���ga�iy!�ũ/����H2D��u�;x��c��;N�6�[I"D�{���vԀ�4˄��P$ 7�>D�����H��� *F�zD< E=D�a3l(Y�����Ŗ H�q��&D����猅+Т�!0'�0#8� D�DQ��ZSFJ�1��0KP(0!֧<D���/@(ȵd�����Ԡ.D��� hM�L%�)����	^���@�m9D�Dh�M:0��Ӏ&ɵa����r�7D�0&)�X�$3e�=U~*��!D��(p��yMٸ�T  �6<��2D����	�G�P���)!�,TC�//D���
ʸ1���I���.6��u�'.D�舠bT#'����qV+.ܕ3f$.D���@�0p��J0NS�i߲�1q�,D��؁�]�Z[���� &*�YI7m)D��k��'A�^�z�*a��)7�&D��,N|�>E�t��brEK�7D��3�F��c�>)���²B`�PJ6D��{�ďdP���B�2�m�" D��eX,2�"��1cUz���=D��4'I):,�p#�Ҫ-���m<D���cD�*r*Б��쎞p����b5D����Ό^���4��^)��$�4D� K�FRx��Tn��mg����1D��E�)Ǯ��W��|��R�0D��2W*�V��@Ă�;VyBć;D�� �@ӕ/�i�XY@��D���Ż""OЅP�.Y5I�4�S�ٖu}��1v"O:5�� B�)�x�ycO4"q�Y��"OJ�g�=i+��"w��8~����"O�$��ƕ,Ag��&�<QBT�C"O�� sj^A9A�Q)J �� "Ot�r��OrB�#u��8C6n�7"ON� �L̫]�2\��
�;.e��"O2U��Uy�	KD��C�=�"O �zp�Q`0.ECr�G�A��Y!"O`�u�5�F91�� b���"O���+X�P����Ǐ|�>c�"O2Q��^��fH�vn�>Xi�p"O��ٗ����|�L�]#R��$"O��W@?&(�=x�阄!����"O�šA��E֬z��]W�=�C"Oذ�_Y��*S��2��Y3"O�Ńd@
 �|��B��� "O~ɲ�m�r�� ����tS�B"O�yy�+�����u:d� "O� j���}i{4�L�Q"x:�"O0���'Cԁ䣎= ��� $"O�L1�Ƙ/�pAH-ܒj��Pڄ"O�s g d��؂���Ip"O��аƕ:t� ��Y)I���[@"OB�Z�$Y&C�(ᒀ��	�d���"O�SA�}�H�S6�	Y�*���"O�� �0eZ�K�(��~�)�P"OV�ziT�c��P�����\�B"O�e)�e�\4���R"9R��"OJp��Ƙ''�D��CD�:U%�B3"Op�4)I޴!�1.^�8��#�"OF!�4����좦�����
"O��� ��`"$���A֏ꈑ�"O�x����<P��Ԙ���L�����"O��{7΍"D�Y4��e��u�"O����#��p��y�S$WP*�"O�E)oնI��x�P��/Jڑ�S"OZ��dV�4\*�3'¡P/��Ɇ"O�%�֢O(Ap�PU� K��P�"O�+0AW�yL��B$�by`Q"O܅J�i��U�-S6�I�\�4��"O�UQ"(�
-cAݑA�L�"OP蔁]rJ�	3��U)*�r$!w"OLIR���8DX��
JƌP"O
�qP�V���P�q��>��"Ox)	C��2��y'd˾} �bS��O��(O�'<��1)�kq(9d'Ze��ȓ|a���ՊQ�o��ER� 	F,��)���T.Z�e;��S�&JR���;D�H��C���$Kѯ�.t�TF�������gTuiЁ��fn�@`3`�2!��C�I�eX���������	βB�5�jEJ��G�<��B6�A�7��B�	�jT�`1P�*C�@�3�ɀZibB�I9b����P �:S�*�R�.	�~VFB�IFR`嚆e��1����!�T*B�Ipybp�W�ͥ8�����GE��0C���>hK�*��]�BT�����>�^C�	��x�!D�f�xD闆�e�@C�	(#��rc�ݮ6�f��
�brC�I�D�����8!L8P� �!�C�IB�^M���_8oN�#�"[�2�C��# V8x���<3�O���B�)� ��as%B�[�0�Qƈ
F���D"O���&B�$�8����F�Y`��"O�H�c4 h�`�� �[Hh��"OBP��H�*���Z��E:=�v���"O��GE���<,8���,K�֍G"O,0��M7�6yP��*+f� T"O�!��*�HxH�s�, _��ʤ"Od$��,�v��H�cC+t&���"O�}�cÎ�Azd��� 	�"$ �"O^u�4?V�t	!ɟv�K��yR���n�0"�Mu��ۼ�y�/�}�d:ˁKp#�lƉ�y��6^��(��F.��8�֣�#�y" ɁY��dw Z�)9ix�IŔ�y��	��L�c2�H%�b̹��y�+�6��i2C��8�|a���yBkS����ƙi]��xb#޲�yҠ�%k�T��)� b�F��Ĩ@��y"�C�.�E��R Y����s���y�)M�V�~�ʗH��=4��A��yB�DUH$M�	�>ߖ���+�#�y2��%K��D	�\�.aa�B�W �y���8c��ɩq�0}yR(���:�yb�Â5��dC��X!J�&�x�����y�ͧ$�rA�"�K0C|zԓAh��y2�X�6����G�N����ዦ�y�IڲR�P��]s.��P�ʗ�yr��r��Uy$�� 4�Y�T�S �y"gؗЈ�1,Ǖ�4��#��0�yD	��f�qw��$z	��C�?�yR��kcf�a���a�`xæ�-�yB�[�^��P�
\���3S�J�y�aس�����+6�8�f[��y�I��N���CU��|���3����yZ���@� ���$�1ٲy��u@Ò���7C�2R|�� ��RJJX�6�%hh�(�gN�"XvI�ȓ4�j1� �eU�"סЈ� =�ȓV\�5�±?GnM�'�N��̽�ȓ	��m�q�!O�x���g��E��h��_��{d�0"��0F`�:p�ȓ^%y�\�.(���5N>>q�ȓ�2�I7k3]?���/ֈ�e�ȓW����a��1֖� ���l �Q��x �}C`��V���� |g���ȓ{��d��0��B�K6| ��j��#�:Gi�{���fnP�ȓ2�u���آ����"��N$ḃȓ`�r!!��:=�� ��0wŇ�-6��Ig��)��%"�׊bޔd��-p09q,ΞL_�9�q��;D�D�ȓZ����v�X1=����磓� �ņ�^���Ѫ#a�4�#��)����=Լ����,a[v`�S��cb@x�ȓI�H�[3k��e_����#�T���ȓE l$x�$s� *p�١j&l��C>��� ƞ$������8gp 1�ȓ`�*9F�4�����A5Z��t�ȓ���)��*=�@�6����܇ȓ&���`lY([M���� '�����@j�1P	ܶ5*��E���#,���jِ�D��H���� v�xi�ȓl?��	���K���4�C<e���������I.3n�) �@<1�v ��S�? ��S�kF� ����#e�"���9�"O* ���@�E�\8wB��A�T�a"O�H#ч�Cn���̒t�2)
�"O���%(�J�9R�͎)_��h�"O|M"�oT2� �Z��ܙ$O�)�"O�q3�)�97�^uI�Oȍi9B�""O�|I��!��$ ��%9�t�q"ON�����8XN2����!o���yb"O��xqL1d��+���\�l��"ON��0�ڇ!$Z�:b+�;&��#!"Ob�S�ާp/���TsE���"O�<a�%ޝoZ���.� 8n�h�"O.d�t�To�8�Q3Q:h��"O�E�gJ�� �Z�GB)P8��"Or�9"���ZK�%�C&Ug,���"O�J��"#�.U��%�+���"O�!{��ւ"<^ܫ�*98|��ʇ"Or���
��Q8��	��Xt!W"Oĭ�vl�}�qXe�:��t"Ore#�I�9Cڼjp�J�P�.��c"O8��ώCq�ԣ�E����@"O^5�BÚ�_/����X%���a�"O�qNݦv6�@a4��v���"OࠈW J�T � �1S"��"O�[̊1\(���4`$p���"Oru�v�]5MEP�MN6()�"O��q��(;L�Ƀ�ٜ#�0�A4"O�<��n��JB��"��U�a:�mb "O�B�)��C�돪-�)�"O"���N�!�^���l��sN �"O�Y���R<Z����"�_4&p�ha"O�1P䙲6g4u*jm��Y�"O�I9��U=���i����)�f"O��P�W�x��+�Z@��"O��x�n�+<f�@�c@�Ch$��"O�s1+ՏhL8H5BD9M��@v"O�%���  �P   T
  9  �  S   �(  �1  �7  +>  �D  �J  Q  HW  �]  �c  'j  jp  �v  �|  Z�   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl� Kp8O9���'�t��oŶL��5��m�-qbK�qU��� ��)U��ԑ�C�4Q�H ��Fa�U�@	�?!�I�?]���ʙN>~x�*�32���D�(����j� �5�@L��@u)�F6�]� �������Lre��r����%��Jް�
�"Z;X�P%%Ɉ�?Q┕d�\Hh�n
�*S�f�ɐ'!��'�"�'M��S*�4�t�7~�Òǎ&L���'0V6�J��v��?�U�ڿ�����?���L/O����t��&Y���QU�?��F��Iϟ��������,?�'ǚl�t�ؙ]qx,��#�dz�z�'��l�5"	�f��$�¡�2��ҭO`�U�Il?ѓ� ?r��'rJ�ZՋ�/�"%!3��8|)�	矐�	֟��	럄��矠�O����7=z�T���H����D	I�M2��h�R�m���M�w�i)��i��|l�M�q�iyr�O�}^���b@?<�v�I�K�;md�"=)�I�O��qӅF�QdYHcn�:���cs�\7Q�9�SB��6����i�(7M�Ԧ����|�p�/�i�fB����}��X�ݟP��@�P� �3��˷(ұK&m�zıQ*¼�M��i�7�B��1�m�,0X����a,zo8i�t�%ژ8��Ř��m��4��vi�m6���G�����{ÇY�/�1�v��7iؾ9�瞁Lb����L�n��X��#ʑQ��7M�Ҧ۴\�M�Fg�(	�4`ҤE�TӬt���U�AE�u
�Ũ};�8��0L���C�6N����o�G��`F��(?�d�	a2�@%��#�:|�� S�=���$#�	����Ʉ#"m��4�?���� �	:V#����  |(������?����?A�����kD'h���x��@M(V���fe��1�R�Իr�j �g(��0�'�Aj��H��05�� ]�j6��/#{"uxk�&J����1��jUaxR��;�?�����W	e>4�V"̓0뾴б��GKb�'1���#R�P\�wi)?<eX���E,���Vܟ�KM��D�P�B�yv�4��OV� s`�%§�y�ĉsK���NnDl�9E�-�y%L
i� �
�jj����u	Ā�y�g�v�ҭ�U嘰PI��{UK���yr`B)$����1�f�;Vk�y2�!����J�K��J�cԔ�yg
.*�H�7 M��R�(�ü�?U�T{�������tK?�8!���T��&�s�)D�@J7�Y�K	X� A�P*H�
�0�'D�����ۍL����@�M$)���bp	;D�@� `�Et��ّ�Mu%�����.D��H�ն�٩��-Y&f�k�o+D�l�S�]3)8X(x&�>K�*C䇳<�VF{8���Ü1i�%SV��..���E%D�\������J@j���b��#D�HӐ�3Ӥ R���)��] p�"D��q��C�?�@�v�&;�Ɣ �?D�[fcƚ_:ll���M�-�XiQ -:<Ov`�uEMצ��'� �F�ǕqK�,�cޡO@�e����d�O<��O�1H��	l X��.�S�|��I�u��$	�NC�d�RX�#W�;����$ �@n(�"��0)�Bm����O%CpB�1�}	s�#���"�'04����L��Flk� �D���h���iX	�(��%���?!���iU(�v��rE�~@����F�����O���#�&K���c�B0t���Iz�I0W�Q�!�1�s���;M�`��K�&:IƬ ��9D�JŇ�l(<	�����╘�A�7lZNȅȓk��u���N�C�|� >n��\��7=N`��S=i'p��1b��q��ȓ]Bp|�%�Nx0Q�.ڶso䤄�>
��k�m�4K����G��o��Ţ۴��k������?����?9.O�9�T��3EG`��U�'�Y�"fԣvh�R��惡ʠb�(1 �O��\�G�[>l�6P��F�\��U0iݽG,re�e�O(Xl �j��!�c>�[���)����pN@;1'٫<�����e� �9Z�d��E�	a��t���L���ߢ�&�0�+G/d�@-;�c�Yx����O^�xX��Њ�%V�x��`����Ĝ�Yߴ���|j����d�by ����:~Yj�`�K�xB�A�w'�E<����O����O����?Y����4���3�p4c�;]:�J7�ߤy������(%�T���3�0=y�f�$�����ɕ� 	@x��b8&ixq�{֖�k�I^���0ua͏av�L��n��	��D9���64���Ԧ��'���'�2�'w�?����]���Ì��\m�GH D��z��V���@�+V
y��JR%4������Ly�#ܾyO�7��O��$ ��=���Ø5Մ�QD��X0����Ox��T-�O��$r>!�W�O�b�� ��qbm�
Wa�,¥#�&rp�����'��+���Ղ�T�#�JP�k�<��&F�ax���?���|�oʍl��A+�i��^N�剳'��y�ǋ<_>Jy�`� Z��9��
����?�'{Vq��瀆SR(P���7���I>A4��4����'O�Y>���˟�	�
ׇ�>D×מJ�0��QiZʟ��I�U��]�'l� %�dm	���,�.���'x�)�2��q��A�ejU�'�~������f�P;��15T"}�ϕ/Og:P*P���T@� 2�X~�7�?y������O���c�H�I󈞆UF��J>����0=�4�O+8H�QB�4��d�ŠMZ�'R�}eHNd5Xr��\=r�'������O��$[���E5$�Ob���O���i޹�C�%j!���G;,j U"�<��*�����0<��m�<�x���Z���SEED�M��P��� �� 7̏�|#�|�|w� }R��k*��"�_* �l�Pd���?����?9���?���,O��Dٸ4��!ף߫6
�W�Է��˓P$�G|��d�)T��IIA��2v�-�Fj��X��I-��$�Nf�d�OF��Q��O��'0o�Y2��ԹH����W/h�Ա7Z#.	������?���?!���.���O8��X��Ã��=�4�5�C�$(.�(BL0��ʀ�C��b�&)5)�)��O��B�I	
�k��T#~��a��265\H���OP�6�d�O^�?�	*85h�T!��|���M &a�ȓ.7h��T&�d��afЊ Zze'�hh�4�?I/O8��s�$�'�|��a�%a��x�!Oާb��Kc�'2�9���'��	V=X�&(� ��/F:x��*����s#`ٰiҪ<�7%
N@@s�*O ��cܥ9>�8@�'9>]lZ* n�D�㬞���QbA�6Mt���g�"�'N�I2R�&|H��0򔙳3H�iO���!LO�=���=,�e2dfׂ?/^ [��'���9[&xp#d,��I�=�u�O�Y��W�p�&�X��M����?A/����0�OVL�����i�2-�^�B�J���O��$_��|щ�쉷t�v��$@?�M�O �S3uX@5K�-F,V�xP�/{�P�;��2�Bm��1CE�E�UP�>]�e�&j�(��E�u}R���O��zP�'�����T)�*�h�q@�&d�^TK�ǄW�<q��Y�z1CV�V$;Ɲ���O�'���}�Ef�� �X!�d��	0I9���M����͠lB�i�O����O�ʓ!a㐥Y�w���І��N0��bt�T�<8B���'=������Ϙ'�2�b�B��4x�1�0��	�Z9,��TH��:��'���#m���Ϙ'.� kf�E=�48k�/P�#����ğ�g�'�ў4���!��݀%K��U���V��l�<a�.�-�P�÷��.O��A���hy�� ��|����DKeh��B�F<x2�t�3|o�� e��O����OH�d�<�|gf��#/K�F��3)��D6H��*\��b�IW���y��Q�2K�����Ԡs��F��T��G"�
�J?~���'#�|���"Ġ|��螩p,"b!EN�?���hO�"<y���
|������X`<`��Ey�<��Z/|`�y �+;@�K�Er�ɪ�MK���',x��OU�C ����+Djݷ;�����'�l����G�#Gϝ�2y2dk�'y Գ�ᝨ4 �q;�i�#։x�'J�Аd��6m$��e(�*�� �'�x� h~tzeC,
�E��'ނ�	�� �R����8b�t���C_�Q?=z[)C*��M=ê�����y�[�w���C#��>�tQ�"���y��ˈOr�A��'ր1�� 3ß��y���
�p��ଁ,-:���Pǿ�y"+N�6��(�	O�7���!Eԩ�y"��c^l�1��\��� m���?�*Ya�����u�&ݚL�jp!ӧ����+,D�Р�`D0�|@�5G8(� �2�5D��qM-�9[ �B#W��a��4D���$ �"f�0��5:��v#3D�8 `�ޜ%�
��2O�	�*�*�0D�D[w
�:z�d Y���/���r��<i��B]8��j�H1`�$93�ގ8CXT�h*D�� =�qF�$��I#�Ck��it"Ov�pҨX<S���y�-��U�� "Ol��*�pN��{`.��d����C"O:(��G�T��=@'���^��b�'�xI�'f6�q���.���z��l��L	�'�|�2��܀o���,×]͒��'ʶx�W�@�|�[�LQ(PI��'*td���qAlyh�iQ�t�f�Q�'��ႃ�l,���@�km��
�'D��Qˮ&n(�E�ŒY��M����.�Q?�������!ӌ�^�!�H#D���1o�,�9ڤ/ R/8�Q�b?D��
ï6ڤ�'Ϛ�X�h�Ce >D�8��)?;׎tٓjW���� 1D��KG�8��M#�  2D����O.D��C�M�@�l�b[/j��l�O&9�#�)�'6�,`	@a�;r:(1����iR��'J�C���3���?^��	�
�'������f��-Z�$c0�
�'8v q�Եx��@ƃXF
�0 �'}S�,X%A�,i��m�E�$9�'���S���5�Ш��B@�8Wr�;,O*U�T�' ��j����1߀x����0�¸C�'C�I!� 3z�`��t�	3 R �
�'�Θ�W�M%"XHx�Q�q\D 
�'�h��*�;.�	qd�Y�j32M�	�'x!2%)o������|ݲ	�m4� ��6ή�����83O��لH�h�ȭ�ȓaݴ�G�_�3�X���ʂ`����ȓ�J��AӬFw�u�©�4^�ȓ.��RO��~�bmi`H��a��d�ȓLyF`@F+���t�b��T�����~P݋�FY���E2�8_r��F{d�����(���!T7b���Ř{�j��b"O��0��PhJD,0�%��	͛t"O|�q�jڏ"RZ�P�� AR1�"O��s��ۄqW^�rw釫a�y"s"ODh�&�b�t�L�(N���"O$��b���(�4fCy'��c��'�x�
���F?d0u�Q7[b�`f��	,�<��7ֺ��(�0kvnڠ͏%m� ��|0ݨƅ�s�vh�ըߙ"�f��ȓEܔ�#͘It��th�$*T��ȓK�&8��ʖypls�$�z��ȓ
�����l�j]�`c�,��\p�ݗ'7T�r�Y��=��,�d����v����l�\����f��1p�ښj����vQ���'�:d����oR�g��I�ȓIZ��S%GLPP�F�W��\��cX�: P�1�QA�̛:�����	$Ecx�	�;�! %K�CX�T3�J�mB�	�Dxh��%�DP!"+�*chC�ɄA\�@��͒�u���Z�(D^؜C�ɞ_��Z���!P:�+ ;_�nC䉓����ț����vIR�B�I#4�DlCT�U� Q�L�چ��=�'��E�O�x�"�M�9�f��q��*�c
�'uP���aS1;�Z���=2�JT�	�'�X$��oAXl8�$D~��	�'�pt���мƭ��(ҽ���J�'���)�Fن��q��L�;m��m �'�@�IW�,`)�M�F�H���Fx��)3�n$�3!Ȁzʠ�A��.YC��1:��0cR��X8*�OD�w��C�)� �1��Ȕ�f��%V�$UX�@�"O������gl�X�������;"O�(��/\Oьز�n���h� "O�)���2`�4%�����Ȁ�S�)c�(�O�x9�� ���O�aJ@m"OxQ��C�Cq�Œ��G47��ZG"O>y(A	 �&�|� t��!��i�"O�4sS�W8Ħ00����W��P"O`�G�ܪZY��`��Qv|-���'���8�' �܁��]*{�I�U��8.����'�R���nލd;rx���P�9K�e
�'�8���Ǎ�r�.UJ
�1͒�9�'�HQ�
B�
|0x��  a
�!�'\�	�ՠ}E����Pl�u 	�'��4ϐ�w�����ۤ8�05[���>]Q?=@w,ҵ<c�i�CdͲE���1�!D��B�H��ay,�)l�e�j���	*D���㭜*gyr����_�)�h�3�J;D���
� C�bp�f�+	d����<D����FY�Y��d� �[�L�(R/&D�0SI�Ƭ�'�S	�!�Cg�O�}�G�)�'Wt����?7Z��;3-]8r��Aa�'���jьP�H�K�O�H���
�'x�5[�h�%Ym�"�J���,Xk	�'��� �PVT��i_1�A)
�'> ��e\��⍙v��?Ѹ$J	�'��X��O��s�\M����;�Dm�+O0؉��'�∫V�e��)[�N�9�9�'; %I�ǌ�*�d�)ǨQ�;%Hԑ�'�xi3��&8�1@��75v���'�LXxW��"2�ٕI�:8 ��'�	"4��-+�h��J<N�|�	�e�<��{3ᐮ��t�[��B�Ԅ����P�ǌ�=j\�(��L�6I`b�Æv�n�F��vӢ���q�V�!	ϏO�P���	�A����ȓe�dD
�I�Zp��g_�x�ȓԞ�
U���>#8��Ć=s1G{�C�
ب��I@0	Ȕ&`�峁-D�XQ\�%"O��x�(6on�d��%I�s+恈"Oj��""��(�2��C��#\��q"O�YraZ�g�2��V��%XF���"O�I�d��_���+㟘hc|i�!"O����b9�Mz�"ٮT+
��"�'@.�ۉ���/:�u �i2GT��`��	f�@�ȓ���qNǝB��l����B���ȓ  9��K�8����+&�n-�ȓ?w�=h�wNm#¤��_?���ȓ`�6���Ń�!{�Bf��%. ̈́�A�����g\Ȟ�Bw���&��'��܀	�d>\�A*��r�$�Z�,�[���}
����:�|E� �y��<��0iv-�o#� ��QD�
\>��ȓ*�ʼht�^�1�"ȳ��G� F����K%�|Hb*޼-�"٪�A�)/�؄��8V�F��>U��t�U�¶	d�bb���#YLB�	&k�X��mB��tEK#O�&��C�	�{�h��F�4�ifb
2Y��C�4	��l�W%Vh��*9Z�C�ɏ8Ar�6�LaNy��O�B�I8J��
QD�8'���83��81�N�=�f�Qm�O����A�^7�v�����"Oҕ0g�G�EY��9�"w��@�"O���s�\�>m��{ ▢q�BP��"O� �%��"��iQ�DR�㙪Θ��"Oڼ�b�k�z!����7TO�q#�"O��)H@����1k�1��P�F�'n|�����S�(��9K1���v���"	�ȓZ��$�g���A��8��ʃ@H�T��������V]Z� �En�*)���ȓF3��K぀�4O��SUb�NZ���l��Mkr.ьP&h��$\Z�4�ȓjc�ӄc�:��V��q�x�'��k��%�Pd]�iaH���%��lp�8��;�����6��I�����g2D�ȁv�Y�>4�y���D��]j��3D��Z��ҷPZ~��щw��UÕ�>D�8"��E:A*,,�s'�30��p�g�<�O^�R��O���w,BJ�\!r�LC(X�\ �D"Ov�4�
m!`��G<H�l��"O����	Q�ڕ�"����{�"O�՘0�ͻ5��H��@��Wn�[A"O��AC܈h�0��B9VG��IW"O�p۶�]�oZ��jal��Y����_#H�~��S�r����� N�;�|��%�c�<��c�H���	�(6E�X#��_�<��	":��L�Ү�`�RE��h@Y�<�a͵R��� eBǽh��哗��y�<�G�gf���EZ��Q�U�t�<�sE_|D�ݻ��ل%.`uRv�Q��;��'�S�O	�@ `���'<�(I#���t:s"O|5�'�Vh$�(R ��(�<pC�"O(�C0��dBq�@��n0r`"O��*qL_g!.0�J�,d�m[�"O�99��
�U8*(�B��C���0O��[�NO� ��a��#{���m�O�'�����'�y��П�ρ!�VL���"sv��2������gb��l����/+z�YB��Չ%���#͟���i��ک.�"YQ �%��#>���W�Z���
��G��/�6|RvCU�\6�� �I
S�lI��	N�.���OXc>eBƭ85$b�P(͢�F�<����@�ɰP)�EرJ����	��$���4�B��ɒ m�P@��P#��I�e�氩�4�?�����;q�$�O�Is��H���ΐh�,���O h�ǉ4<���j^�IV$��|���� V&�A��
V7uZ1��B��yb��{üe	0�x�� :s�+T�-	&cЬgA���  Q�>�H�	a2F���Ov�S�b~҉��/�Yr�$���uc3�y"��P�b��@랲�xY�����hO`tG��_
FK�4^V��A��Ys5Oɟ�'P�9u�'4B�'��P��� �v]۔G_4<����7�@	��#��� ��H��`�4Fx#V�R@l9��>����d�FwP�1Zv�'A�0��� |p(�Y̟����gC��N�)?ve���/?%���$�	S�'O�D��n{�|��@%.�d؃�)B�x5!�d���~��G���DT��eA*'��8��|������ʌ=[���(�����c�'#H�t�Pa�OR���O��d�<�|�e���<k&��⮉5%��H�CΔQ"�8��*3��xz����y��ַ���d�� `�#��_���o��s*�h1�['5�y����?�CL��VDUa�D/wѸ�@ա�?���$&�	�6I�&#�&.`sBU.CTp��=g0Tp'��OAb1#�c�A߮��'��6��O�ʓ^��C���Km���45�B���� KZ��?���?��_
��fK	�b�XKG�����H�(�"�ȇG�B�t�)��^��O~���ݿ�<h���
�\�'�ɑr� ^�t�B%͛t�,DD|R@2�?�����O1H��lOW�@���L�b�d��/O:��c� G�Tx�d0��V&^?�}2�<���A%{�ޭ�d��8
���Sy�F�hUf6��O�����O��^"+�4���S�s�jHS2.�@�D�D�,O�9KtN-5�(h׎���"~R �mYʁx�l҇_\�Dub��<Qd#R`�f�����aK��i��)���`�d�v"�(�g�ʨp&���/K�'��)��8?� (�	@�6��\�5C�p�F= �"O,˙
n4�w�F7H�Z|���ɼ�ȟb5҇F�
�v�CS%�3��%�3G�O�ʓ|����i���'[�R��WU�x���'}-� "'�%s�N�ƣٟ0��E9D2��3�H8Fx��.`0^ԻÓ&J���3���Z�fDsu�'c���'NF�T�\a�Ο�|;w�ʨ%2�F�!{�� r�%?���ϟ��IT�?�O*D0��YY��5�<Ӛ���'4j� �ۈDz0�Bp��<�����O����|�'ى@[�=h� �f���(��ё&�J�r�-g��'x����'4ᖄ�Vk�|>�= �)E�1.�Y �'(�ČZ�ޑ ��`k��'�\v����ԢÜX�y��N	��`a��|L�h���'��`a��e��2!`������1RΔ�0���hO(">!���	���p'�]5o��s�j�<)w�����r_
(��Y��IEdy2�w�P�Ĺ<Y��@9i����a�� O.[4,��$E�o,b�j���<���?��>�.�PMz'�h�mV�_��O|1���\�z�D� �+U��l�h��dK7p�-J����9A�C��|�`蚳+9�ĺW_-[�p`��n�'
]{���?9��4ȀH������=&�l1�6K����O���d�3%�Ҋ�P\��q��}Bd�<�� ��qY����*h����d_Yy��'��'2�^�&��*���!�����B_^"���	A�'GH�@%N:�v��,lQ��cí����O ����>DU
����ٸ@��O���غ��O�s�\a�Z7m�P̋�j��l��xC�M
����'��'���N��PJ|�S`����`�!��Ra ��nD!9X�'�`��b��yR@ީ1�UR ]-i�`�Xb�0Zd��N���I���V�>}�|��/؞	��0�cY5g`�h���O����>���IQ�O�F �4��// �� l׬RnjyZ�'���
M���K��p�#<}��u���r��]0p	q�C5�t`��R��5$.}��3�rP�	*��G4q�Ph���N���ep��O��#w�>��y��_�;�"�'�f���ߌb����S@�(x.{���^���Q����x�>e�%�4��T��N�~����P�OZy��'��{�O�s���ׁ���Q�O�y�nY�FZ: 帜��+�O^]!�j����n�3���qď�݅ȓÒ�z&M��d躣���"��'��՟$�'�b�'B��O��a�&
�bF�Q�![� ��̋T�i)�|�'&�����Y�0 �>w�HmK3 ޸ ��2A��(�S�3'p��C
��ܵpp�\pCfB�ɢuCV0��[7`yR�H�/�BB�ɺ%�l��$e�E*<�cT'C nlB�	0JCV�r�F�v��ġ��<)�C�	���)ƀ��(�6%�B��	��C�	�Qc��Z��N�`�s���S�~C�I-���Ԩ�,E��dK�[�ZC�	�'�z@�%�T�HQa�?ZW`C�ɧX%�"�f�̌��"Њv	"C�3P��M"���.P�t��H.:"�lZZ���S�b�D�:07-����߁�B䉒>e��@K�K$Ta�r�ވF��c�h���mL��1� C�+�0�إ�p54�:�Ly��骆��+6��#�B�'s38��'��`�0ɂ�
8(?\�S��$B�HI���1j@0�1E�9OK�=¤��T�d4�5�T���x`�G�T�`�u�C&SWde��24�$E�.<b�Դ�B_(!���BïJ5b���Ql����X��ɠօ�$C`���Ѩ�ڟ����K<�IJ� �!-�z=��-K��?�O����r��K&O�f�hEy��ͰΨO�U�$ �q`P�s�ӁW�*�|z�"\���r��.)�mT$Js��\R|�D�OJ����d�D��;7��q��ʒ��N����d�OH��ďe�<B#�)V0 ��C�Q�~=�x�2ʓXC�F�J���h`�J�.�X����?��cZTx1��O(`h���&y�ȓbS���d�A��$�u@����ȓz���ɑ�/_"��@_*�E�ȓ�f`�$�ރK���j��?
�@�ȓ����r\�OG�!�Q+¸!=����b��CC� 7"����� ,5�����+�&�+E-�#V�e��N�3�r��S�? Ȩp�Qm�RlHd�K�\��"W"O��8F�ω'�I��A�}Z-3!"O��J��t���Î\�fT�D "O�p����7m��kG��vFj,�"O� ����
����9XE��$"O,����Q�h����,L�Δ�"Of�۔l�������<oyȄK�"O�8����@�FE��ˁ\�� C"O��%M��ʥБ�':��q�"Oh �嬖�W���bgc��%�����"Oz\�� Ŕ�<��a	AF��1#"O$�J�$,/�� �	�
JZ��5"O�U�U`��b�d��♽*�,�yV"O���v�W�fXX���J�gF�|��"OB�V�ϲI)�Lcb�yCvaY�"O�����Z�<8��"L�x�l) �"O�����Cx԰Q֤� J� �Q"Of��RKǛ�L��F��y�B��s"O����]�()4 a+]W���(�"O>E���w�Pz��T0\|�K�"O�-��\��ұ��2gfމK�"O2��w�K�1��*i<\X��"O��X$��b�
A�A6��"O�1Tl&��!mӋ&t*�"O6	�¨)D��a�lݵ0�t�R"O2��˜/Tsz̒kX�2�b �w"OD��5F�z�yQ`ܻ�nՋ!"O� �Ǟ�I�iq b����93"O�|�1�T�y���R�1�"O���uh�������.��ι��"O�-��L��t��".)/حS#"O�R�ɢ4bU𰋁�|y�y��"O�T,t�z�D�\4f�a�"Or��p@P�wu���WF��4,:�c"O�=�@�S�}P����H�Z����E"O�D�P��((�^�۴ǌ�	�İ	�"O4X��Q��x���η	�n�X�"O�Dy����,Od�9��k6��r"O>5�'ʇ b���T�0\�;*O�m��' <FFK�mC�����'��T�v�̨V�xP�-��D�'�4)d�L&�V�Z���%2��+�'��\cd��q�E�U$Ap��}�'Pn%8 � �T<���BϚS�&9i�'�H���BT�YC�9����J�d���'��a�'�\X�F#T��,��'�`���o�=> es��Z�R��	�'Zy�,]  ��$�����$�tl��'�j�(��&'�V )�������'����A��4*
�(�hK���5k�'���S!�0Sԙ���'"��
�'`1[�G��l��cDΖ ��d�'�8ya��S��8:t&�}�:)��'K��sE��o!�l��ƲGCp���'�n��b�q��!s
�B�¹C�'��P�Ŭt��Ӆ�*e+f�2�'��xK�B���~�S�"nn����'͞�6 T�D�:���]v�V�K�'\֭9�)���̄�$�K�tZ<|��'⚜	b�K$�B]��K[g�DI�'#��e�J�=�-�sڒ^���'#6p �i��U�V�r�*��=ΜXb	�'�n!���S�\�RP�RM�8;+&6D�X�c�� }�0!I1@2�H� ,6D�� ����Dͺ,)D�M���bp"O�Yb���8d����Rd}�6di"O�0�C�D</$ k��� /ZH�'"O�t0��ڸ\�v��[�r����Q"OJբ�Cә~Rf���
�K'"O��
��5B��l�Q�^&��
"OX홲K[9~^����k���"O�d�ċ/�k񥉜F���Q"O^�d��
ζu	/��	&"O�u�C�ùcZA��KH�"OT�QubBh���,� �&�T"OP(�S��v��h�a+C:�6���"Op 3�O�3�b���6�)��"O�܊a㒁L�N�+��ʌў���"O,��Q>=݁Fj?]ֆt��"O� P�J�k�f��CJ�(Ʋ�	"O�9x,ˉR<<�Mk����"Ov����B"-��ݱ��U1W>���S"O"��'�8t󾨻����*!t0{b"O$x`��I�I`�����G��)T"O�ч��<�R�������E"O�iC%i7�����@��@@9f"O�&��jzX䩏W��(�'"O��p�ԣ((!��N���C"O̽12�v��#b���R��w"O���${�8�U��UyXh��"O^��S/h4��2�Ӌ#h"y�"OD=
��ڼ����`<]��XT"OFXQ��:'�I�d���dj��U"O4�١�#)�p$�U��Zxp"O��1�K[�D�����.K��rD"O��eaX����T��$K��<�7"OF�CU��G��q�eHX!�H �"O�5ɑ�	0Ts@ۆ���[��@��"Ox=��)A�m�4�V�ՋH�hP�B"O���'
_��%"��1�U{�"OD(�D掝O��ݻ��Od���"O6e�cH �N���sm�}��8��"O�`��J�9�2�
�9]D4��"O�L	�$��KI��K�4�q�5"OL)��.V�gj�$+T-V{�(��"O^M�C�O��t#��������"Oz���.@�A�N�r"��
�*�9r"O�{��O�
vd���׫)��%ȃ"O�@��:��QP??�l�!"O�� �>'�)�fP;8�ܨ��"OqcBi�$F
���B�e�����"OB(����X9:3�ӣB���"O<9dF�,^��Vl@� �(|I�"O Ћa�P�p��֤�$�R��%"O���U_@�qaDБE�vɊ�"OP����
��i��N�-) bI�F"O��[4��*���� G_��h!�"O�0��M����SF&S�0I�"O�Ա��X%\�! �ȮT���c"ODA�AY�2��B#��~�օk�"Ot���ms���R-їk�Ę�B"OhaBf+�$��m�b
��MD�r"O�u��I}a6BU�<�����
>e%!򤕥Gh5z�H��1�h	x�/B�Z%!��0!����ކ}r �t.V9:!�߰$��8�K �?<�K�cF��PyB�ٿhȢ���OY�~��`{q ��yB���2�P`�_b����D���y
� J�`�jG��%�f�@m��"O��K�v�̡	�Op�}Y�"O%��4hD� ��!+�0�"O�K�*F5Ʋ���U�#)h��"O�i��I2]�e��័^�؉�"O�qx��ǳ63 ,"��f�Ƽ�0"O��p�c�9�AOŋ[�Jh	Q"O���BE
rXT�.	>^���Pr"O��qW,C'�.���,� �ꘘ"OH�#��ٻIJPйK��}�N�80"OR�#G�9bT\�J�3��(��"O�J��jZ��r�/�=0���4"O̔�熎�S���[��/OČe�"O����	�\�9X ��.H���g"O$i�υ-�m��o�!�(�CA"OƼyM����	�#� &�>`"O�\�k[�T�`��d+� �A"O�t�`�5���"Ad��+�4C%"O��!��:c����:+��A��"O����^�0���ԕs�x(0"O
 B�KZ1����Kߐp�1Ar"O$ B�K�>lq�1�댐)�@4S"O���5" *`7�R��4s���)�"O�aZp��mQ!�2�����"O�%+#
O,>]h���Ք&RQ4"OR�jv#��o1����Y�MY�"O>0"��3UE$$���6���"O����'&~x1��k�g�1qE"Ohc�b��/Y��"˅;6���7"O(%i%�Lyb�=I���?�8p"O���$G�_�l�p�D=�l$�Q"O<��É==:�R%敁gs0�Xr"O ]�	���pq��D�%q\Z��"O�4c5 Թ �"�E ���"O4�*� a�V�`�a_74^���"OnQ�A �#Z5�I`�`G')B*|��"O�\�a���[�2���h��h3�%�'"O.Yj�n���>��AOB�*�Z�"O�@B�D95 ��Ar/�u��P�7"O�鴋�Y	�y���,[Biyu"Op����K��, �H�h4�e;�"O���B$��`���V/֝#"O�a��D�������
	*���"O�1���i��e���C<@V�hV"O�T�fT-Ct8k�@
�l2���"O�����D'*�-����4�j8�1"O,�Xdk�Cc�\b�e	���%��"O!��ݪJ�Y�u�Y����1"O�����4#��#�B�7�-�3"O���B�U���s�A�'2� ��"O�Q��C�^���B��S��	J1"OPepČ2y�5{�������"O���MY8-z�j��Պ�s"O&������h�%	$uy!b�"O�`�S/҈$�h�`�'�	@u~I�"O���M¨1F��c�戣F`��p2"O����"Y�(�&ջ3��@"O��ۇ�ݧrQ<�j�CжP��psT"O�*bHFe��s�Q�_c�=�1"O<t���'�Ν�@�)��$��"Oف5�2 �1)���8W`��d"Oh͓vkۄT�<رW�	+F�Z�"OZe��cP<S��T;��a�	t�]�|��2��F��h�T�&<O���0���3��ܱ��,�(](�"O� �!&���}
��q���"OĘz,3�
�S�	�q���""O2}��Ŗ�ޱ{9B�Z��C"O����喋:�������|%"O�e��ʟ|k���DFO#�ɚt"Oj-��A;+cL`q&��>�ʴq"O��2'��!��-cE�_'\yF"OZ�#�10�E���Y,>�#"O(�,46}(�hc�A�pzI)"O�k��0�M����h}
U�"Oּ0�B,-&��sg	,OW�ZV"O��Ā�%r8Cs�[2%���'"O��A7�[2i����?F��2"Oh���˧#g,]:�cM��E��"O.y���״^j��p#A�{
JU�B"ODa���G}���En����3D�h��(�	G(vs���v{��.Y/!��_�{�L�Nߠ��R���]!��>b�i�W-1> )3�\�8!��'BJq��������6!��s��@J�;<��K�NB�!���&@P|!s��;y9� -�{�!�$S�{��myC�U4o{&�{��1e=!��U:+�$�u���F��8����.!����\\c�fӯd<���Cَ#.!�U�E`$�E1"����L?IL!�N8[3.�p�+��s#� @�k@!��үk�L}��Tx�a�s'G�o�!�DY)Y{�9�7���x���$���!��
5.�h��B�-7��lKQ9�!��C}�X��e�2hhM ׁ֜I�!��"
����%j��CLR}�Ӏ�+�!�� ��	áH���Ub��� #�!򤓺%�
`���1�6]��^4)!��X&2$�圹V�;�c��	�'���f�м.�}�@׶IR
�
�'���A�R�2��@�g�(�f]�
�'���i���c��`��_C�q�'jN�zEn\X�9#� �wN��h�'���ȦM2!�1�KEB��(�'��	�׬�t�Mp���i5�!�'�0Y"���1x�C����VJ�
�'���d�*rdQyW��>%{����'�(�3�@]01v��lٕmyz���'Й�#.\ $N�L��)c�a��%D���H�;f���GLC�v�����"D�J�k�j��=-�0"w�.Z9jB�I=U�y���_	(��,����/+�<B�*�P�aۡ"�܁C�ߎ�B��D_aP��� \�1��3NB�ɦs�x�aq�����	R�\C�I�<'��@u�ĵa%���*`>C�ɒNH`�bA�i��2��^Z%>C䉦
6 �a��1^F�E���8?��B䉐Y�-s֬E]شգ�"�>LH�B�	`cڤ3��ΰ��	+a��3B\B䉝Ġ	���u�-ZST��VB�q���س/���h��%��B��$����T'�C�rpY�A�g'�C�Ɋ#�D��h�>;�-35Ā3vgjB�	�=�HtR����:�*͑�O&��B�I`X�����_��*W(L!)��B�I�9(�sDEu��0{���@zC�I�$ t�[櫐�y�� ����NazC�)� f��I�&`��ޟ|���"Os�éH���b'L� ����"O����4���Z�Dc����"O�a!W'�N>�����8\����"Oh8�G"E�B����WL���G"Od�t�� +��t���CZ4�r"O�I���'�"� A�3	Z�$"OpU"��%+�t�W��4L1Q"O�(���|]�I��E�h���f"O��r3��c����� �{Ő��'�H9��
ٽh�Д�F���)��'K.�)�@�*k�8@�6��/Ϫ� �'Y�EJ� i���S�P�����'Ό�Y�莚%�=6M[	�A�'����Pf ,.��0H�-6�@��'/F0i�R�|K�E¬&��b�'�*=j�ѵ��;E�ٟU�4r�'GM�b���7[PŒ�!��RH���'ښ� !KT	N��-ش-�Sd0���'(�æ���M�Բ���"��$�'��%J���2P±�^6�:�'�N��ǻPc�c 4o ����Ѻ�y�g�!?L��3#I=-�HP���ƞ�y�(\� �*���D�,(����7��.�y�k�$��a�(��m��� g$2�yGP5 D��5��"�810&*ɔ�y�AӷP84��WI�0C*tA*f��
�yb��:��FJ�:sr@|�A�
�y"���
�4��f��kU(X��!�y�P�D%R�JJ�y;�*��K��y��4&@� ��I�E�y�u���yRKF�q��P�×#p:�ur���8�y�Ţs��4�Y�q�A�vR�Y	�'�`�ф4m��8��	80.5)	�'�DD�6�I|�F�IF��7��k	�'��]�!	��+,����LW0%'��*	�'���do�i���[A��^��TH�'54)rU˃�'���g�T9Z
@��
�']�}��*,�Us�ƻX8v��'sFܑ���0<�~h� W�f�z8��'���֩ME*T)Ѕ�H5K���
�'Q���3�J"1u�u��,�wFJ���'?�8��ꟓs�~�
4g�?p���b
�'>�HT���%�$!����jJ���
�'/r�5e��U��LB�`	����'�iR�E���V
�Cf ��'i�(� �{xR�x���3H�aZ�'LJ@���n� �[F�^�&V��	�'�|8��,K���9�d�R24��'�=3�[�V`�]WoCӜ�#�'�)�tj=-�E��T�z� H�'��}�u��z���NL:�xT9�'����H�5W�ZD��cI��'�
-"�hQP�X���(�tN�[	�'��m�W�U�+@�t�O�$(,�	�'����1Ƙ;J(H<)獜+U�©�	�'���*�)���^$��!�'�
F�M#���v�X\8�1�'!j5Xt�Ɍ Y�1�3�H�f����'@,)�񯂟Y����[:�V���'i���	�2aż,
��߄;�}��'R��eE�b�p*�eG�d��'��%��X%F<+0N͹��@�'D@Q"RB�v�܌s��5�N؀��� f�S�غw�^)���!p��!p"O��fAS���w�Ӭ;V�Q��"O�|�6��"8@��E�̀?KT�p�"O�4��l�9q����ĹD"O��Kv#� lL��QkN%�|E2�"O\Qs���	yD��%��e3�ъ�"Oʘ#0Ĳ>�^�����b���"O��xq��[�5k�� y��z4"O<������wĮ��S��bibX{5"Oz�c���~?6Ղ�B�)��$� "O� �B��x�F�����I��{7"O�*U��E�6Pf�CO��"�"O�$;GG׍x,\2��[�p�1�"OR	أ'��$�r��$
���"OڨY�G]I��x�0ϩ�|��"O�D:g+
�:H0r#�+^ ��7"OL!ICH�(*��`t+]�� ��"O��B���7R޽�dH�W�\1h`"O�j�H_�)5J����ݶ(���'"O|,�E�
9n�ܨ�aoՄ^���W"OD-����.��@��"v]c!"O�gA�4)�P��n�;䲤�@"Ohq´g��-�q�fS�Hْ$"O\$�D,ۄ? ��f%͇1 �"O��
W!Q�5jE�S䗊&���q"OT�8�*MXA
Tj�$t̴(P"OLq���5_r�y�*��cWLl��'l҄�tJ�*L��S�S�;�*��'d�tb� �\*����;�ޔ��'�(�ˡ�Y�U+"���)��x�	�'��tG�ޮnw:�z�C�\Θ���'��y�Wl����Z#�1Y���'��ȳ��F��A��>��1#�'4м8�X/_�rm` G�'����'S�����Pi'������Y6`�A�'3�803 �99�($���O�P���',�eR�H1~�( DݧB�=��'�`%[��D{��y��Ld����'�$\P�#� N��<���I�rR�Ԓ�'���B�+��{��$QRN�i�*�'v� Z�"/#	�l3c@W��H�'d� �Q�ZD:S�ҹ
��͚�'�4Mrq��)x�cM�0
r�d�
�'��+RƖ�-��]���ʧj쐙�'�`i�%O��+t�l�b�.A�0�'�X��U�f�r�eК+���'����խ[
4I%�Ÿ(#��I�'����U��|B:�SU *Is��'j��!���;+���r%�9�.	�
�'y�|J&N#T�̅�L��.��Y�
�'�`@�qM9p��P�˄(ސh��'h8�S�jǠ^6d�H�BR�7��L��'.�$r��+�~�2��Wd�ui	�''�캥f�A��	AC��M#J���'DZ�+̂�ZE�"^�A�.�:�'6:8�`�,5�6�(���H歫	�'4����#@�$w�ȩ6�d�	�'ĸ�b����`�|Х�:28��'�PYu�PW�(�A�Ȏ�`��"�'�8�2q�!�y�#�#:`Mz�'.��Õ!�|D�bN
��X�'�^�K��[���Pk��3>���R
�'��@	d��Tz��`��P�
�'<����	
3R� g��������� ^M������k�e�$�"OP ��� R��4�"
˄}
�ۤ"Ot8i�$[ ��x9W�7=L�`P0G��2cc��SŰ}���$<O�|��V0�Z4��KRs��cU"O���b���dԸ�)Aş�n0PE��"O��t�UW8��S&'�8(��[�"OnmSÃY�u�D+�.s1h#"O�#��S:V1��N$�:]��"O(=�EBC"c��ԑ�L�D�Kc"O�<K� �+Hx.e��fG�*�=�C"O�#iɱq̝�S��?ʔ3B"O��2J
���Ĕz%�9�D"O>My'C�B��)�cV�/�]B"O�a�H�!h���� c�� ~����"O���e.�*.�맡�<'�����"Ov�)��	�Uk�ݹaA��:O��b�"O`0�A�	���#'(M�L $"O���+E0����AG�9�"��7"O������z�5D�&a̸�rF"O$e�c�Ъ��
t�*Y��г�"O
}�	O&C�� �� 5�f�H`"O"�`#'ްJ�<qeBV�e�����"O��ء�˦|[�h ��ą?���1�"O���o�)����B��1"O��/��R	����#P�7v��"O@����[�&����\V{�58g"OX��Ǐ(t(��WbZv9��"Oډ*�l
"�R�ꤧ�bI����"O|���$<DDZ�(94"��e"OT��ed��0˰izs�RK,���"O���!��3<�^�;ń�j9��9�"ObT��z�� 0a�Z�Ϻ���"O*-��J�� "��#^$���"O`����T�:=��q�֕v�h���"OX89#ə�x���Pa�)H����"O���b��U�h%�T�V�(:^���"Oа$�cT�����q���"O�0�m�m�vY���^�ޤl�2"O�\���\��x�j��ăTivyʓ"O𼚥��`���G��#S~u�"O^ ��)Ż:�4nP�8ZuB�"O&Yh��
�!J�=r&푊����"O
��&^�9J����.ȋ�"Ol�����9�����M�>��tٗ"O\\"�"-C!!T��:-**��"O���D�[6Rt�"G%�t�YS#"O`r�͂�UsW!9EF���"O�����=O$���o��q5x< �"O���P)�r.�·�-�h�"O��b1�RO���!�����6"O.� �߰	�����V>+�4Y��"O4��´`���FI��r�0(�"O��HFn�/TN�󈎷E{��q "O��R�ڣp��L*G˳`��#"On����@�N�{ D�>'O��A"OL�ː�41�� Jr�Y�F���1"O����N��OT�H '[.8q�Y	�"O`8�VoZXfҁ�p��"
t�L۷"OZ=�˅�(��i��f[*�(�"O�q�p��V�b��F���n*2��"O����#߽6٘�hH��$P�q "OZ9;g�G�,#�u*惽Jq<��"O��B�y�&����5Wtő�"O��s�2^5�$L�\ߜ��5"O� d0Y�HЅ"�6�s� X��+�"O���A@A���S2���N��<sC"OlTCuMԶ0�Ed�)�P��e"O����fY�B����ᢑ�d�� ��"O>P��*�#� �woVf��H�"O D#\%��Yb��͸y�xQ�t�<�Ĉ�?6��������p�<!r��fJ6BC#�?�L����PG�<	e.��Y���shW�o��=�@y�<���>�zdAAL���δp��x�<�F*	&&�Lĳ�#��Uֈ�a��O�<��E�Ma��� �%����'LA�<���]����뗱4p`�1P|�<ٖ ��![��P��8�lQ*�w�<�'�L/L��u��k�>�t�!�Po�<�cV�zq��Ө�4i��Zcg�u�<9�N�hjY3��� Z> �a@��X�<�`"��P�pe�F�#����"AX�<)b��Q�9C�����6��m�<B%��8���Q����M����c b�<q��=x�t�h�T̤QbgLy�<iDh'��ɲ�TX��YPp�Ru�<I^���2��N��5k� &vo�C�	�A����a�(|
+�Rf�C�I�3-h���I�NL�9�jK��C�I�*�~��fcC*i�N��@	2w��B�uKԁuǉ�+�9ZU��@[fB��>(�f�36".�|�C ,V�0B��&|p�Y�L�#h�˳���Z�C��>Q��� ��	�Z�
DiK,C��C�Zv�	�AeX.]nK�g�"��B��?@�����(?*�v������?W&C�I�ΰ�Kb�٦B�r�#�+>BHC�I.�l�X_�`8��B�8iC�I;+���'�1\� �Pe�B\�B䉉��pf��/]VH;��O�lu�B�	�{�j��d �q�B�1`%�	@��C�[��y10)�MH�I�[2�C�I�T��Q�A"T98���'�S)ƔC䉦���z%�T�y�zx��n���"O��R�۞D�
4:W�\�	甘*G"O�s"�����)6���pu"OE������̌�"�<
���"O�=p�%O�h�����
�n�:��D"Oȹ@3��(VvНJ� <� �ɰ"Oµ�W-��XH��h��3l�8�"O�e��V�>^��Vb]�sO�q"O���קY?g�d|�9f+��D"O��ODG� �ccֹ|�4�G"O�<�L��*&���`f�>b�`ś�"OH!�'T�1����dƧt@�%"O�b%w��ٛq�N4oe�@3�"O�qcn��T1+�	�.I�M�"O`l�T$]�\�
aȄ��E68���"OӀd� � I�JS�BB�� �"Op@P����"��T�BA��"O ��
8k���E��!��P"O:���)ȩ|��l�A�_}R%��"O��L�$I�
�GlZ�H5"O P:�e7P�� -��,� ��"O*�
�)�z�F�+v���"O(�Aw�]��DI�%��x����f"OR��AE�kU-�	_�r0��"O��A�% tԝ�@@�Bp��S��'[ў� 
��QV!�,�`�3gv\�"O�D�"�����-�!3N.��"O�B���{iL�����3�q�#"O|����(M����O�F�"O����`Y:U��J�ע���"OZ��JF��]�p�ߔ+Y���t"Oj1X��H	B7�JՋ]�z9�	��"O~PPAL��ӺÃaމ:j��B"O�	�焎O�ʘ���< d^�;�"O��!q&�eT��B����as�"OȘ�Em�*x�vm���&C���ZC"O����e`z����
����k�"O��x�hZ
��l{ӫW�F��I��"OH�3�!8�P�7"٠L0"O��%)�>P��e"Wʟ�(�tH
�"O���e�Dt��"��J�ޠ�4"O�H�To��V����E�.4�!`"OΙ*@Ǘl��bREg*�8�"Ol����w� ��O[�"��"OfJ�e��8���ĪOh�"Oh�B˝��4����%x L=�"O�9�4��*P������ �;�"O~��Ā�2�Pv�5���c#"O��
� @fߦ��U�Ĥ+|�=�%"O`u�4�B�� @��G�Pj�3Q"Or��j^F��l���+`��"V"O�,�w��;!�i!�^1x9~��"O�5�>DCGe��xʂ��T"OZh1�'�'w��� 0�xE"O����,Αdi&��A�f�*��"Oa� B�'�^�2u S5pd8��"O�a�ĩ�^t�-	�I�	e�#�"O���ʼ"H@h��P�WF8�Bw"O&��-�03����GE�@=,А"O�jUŝ0cBj�맣=��+6"O�}���M�KN���b��b�T##"O������,>���`37}���"Op�kQ-�DU Ya$OW�|N�()A"Oy�%�	2���s�͟�IBK�"O�s��gZH %M�4c0�"OJ0Vb��2j�kP�c(�K"OxźV��16�V��C�Ι�rl��"O0q���	y� -Sd#��H�#'"O�8��^�QȾLYbE(y#��җ"O�0Ƞꏀt��`��:2�&eJ�"Od0�B��s �Dڵg�|<e2�"OмH�E��)�xeZi�4J��$"O���b�:�|�0ը��G]�Ԁ�"OƩS��+��8X��ZVl:�"O�a����m.^�[@�:p1����"O<�``\$z�0u$){�͛A"O�]�,�1V�T]�c6�i±"O|�H��0S�p�R�B�p���r"O��뵊F�vD@Q�G�(sdT� c"O\��� I��`(S�)yx5��"Op�𤧔0}�x���ti��"O�#2C�.,�9�懚�
� 5"O��rc,��k�x��UB^��|�f"O>T�f+�.n|�#A,���hp"O`U���J���J��/q�V�H�"O @�:3'f!���يi݌��"O ����d(���5���T"O��9�B�$��-�d�̐0`����"O����kY�E�)dW�4K�,�b"O� 3�D]9g�@���+X[�2�"O(�"���W�HU �a��Wl��s"O �ѷ�Z?,�q�FD�6X����"O�X�%KO eefL�WEF�EX8M��"O�Hk�͝�"|��fL^9D<�"OB��gP�s��L�ш00+!"O�̓ ��_��x��J:���$"O6�B1�́,��P���"Cbxb"Oa���C4̰�ņ�w%D���"Oh���=؈�� ��bִHc"O���dT1Wp��bա��Z�"O���I�n��%�eeڕ[R�p��"O����oȚ1�p� n��J��"O�!�՚?�V���Ԫӊ�a�"O(�
��)0��#儓C��	"O�)cc@[�k*��壒�%��I[v"O�LSG6r�dYQ�m��n���`"O���c��0i�Z��M
|�Tc�"Of#��%9�1 ��S),��B"O�\B���y80���I,. ����"O�A���T�/N N:J��"O�P���¢h���09b���"O��w���P�|�㐕	dU3"ON5�Sg�\>�p��b�*IV9`"O���KˬWK@�G'ܫ7G��"O�qK�dM��JA�%]�@�)�"O������1�H� ��Q_�1��"O�{u%X2 -����4CO���"Oz�����oA��Q���'u&d�p"O4�Y�h�A�n��th�� u���s"O,����;����ħ_�79���"OrTj�M:+{�8��ƒf(�yb�5[������Kw椩U���y���+��E��p�"TZtj	�y�G�ar$0�ϗ*k���{ҩY3�yb"�z�Lmt��K<P9b���yr	q�"q0"/@=Zm��yk�;vLV�!�Cр5�xj��1�y� Y`f���.�8S��-ipϒ1�y"�q����,�L�H�QQ����y�Þ�q��Ĉu�Ju�@��A	)�y�\+>T�)V��`��� t"Y��yB��`��BE)�fQL���(��yb!U��Y*�Ϭc����gd��y⨓	c>H�����4E��(�<�y"O5ay�8���M�,z#����yᛱ�,�e�N�FyHj��y��]�d����	L�%�u�I��y���`Ր�vÛ�?5�u���yZbX���ԈF3�!8��c�`��Rg�B��Ef�8��@�6��чȓK��y�3�
�48Y��ĿtW�M�ȓ �	#��Y?JF�B�h�vH�ȓ;T���B)��v\R�Ї��J��=�ȓ.]�x��OF$`�Ԃ���ȓ�T�:�$W/5v���S��8�ȓ[1P4�r�]�Ľ�f"+3D��/�� a�]�ԅ&g����<D�h��C�gVt��#�n~(���!%D�T����0Q���#��ٴ<��#D���'Լ �d�E�^�[�����=D��$(��{���b蝵C�z<��N>D�TpC��w��@�����."�r�")D���aa�*L�xâ���f��*T�2D�� v�	/Q�~����h��l����"O��9%#®S���������
�"O����B�.5�؁i�(��|��Y��"O�a��\�>����)�.0T"O�� �	چΜwhÏ�r�rs"Oh��s�[�]
�:�L����Be"O6�y@�ʲR��<8���e�t�"OܙK6� �����e�	]�Dx�"OL�1V�8u�QjD
�=��h"O|\J�F�U��!��$#�f|�#"Oȥ����N��8� W�^�6H�W"O���Mݔ	A\0�%@#��@x2"O<�Q޶��f�������"O�x��E�'��`��Z�!*�"O�\Z$&�n�x��r�P2�
�#g"O�Q��_�+z�%��n 2��xf"O��4�Ӝ2�I�`�:��P�"O��C�O؃`�8x��C�U��]�2"OL�� �� �x@stED��|Z"O�г$��7^��� �'Ŗ�R"O��˙$,&�A��ݓ]���
6"O�zƊ	�P.�u��!] 4��ɨ�"On�*�$��� � [�D�4��"Oj�_,Q>��ǮB�R{��AW"O`B�҄a���$�!OPt�$"O��t+W�,�N��eg��'�6@�"O�i;�B��z�a�����Is�"O4���oD?'��ċ?C�N��C"O�%��f@�/��$hb#�>}��A�T"Of��ٜ%�py �6Nf�!
�"O�"��e������5�7"O>d���%i��cSkT�z�C�"O�Q�U��#Ja���Ӈ������"Or�iA�� q��x��ԂY�2�pG"O�]Z��!Z���f�Z��,i�"OU{�]��Rȩv��-@��xI�"O���#�^n�!Z�\��i#T"O�$���J�9*D��D�M�"3u"OJ�q"nB5g>P�b�l�-`����W"O��I(��Q�����j�"\s��Bb"O����+9{�I�wDA .MfH�"O�)�`$H�nd���+7�8��"O쬡�L�>����6�F! r���"O�8�K'n��	Ra[�y]T9pT"O�!9�� (m��d�R�m>�`3d"O5sqKT�,R�d��޶m��Q1�"O�|Z5#�3%5�q��B�X��q�%"OP̀ao�U���*Ҫ+��!!%"O�I���+3��)H�	3dM2�"O���գY0!XU %��V�����"O�@�j̮@��%�ĐX�� zg"O\IȵK�5�҈���A1yQ�|�p"Ot��ՋġrN�ѻ%�-�����"O�����;���C�I4��A`7"O�9�b_L���B���w��	Z"O����l�$EPH���q�4X��	]x���i��
�h�1�d=�6�  �.D�T�`/��lb�
R�i�@�k!D��xe@/Dr�Qb�d��NF����:D�Zp��P[h�;u�L�c�^����8D��a��&$�F�p �L�$V�!eo+D��j��/iP�IF̞Vzry���(D�lgś�5T�k�	�S�`I�g+%D�K@c�8|p��G�~b]��!D�� ��ĩԒ_��	BW[0��q��"O����Ի-�t9��ž1k�t9�"O����lޮ5�t� !=^v�)d"O(I2Ɯ L�f5
��U�ixP�9�"O��'��/X�\�T�4u8�G"O�e��̆N;�T�@Hkn)a"O��T/&EP�'lޢB_Pt{�"Of�b�g^�s'���kH5\(ҙR�"O����'9;L��q���B�X�"O�����Y�a�f	A2JD�୻�"Op��bÕ?&���1,B>!kJ��Q"O^8g�هd�~�:��AS��v"O����'[�	�$��r�H�,M佐r"Or%���?K�T�� W84L�8�"O��:�4	��!r�UyDx$�w"O�����t����@n�<@/�yI"Ox	'I�R'����- z�""O����a�f`����k�����"O���
+e��4�deâC>��"Od����O1	���j�� �MN�ȑ"OH�+B-�8-x5*U�и+̀r"O���CǶW�Q�U&��/4H�"O�-��̏�W�DI����6ܸI��"Ot��M�/���Q"}�ޕs7"OxH{$(J�'W u���t�څ�w"OMz���2wz5��L2��2�"O�]q�ӒO,�-���7b|Z��C"O��+%-T�lN�BE�yd1q"O^��G�9[������4Fl�چ"OJ����c7��A�n��(��D"Od�W�D��1�G�ޠ��j�"O�u;�m^4(��AT���\k�"O��ؓ�I)_k����M�a ��f"Oܠc�@U�?��cr,Mi����"O�h���Q3H3uk�9��K�"O��1�$�~�@�sf�K lN\��"OVaq5��R��0��|,��t"O�����A��q� ��<fX�h�"O�!0��cJ�8��;7HX@��"Orx�!	�,^�x�ѰN  �j"O@QkgM��c���D�6i,Y�"O���Ɵ�	�椸cW;N�D	 "Ot����M�`}ˣ���W���{�"ON�	�.P�2!2��J�����"O��%�ۼ8�t���J�&�@e"Oċ&�u��p	/�>%� "O��`��^.��
W.\�-5� [r"OtY�-ҏM5{�MG2J��9�"OvhR�Űy��0�w|-��"O�E{Q&q�T��w��59��"O��b�l�Pb@�q(�.%�uXq"O��ꠀX�1�2	�Dg�u�$}I�"OT�
���4d�"�A&4�xDQb"ObM�fJ��0�PČ(j��Dٷ"O$bG	I�S~���`ƻ:���"Op��XI� x2�J�s�� !"O�Y(�F�&+�,r6/ �\���z�"O6��h���@�qNB�P "O���R+�!�ƅ��c�8TD��0�"O~�fn��a0p�a�Í|3��`�"O����۹ r���nҔ~#ZxS5"O���B�<vKP�R��"2V�b�"O�pq��M(t��+\n�L: "O�9{cC�1���$
b_�@qB"O� ��� �8�6���!�T7��v"O��4 ߚG+.�2Aߖ[F��"O�=�S��U����v@@4���"O(��"H�y.r<���"]c
9c�"OD��B.��Q�n�h��!]Im��"O�#v���v�ؐa��F1�L�$"O*0�ש��U6<y�CҫE%�0�"Ov`QD�݈@�C$�����"O���W"��X��e�ƉE���pe"O�E��' G�ʤ��aK�� �e"O8@{�eʥ�����4N\�ZL�O��y�
��M��O?�	}�>�RE#ݲ�B���KJ+;b��7��g4�a22h�;�Nl�p�I���>���� @f�d�@�ٰ.
�d5�k$�i���"���8	kE�`jJM��!�j�*� ��gP+����� &J/�(ً�GD7f�ڗŁϦI��e�O����_y�'�����y�0 ��_N�P�d1�x�D�O��O.#?� ęS_��J�B-u>�dTL�k�'�Z7��O��?�oڽ#[Vl����.���ό�B�[��?DяB4 �H���?����?�t��p�$n�h�;��1()PP���SDp�� `�༒�B��,���f�G�h����F�X�p��v� ��f��/Py"���.8�9 -�lH��J�f%M��P��2�) ��	�R��|@����&�9Ї�s_� �A�b�a��|�f��c�,O���>�bhɛ#!r�ԗ\�^H!"��\�<�lP*�dD����@�x�RoC`3@7-�O8�O��	�O4˓J�Z�(�+��!PK3Q`�+aKN� 3ϓ�?�k& �B�"ф"�Fy�M�o���%`�����)��:3��@�e�"��"r���Vd�e� sD�5�Q(Pq�˓�h �� �j��!��������F�ē*��I�=�4d�J�@*6���7)8	���3D���'��Işp�?�Om�� o�p�2�)+}����']aR���Zep1� �*�\�������I��M�i�剄$�x ��4�?����ID8Cbr��a�UX�,�V΍	?Dī�)������ʟ�H�dI���<�C.�lXn�UN×+Q�M�]���A�=�WƼ	7�ɨ����q)ލcj������#^��X��,���[�)P/�����EW��+�
$L��c��)�O���PA�S�"P��[��hW嘦f7x,17�G �?I���T�xbC���`l���%s��h�����p>�ӳi��7-k�ޘ��ij��̳"�L�8�Ḱ�O�فPb�צ%�'�ӸB�p��ğm�2��` 	{�B�.�!(#$,{�ć�6� L�#A�:f�ڽ�AD¯#uz��D��O.k�q�����N����'<Gp��$�3Zp�C��R(�8(��s0$ cC�,���kl�PF�B�DT'F�����G	�����?9�����N맭�s������(W��:Sa��6�m{��Ot�D4�O���/(x.���	hH@#�ɋ�M�i��'�����0��N� sȥȵ![=_����ƍϟ��	l�СuJY̟P���� �	�u�'���Hg�H�p	/W \,���GJ�R�p�f��8d� H*s������L���d��x�d����(��� 2O�v���GP��C�Z��G_?�I�J��hx�p;�OL�(�B�>H��d�P��C��7_�X:U��O�nڜ�HO��	�m����2V<T2C�(-HQGy� 0�S�$�/�zؓA �?������'c�mZ��M�J>�'�N>iڴt1� @�?   d   Ĵ���	��Z��wI�+ʜ�cd�<��k٥���qe�H�4��6X8$<)�ih�6���#�t�`�ÞP�nѱ�%��>iD�oZ=�M�!�i����B5����OG�wo�[)Ն �eaB
��M���߆�O��#ߴ7��z�fU�_��d�!�^>*b�]�'���2#O�)q/O��2�����h�+O�=�v�.)��(u�u��n;YzRp�/	�){�f�M���M�j1A�4-��7����T*��[Z,��/s@�I��hΏD2���E���F�;\ �u�i��˓��I�1)�~?!p	U43���a��;?�̘��NL?�$Q����<yP�ܑ]Xb���W*B�4�>9:0 �T+:���`b��HS�;��hq��� v��	7y��aX �O����[���$X$�d5���W	�R�"jE�Ml"<��=�	:^a 1sAہ�d<�b�S��6���O�x����0��񥁂5`b��WB�cn2�Pw���O���O �Ym1�B@���VK���	�T�h��I'��O��]����@8x����+E2\}ExRGFT�'P�4�	4e�b)�P���q�&lk�$K�<�c��ht�	;r�'��|��g �4X�Ǫ^ ��(�'t��Fx��h�	��~� ��\��JX�t�z��@.��?!b���⃋=�,6�(}B��9k�$�����t�v��<�R�:�*V��0t�'@��Q�����R��xY�lk�IRp0D�ǰ3��ȵl��K=�ɠ�o\CB�b�D PG<�Q�\	�L���4�r�AU�f�TZ5�:D����)   �v��요�C) (jC�I-5�:��$͐%.~�Q�k �w>C�I[�|���u�\���;Z��B�	�aRDl�QF](C�*5�PJ�K�B�	*!wN �6�R[X�0թظ+�B�I�F��i�EQ
~$R�0�ɷ�lB�I�d��H���'H@(G�GJʖC��qt5ض��w�`H6 �7`�dC�	3��b�Ď%��Q�q`I�4(pb��QrJ�r��R�茰5�xCgL�/���ᦏ*z
<�����b��V�J�Y��t�`%�a�0hȖ�Rg�D�/A
0"���5���V�����E�e�:���#�U����S�V�r�Tl@W�|x�):3�ޯ7BE���#K���4'�>� -�p&]�v�[�&Z4J
!poq�ZLխn��P�J"h�����Uҟ\��/)dd���h�S�,O��PS����	a�V� ��!r��x��5�O���3Bڮv/�tw���1*%Y��x2�L5�?a����'�ħr��1eJ̾n���9�
�=(3*=�=Y����<�T/�v>"���@���Uؗ��U8�s���5U�J	��#tWr�#�/P���d�Or��D_�٘��~*|k0��"�!���<��!�S�L�)&�W�!��ݏVC����̀+WҮ��7���m!�$���Ԫ��0 �ݢ]!�Ӻ�ࠚq�C�z��+��Ͱ�!��#ж�H�-�r�L���
9!�䋌ac�5Rc���.Sԁj�-C�S1!�� 0�`�DAz>�j���jל]�"O:i�0&�6X��C�W�4�&���"ORaf^tռ���.h��aS"Oыp�72���	"�����1�q"O��I6��	z��3��2"O�-)aj �[s$7�:m��0"O\%�u�H��ZH���Ƨl�V��"O��j�?dM����H@����1"OB :��F�2P�1'L<�V`�t"Of���-r��j��J2U��rb"Ob$��A��7�v$��g�^�=)�"O���8 p�$�]�*�S�"O��S�>⸴(F��l<��"OJ̚���]P�@��A�'���"OH�ؠiٝ۠k�	�,-��XQ�"O�4J��:�J| ��\�����"O�I	� ^t���%�V�8�qJ�"O���Ċ o6��C�v�f0�"O� 0�鞖U����"�Y�J<�b"O��[��߁g�L�!�
}��"O�$�eo�E��%h��ݨ�ąsr"OޘQS���>��Hr��!3@`2S"O�\���	#8��X�=A��@�"O�}b�C�)p�br�5P.JYV"O�)��@�]�L�	 �ۤ5�����"O��r"�J�<���Ԣ8�� �@"O,�PgF49�=�$m�������"O�-��8P|���잽��Ի�"O��&EM5?l>��lǴA�00"Of�C&Mx� @*�
E�VT�U"O�1y��8y�n�ÇI\�b,�5"O�y`*ܲx($�0�n����	�"O�ԑ+�:b�$m���"�s""O^2��6G"�@�G��	�@"O^y�'/��J��0J�D���"O��t�/S����Hӎ>�8��"O>%�'���~�����͡F�2F"O��!vҎjN���cm
B%�a�Q"Oj���L�ț�!���Tq� "O>���>
�����P$	%�"OV ��E�*;���dL�a��d�`"O\�Q�Zv�>􀕢y[�	��"OB�����*R�E	��E��|I�"O�Й� �������� "\�$��"O�0�D.��-n$�2 �zYі"O�q#bD*j�X����$�>��"O����a�.'����S ^�S��]�V"OpS�E�$�� чB�py�Q"OJmx$��D1:�.էC���"O*�z�U%�f��q�	�+V�ɛ0"O$1�s�r�֤k�Kn���"O|u���3�L`� ǒ�q;���"O���兤��!���+V3���P"O(t[�� m�����}.H��"O|��'L)~a7�H�Z��a"O�qg��࣏#tt�6d�9�y��>��c�l��9PMr�����y�ʏR� ���˞�.ʹ؃�h#�y������D�,�6]a�J�5�y�,�gt�27!Z� ��p�Ö�y"��u<$+2�G�����3��y�Kмm2l�(E.n<�A���yB�#s���3V�'~+8�ZV���yh�V�t(��I�y)HH������y
� �qR�KT-� 	�Ǉ��v. �"Ova�r�@?Vb<�4-ӯ	8��6"O|9�$@)zj`A��K��L}j���"O$ ��ڢR��L�3���Rd�m��"O]1w������]2��8T"O$9k$H�@E�sdFγ\uh� S"O�y;e��0Oov#���N�H�"O�%ʀ�$@V�;&��88=
c"O�yX����L���շ8�}!�$�b����k͇_S����:-W!�D�9x��1 �K><��[�J�~M!�=wPف	�~3�da$e �}�!��M�FJ�UZ���')�فtd]:�!�$�<a'�0�e��w�`���{8!�ā
b��1�f�94 m��-3�!�D�*H� �q�R;\Ձ�BT�4�!�D�3+nH�8P�ڼ`�N�X5/M�_�!�ރH^���*$?��,`WNM$P�!�Dg�nܻ0���:hl!HH�P�!�Ğ�w�.��'&>²P:Vh��u�!�$:>��u�T*�Ҁ��-Y�!�$ݺU{��CBI�}
ޭ��G���!�4��Y�GM��R�L`���6�!�Ĉ"Q�r����X�0Ly6�յ"�!�W86[Bȣwf}����[�)�!���/2�p��,�$r�=M˷3�!�?l	8��R����Te�|�!��.H�B\��ҝ2�B�9�CǗ|�!��V��J�I�&�3$l۶�ҫ4f!�d�;S����҉��V��[3,��b!�dā5�:IP2�Jl���ٜ/�!�$�#yn�#�mَ4��0 �i�x���d�P���H���9SQ��#��	:�y�j@�3���#g�"���Em��yr����ǫ ln|�6��,�y2��3��!�&��L2S
���y�j_���I�o�� @&�УG-�y�"I��*� �u�.%��+/�y�Ūv���`G+�l%��ʢ���yR��2
_ځZFҏi��Ű��[�<�!KK'UnlP��M��!�8�kz�<91�D�	�:}����*J�uL�p�<9$,�J#�%B��éB%<��n�r�<��g� 56�����(\����w�r�<у��'�`�nJ�f�m#�d��y�+�����0A=]*��t���y��ʅ
�(w�R�8 |z��Ť�yb�ɣ5��@p�J�|��]`��@��y
��̓FZ<oH�T
��y҅�[�݂�J��N^ز�׮�yb�-d7*�zf�M$P-�r�R'�Py⤇,G��%��-%p5��S`�<QBoy�|U񤨃s��jT�ET�<1���2�ro�
<q�KP�<Ad��[�H�C�����`��]G�<Q3�S/s�`3f�K*�n�c���M�<��Ӕb�ؤJb��K����寁K�<����J".Ti���B�@�c�bJE�<�g� 37a�=&�R>�hiC`gx�<�V)Ã7��r���^�F5⩔L�<!��Heb����fz"A %�H�<�Ό;~g��H�b��~�!H���C�<���X�bO"�P�m]0R�:�ȄCIX�<I,�e�n0�')�+1}�iȐ��z�<� �@11jΝO��Hӊbz�y�"O,dbŠ��7�h���F^T^��"Or9��G�x �4����B^LAT"OdX4��(e��PTfţ���"O8Ipք���2f�'D�2�b�"O�E�eM(U+|t�ʂ�&��U��"OTpa�J\���%[ 	����"O�l�gF�'���a[�B���S"O,DAqGϹ3S�ȫ���.m�Req�"O�����E",1�u&��-�멋q�<�&��=F7<DJ�.�V�(��w�Bw�<��CO�O#�I(�a�|Ą�H�>m���һ?P^�y�3?��ȓP��Jui�5�Ĥ��*ߕg�84��yD���eO*O�$��C�D��ȓ>�<�� ^|AJ�.��R8�p�ȓ����c�"B����	�P���ȓ$LpP�@���؁�k"Y���ȓN���`uk��Fy�4�����9�a��Hq:��d�ƞS�� �ȓN��ŨB#�CL\p���Ʋ|�0�ȓ��yec�9+����!�
�xc�=��*��H�c)�:�|���D�Ǯ��ȓO�����@jΰ�A ��DS�d�ȓbX���僕Y7�5	1nO
/����xLM#hK��Q��(�\.�\��E��A�& F�b�da�g�L���ȓ�f�ba�
�gg��T��-� �ȓ;�֠9�.W���܀@K_�^�jU��-"�\�/�;0S�t���% n 5��5t��h��I�_�N�iU�5%�q�ȓJ�YP1m�#Vr�A����3\�ҩ����tcd@�'�Hp9&d�3;;�H�ȓT�����D�R���F-a��\��)���br��;3 i�ŊX,$�Ȇȓ!���d'I�^�d؀�E�IV�ȓl ]��'�<����ɜ�>���P��q��jd����N �D�ȓt0�]+�I�6`;�c��8<�ȓ9z|�R�L�U����iœw�����[(���5`G6k�L�r���g ؉�ȓ4�x՘��3>�Z�S�F��?����t��E��#�Su�A�o�>G�Ե�ȓ"�{�f�*�|
c@Y=1��L$������e��dR�7 )�ȓkI�]5g!x��Y�h�%�d��ȓ;	`�X�Ι)�<���P
o{z���{�t$��V�+n��g
BU�B��`J��W%��U�h	<:(����d�zC$Z�^�zbκp�:�ȓJ�\-p��6E��NI�s����ȓ_LX*��ڊ+odБ#e�2H��X�ȓ<�B�0v�)ՠMAb
2jv-�ȓt����*ӭ5M,0Q��M,Z���ȓ�`�f� �h�ꌫ1��i��@ж%?m�iK�iQ"8*p���$}��������"KU.x��LW����'΄	bJPAB��+�Hą�B�`��T�U&R�d}��E y~hp�ȓ	8����kz \8�d��\���B� W��h��<����?�&��K`�LI�N�r�$ȓe?{���ȓ&Y���)cK��¢5w���[�e�58���3��ƙl*Qr�����'C
l(�M)�C#s�$���S�? ��i��p��`ӺO�L�P�"OR�
a�Ңwȼl�����"O=�ɇ�J>�M�q��j����"O�Hq&h�q�$��r1�`ZS"OB\�c�(5~ܑ��[?e�HPa�"O�X���L/0�a�h�\%��e"O�л�f�_4\�s���u�q�D"O1��,�#a �P��$���1�"Ob��S*��%3ء0OʱP��0ʇ"O0a�G��e��<
�o�S���f"O�A��LG&Dl,���.Ǎ7�2�p�"O��c�d��G@�! "�Ȥ��T�4"O^	x���z�A�BZz�z$"O�ڀ*��L���rD�UI�"O:�BU�	�Z��`�ʔ�&KV�St"O��Ӵ�{��ͩ0)M�(�U�"O�q�.C
EƐa҆�"a{�� "O&Y�cFȂd{���1�J;z���"O�(����')'�	��>O�M��"Or!����� � ��I�+mY40��"O�m�T.ˎWю��u�]�pP�D"O�Ux�%��h ���ϻ5T�M+R"O����ˎu�� j-E�D�T���"O��K���{�j��Ti.I�H��"OxTR3�¹!����v�� *��]Jf"O�1��)�)Ja���%�~�f"O���&m�DoTu���"}O����"O���S�M�'��9�V��"q"OB ��QV.r��Ph�x-�K�"O��vG��n����,,�H�#F"O�	��I�*KT"�2�eL�(�^�2"O�ٺ�˸H?x��E%T�'��8�"O��H7�ݜ6>M+��dV�,�"Od���E�"+�V	b��Z9M��Y��"O4�2ရF�~�Z �ɀZ��A��"O���FNd`�!�՜o�0��"OT��o]7lA�xXv�6O¨�!"O^��e4+봔���T Fl�@�"O(�֌�4?��2ᆀ�hk��8c"O��b�n�:l|�}��L$�\��F"O"L��@l"�Kg��e�"O�!�+�1FTz�kt��/zbT��"O"}�D�&r�Niڣ��3[��	�"O�0*�����*���O(<��"O���g(��.�.�p��3d�ؔk�"O�X��w�YtO�)P5iQ�"O�|ti;[)�ŻA�C�v�,#E"O����a��[X��F�-��	�"O�B��d�`�<莀a�"Oԭ��oD�x�bUXq�X Qz�i�%"On���9s��0�5�H5s��*�"O���G�Ȼo��l��D ;���s"O� !���c�E��E�Q���Sw"O�P���zŀd��"&���"O���A�N(n�4��B�&)u��"O���R�� K�6a��}`�CF"O��d�[pptE�dΊ.6_�X@ "O2�8'��=i��%�N&m���cb"O2�9W���0�Ь!#Y�ҽy#"O&�`���Iq�����:ۤ��"O��C�놓Rɪq8F
�/4�:��"O\Rp��;l;,uiU�	?��s�"OUrM\:<��C�" 	�"OƐ�#&\h�Q�77���"O� ��c +���80��:4"O�l���m�����
�+֤��"O��S�7Ξ�!�h�@�!�"O�"�BF=>Dp������D���"O"@x��C?3�Y�QN��%�0�y�o��s��� ��r$�p2M�'�y��Du���u�ՙx�����CT��yr$���,����BX1�i��y�Ac�"�Y�I�	݄�h�A]��y"��#S|�����Q�\Jŋ�y̕{ʬ!E�Q'~�� �E�yr@�&i�1�CEZ�}+9p%.W��y"H��.y��ʅ�Vq�Z��4�%�yBK��h1@#E{�`\R�g���yRJ^$#v���g��	�	=c�B�9BFʕ�D��Y���2Słe�^B�*f�ਃ#	I� ���Q��>N�4B�Ʉ!�r]���C��#��){�C�/7�cwg�rl0�#i�_h�C�ɝEKj�A�� ��q"�ʇU0�C�ɡ"�J�#�JՔQ�eS5�I�r	|B�ɀ@����p�D�6�� '�� p�pB��:s�1S�'Q�j��p�NN�4"8B�I7�rdIUƒ��%"AO�H_�C�IDyx�����,P�珟;C�C�ɟ.�~�26KC���L0G)M	?̐C�1dE"�@]l���$�$r�bB�ɂW�6�h�f٪R̀���ٌ�yr���Vz*�)��X�z	��ڦ�y�iϨV�ZuJD�0Qt^,c���y�C��2�;s��u#�tJ�_'�y��W�|��裮T�f�̑�#F>�y��@.$����G8c[��"��7�y�̊%S�9�'n,n����*�-�yr�ս8`��+
�b�J�S��yRƬc���`ee�t#�Z��ybI@�tĝ��
E00�.-��oN��yrL���Df (\�a�@���y2@^�w���'<��ɡH¾�y��#by�-P5�Y� 9���4�y���*b�
��YtD���G�BC�	<&cr�#�Q/��#i�{�fB�ɕe�>�i��+z�y#�G �C�IE{��1u�9�t��g̨e�X���U(��ٕ-�R��-� �H�Is�4�W�7D��P�#ML� `���"�8�eN#�E����.��O�P�Y��S�U:�� ΍��=�
�'nK���H s���=H��bȟX��w��؁0Qy���Z�|ie����K�6>.pB�	�E���qa]���	���J�9�N˓5�vM #H�k���9	ÓoJr��Fʪx;�����3_X����+GN�}c�㋲�=b�!��$�&)��[+-J0a�F�(��I�r��㗀GMk�bEˑ=H�<YԋT�2� ᓈW$��`I|z*Y�3���%ڛ<
�(A�h�L�<A
!1��8c"��I��L�'d ��E�f��� �؄8B`�D��'�:Mۗ�'xg�-���W�}.4�3	�'���+��_��V�����2���Y��˟B:�d��eU�[�p8)�"K������/gآ�uDF�;����G�(vp�{�'ʞ�Ԉ`�'Xz��֥V���ڽy[l҂�׈-�j�'� �I�l��a�l���)O=xɑ��D�<8 ޥq����X���G����v"��"O�|�
ق4"�2�y��Ҧ.c�<�4k�y��I�q����Ìq��D	#	�%:\����^	�f�����
SX0Hl�;?:!��ע"rś�*̉a� e"&J�%X�~,(&�iR�;5D�DD(� c�~Fz
�  �3���#��{��N3$�s�'+�52GI��pw �1���un��� ���N� ��g�'ߺ�X�.LO�a~r�;,h� @S�i�^��B�	��O=#6�J;6��q�.�tS��@I?�k���&TS��7a݂<9$1D�@�v���R��|{']#����4-W
�(��ޗ7r�TR4J˸)[ #~��i�*� k��A;3i��C~Q�ȓ1l� �0,
�0Є�
$�Vdq����'C��
E� rh�C�{F{��2�j��pʑ�}BW�_��p>q�M�>�h��DX�b��:7u6�8%��Ґd�B�X���\D���U눼y�ʌ����	[x�D{�+1*�~�8&g��r#1��qaeɨi���y�(E��ȼѧ"O$Q�B��y��)���/ .>%@6�'��6�J%3���ȵ<E�D`C*��0cu
Y!J����`?	^!򤈻3�@�*ܕ>0ī��KZS�k�`9�S����<1f�U�M���*P��h"��T��L3b�����0��#%�t�z`J1@�ІȓH�P���aH��<�C���^�p��K��؇��h�CF�VKz���yk �6j7��"s$[�'����ȓq�މ���ˇ%��!�����<��h꽲�
�6~�yJ0jX=<\`���w6�t2È��Ť͒�CY�hq$u�ȓ36
�#�̩H��dڄ
ev�������c	��L�w��W��d��D?�H:d-C,��)x��P�q����+��ɺ�'��VA*�a@oM;Ģ���H��q酤R Dh�p5����ȓ�����ڳI����El��+J���ȓ��0�F��-D �@���J�l�<ya�O>��i�JÁ
�Д��k�<����Uk&h1�$�+�0!����k�<���_�D͌Mk�؄X���%?T���7�It��řS�A-#	ı 4D���D_%!.�`�&d��1܂�KA!7D�Ta�C�g���P�$./~$�f5D��R�B�(�� i��N2�
����5D�b��2 L��`M>x���$O3D�h`+0eXx9P%�������-D�@���ʠz����ǐEnm�Ԅ,D��i��޺Yr/F��>��L=D�@Y2�7S��H�oE�-_���<D�DhեX�Z5ʩ� ʁ�*��K��:D�� $O�F���D��q���W�,D��3V��Sm�u�kN.L�̉��%+D�쁂�H��	��]����ժ-D����@�F���ڡӆ��B *D�,ې�ޫTT�Se͟�R���,D��#Įώ4��ACKM�>�$l5D��ӈD6�\���a�<9 �N3D�hh�3V2����
?k�8�Z�!�D�5T4ҏZ�Z�<���O�s�!�d�#��PI^()��q��.0�!�$,�tb���g�N�����(Q=!��P�ϸ[��	<5f�ӳ��&9!�ՐC����*%�h�a�QE!�$�K�Irץʛ1(�'�!�^�BB̹�s��!���q���{�!�Ăv2p�u�� 
l"��U.ߒQ�!�d�$P ���Ǭ͞e�@A�'Ch�!�D����vΜ m�L���`΅u�!�DZA���*ߟDäA6�ҥ3�!�DS:?9c���&87<���!	�!�dS�&	���D�F���E�����H�!�Dє,t}0��!E�8\���R<I�!�� ��;b�˭?wiA0�_E6�P��"O
4(ЉW�Ov�4�Q�L41+�"O�Ր��MLE9#Ȟ�jT9a`W)xZD!�`Y��l9�dE=<OBab���5"fH��L؋^H�Ÿ&"Oڜ���%�0�`�h�Y���"O�|�P�
)���K�%}R�|�"Or=�G���J�F�ށ�"kU"OHi�%�Ñ;��Mj��E3��8p"O�a�C N-\NA��C�)�%"Ona!�?<�|$	�엿
��Y��"O����	�i�a�L �~(9@�"O�� K�;l����EG�s����"O,�"��M��Bݘ�5��L�g"O<�3e�[-W���� L�
�h4#�"OE#�cE�:r�;A�үU��JA"O�A��
t��m�7�ϳˤ@K'"O�Q����x�j\"��vY��+5"Ov��e��O��Y+��˘U�u"O�����M"gE�M
@LM�HB@�"O�T;D��&n� TQ3�
2-B����"O@x�@A;9�R�%Ǜ2k8xP!�"Oj���G��x��j�%Τ9��(r�"O���Q K�,%ہC�W�2"O��a�C֙#|�0��L*�"O+�g�<�=�Զ�+$lzC��  p����2~�!Ѕ�[�B� J�Z�Cf`B13H��� �IS`C�ɁDP>���X���v㟵4�B䉦*>�=:sB7s|���s'�a�B�	�0 yA��8WgxU���Q/�B�IX�t���C$�
8�tfPvs"B�	�Az�$�V��C����v? dB䉋fb��T�71�������Y�C䉜nJ��Ё7��XG㜈|�tC�ɥ0�b��b����(�f4p��C��$h&�9u�B�J
 )���I�MK�C�ɻ]K���H�A��ș�뇄nd�C�I73>�}ʠ�J�x�ZLK ,��>:TC䉁#�.蘲"�[v��q�BzgfB�	2+�@ZA�̯n�%�$�<,iLB䉹R7F]� ᪝�g�N.�C�I�yH��Xb��50�x�;Ң� �C�	"�X��A-G�@�X����DW�C�	�x.��FiA�'����W<j��C�	%g�rBe��{1�	�?}O�C�	OE@Hb��`���r�"�C�	6C+���	�L��@���ç{��B�	�<#Ԉ+`g��|��@��땑1�B��+���q��;~�б��Fo��B�	)�NP�S���yṳ0�	��x�B䉯Qj��9%,�4aɆm+�gˮm��C�*�,ak�Y��R��c�Ȃ��C�I�/"���I��&D��F.��]�C�I�e0�Cq뚺O(Q#��F�n�C�I�kf�}ْh	�vLmiE�H?C��2;=�	Z#o��VJlTp'�ō(�B�/J
h���"J�N�R �,F&�C�ɦU��A��� X�8��#�ߠb��C�	&Q5r�"­�9�p���L?e�C�ɬoAj��d!הh����)A��C�I0ς�т�ã�,�JT��	��C�I5Lʀ�׭ԪJX1��^"#6B�	NiÀ�ʕ[J%1GJ��J��C��I��,['&��?��ئh%�rC�)� ��jO
&��j3h�m��H�"O���ւ�2: IG'��e��L9�"O$=��L��v�P��,7b�XC"O(�`�\?���&��_�� �5"O(="E
P�� Jޅb�<ٳ�"O|���NҴ=��H
'�Ź=�k�"Ot� �))wUh�Ȑy�$<CQ"Oи�����L���B
����
"OXp��c\�`��0�N��z��l҃"O:Qx!/:/���RN��`;�x�G"Onx�`�X�t�kq�4o d �"O�5�5�G�j�n��f�\�<�T�w"O��"�,E:Un�tq2J�&K	ri�"O�Q�%�W�J��!i��[<L� u�"Oֈ��.!������%:$4���"OF �
�R�Uѕ-:�$��"OJ��T�0f�#�Thpt"O� X@CQ�~~Xy���\��K"OZ���덢B�^�Q!�)_? �yS"OD`��,�
G.�Y�	c n��B"OXL��I0*���ƀ���i��"O�PJ�E��n�Ջ�+С��I�"O�L�وu���:���!���g"O8,Jg���L���� hȖ ��:G"O���Ϟ(�DqWlA,�F���"O(X1�'T�<؁g-��.Ę�"O�����q(>ay�J:p�\��r"O޽�r/V�*�L��v�J�[0Jt�e"O*THf��f���B���62�az"OЁy��0J��b�ɱb��"O"-H��l�����ą/��8� "O�9�C&܊`� $	��Q"<��q"O�����%;Y	� Q<v&<c�"O)���˅c@=�g`�4\:�L�"O�e�gA�<��XRr
~'�u"On$ �H��ph�ٵ���nF֨z`"O^0��FC�$����7�L9���3�"O�=P�ƍ��Ҩ��m@�~�>LY`"O�$���+'�j�h��{��TYb"Ot��(M�o��E{�;`�:�{�"Of��g*N�f�0�!5��D�0��"Oҵ��%;r)���.|�I�"O0G�֛ d��q&_�Ch���"Ob������Y&�娧%�`���V"O�3�܄�H|3u��Km�X��"Oԩ�r�["!X����-qe���f"O��S���w�x��UۘOVX�1T"O��J/EZ��QP�K1GvJ1��"O����3f�DdI6NǶx�N5�"O��s�Ҭd0�҇l�Yg���"O��X"n�~�DD,��k\,kp"O�,�I�odȲ�H(]pށ�"OT��ai�c��F�m�Ƹ*d�$D���S���n�Ҳ	��*��k!D�XZt � ֌�"��Z�v��t˳+$D�{�)َ{a�A�%%�حr��!D�l0��#fB�)w��4A���2c�1D��削^[�	(vE�>�X�{!�=D�4r��=�\@b6b 7M 4��(D�tI��%E&��J��^����%D��"��9-���+B���j�ܡ�3�&D���,:*L;1�ځD@y��(D��y"O,1J�=����j(��O*D��P�/f9<9Tpʁ�2Cax��)� �T�D���f�d$��i����$�"O�L�C�"��s���7dJ���"O@�H��9*�5*�/��$�3�y��4s� �u��i4�}"�A��y��S�coT1�gȝk����ȃ�yRn:^�ā�VL�pEd� 1���y2d��i]�8�ܻ27 ]��K��y�.�x~����
�.�^��WO#�yi�;c�M�����
~@hb���y⍈�_�֜kJO�nR0�(��yr��!�lס�"RQPR��yr.R)��yh�
�}bt��+�y�o3wE�T����m�4 �A�y��Θ"��M@�Ԅ65���,��yr�Y[��<c��ǎ,����^�y��q��0Gˇ)Wy��80�E��y�V'p�ܫ6���R'. �bH���y"������;�ֈ���[���'O0����t��D	H�	�X�'�`7$P�%N:l��C�d�ț�'��1A�#���J �Nrɘ�a�'T� KQ"A#R�չ��FB

�
�'C�%S�!� �xذ���r���b	�'��Dsn�8b�X\���6W�f�#	�'�LYۖ�:ix��;� S�S���'*\��G!�wi,ջ��6PC(�Z�'�*<�˛�Z��x{��ݞ��0x�'�$�Q��L	E��vOE����R�'/�y�BAX�z���*�@��;�1K�'`x��T,�|qZu�ʿ!BP-[�'%|廅/��0i<�����FTh�'*�%�S&	��+��K��n��'M��i߾<f��e�8;��ܠ�'�&�K�$�e�.�9��Z� �U��'Z�Ũq�ī n�*�d�T���'���QN�w�ĭs��H!Rݑ�'Į��v�Nu7�1��l�H�'!j�Y�	�w�`I�����&gj��'�x�
��D�1�2Y�'˖n���
�'�2�hď�!,>X8rm�EI�#
�'~���f��9^xq��hD1@��
�'A��4���U�3�|ܫ�'�8Iؗiʋ#� ��m��Yt��R�'5f�ȗ�W�'�� 	s&ĘS"�}2�'�p�aqK7i��y�N�7Şp��'/��P���)�\ݡ���0+[���'*>,���[�Bg�x
�I�7w����'(*i��'�;K r�0`�^�.�x�q�'� X�/ްf��qV-4��'��"q�,3.�,�%��-��R�'4�	k�g;)f<y��0#bt�i�'�����$���S��Z�1�'H�����#_�Z#e�@�����'��xtϑ&k#�kRmҌf�5��'X�iä�Drp�YJ̷K7�
�'�Zm�RK�'?N��PQ�H�Ze
	�'~b�YW�X4t�X�b�:BT���'�l�j��K�AGp ����:1
D9
�'��A�W��%Wڐ#%�V�0$V���'OL���
|���ȓDۍ5����'�:I�!�����F�|��\�'��]:LˤH�y�Ӏҟa�0�
�'!: �E�'hf0U8#a
uk(PI
�'c}"�8�8�y�J�rF��	��� .L�!��]A䀠LX�~ό��"OL��peFb%4�ru�7.�ֱI�"OΈ�BFHZ����J�HV��kC"O�,� ⋌'jh��I�r�d�%"O~�A�Ǟ�9(]��һab4���"O�e��!_��s���\m��IW"O�pŦĆW���cq�Y8{[�0��"O>娲�֦0�yf�=절�s"O(��E����2��Է=�9���ݎc��{��(%��P�Ĉ��y2���_��)T@F�NPE��D���y��D�0g�ATA#�Z\��̎�y�O 8\*�XAꙪ"�z�O��y�h�9*"�# ��2`�NԨ ɩ�y�%É`B��2i��qх(��yb.�?i'F���� c�N`i�e�	�y�cԴ������A�XH�1!�BC��yR�Ȧq���C�~��ڣ�F=�yRGE�3sݢѥEJӞ5SA���y��|P�����?�Z�c�'��y�BA�<��Aˀ"��>tZ����M��y�
B��a%kҨj�F=3�L���y��uz�	y�GYS�r�JR�Y��y�B�2d��! �[�Fq����%�y���l�r(���!f2��Qd�?�y�eD�(��E��@.08}�#-Խ�yr�C0/J@�C#N�20�Re@�y���j��l�$�åx�F�*q���yb��,�h�i"s��J%���y*ߤ�4�妀�d"<���̧�yB���oxTD ��=S<�Z�+��y���0S<�CV��x���O@��y����HX`�L�n�n9I왗�yV;N���PbG�;4�������y2��w�|��X�d��E�Teϰ�yR� }?|�2��(f�<��,�y���0Q�6l�$A#3&����y#��v�Řd�(t�[����y2�B3G�Н(�8~�&�����8�y���1��<�S
M� ڢR왪�y"��V�h���b״$1��dZ)�yAR�U"�ȋr�˙o�@�(ˋ=�y)O�DI|����T�p�"\�����y�%��*(r�I��3��2�����y�Ƙ �F�	�ɇ8w֔"��4�yb�=X9�wGE,8�F�h�Ο�y�%�&�A���@��t�0�n8�y�͙�<6�����- ��-�E�%�y��5L����T�V��JU��y�hĸ+ �As�ñx��0���T$�yBdܐH��	.��w9� �w�׃�y���$a`ѱ��ܱӰ�27C!�y�H/]<���D�l>�#W�V�y �l�G��y���x�I���y�.��<d��8\��قuk��yb��l8PÐ� 2��W��y�fF�}��Bé�.����B����y�-Q�<!��`	N�j�q�a��y�ER.a�%��/@6vJe�a ۀ�yR��;L-z|p���3��!5�y���
/޶�ꡡ�W7b��`/��y	ZB ��IIF�1J�	Q�yҬ�Q��A�����v��` )P��y�.��SR���$�ߌp���2$f�:�y
� ���ECmR``�0�>/a��"OZ��,M�T8z�E�%�B�
P"ObE���	v{��x�F��B�yȐ"O6`��/� 4����\@�"O
��t �YgT<(�* �p�Q"OT]bqM[�l����x��0�B"Onٙ�ܢx�P���D�>}��Ő"O�01�O1G��[&��In�I��"O T����1B0)�%�S�X:EC�"O�����8c�C��{*�1�"O��ZG��|�,1)f��5*��j�"Ot:��	g��,@��Q)8��2"O�D�'��ؤљ%�_22���t"O����<}����0m�'yR���"O��@�L_ Um�Bc�5c\v9k�"O� �4�܋f
�E��f�،��"O��F��L��SG�K"0��D��"O������g��%���:G��8��"Ob�PA��N��b/�[ɂTqD"O��􈈵�젃�m]����a"OZ�r��-^�d��b���v��c"O����A�1��{��?�P0u"O�hP��	{�9�@B�W@ޠYU"O>|9f��� i4��#6� :C"O ��Lh��y���#|��� 7"O������NϜ$�D.ޗN�ĥ�V"O�u�4"�6��-��,�)�ƴb�"O��⧎�(��e�f�Zs�@�"O�T�c�#}��(���6���@""OT�"΁ ;�M��jɛ�X�)�"O*@�G��<b'( �S�6�iD"O�Qiu��(x�"���_	(���"O���%���f�,Qd�U��q"OfA��3	F��s�aL� ��8:"Oؐ�K��F9×m͚[ङ�"O�!�%��9uZ�`��iQ��v"O6�� �.1ȁ��*���"O�b��m��Ð&� ?�VD�R"O�1֍Q.��Yh�$C6:
�q+�"O��`V���c�E�6�x���"O��27B��Lг���j��5��"O~X*$j�e�*=�׭��L����"Oeʢ��3c�\���8"�����'�N�� b�KsPt�U�r�D���'�V�ɁHʮ|-t<��Z(5 ����'�0�o :
zdt���E�+���'g*�J�΍%)pڙ*��Ml���'�FXQ�J'8���2V�F�dN�=k
�'�v��.��D�&�K�x� 
�'�`H�B�;XU\QІ�Ov��i�
�'R���Alͷa:n��@b\�g3@;�'�j����Ԣ<G|�	p�ϴ`.P��'Qޝ	`���B�
��GL�_�V���'4<�l�[@ҍ�ck��m����'9(�"�G��:���"�z�(�	�'IZ娷�܁y:PI�Í.(|ʈ� <O ����V���胄�%�}(A"O�����9D:����G>%��zw"O�1z��?B6d8p��b��-�4"O6��@��%rʶX�t�� UvZ�ZD"O��E��2K�B�iR�q��"O|���_�t4�e�6TLE`�'g:0��JO����0����p��',҅��NG��^0�!����Y��� V̱�L�N�f��"c�������"O���¸^*d���J1 �����"OڹK���$m8�bK0x��᪡"O�T� �'�<�aKW=[َ帀"O �kb�̒q%v)Hd�W�쌴Q"O�m�����A��[%	�l��v"O`4��\�LTd� ���ZD�"O��@ִׄ �9P������B�M�<��³&"��W�w� ��¦G�<��U<#|�)4�U�F�@Y@#�YA�<I�d�%0QI���x�$��2J@�<�5Ł�<��qJQ*m��p1��z�<)tM�7��\0��&>\�x���_�<1��+^I��2�F!8K`���e�\�<9���xUʵn�6�^����M�<�׬-�|0�%fX����eJ�<1r'- fb�UnQ̅!�.�^�<�`�ְ+u&��UD� ��t�)�X�<��2E�����ʛ4Q��:�`EK�<9�CH2���h���n�t�rLP�<y���:�Ȧ	$U�x���g�<��C=�:Xy�+\p� f��b�<AqIɻ~|���Η�<�^͐�VW�<��	M�Y~�J��L�\ًF�I�<�u�Y33>�@�G�B�6j~�0�JQ{�<�%i�YO"�ѓ��I>��`_�<a��܆Q��0҂ ��.X�ЄK]�<Ib�Z�X=� �0&K;jG={���\�<J	0��!u�41�0d�d��d�<�5.�5; ѶE��z	�p��A�c�<�Bj�}����-��y�2%"֋�W�<!b.Խ ~�8h���A\����V�<Q�Ȍ ҜP�&$�P�YP��~�<Y7Y2���ba�+}���q��C�<1��ɪ�vm�pDīL��0���}�<qQ��
���£.�9)M�@I�v�<�&�I���)Ce��{6��"�Hr�<��=$����#�m3���Y�<��.�%$�<8���5&\�D�3�U�<I���R X�K�杜V�l�G�O�<aǅ�	#`<���F� �h��JOG�<q��7(�dy��Ww�4q3�d
h�<96�шY�^ ����4Q���#SF�b�<�	[9(��8;�◇Ec����A5D����H��G�$4�'Z�0����0D�d��J����6|'B}C@M.D�<�`i�YN���O�&	1s�*D�\�7�B-���V@��+%�<���%D���"m��e!(���*L2Z0�d+��/D�h"�i���T�,�,ʑ&0D�����Iu9��ÇBіi�s((D��u#�Au2Il�<BA�}5&t�<!�ĉ	 ��3�6��$�D�ȓ���R���@��k�"Ǝx��܆ȓ0����#R��̕�֢��d&��ȓ*L(��C��)C�4e�&Q)�=�ȓ5�Zez#�P(;�"T8��G���p�ȓK5ڕ���ÞBS��B�� gBR��@�3C�V�lJ>�4��eo�X��lV�%`�8O��q���;�͇� �z�� L��9��I��ȓ@��XA��P:J)bQ�\�D�2x��qha2rg�#��R��ǊM��>�n�@�e�7��,���P ��х�S�? R�xu��?0ܐY�i��X ttj"OV�qw�F?u�t<�T�޸y8���"O<ɓ�Ξ�J�25��ņ�'� 7"O4A�#��SDb����(p���$"Oi��D���De'~���ӳ"O��uH�r�����f�%7����"O4@e��2IfX�!Š�>�:=R�"O ���jN?hl�@XC������"OlHb"�]/c�V�3�G�,?��a�"O�8)�͠q r�P�K3.R]1"ODdC��ڠ�=�c�MM��;���O��B`�M��O?�IT��!��[�'��`҇�a^H�*Q�k�`)y#�A>D��8�b�E�`��>����ްh5��)E�
݈q�G���D�i��衦�ظBF1�	L?B��p�ҪOa�c?�؜&ٶ�Q�őF5�U2ԯˏ�b6M[�6���'����?�D�ܴ�]:��J}Q�U�7CA�
��?����	3oX�ip�(ˤ})F�Y$�F�<�5�i��6�!�����m\7(t�i� <W�ƽjTD�!��IZ��Z�4��<Qǫ� _@ce�[�Ȑ�R��Aӄ��q��2a�r�������ޱS��O^��Fx��˨C96�����r���`'���R(�Ls�%]62c&�:ǎD��8X��t5h@/�`�:�zuj%�^!(�ZT��jzha�c�'U6��u�'��7/��Y���	T}H5A��Y��ƯE�**��(�y�&~�H�*�씂-�����G��! �n3�M#-O�d�o�J���<�PE��u���2���4��<��b��B�$�20�ϭ��<��B��$�s�K=E(�,���GޮP� IՂr\�T���R��p�9+'�h������&�bQ�*�=F;X��3Aށ~#le;c U��d����=}䉉t��$#�^�dӄ}�QL�*t&tS0��	�,�`IX��MS����$�O��ʧd{h�āމi���:�`��6P�T��3>̒&��7��RW�
�]�����N���mj�Z˓b#d�T�i���'��ӡ�^EHQ�иo�
!Q�ힹ"�:�'K�?y���?��l9�M�aeԩU�ޥA.�=I<ڱ�'h�d؈႖�P�����n�vFz�F].LW,�yrmL�uj��c
*]T�AK�E
"�@��F(["ym^ͩS��f��"=�w�̟L�	�M�����鉿Ж��d&)� ԰��,X�x�	`�S��?9��2Zz���7,cH�QK�#�ў�&���42[��C
;����K6{Ո�{嵭gG<��435��`�_�ԕ'����O�'#�t�K vʼP���%FI�1���q���r��_�h�9�\=Wh�r����Ͽ�tON noȄ�7�����`�˙񦅰3��@�j�iEF&̤�2�n��7� (��\c�"$lG2RSś�,R	]��5޴C����IП�4�?Q���i���	��z���T'�,� ���',��d%ғD�Dpӆ	k�� ϐ���Fy2&hӘ�l�~��")�ծ;Q<�l�,Ghh��aPZs��'�rOQ[�����'5��'��a�~*�47�Ą9Ў�V�̌��Y�@'"M; �@�9��mx�n�y�\%I&�/7����Q]�'����kӍ�D�Rѫ�:.���8�JvӒ�[ /_Zn�m[�Z')��O��`S�y�>p�B��ă4:~���lP�T�H�$E�;@����O�0J���	�'�����A�	���J	��QÌ�8,O�����";�K����-�P�1�h��Mc%�i��'����O��'��&�O |  ��   4  �  0  %  f*  �5  ?A  {L  �V  �_  Zi  Yr  �x  �~  M�  ��  ӑ  �  `�  ֤  :�  ��  �  !�  d�  ��  ��  (�  ��  ��  ��  ��  ��  < �
 � X �! ,( o. �/  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h����z�"��h���J���y�Α� &�n@y#Ov݃�*J?N�Z��5
	�~Rdd�Dٌ��s�����&@X�fD?C(rap��'>qO�Uc �G7x�ֹ��,�TI�"O���#^4�H��Ǣ�X�#"�$8��?u�	�͈e��i�p,�`�3�tq ��#D���B�]�Tjh@�$�a�)y�,���>)�7#�)1i�$�6&f����$�>D�a+�YQ���ō�yɄ�Q�'lO�� ��FiL�ZP�N7/j��h D�01u�M5*��JA��H7���� ���<!A��&H�u���0�X��<Y����&/F�{W����0���Ɉ ��C���4�$.W*�zM�V�H�2r��>ь����T
��!�� ^��p����"�!������E掄1J��;�`��{���M��H��H�V�:�� �	G���0"O
P0��z�h `g9�6A��$5�S�I� _����#�6b.u�-ŔKR!�D
<k	l�{�#�"k��͑M�s>!�d��:+d�2P�0'�D�[��$!�Z'=N�(fرK� ���O>d��'�X��<�����S	�A0ԫ�U�)�#���E{��iĀ=+�o��hX�0�Ƙ�O�!��Y�x*1;�*�J�=P�X�-���>��B�->�B$�Εgh�CN�q�<2�;6Uڕ�n֜��(��!�w�<1`˄�SO�����w?��&* r�<q�h��*t{Wh<�:��s�<��B�3��A�*ڽM�,l:$��q��&���¡Z.�H�5?j�����6D�TPd��������f]��� d�'D�8��d�8�RT0CꚥY� �'D�� ���_!!��X��q�T��7"O���&jޤ`�249!��'�"xg"O�����DY0V�o�,�14O���D�G�B���=���6 �)Ba|"�|§��)8r���'����"=�y�-� �.%ȓY?$��d8�.թ�yR��\l���F>�6$I�#0�yR�Wx�����$X1,��뗏6�y"��/A��i���T2"��ɢ�ɣ�y�e����1� @�r�Ҋ�y�E�/d��iǔ�f(���,ؘ�yrE#@����m�P�2$R�EÊ�y�L��x���E\�C������4�y��ڊ�XEҒ��6eƭ1��<�yb�ۯ�4�T�Y5*n
(���
�yBI�$qظ�T��)�!��(M#�y�$�+��xJ���?H���J�?��'0���h �D��Q	�F��91
�'	���I�&X��:1)G�C�(�H
�'MB%鳠�q�,�WmP�8���
�'�X9�a䊂D͢b����U��'�xґJ��~�|б�z��3�'Kў"~:Q�K�w� qa�.}�l�Z�<q`%Ǜ-� #� #_�c�L�^�<��C�\� ]�b� +$hʳ��X�<��9U�΁��N;t�Ȍ��T�<�4-�u"%���7��R@��>%�	���<X�%%@�l��}��a��+p�9h6Z���j�@�2ّ��}:�.h�@j��(���Z��\w�<���ȸD�v`�+	�Z�)��J�<�����A����W� ''�Pᡖ�Gq�<�d�@�Uj�I�Oե,�ԭY���q�<A��)$V��'͓C�0pI�l�<	 ��Fj.ĉ�"N`}{�Bb�<���x:�@�:S_����BY�i���Iv�����P��	��
��8_a@�w`�8�yb��0�ޥ�ւ@�b�4�D3�y�j�% [�H�7��7U���q�[:�yr^%\�v�X�P�L+:��K��y�N�d��p�Pb��yF��qn��yR���G�Ё��O+=Na���ՠ�y�F���UI�NА��ʍ�+���$,�S�OG�P��5	O��ґ�ET� ��"O�x�S�N0���)e�P/o[�{�"O��1ekͤU@2A�W���`�.m��"O���J��UZ�p�@D�Q�(@�a"O*m"wD��&x0���_�]�@�@���O����x�vǜ)C�:(�SH�7Z����D"OJ\�І]{�(�5�Θ���R�l8��Ô�U��I��l��� E9D���EA�b	��1VE�q���d�*D�\��� (:�T�1�ϖ#e|��(|O*c�ػ���R�� �IV�S�\k !D���P!��l\N���o��t�+q�4D�0(�o��D�Y`GΧ_� +4@1D�����]5՘�+���5=��l�@�/D�p��׺X��$�%"R�F���u�0D�p)�#ܻ'��,9`�P.>in8`r�_h<��eS�#p��ɗ23^�C1��YX�xGybH��a/t�õ`ͮ.����D��y"H�#Gl򉓠$�8=�e��o����e��ٴ��S�O� ��F�ßV�H��W;!�9�+OTXi����.��=k!M��p��8q�	
�d@�O�1Q���M;�S�? H9�Ԡ��:cT�q��+����Ǘ��l�����L�0m�*(����͆/e�D�3j�8=�B�?�iA��Y^QnX*��]0P b��o�s�'��'fdܲ�,T>zd�C�ݤn�4����'��#LS�av��#���`->���'O2�З*�5":��&H
�BY���*�S�t��<ݬ��
ƺ	��U�
��y"�H
o��Cge��p���#P�߀��IU���O��	�u+F) ���ƥ��v,P�	�':�h:2i�=e��9$ٺx���'%j	��kD�.چ�c�Өwt8��
���~���>;&����ƐA+>j4I��y-�(*|� ��͵#��h��M��yra�d��j�i�*�	G ��y2��B��H��c���j���y"O�	PRTZE
*A�P�����yb�й;��2�A;���s%�=�~��'Y����ϒ���"����"�R������W�Ia<�pa �J%s-08�q�Ҩq�jB䉾S��yQr�K9u�2��N��"0�B�'s�pP��%*$��VCP�#PB�ɿ;V}B������׈Q'F�C��6VA˦ ��L{D�*Nj\C��'���
P��/I����%N�iJPC�	$	��Ź�"��6E24/͕M5�C䉿=����T�g�\T�@2�TC䉱l~���=/\@���HB�J B�I<\�^yZri�	_4���-�9+1C�ɘrf�aŋ��x��!O�EC�"$)�-�3+Ȳw!�Ā��I^WC䉨q�|�CO߷VrTX �O��=B�	-t3,×��+E�h��	=;N�C�I>��xŨ�Y�f���	�9�|C�ae����J4I�2k�iL�9x\C��"[6ʵP ǚ.D���_�B��C�(&pPԥ©�&I�uޙ_�B�I�U���H���T8噢 W�
߲B�	�x��i"�� 9xbd�P�T�D��B�	 @��"����ZI ���&ƸB�Im_3�!�78p��3(@�^�\B�ɢl6�!Y1,�&"'`��^+Q�B�3z	�3Ev\���j
$#FC��*pq �h��z�A3w�ZH�FC�I�zR�����+�81䃓`�>C�ɖD�����Ǆ�rAk�
CkC�I!�< c`�*ZYA�a���yh�B��@� ��P�ٻW�B}3R-K5�TB�I� �.=`����6A�&N7rBB�	z�)Pŉ�P��{�fZB䉪d8�0�b����adj\#9`�C�I�tp�pT�O�/����#@,J*�C�I�K���&FBxĘ;�D=�B�ɁC&��ʄ9v����ϗI�C�	8��É��s�ݓ�N�<�C�I3O�b��c��.d� ͕ �NC�	���E�ʡv�x �W=Y54C�I�|�B�r�4���J>1�C�ɞ?�R�J@(ה�<r�D�G�:C䉿^��͡7"Z<ߺ����|�B��B\�{�M�	%�,aW��8q�4C�I<(e�Y�"���sY����Y[�RC䉉o������w��Ÿ�B�;�C䉈["��ԧZ:5$�	�5��9K��B�	0{�V`1ǍI;[�҅Z�NF�n��B�)� d��5��"W4��q�N�j�!�"O���?(��)��"]{p�0"OF��#D(8�%33G6mL � "O��DHGq0�� ALQ\���"OP����\8b����7��hR`1��'�'��'���'�2�'Jb�'�)����2����4A^���R��'��'B�'�R�'��'���'��`,W�i��+P��pP���?���?����?���?���?I��?I��7W~(�hģ�49�N��Ї���?y���?����?����?���?Y���?9'j {��l���ͤ0�8i�!Eܐ�?���?���?���?9��?1���?��#\1;è�t��'�8:���?1��?����?����?)��?q��m� ����K��a���۸5�
(c���?q��?���?����?I���?q��`���X���Xhv�* �*h�|+���?���?����?���?����?���<�2��!�[@�])��'*ò Z���?Y��?���?!��?���?	��7�@�r0�����J� �<������?���?���?����?����?������!�"T>+��/�q���?���?Q��?)��?����?��,��ڵO' VX=�� �3a�0`��?����?9���?	��?��?Q�U�QسC�&����r�6T~<����?)��?i���?	��?Qg�ih��'ƾ����(7­K����O���ȇϻ<���󙟬c�4 cx᫢)\�U[��jtK�$%�@�2�[~~�!r�n��s�@��"\�"Iv�% �T%���Q#�)��៬`bf�ɦ��'��iH�?y���ix3H\�q��si^�s��a�D�Oʓ�h��� ��ߔFpz�X3遢pe\ ��Hܦ��..�I\��^%��w�"�iC�B��S�X�<����'��;O��Ş"bm�޴�y�dǍ2.ٚ�@^�a!�DSG�^��y�1O���	4u�ў�ӟp{�"]"d���G�F���	w� �'5�'� 7�܌�1OZ��*B�`89�K��npr�`�,������O����\�'$�0��P.,��̱ŏؼs
��O��䀐Id�x�����?qѣ�O`�R�k�wd&���O�OO��"�<�,O
��s��)be�x(��@$s�$!U��<A��iR���OmZb��|�УP�c�\I�&i�e�����<9��?�����Rٴ��dz>-��'B� 8�lH�a`�h�ūW�>�1b/"���<ͧ�?��?9��?!��B�J�lj��@.#�\X�����$[��)���ҟx�	ʟ�'?q��/^N�x�q톋f
H=�&����ЬO����OD�O1��<�FGO�<9�88�����~���a�H�6�8?��By�l�I_�	}y�T�h�<˲	�S��t;�ǘ#$1���ן�iyr)fӬ�h�D�O�(��E��YZT�h	9�Ȓ%��O�n�K�+�����	ޟl�S�ƺK�4{�)�7"�!ȅ�� !��`o�Y~� *~O���t�'��$@ݝ/���R-��3� ��<����?����?����?9����޸6����'��e��XBǫ[����'.�le����1�R�$�Ħ'����^�`��p��rP����_R�����i>�;�Cަ1�'@.��� 15���A��R� }��HF�E+ �I���'.�i>E���\��(l��A�(ą3a��O,|I�(�I���'�`7MO�L�����O���|Z���)W�P�# ����&Af~rɮ>����?1M>�O�h@�0�IC~iXC�Rc$!pd�pF�qf����4��������O�a+f��+fL��!׊�!�" O�AnZ���`����8L�4A�0&�4z*� g�Kgy�lfӶ�p��Oz�䛶d�\�i6��z~T�1�K�jJ����O��Ad�gӎ�|"t*�?ɗ'˰�X$w�tLأAlO
�ə''��Ɵ�����8�������Y���&C����X�'&Vo�� N.6��#D�d�O��.�9O+��y'ɂ5���9$��2& �K5�@<e2��'�ɧ�O��F�i6�dN�*���*�iP?%j��&)ˬ��$ήH�����o���O��|��\xI�E@�f�^  P)�=�:����?Q���?�*O8Ll�0{��ןL�	#	Z���n�I����N ;�0��?� U�0����,'�\ك
͌a� A)�L�]�<P*3�9?�Rl��F,���P&�L�'@-��d��?9v'��Z���SccE=��툰a��?����?!��?y��9�|EّLׯ>K��+��Ī$,��P�j�O�oY2���'-�6�1�i޵J �D�7�q{bALx �d��eq�$�	ߟl�	e��oZv~ZwZ�4���OHJ�F�Q�J�B)F�N.?� ddPs��Ly��'��'R�'�ҍ <P��Ag�a�>5�m�-q��	��M�����?���?�K~��IS|��.������I^< ��\�����O���(��� ���%*_�c���`��0<��9�M�\^���a(h�{��'���'���'�$�+2�څP�<�S�Mw�|j��'r�'9�����P�4x�4]������U���H�OC?D�@)�kҡ-�X5R�ݛ����~}R�'���'�DM���]#+Mp��!./T��
�"�o�����X�/L�Q��t����� n$"e"��I�z*Y޼u:O��d�O��$�O(���O\�?Y�P�n��iC� ?�:���.uyb�'=l6-��V��I�O�mM�Il2��o�3Քa�$��
�''��O��4�F���~�l�.xd��Mq"�%�!�6#��;�("!���^�����4�����O2�D�e���a�M�`�\%:�m\�T�6�$�O�ʓk9�6-��Y��I韔�O���2`ܷ(���c	3�2�Oj��'�R��?Yy�`�h��`��<y��H�֕'ʘ"�D\ ��얧����ӟ�#�|�T�];w�ת ����n�!�xB�e�$=��JK6�Έq��A�Dƴe�Mٔ�����O"�n�u����ڟp� ȏ')b�8r��o�4�����p���l@�o�Y~Zwsb�(�O�4ѕ'
��DL�r����`g�P����'g��ݟ��	ϟ(���h��o��"�2,�R�RS���8�B�:�6�݁@+��d�O@�$�9O~Qnz����ȉX,�� DTzb��� ݟ���y�)�7v��l��<�e"8YT��(DlEh2e��<ِE�/{���	A�	}yR�'���7Yv����\T�0��7��B.b�'uR�'�剘�M��L��?����?!Gd�$��y@KK�J�μ��o����'���?y����	0�,1�[ 	.r�aw���	��a�'\���ư?SvE#������l#3�'X�p��R܌�aTCI�I#����'�b�'��'%�>�"p���$���栮=��\pb�'�v7M�<HrT���O2oZf�Ӽ��o�5^�(�!d�KiDФ�)��<���?��.蘁�4���ih"��,�\Ayd��~H@��+.b�82�5�ġ<ͧ�?���?���?)��	E$�1QC�� a&���%I���DBߦ���^Wy��'"�OXrB�j��aUg�W{Z�*w��G����?�����Şw촤W��z �P���$
�a�Q%�P���'4��v�
ߟ|!B�|RR�� eJ�u�脻T��z�hJ��Ɵ0�	���I��yy¤w�zTz�K�Ov9���
�%�\�&GP�@�
�O��m�y�|\�	П ��s���
�D8� �*G�|�"�떫�tl�l~"��[��}� 'Y�O�G+H�v�����&�,!�ă�y��'<��'p��'��i9Oؙ����_/E0v$���^�$�O���W֦�Yb��Jyr�h�t�O��x�&E�g�ġ�ϗSfr��k8��O��4���4�r���Ӻ�ݴI�)��Qr���"rɋ4�'��%�̗'}�'�2�'����!U%u�;���� d�']�U�P��49K ����?!���I߮)`Ȼ��4( �A;2o�*x������d�Ot�d!��?9��+	*0�fC�O�1P�d
�bփ~���h#o����$�M|?!M>a�
΄&ޠ���s�:T(b�?�?a���?���?�|�/O�o Q�踋�`\�T͠�@vIߜG��2������-�MËB�>�R�~!�g"@ZR�� �D�8^��#��?����M��O�������O?�(0g[��(��A2��"�}�<�'1r�'��'oB�'�� UlM��N�5y/&آ��XT�Q@ش�p���?�����<Yq��ywV�F�����	�:}b�+`�Z�w���'�ɧ�OU�]���i��5�x� m�&~�p8'�5:����%�r`���t��O~ʓ�?���O�R�&�K�<��l�!I`+���?��?Q,O�ilڒ
�y�I�$��;H���uS-dt�5�W3Q��?T���I��d'��I�`D�L��S�D�hO�c�0?y��g���6�^�'l~�����?��J0��LäA�>!Ɣ�G�c�<��II-x@H�fýf���!�A��?QU�iqh0���'G�{�L��$~�!A��-�>z/��������ϟ����N��u7(�;{(����i^ʉ�$��Bɘf�Fh�$�Д'<��'a��'�'�Z1[u��1W�l1���(|�6Y�<cڴ+OF@���?�����?�6�����9�.N����S�_	 �������k�)�S�l�j�H�h�Tm�6��/X�m+ BD�t�n�a_,cF��O��I>y.Ox��&@ܾp�N�B�Aɏk��8+�`�O���O����O�i�<Is�i�c��'v8�Pӫo-�u;��@� �!�'�|7�%�I����O2���O�Y�mTDC Lr欚.dj���OV��7�7?yb��?vD��R�S��}�$�ӳ2G�1	c�=;�z��0q�8�	H�������⟤��C�V z�.yf���}��da�U��?����?1��i��I"$W�pٴ��|�$���ʔ�B�Pp#D���U�O>Q���?ͧSb<�ݴ����6��`r � ��$C�$fF�ÁoL�?Q �-�D�<ͧ�?i���?�Q)��K�|����7���V`ո�?A���]ӦU3�f��p�	ٟL�O�|,뒯gpT�*#�\0�����O�1�'���'�ɧ��ɓ�X�o�7�RI�C�u�<i��	�x˚6*?ͧ"���	j��,G	8�sd�;\���8�	Kp��������ҟp�i>���#d��'�7N�ڰzu�̔=���kbň*8��7�`q5�'�R�j�f�O�Q}2�'d����{qhqpb�:!c*=���'�,=��;O���^������vBV�S�? �1���A�D�}a��ɋG
�<�37Oʓ�?���?Q���?Y���IL�5I����pŢhi�O#&Ӭ�n��`\�I՟���Y�s��R���#V��NH�-�0��4��'E�3�?����ŞVf�5��4�y"�5L無�"�[*?�@|���ybN�1,��������?�Bbe
�6}ؔ O�Pfn8��O"O @mڑc^�t�I����9[�4@WIP>T�=�d�@�L���?��[���I�4'��`�6	}��c�y��ȘA&!?!�Lۭ$�0 5�M���'/�>��L=�?�������Zr%��bfT��-ܽ�?���?��?�����O�a&���6���#��L#S��<ɰ#�O�n)%���Iߟ�4���y�`H?I�$ç �7˨�����y��'���'_�in�	2*���I�ן$=�%K]I��c�"� ���+�b;��<���?���?���?�"m݊ �����
i+i�d�G�����y��n䟈��̟�'?��I�g}���V'�� �.��6�W,v�*8J�O����Or�O1���9p�@ (r��8�FÓi (���6�1?�`���{�L~rʄ�>2�DXB`�<u"R�BB��?���?���?ͧ���ڦ10������Z�*|�<ZA�]�A�V�x3�}���޴��'����?!���?qu���{S�)��J3 ��P���ޟ8=�ez�4��dҲZt���Oj�O�gN�'Z����pf
L�DyĮ	��y�'�v1��Ӧ+��q���":6��8R�'�r�'a�7�*6F�S��MkK>��$]9$ z<��d\;~={����?y��|�&����M��O�nV9v��)�w���G�1hй�׉�O$�AK>�/O����Oh���O����rm$�bt��^Pڶ!�O��d�<���i����'!2�'&��|�V�sE�˜7���9�FU�(D�pI�I�l�?�OP�šaJ�*�֬"�hІH.�����F���i�+|��i>1��'��5&����!��f��2�/�!�
�@C[�|�	�h����b>��'��6mӠ͉^un����mٜ.� ;�
�4�?���5��F��v}r�'tʁ���ǜa[r��ee��9{(�KE_���A�Φ=�']~eW�?��3S��8�a]	'b�#ÇS*���&,~�ܕ'pB�'�'�r�'��Ӵɪ
 
L�y\hh�S'^2�K�4�ƅY���?�����O47=�Dґ�Q�	�dy��a�,�$)���O^��6��	�4��6~���.˅\��zd�SV��p���b�T�� -G��OMg�ly�O(�Ȑ�ϖ(q�Z�GW� f4x�2�'���'\�ɹ�M�FC���?����?���>fN��=��������'k���?�����>U.�I��PԲhr0dԜxH��'��%�4*m����Pٟ����'�&A��.ߚYZ� y$m�{�A���'�2�'�"�'��>�I��^��� Q�hl>5�D́�
���I��M+ㅧ�?�����4����(j����)ףdb��4O��D�Oz�$	\�7�??��(ӁR���) t���̊$="1�scD��<%IO>�+O���O��D�O8���Of�C��]V���C�)	'�2H+b��<iw�i9�=��'�2�'��O����8�>T�E/��J<h�����Kb��?����S�'��Ly��M!�n�I%$$a4���R��M+�P�$	�� .��d(���<�B�ZP�SI:p'l��[��?����?����?�'����ۦŚ5���䐔h\�&�,5��i�h�d���{��[�4��'m���?����?	��M�U���	f|����j7
p� �i�I0<��˰�OGq���N$v(%�f��+K(��� �Q�}����O��d�O��d�O��S�']3���qmT�fĔP���������?I�.����0����'��6�+��%$G���W��#d1qaAЂ> �O��D�O�3YE�7�;?iD	��2HN��BN�/?��٠FѧA.ě�d��X$�ĕ'��'72�'(� ���
�
�3I�}�4H�'��_� 3�4JU��k���?����I�6L6����θ^.��g��9aq�I�����O��$3��?�cD!d��x`B�}���!"��0|@ЛBꂛ����D.��X`��|�!]��uk4��q#����阝$P��'yb�'��O
��SL�j剋�M��MP�h�i�d˻_�|�R��
o,d! ��?�ѼiZ�'�B˻>���r�(���&H�D��o�8DI�)���?1��7�M��'�2�[,M��1���q��vU��a��Ҳvb�����61�E���|�]��UT�v�C�a_	["� 6�׸b$2 ��8	��P����4f��+$i�j|�a��~�Vh0�X|��P87���l�����È^:�&�D�zXh��˼��H!��y.$�Fx#��q�ĆB=J�8��A�n8d���é/�\	��L���A�IN=M��Z2�˒~t� aD)B��s�ƣ;?��I�P��P�DJK7Y�B��uE�.Ci ��%�`���E�b? �;�krӎ���O*�����@�'��y�ѓ$���~4 �ǰhV�9�4W�����䓵�OE�D�/�źB��%.��!��SWl7M�O��$�Ottjb�Sm}R^���	o?�a��ƈ�v�� К0�
��'�����|��'��'���Jrk�&kK
5���JW�:�h��h�d�d�9.5v˓�?���?�L>��x�x�B�M�_�썂ԥӞ����'?|ٚW�|��'��'��	�� �h����3ΈR��D%i�h���&~#��kyb�'��'�r�'aV���)j�&\%�]#!vrȖ�X�L�'F��'t�Z���[������+0{t	�Ȉ� � ��Q�_=�M[-Of�$3�d�Od�dN�4���ɇF�6H��!�; �I��A�L��?���?Q(O��pp�{���'�6d#p�_	2ؼ�� ���PZ2\qc����d?���O����*<*l��A)K�g���.GlR�RaԜA���'�U��.����O��$�he�FOZ�>NX�Fm�bdB��&b�K�ԟ��ə2M�?A�O�����!J�ٱ��n�L(�ݴ��$A=-Ʀ���۟��I�?�OkL7x��yjF�4U��b��Y�`���'�"fA�W��OR�>�1�)өf� ��Շ�	�.������ǌ��9�I����	�?Q�O�˓ևB�O����J\�V�d�i!����M�E"��?9I>Q����'>�*�Oқ	�T�S'��I���(�,~Ӷ���O����2��'��埀��w�~iPSȈ�Z��BΎ#)���>yϚ����?i��?�I�wh0
��D��Mږ��/l���'���m1�4�0���O��w����n���S(Bs�6�<�����O����O^�7�P��I1~ݮ@��Ƈ�=�T5�4�A[x�'R�'��_���	uB��o������8{��������Iu����	uy��_�����^�A�!C��L(.��`������D�O��d#�d�<�'�?�7"zq:)ze��)F:&T��aP����럈��Ο�'�ܵ1E&'�^?:�X;я����@���6t�n���|$�(���t�'��ZJT��9[��9�f���aJmn�ݟH�'�ҭڰ$���L�I�?�X�8q�%ʈ~�p�1��r*O��D�<Y3f�Q��uG�Ѝ[�B�*�).E�(<S!�ɗ��$�O��WA�O����OZ�����ӺC�Ǽo��A���9���#�Hߦ���uyRǚ��O�O�x�R��1X���v�ܨ� �+ڴh��|���?����?I�'��?�R���O�=*CI��v����\�����5��b>��	O��P�JV�F�l�%���$�H6��O��$�O������I�i>���M?��I�9��Лt�B��(Bg�YȦ���S򉸐������w?�K�&,����+�$�p#F}��X�t���xy��d<%��.2Ad�	�jW�-^�$�4��A*�����'|bA�T��pW�yu�Hw�[�a�AZgUay"�'��d�O��ɄI��4�uA_� �!ܩV�7M�.D��ğ`�	ԟX�'�cUeq>ٰ���'�M3p@P7M?�����>!��?������O��'�?��.�F���Z2M�L�33��f��������ޟ0�'s%B&'�~"�.��L�!��p���C'Ğ�㔹ia"_���I矀��p��N�ܴ˒��U7Ԉa�:n�t�n�����Zy�$e!z꧱?�����^wZq�wO��]T��0�5=�Z��'��'�r�]�y�|�ҟ�x 6�U�1��Usc�Лq��`�d�i��	�|����4�?q��?���f��i��0oϱq�ڜ�ՋRj�*h)Љu���D�O"̫�>O*��O������5�� 0�l-%���O�r����� 0�7��O<���Od�	Yr}bQ�Lѥn��P~��kv&���x����<�M��eg~�U�4�Z�9��08�����<;�!({f�:�i�r�'F⭊_�������O��	p3\�S1��D���R��&5$6M�O��d8��S�$�'��ҟ�@����<*dl4�1�وf� 騴�i��g�ʠ����O���?�1t�t�9%c��j�F)	�X78� �'�2ٛ�'���'2�'��s���qھ�
�:��: K
�A!$�M��ЩO�˓�?�(O���O���˞"��7ً(.Ȩa"� ����7�~���	̟��	��0��JyB�
>=
��S$O�\��e��EZd��Av!�7;<!�����On���O�� V<O���
��Vʚ�f�O%�|Cv v}B�'B2�'��I�N\R����$��&��D�PiZ�"i��(���&�n�ş��'h"�'������Y� �(X�����U�ܰ���v�����Opʓ㸄�5U?��I���S(��H��,[���JU�T5fd��Oh���O����3W�$&�D�?��'�DS�7�ރU8�� ��m���	���b״i���'R��O��Ӻ�EJ�k���Eㇴ&Z�  )�ܦ-��۟�@$�a�p����'�!4D�QGL�%%��z�*Č'�6�E/�$DnZџ��I��T��:��d�<�!Jӗ�܍�s�R&3IF�:�!C�v@�l^1�O4�?Q��	VThs��G���xACO�v�j!��4�?��?i�K-88�	jy��'c�d�,0D8���JN��@�5���'�剔&(�)j��?i�,0,(x�$ër�l3��̻Qh���i���m����O��?�17��)H�*�`��5�4e��A^��'����'���'�R�'��]��b,��*�9[5L��7�d������ ,��O�˓�?�,O��$�O��dE�ML�-� �,%�T���6��A t0O����Ol���O��ľ<9��F/��;K6����䉡jR�ɦ�i]��Y����ry��'R�'wY:�'�l�5��C������b|C�D�>A��?���$��9�OB"�)� v�ZC�&2f0�Bc�,�5��i
rW�d�I��,��7e�b��~�l�t!��kǏB��m[��+�M[��?A*O�	'O�z�4�'�b�O
��R�ɛ�c��:%�?:ԓ���>Q��?��|<����$�?����	[�l��(��P�r�!+qӰ�~&����i��'ZB�O�r�Ӻo�����;q����W�}�	��DQW-��$���}�1͏�z0m����V�ڀ&Hܦ=(�*F�M+���?���J�Y���'Fd����ү[�t��e&�I�1�l�2��<OȒO:�?]�ɓK�\��h��E��E
��L���ߴ�?q��?Q�LJ5���Yy��'�$��|����Q�i醹�wH�?����|��Ҁ�yʟ����Oz�Ӏ5���i7���D����+E&s�6M�O�m؁hOy}�W�(�	Zy���5�@әk��ݙ��ڱl*��5�P��Ms�H����?����?����?y*O��h��I�Q�()�.�2-,�ղ��0�l9�'��ן��'���'_"ǎ��(�Vz#�ic5��[�6i��'(�'�b�'��R�l�7�V���E�o��0 Ȇj��ٺ��<�MK+OF���<A���?�"���7�F�����7�J� �m�NVT[��i�b�' 2�'��ɉ_|j�뮟���_n��Sc�Մ_��9�amV8t���lZ��'�R�'��i��yb[>7���q1����	�s��Y�'�վ���'�b^��T������O������h��T3b����@T�
v�����Yp}"�'�B�'�x����Ĺ?e*reE|�ޑ{ �X9�d��(vӬ�!:����i���'���O�d�Ӻ��i�9%N%*eo#e�"(�w�T馩����qq�0?Y/O �>�8u*īp��IC�ϧ5���6�o���8
����'"�'��Į>�ɨ� �ّ�.Fhҳ��[�2�{�4'�d(Γ�䓽�O�e�5f�2="��@��� 1��|p�oӜ�d�O��ͳ-O$�%���I��L��B�ҫH�zUyw��`�&�mI�I�t�I�K|���?��>H`�E�!:�t�p�<)n�f�'*�;�.'��ҟ�'��ث\F��zF��%@$�XC�$X�=�DEb����d�O��d(���dDE�,Ν9.B��L��x��9RF�t��?YJ>����?��놧K�epc�JL�j���Gxt�����$�O����O��^���P0�D���&��TH���x�U�!D�~}��'��|��'��a�$�­�b���&�9M4!Q�	L3)[�듷?i���?�*OD���Tf�Ӈ�=��-����ȱ�B�$��P��4�?�/Ox���O^�$��]W��'}rD�4:�d��
�oN(	��U�M����?	(O���0B�]���,��0:L�ks��D)X��2b��8�J<Y���?y��D�<�I>y�O �$�$^-�]��l]!Y����4��$�)O��n������O��)�l~r�^6&�LxV!Q9f� h!5�O��M���?�Q��<iH>!��ԃ�D��06"ɦt޲XB	_��M��rś��'B�'����8�ɺ�v�����!�@F��ew�X�4Z��܁��	�O�q2����:E�Ӥ������4�ަ��I��T�ɑd¤�ۋ}b�'��d�e3<u��F۞1��5z���^��|���e��T�'n��'�f��g�	�?X��t*���<��jvӄ�]#\���%��I�8%�֘"��i���<.���
�.��V��,=XM>)��?�����DL����/�m�����=���2I�}�	�����n�I����ɓ,���zA��[0p`���y��M�Ǩ�ퟔ�'k��'�BV���E����$�ޓi�Y3"D��iU���g��>����Ov�=�)Ot�Dδ\_p�[���#Iȵ��T+�8��'�"�'��Q�x24	�ħ\��\�A��a��%K�o2�����iў��'5�~��"��B	�a�dD	;e�P��.�̦M�	��,�Iܟ�u��j��T���S.Q=8��#�������z���H<!����ȡ>0�֝�rzxd�PX8.��I��FO�1TN6m�<y��@�^y���~����*���h��\)l0���C���!j'N$��b{�㟨�3�.2�ڼ�&f9 ����+�	�����W���'^�'E�t�'_�U>�(�G����!zT"��Lu���IБ���m>�b>���hF��Č%&��$�󤗅wȨ�4�?���?q!)�eV�'���'��$( _���砓0�������R`�O�-�T��O����O|�dE�k��8a��#/��wWԦ��I�~�a�}�'sɧ5vL�F�̤�5�=NDa�'�A��� �i1O���O��$�O��đ���H�֯N�~5���7O��h�I�<����?�����?��'L`��$��`1��츳�4}�''r�'�"W��p�玁����ְ��]�u��\��TN_�M����?����?���'f��R�Pԁ�d�>�l����I�|��ʟ��	蟐�V��A�4�'� �S�ź|�r��C��zD��bӈ��-�d�O��;��H'����V8�$�
�'��#et���b����O����O^z4h�|����?���\��-�'���e��1�d�u@����xb�'�剂^�#<�;mT��8�22_�M�܌���o�syB��h-`6M�O��d�O����L}Z� �%�#d��K��E�� Z�E���x��'�ў(�Oj�(�FjX���cm�|8��P�i��1�p�'+��'��O��	~��� m�*t�Ǭ�gF�Iz`)_�0�:r�Dx������|o����
~��i���K%)�kIH8�iqq�4S�a}BaۛpC|4k$�Y��\u�ʘ6�p?I��̅oj�	���>e���PG�(�>Di��'wh��3���!�iCiD�l�F�0y�f`��B�<�n䩕��1[0T��c�<�(1"AJ\�njr�0�@�#*�0�r(���
g�P9~h�ss��#�F�j�HY�zB"� ���Mw"$
��6.��1�� 
3��! PN[某�I���	�i�!�	����'�T��5G��s��eqF�I�%���J�'�&c�~a��%PE��*��C7��X��,^���+# �<^~���a"��3���h�L�;\�q��'�+
@V���)ڶ�D��P�"�'
>x!+��q�&���#�B�����	N�'�J�Y�K����҉e��9��' ��2�I��e҉��`D�o�ļ��'eZ���d�?IgȰnZƟ���~�dMP�J��9�aU�^����JIl�&q�t�'���'� ���_�s�|���.Yj�T>�11LN��\��U�x�	V'-�A Pb
@�+&.������ħ.\IS��� E�uM�- �YEy�?�����'�?Q�h�A�X�k�n�!}��Ppb��?����9O�t�.��ބ9��͞*�DҦ�'�O���`�}x<����מ-t:�7OX����h}2�'c哏M�Ұ�Iן��I�'��!U��9���2C��������R(f��p��_6 3�S����'�*}I�dZz�^���$�=(���ɡ��#xM�,ɕ{- h�a��O?�DV�O�l�`�
�"Ԫ��ԃ��Md�����O���,?%?Y%�)���(z0�f��6[j<���=D����&-��`4�BF,`X3�:s����'F�J�h�o�:MA^� ��	2_�0���?�A/��c����?i��?	������O�B@��|��@��
�O�رbe�O>\�5�w?����HXs8���eC�t<"�k�ԯt,%x'����R�8@��=�M��p<Q�Āt��`ʡ�&+�  #��`?�w�ǟ��	l�'��I�D�����79���UF�=��B��'{�\�:g��
'>�|p�b�1��I���?͔���A��6GXw�L��M0Ƙ��!P�x�P���Op�d�O"IKp.�O>�{>ٸ�_�3Ǯ,���q��*6���K��^DR9�R&�d�6��1T�X59ԮǰP �D��a��8x��S��t�a{bg��?���Z&@��&���SQ����9���0�Y$¼����%oq�1�ւj�܆ȓDHxy�7/S�86U� 	�8ւdΓ �IBy���m 6M�O@�$�|�dbD�
�<`0K�7h[h���7��(���?���X
�̢�Lߐ%}ɧ�i���с�Z�xF�(A!�<?�Q����+���D�D�C:9<n�(�-8�� %ʻ�(O���%�'XR�'bU>!���:J�(��
L�L26��џ��?E��'�N�֌����]���C��
� ˉ'�<S����g�:�A�ǰ' �9��')Hș���>q����	�F(\�D�O,�j/ΡڢI��0|���e$�2D`!ص�ѱ��
��W6kf�YP�|Z���>���A:.l��
S�DD\���Ġ+�\Aؐ�F' ��E V�p��?�R�J����y�y�Z�X'	�+r��I����z�r4�!ǾU��["�!e����`��x7g��l1��GN��DGx2F"�S���;XxZ��S�6&��r� 
�q��'GN����SW��'r�'���ß���dčچ+&=��P��*Q�}��(Ly���d��>Oh���
ٚk��	1N ͠t��,.����땍)��D��ڟў��٘N�@��ճP몽j�챟d�B�O���%�d�O����<��!Sb�a�tj�
Fda�'��J�<9����
�����0k�áFD	Y��']ɧ�D�'o�I�Jhx��4N��@Ԅ̀1O�q��ݳIJ�����?���?�[�?Q�����.+TrrM�d
�n%�\��۔3#VA�b-|hH�$ǈXXH��D��k����D54Rd8�(�I�I����X;�D �ɝ9�$��I&p�����O���9Ķ�Y�����F�(E�2���OV��0�)�C�)ɰ�˥�O�C>� p��I�<i�$(R���0�_7qH�[�O��<٢T���',j�C�ei�2��O0�'x2|�� D}�(I��J=N��P@�I޷�?���?a�ʁ���T>��#CR2DF�@�r,-1����  �`o�0����Z=n���G��o����S�Q��3���OV��O���|b��4lE���\��f�N8�?����9O��kX�H��d�!�R�	�~��'h�O� z�� -rz�T3�%܎#)��g<ONI�D'����	ܟ(�O������'*��'�,Că� Ҷ1"Cҩ��$��*uN�	���W�-s"��O��t�矐�@�>���!c�M�0�PA��8�|������ه.��?E��{l�� ���e�gd�|z�צ���?����?������G��1 !�89�h�"4ϋ��yR�'��}�˸M��H�� ��D��W֑ �"<���U�T����=:��Ќ_>�2�P/+�r�'��	Qt�/-���'���'?�'�?���\�,�Z�b��u�~ ,������'��y�R�˟B�> ��@�SF{�
��8��̦'NM:�*�8/�`����28lzC'ج�p8���hO`X�M��B��Ey�R�fɼͻ-�O�l"�o�Ot���O�Y���IVy�hX#u ��cŚz�r$�Jڏ�y����Z�u�C�4A���YF#=Y/���O���{s�yJD�ؓm�nu�F��3:�!�d�
}d� R�_�[��K��_c�!�d�"D��a�d����^�p��"O$����ˢJL�d�Ǯ�w����"O@P���R�vL�@�l	�.]v��`"O2E�Kː	�l�H�l݌VX���"O��bg�|%�Г�ň�[�0xE"O\��-�$I�z���t�� YF"O�8�w��(-:6�рf[��9J�"O��x�� {���$@I2o��M�B"O�|���}�~�S#
�
D�Ҥ"O��%$ܓ�d��-7�=�"O�y �Jwt	v�U�^�F!��"O�	�W�$����I�21p�"O؀ag��;>N5��"P�V�T�K�"O~,
��VjN���QD����H�"OFlzD�l��0r�	[-n9��"O���#�^=I^��;��T}�@b"O��6�G�>0�T�N�b�����"OH����F̾U"e���lul͈"O�u��$�UR��VI{X�UcB"O�Q�� �(�}�@�ZD�zL�6"O��+Շ@*�.��6g�#sq�je"O\MibΥ!���&5^� a"O����ĝO+D�i1�Ҁ&��١�"O����ᖧQ�ޱ�b���z2"O�\ ����V�d��%㌶o����"O�`ѧ� wA45 WD��T����"O�}����=P�퓲��AN�\26�ȗ)}~@���i 8�8�#���էY8k�ǔ��0A�	�	��$H&���$X�9z���BS4���P �$x�џ�c��
(Q0�'���O0>�$@���R8B���Tj� !razb�<a��u(�G�0yZ���!W0Z�$bn�),F��u�ޱ����e',�&�<���^r��#�"�B���2�\!���N��i	�"��^l1O�h�*���(�*���������䘟E+�L�f��b�~��灖�}d�ɺa���'G�-XUl�x�'��M��'N(]WRi���GZ��qbʤX���q-�������ɻLѰ�;q�;7dA)z0�ɰh-�ȱ��M��0=�1
O8dP4"��M�� ;�#�͐��ƓLm�`0&�J�0,>��/�#l��|�˓r�X}%N�X����]3LF�Y�,�p��)��ECBl���'�(��(�Bm�����I.�W�M�`uX��R�
��I��x�T1z����"̥s`*���a0�<�c�P:?r���� X%�� ��C# Ykۓ|�
��)7#F�h6D�,!rhݠ�Z%>t(:f�&����PT�)�;��D�<���(��',R�g'��5bߌ1���3�:B"zrJ�����*��5&͙>��E� ��Db��R*+R�(�7�O��~/�URX�}&��Z�$]�g
�)u��e�R��sF^LX��W�$qK��P���<A���)!`)��BU���I�7��3d���
��l�T�Fy��E �H�3��Ӽ{ϛ�QSZ�#d�B�#���a�HZ<yǋ�(����:�2}HgF��&�|J+O��0C@z\���H?�I�I/�8��V&`��T�<P����=52 !c���"/����'�XaRe
g��4�
�.�Ti�'�6�rB�Y3~*�����'�Du�4@��@y�D*�(�G�Zp��O��PFA"s(��M����3��#� �svᐵ�v�S���2���%!4��pR�H6z"@I��U�z�*���)�(gŎe�,O�p���>��>��!k�i+�g�������+h6�ad�5$��[e���U��ԡ��D`��bŃ�9K����I~(�aJ �>�5"E�~|P�>7MJ4�d-�7n�6u&�r�B �ayRg� Z��m�a����$��._k��D��a�e�/��I4�|%����m��y"oς�\iR��-c�t0�vf���ēNn�"���i���|b@�� a��[�K�C��q%�8��T���4.yB�	.1&Ly�!⊍bXU�F��>.)�P�ʅ���9�B�!Δ	o�D]�M��:�wdH���ed�xL��gH�Q��tI�'���!e�Q<<,�B�8F��̢ڴ$�9ŉ��e Vӧ���E���K?2t��+��N6�83�&D�dJ�E�G����ӥC�4��%��K�>����n�J�#"&!<O�Y���ھ�D!�(�).�T4���'��j&��kTpm�ӈ�:Pڭ8�o�*�~��&L�Vh<Q5Eʋ�	S�̟(p�� ��m�'�n��&�U#;
������@�x�A��2����0$t�<�� Y%:�T
���VGJ�M���%	�L�
���֒>E�ܴD�l0T�3A%��(��$�LE�ȓQҭӴ ۖ R ӯM%@�i�'Y���
ȸ>��)��I�C��c��Оl��}��� W"��dL��E��i��Eav�#B-���Q���ͣ��X�'�:� gX!�<Z6(59��l��d�(�	�7� '��O�l���aI�7/�1��� '��L)�'���4"E�'�,H��S8#:���ݴF���L�%	��ҧ����G2͔09��3�� �I��y2F���`�kv�L�O���ao����֞&��e��I
=_v&���hO
�*��̀=������)�@CE�'�P �6��
�(���?f���r�G�K7��%�ɋX��a�ǘ�p?���E�4P��_�oJ�D��0�q�ċ�h�2):��ß_�ݥ����	 �lawʆ%�¥�"OX�p�51 r�
��ҴUs��)ֆU+'1.Q(� (,LY1�ݾ"��>�	.?�P"f�8%���!C��:b��C�
NX���k�!�ڜ�Q��o�¨�@��->�F��9_��h�2&|�QF}�+O~i��A��m���!$ʝ��=����C��E��G�v|�`ዝ\�p9냃Q�Y��� ���Q>��	�� �T��Qh�"���0J�(8�=-C!I����������n���Oh4��n��m{Aa^=F"�D��'QB8h��R"'J�		�)��q�F��-��	($p�̊� 2��i�Q>���'�ɀ�W�M��0�Ł$b����$��E�#�2�,򶼃D�
`�H�(ҡ���\�&g��`�T�b�|�6)�E6��R1cG��nիf�&,a�[�#�);�O��%77�T�u
�p��,����xTN<h&d�h���:��˙¼!�C�ԣ&��~�����������>A��9]'�~b`�/a��lX�c1�t0����ZX��!����?���cS�B]�,�mJp(��p�')Ё@S� ������VC�#|L ��+*���A�(�T�3Ư�O^#|�"��$)D%�2���R���()�6p9e�8ʓW�i��	��T@�K�@76��ё��h*���t� ua'�>]	Zኢ
����Oح0�l�811r� d+ٔ��i���'�f��d�.?F�H��f�1$nf�91E�Z~�0��Me2��2�n�Sӄ���	��p]��b�+i��%�>L�c���!�~̦ph�Ǖn����N�O�;��[WHJ
-bU�T��Q���/qh�`�J�	��U�G��9Y6  ����Hf���GJ5=��	R�O2lA��l�f���!_Ҥh�7��]��FN@�R5�O�m����8O�f�������b�11@���a��@">�A� 8" ��8R�b��MO�+�9X�	�!zў�#5����Fe�W�Z���j����1��9U�Lrl2�����G�I�?��"I��F���0Y��\�v�A�2����fH�.(ZLb���b@�h�L	�A$�-��)�@�O�8e,d޹�ĉNxa��D�JhAH���?��ƅ'_���f捰@�d�K��
 �\y ���-��		`@�O�"|��L��|���a��q��0�~���%�%(�(9YN��P�gJn�g����� �=)��T�;T�"���A �ё��^%P@�Aq��ƈOt4�D$*��PѠ(�=�e ]1k@�a�b�^�HO�jT+Lh�0���`r�����O���2\pB�\�],�����_�ՈO�VЃF�K�O� @��u��[R�����v�"w���B�d���ōfܐ��}N8�n�C��O�	�E�0v����|�E�2r�Ăd�W�O$v�AȟT��9z�e<^d��b�4`�� ����ϼӧ����D��O*�t#j�v����<zET��$[�p"��hC@\`��K~�O��0��g�L��C��j:5Y�AB�o��{��~���褮C�U�$���ќ�J�K��:Kg������Xy�%�Ž0DN��pN�Z�ɝp�>=a$�`��ĥH�	b*��Ua�s��\�V,�$q�ը��	i0V�KF�t|�Xc��58�6��>�B"	.�^l�K>�F*)nx��K��?I��Y�"ݐ`"�t�Ug��Y�N5��=扡N4���e��"�X7�V��-,���n�=�r����~ �����2r�%���	��r��Nׇ��)�� ��x}0*Pe�;Q"�(cum�Y\q����Bզ�!ʛWF��'�4����U
��ֳz~X�ȧHL5�JH��J�p�j<��ů<
�U�Ԧ4<O�a7 R�Q4x�$�G�
�@r [��� �J6	�b�"}�dЂ/XL��W@T�|�-������<�SHD�<q�,����{�,j5��"s��m�0Gd*%�����A �	�$D�2t��Y8$Y�0�赘CCAW�T]����*���3u��-b��c��1q��"�ds�C�%|:� u�l�N1�C��Ln���"";4�R�g�G�n�:aZ�L��!���I$��i ��f�'�h����0a4�N����p�F�\P
\�Q�!o�)��'�/W�����5P��5��s�|����@�u�W���D�+ �DIu^����T�`Z^ �!�'VhU:D�XM���;BլL6��Bg�N�#D���MB�3a���f�'�hT8@�X(��9J�~�h���:V�yjR�m_8e�:�
�=a���d�	*4�P)C�C?Dz�pc��6��ؠ��O��Bv�_�k�vyj�ÿmj�"=QǎZ9R���B>L������]��d���$ە��c)��I�Ξ���\9��,�4�_
|�Rچ�Y�$Y!�dS<,Y�L��U���s��T���-�	`�tS���4�@1���F��M#�.ȩe�ڄ+P��ٚ,O|�<��[N^���m9�D�m��/�^�����\��L�v
�3ғXl�Ӕ/�? ,�pS�[�n
\|��I�.�\}��F�p��r�-�4�i@�C5`Y�KGZ���ɺD\��{T��9���GOI
&�b#>Y�60:�|ړڽDn쨂-*C�	��l�k�<����D�����+U.�Ɲ�<I�CN;~�ȑ�<E�4�Ur���gL��c����a䙠�y�
`LĨ�揟�p�M�����Y��%��'�Aˢ��uF4��&�&�, �����)�K�$'b�;�
�d\x�� ��I�$���|�ya�@�+C
\�9CB�uG|��k�);��i�`g�p����81��Ę;hq!�D�) �$e�:���-B�`a���V`S����	U�D��O�'}�>��gK,s�B�I.(�h=X��,.,ܑ�e��{�B�`�Ly����T����Ԣ^�2��bM87>@��`,�OhZ�`�0VRH5b�Gћg
�M���lx�
�'�D�A�L�w瞁�rO+}5�l�����c�v�G�T�J �U	���(�XM�&��y2Y�H2tL��k�p  ���G!�yrX찔B�/|:q�UE+�yi�%�D��5�m%f���y"NB�a��I9F#�;+�*�(ԅ��yR�q{�#`�6u:����yB�
8i����j������y����-�6��aA�!]l�1�B��yB�X�&K���i%@j}rq�E�y��M���A���v�b��/׉�y�j	's���%�q�X�A�m@-�yr20
D҄�
bI�рA���y2_`�9*d��0W@���E���y��I(i�D��fÍ: �s��4�yRaߢX�`���#�?*� I@LK��y"��>/ЌAiX%�"A��y�FGi��ˁ"\�O��H��F��yb�72ͪ����M��!Pa��yn�F2T�aV��D����Tl��y���'���� W�$R$-ؓհ�y
� x�[֎v�j���#A D\����"Opջ�&�`�>� Ӂ[ yWd@�b"O~�pFK�Yf��� Y�7r�̓�"O4�t$�= �J@�aEՖSg�� "O�ـc�4t0=8q#�8L-� "O������5$�Y�P"8��T"O����0]��Y) ,�)��Z"O����cЍY��}R�L�H5�`c"O��[Pȍ�7|lU�CKP.*D�K"Oj��-j�n]	6�I�� �ɴ"O�"A*�Ep�#1�I
n�p�3�"OX$B�
�0�X(���F�Z��"Od�{w/W�O$�CF�V�?�h-H�"O�����͗(�I�!h$�@���"O�w^3N"�+vE���l��"O�(�⇚2g��|Rũק�y "O<͊�l-(!��2����?tZ�#	�'�M�d���%~ 9�n��ef�-`�'T�		���:]�u(ËQ��b�	�'c�\�Wo""z큲+.}���9�' 0ȥ��>p�,p��F�t�pm!	�'P���&Ô2Ċ��kS�Bp0	�'�֠�DlSp���k�+y��i+�'a����jI3eX|Z�昆p��p��'�L5r�#�3{<���� o��EQ�' �]�H؉m�v��e��S��}��'e�ź���~8�}�W#[P�hа�'�����3P�5��DW�v�R��'��L� �:jH��r�gؗl�2�	�'�ĜH��^(>ȑ�0,���p��'�@�r���K�Y�T��P�p8�'�n�s�	P�G�a�ΗJ*���	�'<r�R���0�(��F�z
�'>�ȑ�舚��T��Ĉ�7�~ ��'t���r�D/CN� �1IS�D����
�'�ԝ8u��*A�:1�͂:���	�'D(�i嫆�)�V �C��<����'�L#j�-~���b	Ékz%Y�'�yjBhȺ[��i��fν|_���'���Pf4|�\���*ץ`s`���'<~LfC�2:�"BeN�O��3�'���L��!���
\U4�r�'�x�3�F�"#�����$��5��'a,�z�&��,���Qn�����"O:��돃4j��֏<M��1"OXl�u��>P�Iїm�b���3"O�E���Y�!��	����tYQ�"O8�POڶvΡqc
ߚg4Q W"OTT�D���,P�QI� ]j�+"O"�0�c2{�2`R���3u!��"O�e8�"���!:ƮJ2�-j0"O �S���(W<�e��;��X��"OK^�*���ҌTJ������y�AӺq6�1����9�1玲�y�[1<*����lU/C��0�r�;�yR`E�z�N���H9�|�����y�%� yâe�qF˃ �q�qˇ��y��4��%�+�49���y�](t���g�D�v��h��eӏ�yr@�M���ȶ휬���k��(�y��Y�8�r�������1C�_ �yb� Cn�K�.Ѷ
=�xe�7�y�"�8mO�y�6+�9�XM�!�5�y�.Z�CC�`qF	�~���a����y
� $0�'��8�h��Ez�"O��h"��to(pLہ5�r�id"O�ay��()����ȓ�v�����"O
Փ�B��XU̠8q�]�o�U����-ړ��v�1���gh��1&��cMHA��� i�Q.ЍE�$r&;M͖Շ�cF�k�"C�L$x8�E�� }�b��__���.ţE��:� X/�؆�%�,�9Q��\/Эٰc֧fz�H��ov8:�^$l 8���O?Y�-�ȓ9i�=�d�� ������]%*��ȓ	����S#}��M;���	S��d��U'nM�6d�%i��J@���TC���ȓ0͘2�� ��tҧ���	���ȓ!�>�{�Γ4ttp����0�Ć������l�n�H�J�[����ȓO`$�Y�e��]���Af,̥r���ȓ��8�d�;Sv�� � 0����r�da�I��C]J	�HX[�$h�ȓP0��('̭O�$�C(�
h����ȓ���@%Z�m��m�n]�3"U�ȓ��py��R.T��T��IN_m�؅ȓ/���VD�Y��D����|�T��A@b�[�E\H+���9S�4���G���5 ��(f���~쬼��J����V�j�m�'x�楹��-V�ɱ�9D�X�Oш�Ti`X9-%lRe6D�ѴE��ʮ�'`A�PDI��K:D�4�ɘ�6�RF�@0�*=��H9D����AH���9�`o�E���q�7D��!F�W=�@KG#[�$|[��:D�hU�N�"�-��h�)�~<"�9D�X�t@ʴtj,!���V��G	"D�8ѥHG�W�Z�b�X7_N���e,D�`��k����@�R�I��t��)D�h��?�=Җ��
�)A!"D�ܨ����`����*O���`:D�`Bcc ;���"�̈�}v�o<��s��`���I�|�H���!�1A�^���+ D�Dk��5r`�0�C�_7a��v�;D���U$Ng��ѥ��P�0���5D�t��-[)F%�Ѫ�� |X ���>D� 8�I7 !�h�MAu�7D��ʓ�	l���4JӹP��)��3D�d���pn5�����e��d�&D���0gK;���Ι.Y��)[a2D����"]	�P�W������Ũ#D�����L�]@  $/��=Щ�f� D��j�g_h�RI���EN���b"�È��pzS��7v������ڔ�9&�|��)�S�kۆ�y"Hm��Ոŉ�K��C�ɬX�:\c2e�(P`P�!0�W���B�	3t�0��
e�]���[�AB�ɿL�uZ@��+�u�Y�v��C�	:�ơYO�	�~ɸ�*�~=�C�	�h���q�΄�8fj�)s��3C�vC�	�AL��b��MuQ.��"K�NLC�	2
��V�U# ���F��A��C�I0	�Dc7➺4`䴡��Z7y"�C�	�j>`���\�q(���3;�C�	2$0D��w�4{2�A�<O8lC�	�g,���G�%8x��'���B��7!�����k�.{�`�D���D.}��I�\��q���rU���ڒ�y
� ��r
T
�䑆OX-*l2�"O|@��
�>��ӈ�'�Ҝ�B"O����m�z}
	rA��v]�%34"O"��g�l5�E����@v�)a"O��cwF�%B�4�#�O�hj��"ODa��A�+V��D�!ܣ|b��e"O(S�'�������J�>'-��G"O��HӬH��b���I�}!����"O>K��ȮV���4��k-��h�"OF��ԧ�0U`�h�&Z���#"O�@ o�|���z� E$/iʥb�"O��p���_�0��1��aG��"O�A�D��$(z�� ;&�֨h�"OR��J�#bY��b�L � ����"Oz=B�E��B��\��;V+K�u�!�d=��� �ˮF�,y���͠o�!�$�2h����醇I�j��-�� ړ�hO��HPm�_N�!3��k�H�J�"O$���$�<\!P3�Ety����"O�%�6�^����r%���jp���'�ў��
`�(D: �a`�xK�+D��W�A������,$Ҋ��/7D���&�['W٢A��N5�Xɺ'!7D���f���|A0)�0��10 �]�� 5D�(j
Q�x���f�V)B��R�3D��j'��,0�+W�� k{h�a�0D�Ժ��J=_�<�G��fS4��h9D���B�I�&��U{�߬��5��<D��ha&K�vL�"`JR,&��f�<D�l�R(�0HI�|a�H�F�
AZr�$D�L�T�M(gF�q�cƞnpF�{��>D�$	t�G+u���n��=3r��n=D����S�o����eǟ9���P�n<D����"�<���f��<{�H�be:OR�=��L�r�P"��CNAٳ��F�<񑂙�  <�҅
��F�NY����L}r�)�'9�N�2�%ް#��9��)h���j7Dk` W4,8A���R.8tĘ��]
ʴ�Ee�&N&T��۩b# ؄ȓ0�F\2����!h(�c�("�
��fS�}����?WT�(���N!b�@q�ȓc.$�"��ʝni��#iV  آQ�ȓ(��`��kE#i�2�t$�}E2���d{()�"�^�jL�L�4��w�|�ȓ.��I`S��D ̠�_?A;��x_�̱7&��u4�T�W��q�<��6��2  �c����7�@�i� Єȓ �0��%O2VX�ր��e#(�ȓ��(D/���H�'9y}�5����5ô��x�`�4' 8��-�ȓj�BD R�
�8,8Umς}�ȓ-�<SVCK�c��A��
>��\�ȓ
��q&���0��uڦ�K�����1�F �'B�F�ڝ86l?+H�h��Z����'!&��!IA�C�f�ȓR,�(�씨p*�Ď;{�x<�ȓL����4��Ɉ�ό4?����J����0˵J��d�Š�8v5�ȓ.m��e�W�u)��©p���9|��+W*�.�L�g� �N$�ȓ[�j�j�A�7:�|!�=f�lD�ȓ	���G�D�D��F����ȓ��� !�n�XE��Z;v�݇�-g�u9�к0��Q�ЭC������S�? @`�q�@ ���#���#&5�5"Oj0����S5l����[�>�9�"O�1�+�P�<��7dW
F�,��c"O�(�am8b�jXZ��V�3����!"O�Mp�C>S�R��d±qS��z�"OΈ��F�$���r�R$+L�Q{�"O��:a��y耀:�KK�v[b�i�"O ��L!f-2yh"h�4S.�WL�<9��]Yppl+���R�8���)�\�<��	X�˳�Hd_�m�4��`�<�4��F��f�>,��Y8�.�U�<!��@�rk$e��1[�hგe�L�<���.V��{��ͰzܜH@-�K�<�C҇!��w��6B� VjK�<�A�Էs ^u� l�+*�����DJ�<�r����9�g�'&>V�F	JH�<�g`��,sd�h���,ex<�	�D�<	�h i�T�8ce��$=�q��h�<�/Ú���c�S�P"�g�<9F	:yC2a���D�`	�f�<y��
���4)�ܦ%.�����a�<Y oE;mZ�[�F��"������s�<A4�-iH.��퇟[C0�j�/Xp�<If.M4u��,b&Əqtz�㏟m�<q4���PNP�A*�S�-�ĭ�B�<��m�8l�bA#qX�P(�!bW@�<�X"	b�t�g�ԍ�h�
�z�<y��P�B&��eBn|�Ҵ�Cv�<1�%OD~Ճ��X�Fr�<�a ��9��T*�\���)Kk�<�A%*��@E��9AN���7�i�<qd�_n��)C�`C��h�K�}�<�Тˇ  ���-��`r��eI�v�<كM� k� x�ے�����\u�<�cm��PV���[el��w$�j�<��L�\�ZQ�d��XW����\e�<�&��59�������b�ha���^�<1aO	B��:V^�$�0i��^o�<�d �?��e�%G�{Q�I�v�<IKW?O�����+�l5x��%�Kp�<��"�3�*1�@AĂF��A�ho�<	�*P�D�1��C��W���ia��h�<����1t��5��'��TuI�B[�<���d�\,JA T&��#� }�<�piHV ��7,�
R�l�S�<9�&��	����ϙ�uw��T�KZ�<)Fb@��jHpG�K�< .���a�<��Y|^�m�G�ׄqb��_�<�㯑�+��Z��Y�"@U�R��\�<��l�.!�qD�Z�1�nBB��Q�<Y� W���RF��.x��$�Q�<p+^�^9�w9O�<ai�h�<I
�B�t���I*X�0��.�e�<�7��A!���P V}���b�<��O(��§�D�P�r$��%�I�<!!$\3����b�En�C��\\�<C��m�t�ˇ ۄat@�{�'c�<1b��A7�c�
�&�����)]\�<��g^�8-�Ċ���_V\�զ�Y�<!R�� c� ���͍?��x�͑U�<�d�Ȧ@2 Ӆ\��d��#X�<� +�2�(��ꘜN� 0�DNU�<92��G�V�P�J���XT�\J�<QGP\���R C�6��Q�\K�<� .���+�	X�"��;�}�"O4;Q�N}�|tk�Hu@�ab"O�qk�-P*E�"92ō�"uR��e"O��)��-��ػ��+��DB#"O"%� � �α1q�H!z��""O�y���&!� ����ruZ�G"O�%	3�8���� �
�z\Ja��"O���PJ-y�X�Rc�ʘVnF�!�"O~P#��W M�T�"đXt�Z"O���5pl��x���1 M�Ik�"O�m�&+Z�W�p����$b�b�"O�U��!ܨ,�����&��#"O41�R�H�;�i���X�0r�"O��ip����r�8L+��A�<�W�רҜ��f®J���3����<�u-��I�ZȂ�4Q�"xs�L�v�<��.Al�>I�4������t�<!'��Xh�}@u!�������l�<Q�Mݛ>��"��؅.LĬ�H�M�<y�Í�~6d��Ac��L:S�RB�<Q���,������ -��I��A�<q0�Bx�Bc�Z�ej �9�x�<$�����Z�˃m�`b�J��ȓ\���%[$_q4�q��"����j�:�P�#�_d )�ũ�.��3���w�C�A�pm�bI��^��ȓ.y����FԤx�i��j_�Z�f(�ȓ�钶���g�����\#@hY��5	t��9%˄@�E֜5ށ��BP~HJ�!�2���C�Z*> ��ȓ|	uB����8d@��z=��S���f��;x�ge%�ࠄȓY�R��bM?L�L�T`��ט����"�*�AK=@����d �<>�V,�ȓ@|"�P���7�p���A6G��e��g<�))��z2I�rhܪr��ņȓi[�����tbjE�|^<<�� �.�3�e>~��$D�(��ȓ
Ć𠦣Шo�TP0��<V`a��B�t����7�MH����&"V��ȓ:��M�n�4/O������4_��t�ȓ<Yΐy #�����F�A�h���ȓl�M��JeJA����d����c��W  ��b��g��	�ȓ�ʭ�'`T}6HH!i;>�̈́ȓH��l�t��0M�ԣ�� U����F"���֬�i�\�\I�:�� "O���$(��[t��u��h��"O4K5�0I��������y�"O�,I�y�N��#U��DT��"ON�І�λ3�Pq�Ӈ/1��H��"OH)���!=�M+a��4<�&"Ol�����60��ń�_`1ӕ"O.�� F	)K�ڈڀ%F�A�@P�"O���A�;P�8Qrģܡ��S�"O� 1�b?H�+b$�8w.ۢ"O��K0�ϧ��X�!��J�B�"O��H���L�x	y�����Y�p"O��t��k P� AG0~z�H��"Oh�V���( ����a���br"O�p��C %)�Zyi�Є*z08(�"O��P��P�(m�7)Y�;|p�it"O^�#��[>M)�K�g�8v��a�Q"O
ģ,�/u����?�����"O� FTq�-�������͙���
�"Oh @�<{��lKVMFG�P�"O�MZ�Ğ ���*�̈́�k��T�#"OD�"��H�����x�6"ON�裯Q�!�X���V��j���"Ot(y�fZ�?$HQ5�"y�bh��"O���i�2#x����;:�)�"OBT)����v��,�I��&��\�"O^M8�G��d�Ps&�ڽg����R"OR!����5�a[��v��q"O�]r1�G%i�U���g�d�zQ"O��xÄЈf�^h{�ai9|�B�"O�T!�ʙh�i��R�h�$�#"O�ɠG�W��
pJ�mR�"O�(�Rh��(\ҭ���Ks^���"O�c�"�	j��Ec��Xm��ٳ"O���C�h��}�wÜ�e�I�t"O�h�ã�e�0]i��?\D���0"Or����� 3)PA�'Z0���"O�1�
�]�$0z�≐x�\I�"O���G�xz�MFD�%���� "O<uxb�	�lUȔ�! F�< �v"O����?2�+ª�z����yRي,b|�/[�b̌A���yBNY�(UVm� T.�+R�ݝ�y���'k�f��r�à2��`��Q=�y"l�}�>��%o��M8Tk��y�さu��l#A��3ڬuT��yr���>7<�tk�2�bQ�K��yR͔�N�5� �R�3�J��3�yR.�9g�4R�cP�S�3�k#�y��X6t����Y�
L���ꂤ�y���*$W(S�}�X�r0"���y򦖨)��LK��	(�|���&�y��Y>3G��Ʒ&�^<Ip���y�ra�Ŋ�8��x��,\���'�����9�@0��j� 1�����'-��)A+.D�8��Ah�0�`x��'#UZ0��ʸ�S�(�{w�l��'�Dd�JОT�:�{$%��o1���'2��&�Ϯ{`����bVU�	�'�t���H6s��t��
ø�"Q�	�'~��J娅O��0���:�qR	�'�4�0�~��#�"y����y�h\�&vlRCUN7����P��y��Xv�䉲gCU�HHp�{�FZ:�y"��/b�2l˦�]W�`(�B�E��y�]�u:`3� l�(�G�Ւ�y2��@����L=B�X���A֘�y�K;[T@�u�I�>f��ё�N�y��û"oT�q�BO+5\0uC�Қ�yR�̦9%�u��$C���#�ԃ�y2�ŇO�b���S=fu�,C�iX�yRa[�k��0��U_u(�"��W�y�Ţ3٪T�pꜾF��G1�yjS�p<Ѐ5'�%;8<�t���y�h$VZ���`�ÎC�~������yb��N��@'7߶lh�B]��:
͢b���
*�4ϛ�}�tT��2��|�#	$#��z&ˆ0<��0�ȓQIZ<jW�N0����g�7C��A�ȓJ�\��nzi h𧪜��x@�ȓF HY��ۦ0�l�r2�Ҭ~2@��{��%���ц]*�M���T!U�T��S�? �T�6�*=uv��G&^
B�FE�g"O�}ӤoҠT��3&^&.����"Or���M�� ~<Mb��G/��q�"O���`��& �2�˚i=��t"O(�pc鏈3*�͌-0$�!�v"O���,J"$Er"��U8ȩ"�"O�d��ʝ1���`,l�b|4"O�(�V���\���REظ6�J�?�y�É�?z\ٵ�Yiʶ_7�y�b4n��r�	}���HV�O9�y�B�(w������_��4�f���y��'w̠�ʆ�YFu���Ո���yҨ�`�f�a5c��DW�8˲	�����hOq���
�T�t��m�Cn��z��-k�<��_ 8*��(B2}�I1	f�<�ģJ�y�*t��ǁ1]�����i�<�D���lu	��j��`�r�0�i�<� ��m��t@�eZ0yZ`�P& d�<�Í��}��5P�H�$��𒅂
]�<�B��L����E�ܤd�")˧k�~�<�n֨H٦]I���$U�L�*�j�t�<T�y_��#0kxxU�O\�<�B_�g~��c��%*���˲�Y�<Qv��
 	6���Ɣ�])�x�� o�<q�b01M*���&��L����7
�h�<i*YJ@��r�Ji�F�(pg�e�<y�Ɍ�8���Q`�ѶM%:�;��i�<1�-��ic`��6.V���]�<QW+�4!�1�,$b��,�V�<���Tn��
`LT�
f,%�BfM{�<����:]q���;���Vdx�<w�W�YHD����U�\r21:f��v�<Y�H�-Gc��x�ݬ0Q��"#o�< �ҙ~Dxaz��H���!�Dkyb�D.�'C`<���+O))�,�'��B��܇ȓ[,V�#�� L�@ə��d�f��
t$R͏�3$a��)Î�*A�ȓ+k�(Ѧ��6\"<�@�@#�f���# ��r��#R�0�?|�1�� G�]*��E�\FP��Q=MN����m��Li''�~5�����wd|���Kp��8iD�%JFO\F��ȓO�TYUK��W�]H ȉ�=�<����AR�JY2gL����#C�$Ƭ��� �DAfivUtYR.�9���ȓ:�<��-
5d
"�9��G4:F��D��<�%)��3H��0��P�rE��FDcC�o�2��A�'1���r������4a�M��	T8�BԄȓ���yŤ݋,U.�3oE�b掔��M�5���'ai��#6�T���qY�#���j��ءeiV/T9X%��`mͲum���.@�#�d��K�h]��I	dR� ��N%9��0�ȓ�6��)2Le
`� o\Z%v���]ڼ%A3�\gb�u�Ġ�D(>I��Q��Q����g*�a���r=�ȓ�� ��O�7�����+�����[��}zlN D<�OO	�݅�N��I�K�`��p�Iшas��ȓ��0O��x�ppp��@�
����Ɠ#�6aPZ�d��؀U��.V��Q�'�1i��A�Nk�![�a�����'�B�F�f�,l+�G�Y<2R��� �L;�0��IP'2u>�T��"O���̩�p�R��)n�&��"O�p���Qp"��a����e"O�8��^�u�b@���I�t����"O��k��ɫdJv퓐�ݜ��c��|��'�ў�O���B"y��� ��?Oxl��'-��4�Ƙ,�����n�4�����'�n�`�@ 0(U�fFɜ%����'ZBq.�u�Dt�ebP�\�pi�'��;0+4�|
�$�Bh�I�'�X���)�=�p%���աk�Yi	ߓ��'�X1��F�u���0��58FX��'�L�����D�C n��(�t��d4�'$�xU�V́!zh���Z�0���?����j_H�m��DN�ar����a��[:m�F�|�p�ȓ?k8�'�_�f�.ǂm-�����mK��]/�r ��i�O&�ĄȓP�[�,��4��|06o�Gt�|�ȓd��Y�ע��1_�%�BF��4�i���Ɂ(�y5Lp���0E�za��	��,����J��DL/^��U��]�Xp�&�2�Yb�Q+u�0��dA6Ȅ�]�"[�	JDL�I��ч��T�`f��'k�`Uɰ(�|�d0�ȓN)���[>J���s�%��Ѕ�ږ5)�,�0������M�l?4���	R~���C�$i'L�U�v9�˔����?�
ӓ8%B(�gI
�c��U˴L]�_���}��a
Lr�&!s��9Qg����Bh��,�(g�F̢�j��p�f�ȓ^T @�������/1Z���^8T��p�#�XC�4
P���@�u�F�/ɬ�"%E����b��G{�����4��LY�)!�XCbF�y��J/t)d�	���C���y�oS��$P�'.�9i�pe�H׵�y��M�'�����)P}�`*Ō]�y�R9J�9Ǭ��^9y%����yf��:o�Y񥖘 ������<��͵
�(��BgW VQRF(�
����3X��ɩ1ǔ7X�Bm������0?	�ć8f��
��])Tɬ݉uJTZ�<1��^X�<X"�ӊ,�2E�]�<�"BF�L�����V
e��`s!�`�<�w���U������D�3&��F b�<�'��4�i�%g�O2��	7Qߟ��'ў�>��e.�&U�ܤiPj� D����O,��2�S�'@ ��Ғ&:v���YZ>��Rui7D�$@p$|�@�%J�C��HFo9D�4ʵ�I=?��3!��M�����A2D�8"@�Cݖ)�ސ:���S/D���_�(0h�eJ^P�
$��+D�����ۭ
��]��c^7#[��� �5��刟rqȱq m�E�rFx�{��|2[���
`$�-�cV�"��#��-�&C��'&`:,0EL�~Q�hRq�� �C�ɽ}4�I##ҼO�����M �B�I�>j]�@晩P�RA1�a��~��B�I&?T�!cqɏ�
R ��!���,D��:�G:���U�θ)EA�g;D�����֒,S
�3��K�vV�����4D�t�&�MlF`���#Y�U)6c1D�4���
Y����SI˪i���F0D�� ��{��������;�`i�"O�����2KH�bD�� <�&��"O��JL-Q��DJWJ��3����e"Od\#T���9�pК���|���q"Oи�u�IvzБ�I�zn���P"O�)���	?p�Z`.��&w���#"ORA���(����3�eY�Œ�"ODT�A*?9~��VN�XH���"O�X�6�	.�TY=iDe��"O��J� �<<��P�K^�}�"OάqB�6F���5��!c�} 6"O�͹�� �*�u�ũ͜iU��"O�=:�ヿf^��G�7Wb��F"O6�p`_	�PR1_N�A�"O�аG��v���ڕF�%{��!RB"O���5�� @�D�2��.�ع��"OF�{���"�ޠ ��
b�`��O��X�-M{�*y[��N�S%8D�dS�ZN��F���W�࠳#"2D� Z��P8.�TA���"��;��5��N����*<8��v��
 /�Cd�!;
B�ɞN��e0�����x{.���B�	yw�=��*(�j��N�S+�B�N�6Z-*7��X�$H�ܔ�� ?�g�m����d�A�T�P��Q�<ѳi��PB�ǅNqڇ�K���̓߄0:�Zby@}q��K�l{�I�ȓ�z��&��j�����T"W��E�hT(�I��qTrpӗH�(r�y��=��T+�)�4�1�6��D�ح��R؄#��:�8�ӱJ��[� ���������.$�|5�W+E�	��uۡ��(�B�	�23��G�W�HĤE�`��6�C�I�-�j�(gO;~�1��+��㟈G{J?=aB�^|v��EU18f��jU1D��*D��(m�Ĺg��/[!�(��/D��q�)̀:��ٕC��`nnز�.D�x�e㉐�"XbgOʖ u|԰�/'D��A����5�2��"L�r&D��9�ؾc̶���� o���%�$D��q���54�q��(��R:A��E D�(�t�G�y���x�L�}۰�=D���eÂ5>}r���)F�����k.D�<¥��i>���� 6rؠ��h-D��cn�`xN��$�]5R9�\Y�7��Z���ӎH�Eb3

1��5X�(ىr[2C�	�X4���G��nI�gd 
C�I�t�B1��&E���QC�4b}2C�	�\�����x,�DIA�<JB�	�ܥcwad�P4³f��B��]|E�%��iqVI�kZ�T��C�I�X����%k�@�"�x0FM'kJ�$7�S�O�����D��q:�Y��(A)FL�`�"O�� 	o$l��ğ-DV�M��"O��!��ڡ-�aذ��;K��#�"O�(�

al�ݢ�jA�C�2]� "O,��UY)Ӫ@I��!̪���"Oh��v��r3<�вgB�Ä�8C"OP$ɤK��,D2p��%�z�V"O2\Q�Q�lj�o��� ��"ON�`IL�<8Is���=c$��P"O�;`��zA���ѿsVn���"O�i �ٴR�(AJF,&C�	e"Op8�b�̵8G�aKc'�8/8m8�"O� Nձ�FWnnx�G�Ha��ȴ"O`�,�5{zH��5�ȳOX�i�"ODA
�α�mI�n�J�rU"O�]@�#�9@��A��2<��hv"O���P��(K�P��"P�;��5�@"OD��aڭ�� ��b<}����"O�	1���U2�a�^���"v"OT��,�<�E��"�'���`"O�l{B�d���Ёa�(������w>}��.s'�8���6S�ݩ3C1D��J��-B`ɪJ%�xQɒ�.D�dH����9�B	�Lꚍa���Od�=E��'V�%�,�â%����h�4��7K&!�$|!�\�ff�8_���%Ɋ%3!��W&.8���D�"6/�y���� !�$�	^�<�X �/]u2���&U�>!���r�T�����-o��s��W <o!�D�$�¤�"�P�k���x!�7U!���-'�<�x�(�Ov��z��� �!�DV�A*�SU�B3fE��P�㗩\�!�Sf:�q3�ʄp�д�@C�=�!��S�Z7��pU��T�Ĺd���}�!��
/'��B�
=2��hSa/S�2�i>MExrj�<uP��Z����:�,�Hi��y�D *�$�� �4�\� 1�޳�yr�@!*͔i�q�-3�`�̳�y��#�0�J�f	�#�<HG����y፼�F�Y��M	'�x-�iڈ�y�dS���ZD�وP��5����y�(�/�tA�"�#V�=�"g����)�S�O�V� 1�"q2�,+w�ژ���'�$��p/{�Pq�@9�8��'D��{�]��Id�6��X�'�,F�ǣ;�8�� z���'� �ە�M5S�䴀�
��
5�'* T#�%c����4R �t�)�'�6\a��=
�����h��	�
�'�^� ��y�p�3�ԩ]�Q
�'m���4fI`������>l!�8��'��dzb(��uG~*�BӒeZ���'�t��ǀ�N ���5C�\ �'�J��7 �Cr����e�*�i�'����6�Z|c�����k�.
�'����Ô�pkb�y���a���	�'�݁g��6ܙ���'*����'p��6fѹk6�P���(h"��'j�d
�J#p6��7�"/�9��'h�9�
,�@����"
:D��'\�m��,L����g���20�'(�Ͳ�ʫU����&�ZJ�uy�'o~��s�(0�T��FL�xm�
�'�h�A�'Z�6(h؊�(H�8֠��'����Ӆf�ҍ#t`��7�7"O�=B$�W%7p�'�3i.)х"O�Hqphܦ~9��B�X� hV!q�"O���Զ?m�A:�8q>N�j�"O\�2��7d ��L=W��"O�����������?`���/D��R�!<����% ͚:���";D��3�#r�%
�I�@���8D��(֦�!k���3ƚBY��aa�6D��֦�y_�pAEЕҮ��4D����\�����E��/P���0�7D�D1��&D)`IiR-�&:����q)D�� �e��O���l�)�Z�:2"O�X�s@�h-4QzR���;��Hs"O����q0@q)D+͕|⒉ �"O�Y��Ϗ6t(���'ʬm���'�!��&B��!AbC�Q��q�uA� �!�C#8rB�"ǭ��00��"G!�䀏]�Q�!J�+�"�Rf �x)!���a�~���O�y�1�  B
!���|�^@Y�ĕm�B�U�/�!򤙿8R9��&�2|bm��Ü�!�D\�@G>�j�M�L�N*ԍ�A�!�$	�-тTS��ƥ����0.�!�D�*nb�i�f���P)�3mw!�d��� � B):�����M A!��-}O>�r��+:��e3s��9џ�D���))��e�Uf�1
�P"9�yRā�#��`;Tɟ�kwb�(P"
��yB�ֆj{Y� ��c1b�#0'�.�y	�< 6mOW��E�'�̴�y�lR�M|��9PL��Crxx�蓶�y��H�+||��WN�:�RA�雼�y��<� ��R�?���s����y��h�rN7�P)d �y�f�7w1���
�<����CEȣ�y�M�w��y����
�DiS됀�y�ꏽm|�r�,V�Qֲ}K@K��y��
1�J)s0*ίEb�����y�Kޔ����6�ȳ>P �R�/���y��� ���FU�lZ.�(g+֤���hOPc���A$�݊uCX� ����H#D����I5�8����T�r�����?4����hƎ}�^�AP���TT�<!pI�[�Z|��ś8�"����SN�<�A獺m�V��e� 5x�X�Хm�e�<����e��Y2N7`��w�<���ƆF��y'/�0N�Ӑiu�<q�0;�2)�I����3�MZf�<�N�'D$��*<Ě��d�<a��X�� ��0@�;OC��S�U�<���D�����ĺ.z��Pơ�S�<i���stM\�a�&"�e�<abgò8��K��5�8� C�h�<���ԩ>�`@�Ő<��F��O�<q��6E&1�6��` �tR��q�<ٷ���RѴ(x$*Z�J�q�ɋR�<	qoB/P����%�|��!!��f�<�����D����I�]t>�@N�a�<��N�o�J�*�� �]���^�<9u!I\!`w\e��頶��]�<�F�3��,�rX3�R �q�P�<�A*:H{�)�*)pt��
^N�<��Z8�:���&J.��@��\Q�<a�ۋ�v� ��"w��!G�S�<�@�٠^.���&ɴWIX-����s�<�F�� `t���@���j��Yt�<Q�./�4$���(D�Hq�<��C��<m��g����9Z� [W�<�ga@�-�>���g?������GR�<�1NΌ/�*�	�`E�S��Q�Vr�<i�����l�"�G�o�ry�k�n�<ᶣ�.$�$8a�)C"7��a��
�_�<�� 7"�=�W)N_��,��q�<	05ߠ��J�=��l��y")F!8�I�B�:�Ui����y
� ��A�CdD��q��#F")�"Oxu8`/�"��5p��	O�D�2�"O�����~h֮7*�@�"O&<�2@,E��E)��9K��[�"O\�2%�P����QwB��i.a�"O��c$CE�K���0�.X��"O-hӠ�   ��B7@Q.i�N$��"O&L���v�Zģ��AK�U�`"OV�aP�S�m�L�@�:<����"O����A_�s���3^�uҦ"OH�r�o;/,�H�&�����$"O$H0l8H"*R�N�D��`�%"O�TQ����,U�UGf�4��A"O 2YG���8p���T�thY"OA�FP0wS�����%���"OnI�ī�g�4���ދXr��
�'�b�w!�e!J��C�{;�R�'о�v"N(@*83����B�d��'&@Q�,��J[���=�T}C�'��5�a��5T���둅�:��Lb�'h.��sH�'_�69���9�pls�'��-{�E�2u��h��g��$z�0J�'� "�E�	\/pa�ǤY2!_H��'��=;�'��\r8�ċ�p�ȅc�'���š�C� �W"4x��'�*X	�Œ/vp��ƪ͔@��=�
�'�l�Qv�ҹE6�)f �=����'���ar�Z��||����&7��	Q�'��mw�� &ѳ��<�m9�'_���t+{�q @
 ��d"�'���0G�!''hh�.��A{����'��Tm�)�4��cl�!g�4�B�'1laR(V$L���3�H,d$���'��up�K/'��=6��;KFb,
�'�Z���l~u�	�RlT0�x}b�'`V-���J�H��1	R��@[�'0����l�0~�����H(C�����'VU�'I%V�����%T�Q����'�d���/ڧe$l��%�ܹ�	H�'i���:2\yD���T�8�'C�@�q	�=&�3����'��$[�!�>f�nc��H3e/T��'2�@�aͦ�6̡"��'I&@}��'�V}�6o҃OC���1cމ��L`�'Ʉ؈�"%q�b���O�b��i��'r����煈"�:us R'a�^P�'6���'' ��9B��?i@q��'Wt(�oP�ѱ،g�0�'T�y{�B:Zћ�l��d��'�P@!�O׸\!�<��E?X����'d@y��g4�@�`/[�?�$�
�'�J����/���G�O�<%���
�'Cb4�@(��bgX�:��DA
�'K��ЋH�dshݱ��6	`��vH=	��0j*A� %�������%����J�_JP(�����ʓF�\ժq
۱$(��oZ$7��C�	�l�4�����I�U2iRC�	�<��ʳ��
p�	b"��t�NC�~��-#�លs�¹���N4�C�,n:��ʱn�>_6�1� [��B�I�Uta+v�A';\��C,�rC�	�٤����َtaV雵�U�
0|C䉈�:sDْU�ژj�H3 �B�)� XX{emF�]xh��́@�Q�d"Ot�(��)�
��"�*`"��"O���BX��]3F!]8%�Ve�W"O��(@!T g�
��#�;�tl��"O��r���'r��9�g/��!a���Q"O�5s��8�<�@�/�RS����"O�0���?4戜Q��[5@=K"O�����"(�|�S�Tl �y��"O��Ks�+^n��yblU�O� rD"O�����; YhA�Jф*iz���"OZ�
qK�!� �Qj�#Z��;�"O�$��hϊ������(?�]BF"O�yK,��B�\
_�
�AѡեR�!���	v�������c����4	8I!�  Ԩ�P肅_v������U!�K`��1��E�nV��1`�/�!���*w�c �X���� @H
�!�D�6�@P��y�eU/�Py2GMed�Gi�0H��}㢁��yRe䝑#�ф0ެ:�k���y��*#��3 d�'��X���<�y�Fd�n)�4	��!*:�!�#�y����<��Ⱥ�� m�l��DW�y���p
�u�t�A	q����y�m� #Q�-Q%��^��Q(���1�y�f��9��+S�X9Y�&�8���y��PE�X8;7D�Gn:D8p�A��y��1k����*��CSn]��L�<�y⌏�CzXid�
!��H�yr�H�CƄ$��G�]q��eF�y	�%L�A�P�\g��;'��yD]�M���В�=3̝�aǗ0�y��͗���DOt�~�@�����yr�L!�L:e��$i��eA���yR,��//�T��ʣ\rHR�ၔ�y�ؽl���R���*gw�@���"�y�� Nr�0����\j`�K��Ж�y¤�*:@>l���
�'-B����9�y�H��5v  �l�2�4�hV�y��ч`BI�u�
>��3�ѵ�yR҅L:X�b!g.��1� �yL(�`#��3<S�pRQ"۷�y��t��A��ߞ`2�@�X��y�	7T�Ի"g��Sx=�0쓗�y���w3���K�}Ev@p!m���y��6s̢��I�!#�ir�$
��yB+�>s�@��W�$1����G�	��y�F'~.:r���'��y`L��y" Ћ\`�A�v� /�\�����y��q��`�Ĺ�Ȱ�G�Y��yҎ�o���s=P�׮���y�+�7j���l��w��%��>�y��
AdP*�.Ŕ��ō�y�CJ�� 
%�a�l�[�yBPrl��A�FWj.h�T�0�y�&ыbJ�da3˟274���B�B"�y�"B5H>L�15Gř=ft��R@Ԡ�y�*֕Dj�`& �;ǌ����y��=��Lہ�_�15�y��b���y"�R"U1�9��*�1y�k3�T:�y�J�>���BLܘ4���Q���+�y��TṈp�A_(*���� �y��T�.��g�!�0�cs.���y�`ۉh�|�b����E��j��^��y
� �h��-H�����CJ@�x0��"Oށۦ��$
:��S�Ʉ<~zt��"O䵢(B�S��PA�	���S%"O�͹E�Bd�srA÷-���@�"O(i �m�zQ�� �O @ 
�"O�a���j������hu9�"O���&��(	<vm@'+K(>f4yC"O���raZ��@�I��_x8z�')`��p�Ŵ�Dx�nR�����'�X���ƾb�~��,B>$.���'�:3h�<+��<��&��FU��'��18���)O��;T�ȧOy��1�'A��%İ:7��BV�C6F��
�'،P��!¨X�Fx�p��+F묐�
�'	"�	���9V�As��,t*���
�'�΀�aN0k(�Q�R��Cw&�c�'M��Q���)\a�l�$�ln89�'j��2B�DP(<�a�@�,����	�'E�}gB�U���6%v2�0	�'!�d�iŦ��P!U	&I�y�'2*����0m���ڄu�4���'�����:#u`4G�ȿr� �'������<�<h���_�( ��'G�e��Z�� ���'M1f�r�'�ش���_�+G��Z� L)P�2�'����V��8��lB��F��P��'��MIa�G�l/ ��vAW�UP�S�'�h����G+�P���m��V�6iq�'�ȕ0�Рv�����)\!A�'�m����H�b�� ��9yZ���'K � �����P���!|�E�'��͸։L:*�$��c���m�'g�!��Ȕu~�p�ČH�^�"���'�d����x�&y��A�3'�����'I�ݻ"�YyV񡐌ƈYP��'� 1�b�����l�	�@�'e����%�l$tcULW<�\#�'�J����U�.H@���#�<>"���
�'�$����R=em����B)6m�	�'a`���
��D���O8G,j�;	�'��X��O�9�Јi[�F]����'3�@0�*�3HN����fK6Ix,��
�';R��4�*��մnBH���M��y��տOC=!E牁�5KX�}�	�'u�@r�gT"w�$:��� �`�b	�'���AH�'���@g��"�~��'���B�jԛ[u:�!@��v��8�'�����\�N�{�lG+�"�H
�'p��ZѤkC�	[�G!/L��j6"OBЉ�I�>�^q��jɗf4E�"OR��֌V�`�b�J$j'D�J�"O ��F�)�~x2/�&
���R�"O�y*%c$6�f/5ªDA�"O*!C��78n<}H��92�B��S"O������.@�}2�Æ�y��"O�$밦�g��������"O4X�R,\�v�:a8��U8f�y#�"O>��냣P� ��E��A�!"O$�@�dǵ�����,�riXT"O Ś@ �#D��M _d����"OF�$�5.@nТ��M���be"OV�b�!4�-��.>	�h�"O�ֆ�}�<Y4�y���"OF�`p
J;��Q�My(�2B"O� , ��o��s@�c�]�r�l0B"Ov�p �/W�v89�v�"&"O�E��l�w*�\��j۝H�,e��"Oȕ��kԆ|t�ɹ���XfFA#g"O�� �U�S:SD'D2�eX"O�!��D'�| �]�`8����"O���N�������7��� "O~�awN�*q�UH�D]:���
�"O�Q�G��5K�9�dT"h�%"O���
�L9F\c�bV6)BޘZ�"Op��A͏s�<)qcB�a��S`"Ol�R2��+q����∪�0m@ "O6� Ä�Lgν2AS ��)��"O�L1F��!iꙐ�o�\�R��0"O��OA2n����A/J:k���s�"O� C��Z�Y�L����N���1"O�is�m��_g�y�&-�4o�IC"O�-RG�Uߢ� �־��l��"OfTy�3�$�JV��+a㬄��"O���'���0%�t��q$4M�"O�JȚ91�~��u#�.v���"O�髶��,!2$��a�8�l=��"OvTc�%ՑJ������t�f�%D�\��A�aLy#aʇH�*}���(D�D:6k0�&|k���.�	�a'D���b"�m���bS�C _��sVj*D���g��92M�i�Bn��M�B��#(D��#��[6w�D���/x�tyD+&D�`cɅ/D{�(`���j�,�b��&D���6�?f�U�n��(:,ܓ�!D�PR�/Z�O�����G�V��]1R�=D���� �70��12�őf��}"q&D�����v�p�vȞB2�Q*��'D�`�v���H��xs5�ں���3(+D�Pq"#	�W� ��m� `�e,X:C�I�$�8a�2K� X��C�v�"C�I�~W0T	���"X����曊#z�B�	^�tR%���&
�]�7�֑e?�B��,;ƺy �d�*}�-�����+�B�IR����!��"�����		Wҡ�$�	���[#*Ѣ(�j��t��<A#!򄞌5�,I��\�ڂQ�����.!�C� � p�3 �#`�H,�b!��pe!�L��1�һt~��NQ�Z!��&Zm
�)�,����v��[h!�Ę�6)�YiB�L�8�ԝ�^+4�!�<��4{��NnI�׀W#'�!�$���(�(e��_��j�@B�<�!�DGm�-P�o��,�V��k�!�d��z�I垛W'Rj5�W!�d�+�@���g�	>VpB��_�R!�d� %��,�n��c ؤ�Ǫ�!3�!�X� �B��J
@�6�W�c�!�	
�IH�c'u h�AE�9yx!�DſJ�b��o\�T��S��C=Pv!�DH[�T��t��G�Dq�+N<cy!�*�D@�K�����ɂ�3�!�^"r�&��1���(��I�D�!�9DTQ��B���pZ5�A��!��$t���d�Z�n}{�IK!9k!�ć�d��	h��L2w��cS!�d�?"58
�c�_mcA��YG!���/���3�kʍ�nᷨ�-4!��`�<|Z�FԴC��d�㧎~�!�� 
8��ڞr"�rS�܌|�캲"O��i�G�L��-:&��)�|a�"OZ���!�g.��f\�$��9;e"OСb�j]�f�������Sњ�s�"O8��U�C���ps�ʮkY��"�"O��z#%��B��[�aBMR"���"OU`N����	`��3�pyr"O*�5)D4
��Y�[�f@p�"Oz,s��5T1F��\6g�b���"O���bn̜C�t;���<�3"O��+�!�P���G &'X0k�"Oh}�C�N�ęQ�N1c2�9W"O��ҭ��a��H��P�)n,ʐ"O�Dʗ�
�G:,����=Cݴ��"O\�'g�������I���G"Od|b1�Æk�42�d����h!�"O��CGO�/�S6��Y9���"O�Q��-|�����zl��"O ���K)z�<B��ݦQ��9Y�"O�,�cl��j/���Q
,�& ��"O�����K�9.\���	gx���"OR��S�'M�X�˵^svF� "O8|K![�
�:%�&��
Ndڡ	a"OY#e�tӜ�[�G�FP�AH�"O8��w�[&`�u�f�ۋ ���3D"OP ��Gҝ!QP�� ["�9��"O�Xh��	�3O�c��U4wj����"OPH��@,5V�\�#
r.@�"O� ��-�%t ����i�p�	��)D��!��.:�"	SЬ�x�!x4D��6��	bۢ�+VA�8;~�/&D�x2���0RDT�(�l��U�d}kb/9D�H:%ɇ�n���Ka���d$�x�e�<D����O�Sod2A
N����q�:D����G�>�h� ��Ivִ���4D���$�U,����@F�c|ܱQ��>D���e��7v��l�se�*NU�Չ��<D�$�`���z����=�0���F:D��9N
��2r�ȕ$�����9D� P��Ex�$�D�E�""�!Ȁ�8D����*��ut����A�0c�A	&G1D�@�j\q}\b�Y���y��9D�����f	��m��Α
V m�<�t�Y�{B]:�6U��jtvO�q��P�B���[ M>8��]�"Ob���͘7m�dq��A��%{w"O
��	7k7�����Ʉ�|0�"Ot�C� ѸV#�(0�ފZ���"O���P�D���W�܍����"O�!���ˣN��($+��\�b���"O�)X%Ƌ"��ܓc	#GP�5"OP��sn�;��"鋆Q�|�Q�"O��j!�)	<(���qۨų�"O����Z���f�+ir�`��"O�h	`�\�t��Y`'�	���pG"O�y(��J�.A�V�arhH��"OH"���a�r����XU`iw"Oj4x�Iӆ.W`8�h�
3:���"O�٨�Ǜd0r��tC|Q�s"O:�1�@ɀk�\��G�[>x� �W"OHCM��%ն�����?ST��ȗ"OR�DP�/���yg�����b"O�MQ�	�cm����
���j�"OXEb���+n��}�դ;ȵh�"O� hd�aм9�ik��F�:�^YY�"O�ű�#U>2�����bK&�TH[$"On���̺y�LcG#�q�p�
�"ORd�RF��h.j0���C���Q�"O�A)���(w�ڌ�B��?ID��%�i�铉�)��d]d�,�kD���t�if$\��a~�Z���uL�HZ0�B�Z!zT�5J�>	��R�z�ѸRF�뗡P�@q���"OL�sզٮl*Q�f㚬9iƱ)""O��d�	�,����!�$g����x��'B<�"�B/p��J`FK�6�H�	���~�cO-d�"����7r�L9�RjF	�yB�2%N @�@�M+VRl���R��y�)9,���)RO��SΆ< B��y���-��ͱc���L�'��y�gU��y���3G��&)�.�y"�G!0��23m��>���f����O�~ʖ"�"�u-�
l�1T������cg�TPhM���VD.D����@K(8��0��7+�`�B�L6D��A�bO #��P ��k�rXX�H`Ө��IyGqO�">yWb�",(1兓3�`��Tq؞tnZ����c����/�%R1�p1���9�|C�I������X�H�Њ[�v��b��Cő�ʧj@`�4)Z>q��D�f�\!���,~ �d��4��УG�ݵ1�P{�Ŝ��Q�\��j$fQ!G��<$�LpBKK:<��"�	=
3܈� '��4`�[f*E�!��7-���?)e�Q�����$�Y����x��4����<<4	��B̉b�d$�s�N*�JB�I�3��k2�&r�Sr�L�e��E{��9O����f�|���3��<[v�	Z�"O��SmFrZ~�h�-�.b;b9�:O�b�h��43�M T���P<��0��":��C�9l���03�Ҷ@���� �˒M�C䉀�zT�冑�5"����A�-��C�I+p����Th��ʍI���I��C�I�삵�b)	�^�L�%F��gH|C��.#Ct�z���X�A�Ӎ�"@<C�	� O�m�U*+e��8Ql�@��B�6PK� `�03�.=�B4w�tC�ɘ\wN�V��[�ͩCj�M�@C�	�~�01�MX"�8�ń?.�C��"0 �G���,��I�_Vv�I�'B- a�J�*8��*��_�{�4�hO?7��9�� ���%SӰ�ؒj��_�!�$K�B8&јQJ�0�r�$�ǑI���HG����&7s<�p�@� M�6�4aF�ybI���2@Z�'S�4F�ԡe����~29�S�Ow��@ �#_��8Z�*^�M���
�'Ҩ�2�NĮy(X�2L!F/,�kJ<�}6sѠ�k�����9�"�Fx��T]���)�Q��А6Ƅi<�l�!�Q�!��Sr���/L�d%"��T�t�Zi�<��Op�E{Zwp1f�)A�^1��E����lÉ�$>�S��@���S L\�0�
0Z�LX
�y��9�= �o��^5�6G�~ˎ�=�S�8�?9�3���dC��cC�m�'�ax�bǢ0���a����Q��ԧ��=Y�y�DNq�֍�3����E��yrd�Q�L�BD�3in=;�JI��'G�z��
i"���#+>$:fe��x��5 �9��5����-��֦C�ɼ6�.u`�X�s�p���N-+�zC�)� �EPG��<\�T��f��"`v��`�"O�eCe�./Apy�5��Yt:E�"O�0����^HqZ�(ɦ2�h��HRH<6�C�s(QH�̗4Ք|
�l�H����>�U��)r���"��N�fd���G�<���)G`(S�H�y��иs	V?��{"�O8"=yRɏ�w�h��Z�H�t@`�lHg8��&���e��#� I8�iDIkX�2D$}��'�V� �Z|��䍆M�x��d7�S�d#�&�*-ғ��"�0C�-�
�y��@�v�HR! �n��O�۴DEz���'V��EHI���1�ԭKM�i�'o��s����~3�EaaO���q�O����K9N�T�ٸ�n-�ՈQ�.���V�O�2�胑j���c s���"O
�ɔ%�f���"����_��(O�=��r~�%�r�V$Z�����kꜰ��n� l�a F�`Z���/dC��ȓi�L-����
#
|Yg�A�R
���_/>X��а7�ư8����d��ͅ�cEtx`s)�`OV-²i۠[�d�ȓ,�X=t`J�]�x�E�G��,�ȓ\Q�$�G!��K7r�Q��Y�m��+�~x#di.��-�RI߂����=�tpw�D�3�&�k�cPdc�	�ȓK�(|)c�8uQ������;xl��ȓ\�N�7b�o��y�s��55�-�ȓk���#�%A��rh)0�����Un@�%%��h�@�.v�� ��m@�ď�>G#Z���	I�����ȓY����Z5/.�h � C(` ̵��r�J�����| iP����^���;���ڣ�+q6DD��>B2��ȓb��HB��?��E���H�V���ȓD��"���;y)�h����.���>����?m��$Z�������^�X!�^�<1k	�'=���@��,V��@0�)xD�ӈ}R�Q�Q�P�'O��!�͞�{�!8`.��)�'#�-C&��9h�x�XǠ�.E��'�ι��D���#�jJ���(��'�����A9��!�uKE��>e�'��@�&��9t��J�gخvW�H
�'�L@��2�^��&[�oK$��'��4!�˘A���x�噠c�`,��'H���3��5�1IE�P&�h�'��IJ�I҆����/ t��'Ԧؚe��������Պ(�Y ˓�(O� "3hf���a�Q�=)9X�"O\ũvj�,5N�((�!�22�
��	T����=�q�Q���h�P�P�ޖ�!�D�"	�PȠ�f:(\zL �#ѐOk!��	id���h�`?�u��Et���Di�&�8"��)�cV��b��ؒ�"O� �!��N�$�xRG� W��E{�"OjuP�gäY����e�K4��"Od���]oPTG��*�Id�O�=E��(�n�~)æ�T!6o��5�ރ�yb#�.#���bN�,�d\�u͙ ���BX���f��1\5ƌI 	!��H���?�OR�+?�)�� �t%OH�V�$�ȓ@t{Ee߭_nĐD�Ǉh���,��J�>yŀ,��
UN2�����0�%O����i�ࠊmY$Q��9�앰1�.�,M$���}��4��S�? ������,:�^����41\lM�"O0�(҉
	��J�N9
�`��"O��(G"Z#-�Rlb��@���2�"O���� ��$�	�R,xT"O�CUf�+���j�EǾh�\@�7"On$�g'�4r�ȥ�Q#Q��j|"O^IiDa�6�����W�ܖ�$"O�pX2�C�.������v9��"O��Y����*^��0���Z�""O�MpTj�=}�I`�/�2�-�"O愨��L�>�$x�,Z��Q�Q"O6I�Tk�!5��\�Q�J'����"OK�Am L���.��1�&�y�ȅ�&��cl@
WA*�pe��yb�\����M]�@��|Z�,�yB�t��S�OX�=А�He��yd�mH�"+L�%D�ȓ֯���y�BW�S;�+Vg&��r�,��y�OT��<Õh�8'����MF��yb�4�`��E����f8p�Y�y"�?3�V ��nK(/�n]�R��-�y��9�Q�č�+��(Q1
 �yr�T�n&�$C��G��<,�S��,�y2�Y�B��$��\!c�pc�0�y�BH�G�r0Z񄍬&��L�"��6�y"� 6hZV�����$־-����yr�9J�b�Sbf��j��E#+�yb&��<�\�z���8�b��*�5�yBfF,%|�9�Ͼr���y�*�&a��I͆!w�eza"Q�y�hP�1Čȇg��.�4]� �R��y�iј!�0���gΎ"	� C G5�y�%pz!qC�� ��a�����y�h߿yi M�@b_�
R�(���V��y��_VC������-s���eL���yR�^%�D\��eT���$�G��y�AICyl=�ga��LO�Ԩ�a(�y���.5opmi�K�jI ��ӆ�y���
�dJ���[찈PMУ�y"@��^E��IA#jԬ!��V"�0?!��P�}"�Z3@>v�>��%�ֹm|8���Y�<AV�6d���*%��9J���"v�0T����K�3ʄSD$�=+z��<D�<�S˗bu���U�\�>G�H]!��,:��ӊ�Rg��<Z^ʍ�"OLU@o����vM]�3�u0�"O�5�'���n2�Qc�=M�а 0"O�u(%�ʷ(d,$�lD�G�K�*O:��u�w������i�����'��\�.�����"X���8�'+��s e^c��� ���,T�� y	�'�ܡ�C�#m�8)�o�Yd29��'4��I@�/F}��R%ͦec�'9IY��f�h�ѣ�
�x��'���ˤgޣmlh�
�JY��'�h����^9���6^�w
�X�'��yvc[\�sf!���n�r�'�8��&���9���{�'4���/ŏj\�ď�V�Ei�'��Ș� 7<~h�yc�L<K�A�
�'j�:���#=�b�zS#_#<q0 �'G�a����\�dMysEϨ4'^��	�'*��`���Wт�qB��!�^�Q	�'��m�i΀B�<U�$9!�hi���� ^aR���"�Zɀ0H�:Ф�SF"O�tXu��nB� X���X���0"Ob"V%�$h8�8tF+{�\�e"O�Ԛpa��k5N� ��{w�iSU"Op2��Ϫ=쬰2 k\�P}��!�"On�'bƌ;�b���;cj,4*�'����烶��U"$�6{��e��'yp�E��%o��RM�z�$z�'?��уO�3�t��W�BKV P�'���Zĉ
(Î%#�oK��	�'���[�K�x�� �w��8<��`�'<1�f�m�v��@�L�pH 
�'0L|�%N�q�\Qp�F0`z�j
�'��3�ŏ���pу�x�r��'�$k���lW\mP��h��x+�'F
@;�e){B�1{6��Zs��<��I�=�(d�s�Ȯid}��b�<��j�31�Z�ʠe��f �:��@A�<9E� �X���q�%��r �]�4��B�<Ɂ�ԯ1�R�KRǛ�K�pQ�CM\[�<	P*N�x�lQ�V�X�cH1SAF�I�<��H.P�([5b�<p�L�SN�|�<�'G(x���0�Ð/��+v��=jsv�&�;V�}�g�䎛O,b�bv����[�!�ēL:I�CͱK�L5 ��S- f�Ӑӥ{4���J��}�����#��d� ��b����I�W��T��¥�6��'�)�ĸ4��Š7";wPM��'\,��@	=E4ep�DP<aR��L�`�H�}Ȱ�QE�O����!D�S���y�aIt�fQ�'4��Xd�2)N ���=���c�vDB�1��p�G:�3�d�,U^�$
���g����D$�@��֫,��mS�HH�)Q�I���4i��M2�J5��l�B�>�O ��j�&�ԇ�	y�����'L�8b��Q@+���[�T�c/B�F����䍦r��ҧi1D��"ů
_��Qb� ϼKPνi�K3}�D��}���+s('P��?�)���, �5�@͌f$����+.D��[%�hP�0�fi�Q֎��ǐ86Vh4�.ODQ2/������-��'eN��V�*l�Nh�ēD����r#P��h�Fi�^0s�Ύ�.2(�	!e,�O�(; "u�0L�e�ض`�\�e�'�4D�E�X�a�(�$���Ҙ?ǖx¢�6��C�	 g,"�Avf�Co�(���Y\�lB�I�SF��R���F��a4�V�sBB䉄uΪ!7iF�4�8=��-h8B���ƭ���]eZ'DOv-B�I'5�6Y�r!�8-��x��G^9
��C�I�~)*�*T�ܼ�����(YB�I�|�`	����=��@ЪV��C䉖����!o�k�������"������#��a��46��Z�AR8@VD��eU�=����x�.�0�+�j�V�A�Ę1���Ez���NR������ �J"��ɚթ��~�������)AP�˒���S�ݱ��[�b��F*��3[%��h)�i�M� `��O�Up��X��x�ĄS)S+���$�ɴj�Ty@��-��t&?����WN�� &�H�Π�� ���R��5#p]*V�'���JP�[��j1C@�85<)�I�`�I��iֲ2��C�O�O�ؓC�I���b�M/G�õ`��F�f� %-K�<ـ�:��"a�Kư�)�����`�tbE�#�bD tN�]j�':���;��	Y�νwZ*��@Oֆi8� ��Ik?��P*��N����皵2�E��+[&i��(��m�0t�i{n�t�d��b:��?�m�N8:v_
Ry8é T8ў���,��-�W��C�O���, 	Z���N��;KR|��'�P���<rԤՅ�I�'haIU���z�����d�e����VW���w.��KEhi@��'MMleh���% j��#�����p�Z]h���1D�� R�:�	�,���!��}�|\q�Eo?q�eت���E���9-t����V�Ɋ�ywF������� .�P�+W��>YՋב0`���!Ƙ�Q~�+v=�� rt��/3e��8Ձ�c�2㞘��哩���A�:`o��QI�.^ �E|�!_�[%B�zWL=�O�&���ٻDW��r�O�7����'?���3h\YA.4�wX>;�p�'���R��B��ݥO�>A����C�`tR��alj1H�?D�,؃��c3V|颢H����A$�<D���w��1Ndh!��p�i:E?�O�a*5�/�M�!#(01�0��^�YM^�:�HCz�<1���( 0�h�n#o��ZAD�;b�'��Ja$�;a�ɠ""3����e͚� �&���a�h�xe+�w<�EM�4FE���H:&������7L ks�T8��Sr)Lq�Ă)
~�~�I�d�d��FK�alt���:{���?9�Ϛ.z���E������ƃv�
 -T�x�x��ެj��D	k�^��S�*�0=�#Ō
�j�j�D7j[�au�A\y+aּEY��T�sq��cjـ>(t�� ���H���4X����a	��y"�T8T��l8���_N2@a	J$D�S-Oz-�P'/L�`H�?%��'\�ͻuZ��Sc��J�/�	�^=��Iw]�(�$��.e�>�Q�撦-	2!*ѫ�N>�RV��`o$a�Oh�,�����?)�B��,��P�Ng�(�!GJLO�'(�h($�C�<e�u�@�?i�a�j>�i¥���	VI���p���+��-x�'Z扠զ�4�%aD�{*��a$ZyB�S���=�TO�jq�\��#��7\셰5mU�!8�3(�*d��_�r���O��b�ŗgR�K�'[�l� ��뀼/��ɟm`��;����Z�e�����V�|��U��]H�,F~��SL3a�^C�I�T��	;��: ���K�
"�n-17 �1p�2�;"����8��ҟ�K�;!q��d�	ia�ia6����]a�j�q��x��Y�k`
�g�x���#�$�9BEԧ-<~��B�S��/R�!QHe���9}&� ����L(�W
I��j|Aq��oK���t�n3؆4�t�Hz��Zc�1[�~�(cKH�.��`�w�ۡ4���իǉ3�a{.ݝ,٘QE����xIR`���'K�
w�\8?S��j��"~���$��p�ʭ��e§n���A�	�jT��"�W#3�!�dȫ	�fm�s�#WQ@���`J�ya��� k�4=��"��(:��g�*
�jy�c��$olމ򅇂�2#<\�Bi�IK�as�-D���E�7
|�Y�Qʙ�Q��	(ʑ{X.H� g����zuX������"�I���+�'��h	b/����ԛ�FO�Y"�\3
�zP��Q�E�mK�e���592�Chѭ?V �!�@�?��hã��횣E�0az�䏴6M�h��G�6L��j���	��'��=�:��qc�[)�:%Z&H]0d( �s��S"D蕣8T[8E��c��h 
B�I �bEX��u2�蠣'Ae$)�+� #zd9�я
=�`
��zm`�B&����[�d��~,�:P��{7*��.�j�<����%�H=C�Ax��	����m4�9
U�tZy���m1�ɬ;Os��u,��T\1O��W�'��f턍~׬��p�'¨����7��Iҏ��Hs�4₨T�"�5 ���s�ɳTg�#/�@�rQ"ق�����&G�Х�D�D�+���#�&ω)��O��aEI�����ˈRj=�WdMVbm�􈛐f��`k��!, �3�k�>B�	,7���c���6=�]	�cΩC6Z�jh�eW�H�c�QB=��2�6���k���2�j@@C5��d	e ��>o<�+"OĈd. �<�9UN{��3�J�O lɁ㚑P��쀗G�?A��?i��& ���H�.R�ze�(AR�f�'	0=v&S@yB$L�5���OD�`�O�$� �(({�a�� �
0����Uܘ9�@L��[x�`!P�>�x�-�2�6˓HG��j�6d�.ô�6���{�,9QbGŶEy��J�'�;Az��ȓ}���q$��150����A�c������F��sC#�."��?����憘\F�Oڀb�/�"ou��:U����HC�'� |�f�kH9���[�/��Y6k�Ojx�q��=��.1������'�h�Waϩ����C���U��1
����E<�0O���(�H�Z�*Ƙ|����Qfa[��՚1"O�(�g�+h�R�h1F��axlʣy�0��"`V-��)��<�󆁧W�X�4NTR̀�qL�r�<�(CD2�lP,�8��m�p���<QtH��+@�?\O����: 䱫3�)��\94�'�B%8�ˢD^A��o��������9>���7�y
� ����"Y.e���0�/�BTjC��"Aj����3^�Q>�8��&Ҍ��2��<FO.D�HC�*6w���!�`�(�0TI4v�H#wn���S��y���h6���̻X2�TI����y��`k���"+��D�TX�bg���y���(�l�z$	�e�����?�X��&JO�r�|(��)�O���e ;$'F7-�,n�HP��էa��!i�X!��)l�>pz֢��{�� !��ދ/0��x�a���q�>�;�$G#xb��󊑞<�$D�t�&D�����+��0�K�3eN�4�$D�Ы�*y�4������lL� D��z2*��c�hHbPE�E`I�A!D�P�䪛�N��I��+#r�S�A?D�0����hd)Q���B�`DЋ?D����ě:�����!��I�^A�M=D����fJ:���a�� (�h�R��=D�p"�*$x-�p	�t����G�8D���蜁b��H�����(,�I4D�lC�˄";%��;`)��m:p�5o(D�9���u�nH���I�1�<��&D�\9U�A'W(8ɠ-8 ,��p"%D���S��qP�pj��_��� c/D�4#P����3FEޚV=ָ�ӄ0D��bq'R��4�j A��1�����.D���R�]�4<�	qKP+EMF�I��,D���@�L�Z$,i�&��\�4�K*D�dHd眩.����HM:qYڴX�2D��zs��'�6�yiL�̭�*D�x+��D�"�X��P"��9�(D�ı4���;�L$ �3�C#D��(�:���MK8e�@|Y@�2D�آ�E��T��"�I)E|���0T��2�'�~��ī�W+"���;�"O�Ļ@)֍-.�9�֢ߢ?��5Ap"OF�ɣ�=� 	V�Ţ'piؓ"O$�����qj����D�i�%�"O<0p� -��|��4vF��f 0D����B�� 	t
2%^�9�5��L.D�����T�NS��HDk�/ux1G�/D�1uč�-n� fĂ'l��+d&+D��[F���$�4p
�d.E�IS�(D���(D-HY^����'٫�$=D�@�@�]:$n�}�Kω��1�%D��Q�̛+�^4�W��c��ɸ��"D��Se�?U��|�SG�2��°�>D��@��/)�d	�+\&��9p/?D�d�SƏ��|E1�Ț
�fC�B=D�����I�_��|!�c۬=�Bx�&
?D��"�� �J��֡
��!!u,(D��8�I8b�.�S@�����b�y"�Ƕf
�=��@E� �\peN��yB�ұ	�l���$�h�,��y��3�BY���̂�Nb$�8�yb���*�[�d�۠9�t���yB&�:"Iw�UK���d�M<�yr)�> 5c4AL��s��	�yr�P�t`���1,� 8ӬPR3����y2��O.�se΁0����"K��yR�=KS�u�)�*-�5
����y�ӄB�]B�I�g�D;Ņ��yb뛭8��c��Ņe����W��yr��$��c���%��Rtc�y�[�mLf�Ȗ�~��)�b�Ҩ�y��ۆ8��)�J٤k�Z��%-�?�y
� ����Lj9�(igf�!�B�1f"O&�
ֈ�:�
$y�c� 7n�aA"O��i����@�x� L�<�t�q"OJt��cXXsvO�9#���"Of�+��nqy�/Z :b��b"O�	Ca%�"f�
9;�N�c�B�6"OY�P�@�On��s�K<!�^�8�"O�Q�r��"B�^ 20K�,@�A�"O���L�T`(�*�Y���D"Ov̈ �)C�U�wJ�$�"O" ���A���Y�`=4 0#"O�ɠ���-h)"���n�7+)���"O�����ƙ��q;,�"!ʀ:�"O� '#�8	�,9S�l��CΉ��"O��"D����Y�3�
�p��"O؁J��ʟ,�����d`�b�"O&D0C $q�����bD�*۴`�"O0i0�'G�Pj0��!@�a�b@R@"Ol��T`ATʰ-������E"7|!�Y�**�SR/�M�x�E�J56!�Y�/�t�S˙K�D�0�,2J!�$ުD@��� 	�41���;t-˲K�!�䞿W��\Ȑ�T���5� ��5z�!���;��`j$#�+<�p󵄊�>�!򄃾I㪹�2����ԃE�N5]!�D��E�7%ң�a{R âq<!���"�9�`˙G�`4ó�]����1�|��B�\���rRhz@l�6jb����"-D<�ēZ�08B���[�MJ���~�H��sJA!a��U�9�O�8)3�C/)4d�F픧M������'��ĠՊ�4P�:��Z�P���ܙ��|8��M�-���B��=D����ʛ nT)�I�'?� �F'}r&K*j`@���_x�?�YT�P;	�j=�$!�N�v��G�'D�Թ1@�XO�J��"{R�V�_�	��-O�p��Z�����g��I��i�)ha�asoH?:�xi�Uڪ�ɕ&��#I��ۄ���X��1Ȅ�̛Zf��Z2���̰>)p�SMbp��PfĬQsV��k[8����B��^�	5�l}r/�57��#��N�]&Z�`��!�y2-[���y�9 z �aC���p������mG��e��RI1�R�04�+�bć�y�ՖE�R-
�F!h涍Z�&ΉTuq��<��E; 8�>�O�=����A�
]�ӭӱ<."�ѱO�9@CP
R�85B��ȅh=�} ��]<&5�%	ӣ��>!�ȐY����	�C�L���k�Vx����I B�H��'�b!ص�C�L�� ���L1H�0	�'���4B�9��3 FT�W�jQ��'�L�" �u|:)S /ۀ@��
�'��0��-��|����+V<���'o��Cr�6�z$�O��V&�0�'�JA�8�����@0��$:�'��`��d ^� ����}K&��
�'�N 䂌=i�F��#��@S�$)
�'�zx�L�QעIS`��=e*p	�=g.x!�g��Q�E��x�~�9sG�z��� �"O���� "���-E>v��9鉱qÌ�)�.PQ�O���Gn�'($�rV��>C�`�	��-�v��._�$Չ4j�-�@�2A��A,lXQ��K����(4}���d��?94��8��a #f��A�4�[@�'���JAԳe��D��������0�-�8>��i��
��~�e 0h;������k���Z�����L����0H,2n�rK�[V(��&��%�"��Sⓤ�2�&3\��m� *
�s��j�G�0r�6�"O���@�Ĺi:T�\��5J�,}�����m�ҠϪT��Q�#e4/�Y�H����7�l�ա��������I!�%��'#�9��FW�T�Y���r׾�1���&z\k�XvYA��Z�-�<�Ҋ��S�? &�+���� �`��F�.f����K��Q� ��q������$��9uN}3���i 3e���~Rjp��eCpfi��<�@�E0���;�eZ�����`�OX��n\�V��a���~J|����	�$�`�	7:X���[�E����!�Q�C\C��\�L�"Q#ƗXx�hRq���`|�<��'3�܂��b-���A�|#n��I>��7�p!)pĉ�m������Ԑ;�Z�*�'�^�`�ד@2҆�J2,�D8Å�;LH�H�Ń!n��(Ӳ�AܓFT��|jt'E!�$��u��2'`\��j��O�� �1��rF�$��		/G��`��6PS���Qh!�$W�t0߅tJ��`<!k�D��8�*��sBĿ��)�'v��:�*Q�W�	�]!���cRFUˢLF3}����S<A4
̈́ȓw&̠�i�� ���ܻW��(����V�� hw�i5DM�r�b�|r�ύmCZ��
�'��H�ĩ� ���2�8С�(��
0�4���N�^�$�0��w�r�)#�� %�� jò ��(�	�'�vVʎ��-B�LԠ�y��iD!(�lH*\�(<�$����U��M@���(R���(�$bdda����5n�RXD"S�g�����O�b��Ӈ69FT"W�yN*0�n�2���)r�b�#��(u!az��I�hT�S���|4��;�FK?������0F��.���>9���x�n%A2-އ�|fДR��)�"�)�!��6z*0q`(��&���,}��H�W�䳠�S�4��=�7b��K�Ox�C�w5�+�@�m����&����@�E0�=K��G�$9��E��;ayu��&�� Wd\��<V^��N���VdF4~�q��&J�":9Ƞ(ˍR�Vܘ�����O��@D���*;Ruc!#>��
��7�0�k�cF�.�1+E��y?i�A^�9V-@��9LO�y���d�n���-3ox`��]���U(ǦF�ؔ���Rw�'[d���B	�-6ڔ�$��	HZ5�w;��b�6D��k#�N�!}�QsA�N-U������84��ʓ:�L�&�J�U����%_�	��yg�߾b�,"�C?]�|ҥaP �xr��?`|�XTmۼ]|Ј3�a՘S���X���GӶ���'-h��#|r�.>5��1@IW.5Mr�ie���p<9F��%\��<�M<9�i;,�<��[eı�qf�@�<��nQ�����1G��V�)$�@�<�v��J�n�Q%�
0�&�POCyr�*� ��I�O�%1�iǙQ
L���0���$;b;p��	� P5����F�t�ڴ�q����e�r���;.��cn
dg�$Eyb�f�|��ՠ]G�O6�*��^*E���@/ҁ\-xQz�'<Q)�
T��d���P�v��q��q�T= Q�I���)�矌�GLϻS�����NO-�Ni��&%D�X�"��}ĝiV��#]��3�Ǡ��sP�M�t:
���'y,zPΟ�=���Zr�֥W1���[�P���ҜH�(�ԋޭ::����Z3q- ��v/D��rWbʀp* [Ҋ�0�.a{'�1ʓv����Ks/$#|J���K��*fn��h��7���ybHC!f�jq*RU�s�x(�c 9�0R뗥'\�)O�"~�Ɏm�����6Fƌ�ȄoM:U��B�	�~���"unVF��U��c��O���I�r��,��l�>Raz�!�	��ڳ��>#�&��ѯ�9ܰ>A#�q�0�3A�@� 䀧� /,��ò%>x�!�D�K����ڼ'} 3rў�Y��"p�o�`��aH�|����hب"E�B�	h1�ܑR�g�r�Z$ԁKX�B䉅OvR]�u�!��]j� R9�#=i �B':�,�}��/� �'�0T,j�n�Y�<	@�
� ���!��E$ \@�`�� %��#�iCNɧ���BX�=������Տ|����n��yZy��M�h��9S����NQ�$R 牔<��U�[�@�r�m|@1R�nͥ`�Ne[�\�X�l(��I�g���C7<�=�JV5f�4Cd��{�`�S%�#D��Ӡ�ҿB��ɸD`DfV�	��<�@�ب�g�'|���|2�˵	V����)��EM�y�<a���e��������b��S>�r	:��
+}�ӧ���� �)JS
&�ʡA�d0N1Ba"OJ�����?BhH�E�q9p3P=O��C���V��
ד��5镄!z��<QN�#����	
r�R(���	o����7o��*z�/�.B��)-D�P�l��3�0	� �T&q���!�/�~�֨X�rb>�|*��d��Qa�wl��X��C�<�0�_�
 F<sC��8��ѣ�9����"�140^ӧ���d�0�n�sҦ��b�}���Ϝ@{!�DA-6p����j�;kh�qf�(��$HK��}��&V��p=9p�PF���2������H�e8�ڳ�أc�
l7'x	����ol��X��ۼ�*B�I�^�ً�]��,Q�i��$�B#=�4j̯y��}"c�<R���p���kB��H�,�h�<�"��}����SB�U���E �e�<)@F��.��3�ܝ�d�ۢ��z�<�4�P�<�|�`�(rM��a�|�<q�l�D$��r��-5���j�E�<��h�.న��HD��ȉ��K�<y�
X#YgL�(5K���`J�KY�<1R�Ϭ�!�@�ku��9��Y�<A��P�H5	5$�~�Vd��	�<!�L�|�z�˘�m9 ��.��<�5�M>j��S�	w��+��x�<ё�V�~II�"ǆAB&�˱#Vy�<�0m�"t=��^�#�̼�3�]w�<qb��Ҵ��oł1�ʔ���X�<1�IA l[GL�y^`��fMZ�<�у�I�.�'�W�f�����(WR�<!�Tg�j�H�-خ]-h(
G�J�<YO�G2��A��¨	��!a�͏o�<�� \�"�u���]˘%��)�n�<Q��N�dᜫ�v΁����'��q�m_|�vdѫ XpQ�'�X����F����+�U�ru�
�'�B�����'�����.�e�d}��fʈj��t�(-�w�>y����ȓ[��"�>J��Q�?�d�ȓ%��=!A#��l�@A�B�2t�}�ȓ/�>�s�>1�D5��;�b��ȓ9GR%F�E�/t�8LV�.CrԄ��ڱEy��AP�g�]�n���c�X�SP�NzH`��Q�g�|���&�x�����YM�,���C�P�,���#�"E�G�W�Jl� �E�o{�I�ȓ-&� {f��B֨�2f�st �ȓ����`H>3����-ْN�&���J���[%ˈ���08��bl,��ȓ^����@�y�tC��X�^"E�����>ŃR��0Px��6 2jE`��͌i��$��w��AB�<�>!���>E��aXT��d�!Q�&
�<Y�jZE$�O?����A��"�%�p�]�G�\=B��I��������蟌�K�S
N�nq��+Ȥb�����~~"eIĸ�&�g�!Ñ	E�{��c?��6���ޔ�Q��`��y��gD-�?A!�	D�&K�'N~D���q;��9wo
�*r��(Q[
x�F�3��IaCe>$�e�S�O�ҥ��E�%$��D̀�XeV5·	�~]qO�ᓰe^�X��::���ա�<Y��=�@j^,�a�4�W4|:|pAC��:R̚!�ĸ��I�(t�(�%c�	q>a��M��=�$�
�:8��D��~� A�P1��q�e�T���z@�Bt�ٕ�Ԑh��ܷ_���DY�D��Y!�n-}�����(�TG�?IS�E:�gP@�f�G�HtF��$��ȸ5�:�$<��<b�s3�Չ���*�l�#j��	+4��;E�9�X�CӢK
��ap����9�真�#���iz5z��9�T���[�O�8S+�{�r��<O�a��� 3�`-��\��D���O�V=:��G VL)9��̘`9�pbŃ�^xh-O�ӧzpj��|d��3� �@9A��!]�d���ɂ����;Q���
2���]�>-�0�%�Z����  vp���Ւ��Xb���8�}��J��Z�*���aJ%��Dؒ�0|Z�Ӯ#��d8`ʗ�M���3%/0�2"]�\j���Tua�t�&1T�ZA(ˊ@T�XZ����/V�l�cU(��^a��#�&�ԀXV�Nh���������'�0Q���Ol&T��v�v�z�#Y=O�e8I>q������Ou��#�E!ch�Qs I T�p{-O���1g-�O�T`d\�D�XS����'�AXt"O`eq�O܊K������ L�pı6"O�՘������D�#'=w�
J"Ov)���Ry훱kԥtH�*q"OR������[!Z��D��9rr��"O���Eܼ\$���Uv[��W"O���d����%3����F:[6!�ɂ7î,th�)J h�k(��~!��X$a��a��f�˦�޷e!�d�&u�u��oA�v2��#e��X!�d��d��#��yf�qQDϧH!��>��9�aΈ7� y�i�/U!�2(2@ر�t���cSH�zA!�Ĉ1U�`IJ4�5�����5z>!�$G�\��l�8��a6��!��5MY�l*�C��b7����!��B	���[ǀ�.�0Q��"Zh!�W�)В\�eN��r��Vc��y!��Y�}je�Bf��y��P�a@)'q!���E� !��KK�6��׊M9�!���:/DeRr';}����#�!�� 1,����
:A�Ѐ4Ψ+!�� 2p��7b
�.���E��Y"!�}jС$F�*ء����/7!!�D��-�ީ��À�Z~���퐜\�!�XP�
dI���(Ђ��!�G�zq!+]�m�����a�(�!��p$(a�b�È8�(�Ca�*Dr!�B�l���[c	��f�(,��>gT!�I����8�g�7�K��w��t��'cD=y�MK :Â�Fd�-vAd@�ʓlL�%���r�~M��Q>��l�ȓ7^>��r̃��ԡr�l��J[&���9�@�Ais�1S��
���'L�9{�� z�ְ�/E+l=r	�'x&�@ǥK-Sp q�pn��'4��R#�U��DTypHŎn]i��'t�;��Do��$!ܡk:��(�'D�[2͗�"m~X����O4:�8�'��,#j���	��ID��H�'����K�F����Q���9�"O�)i@�2Z��ң_�/ah�H�"O��mY� h�b, N�ecF"O�T�� �r��(ᄬ�<H&l$;�"O�Ma� �?r11��P�{�ZxJ�"O�Y���}�41�C��w�|8�6"O�$r�BA�bHc�B�qԨ��"O*����;Lva��F�/\i@%"O��A����2���)p��"O��[��wf>p)�I�)ϜZ�"O�@��>�jx �8F�� "O�s��%�iap�^T���{�"Oȱ��+�����X�>X5��"O ��cE�oF$�D]�J���t"O J�	��<q�d&>e.�F"Oz�s��K�f��cɜ<\�`8�"O� Vd
%%�"t��e�#��;�d�9F"O�O��z��ap��b����"O�b�ɎeB.H�Dю$���c�"O��;���."�*!���@1q���*7"O���r�ށ�n�
��\�q||��"O�43քV=$���Q��( 0��E"O�A�D=`��l�@<ر"Oppb��ЀC����e�Y�(њG"O�г�N��fZ�M���C�D�`P"O���v����`�s��y�$3 "O��2g�ׄ2��*���4ed,j�"O<��D!ՠJ V0�D��`d�T"O��(���<��y��CJ�`>���f"On<2���s�N�D�
2>�г"O@	�͆�q�>�j�(�=n��Xf"O����-�"r?N��H�1eA�"O��ǌV*3X$�p��|O�@��"O�ł��\�V3@Y��[bA���w"O�Љ"��'�0cD�=|'����"OU!��պZ����s"_&=ֱ�u"Ol��#��
<��6c�%�k"O���A��) ��{6�ԩ���t"O�٢Aޮ,�2��B�� ޞ���"O�`���ft�Jǁӥ
{:�"O�̲!�"V�cEV�L��"ODP�q�Hp@�IH3AY�/�.zt"O�с0U�vv\H95�WXq�"O�4	r�"�@�@�D�WJ�h%"O�\�d�����v��:R�Ȉ%"OF,
� [��Q�N d�aa"O,a���ۧwq$(�sV2B^��`�"O�U�B.N�mg������3lC�y"O�mZ�@n�����%J7|A��"OB�����N�;�گv*�A��"O橂Ĉ8�̄2e�?��[ "O�)��=o����%�*GjZ�A�"O� X�eR�}�����ы+r69�"O� �ԩ\�|�vD�sV�][�"O��UF^4N%�AA�o��L@�m��"O��� �E�����":.��"OTc fU� !`�b@�$�c� �$�yr��f��r�[�օ#B��
�'jLa�S�~���!���3_&0��'� �H�M.]w�U��o�1�����'�Xɓe�I%,��)�u�X0#� ���'~�1S���\ b]�@��!d����'�bX"��R�sa��� �M#~Bh�'��:wnF+�\�a�DQ���<��'�A���؞ #'c�� `- �'^n `�
ig�0���zp`Y��'|�1����ht�]����J�NA�	�'��@�i�9Z�R!���Bs����'�X1�	�_/�U���6ܔ��'i|x��N<:{Ƙ�B����b�"D���#�D=A�����Ӟ~9�e��,D����KҰI��`X�hQ�"n�kR�+D��#��F���H��I#\"�h)�)D��F.�p^`�`t�L�s���ҩ%D�$AD������U�s�<9a� D���%�B<:�
8���8����V�!�/3 $����(�0�u���!�$ךN�����Q*���Į�d_!��T�&�i�H��@�<�|q�"O.�y��ݘ}�΄���@��@�V"O� �a{ -F$~;Z��7,�q8C"Op\3 �/T9V��$ʐ"@�[P"Oʔ�c끌F$���Ϋr�1�u"Oj�H���V>��ڵ"5Ԭ�`B"O,��A�U�M`� �f� �1�"O|@��M�2���4�K�k�`��"OZ4�$�y�)2�D*,�c"O�  ���9�j��ԣ��ڜq�"O�\�d�Z}uPA��ВA�N��r"O �dkC.&a��;B�[�[ߪq"O0|J4 ]�p�!��$j����"OXɃ�G��m�n �᠘;3!hMQ�"O�����x�-��l�Y4"ONp� %(�.	�d�É$�R$"O`�ف�(q�r��
Mp�X��"O����ۗ5%|0"�/	#���	"O�Ŋ���?7��+�P�*�� ��"O�)��)�%+C1Y����Q"O
�iFn��;�p�թ	%L��4 �"O�({�j iD�����ˈ8�f�x�"O(Ț�@inܜ�F	8t� T"O�M���ۖ>��@i�j�
Ah��Q"O�D��ۻvBp䑁�!+Lp�9�"O��Ħ�tq�W�֘]Cm��"Of=xՈ��a�t�aDmRP�=��"Od��E�� ���t��X�ҍ��"OFX��AG��^�K
Ժ\ǌpá"OP����A�i��9�i)s����r"O@:F�^(�@k!Iw���T"O܄Ib���Gำ���#� ���"O�u���]��lA�iک^��=(�"O�A2o�2p���SN�9U�^,Y�"O.e��eP(�]���Wb�e�`"O&9h��ͷz��̈��O-6*��"O�������S��L�S�^�e$p�
�"O�A��89fA�1>�����"OD��J
j�02�N=I;�}j�"O!���L�I^b�P2�Y�f�aE"O�<ZC,A�g�2ayu����r�"O����d��)،M�׈Y:i��Pi�"O^��ņ^�=�B=�&څ�:��U"O�ũ4l�[�͹�f[",y��C"Olq�Ӧ��[Im��f��s�� 5"O�z!��I�lh���!Bn�p��"O�=�*�FhH�cʼ]Z�`7"O�˷jz�3�Eòh���*6"O�`�ė%*�)�ď_�\�	�"O�H��)��`�:%�� 8ߌ<*�"O��7��9/Kx�#7�-d��9Y&"Oxu	`���v%`�U1����r"O�j�&G�dqH�eN�h��"Ox���܃v#"Q���ÿ��h �"Oґ��(�B�����a�Б""O��QÁe���KgN��Z�B�"O@t{g�L�8�qڔ�˻?kz �"OZ,��#�� ��I�Z��h4��"O�)
�� ig}s��^�j����"Oh�3��J�|�*��-{��p"O:	�p!��q�ڨ8���>~s�,��"O�q�%�;"�����_���j�*O��Ŋ�+VZ��.@k0	R�'�H��Z�3�~�  !A�&�)�'�����GH����2�]�% ��8�'�@-�F�Y	���3򨞜$i�u��� ��O@�?�\mZ���t<B�a�"Oȭ�ټ]���BO®>�Xձ7"O�yj�B/u�H�"���)����"O��L*OMԢ���9�Z� �"OE��范;�L�K�(K�E��� W"O�SC�Ue�� h�K� ��"Op����+b��I�G��N��B"O��R��Є'��x��&;����"O
=SP��I@J��`%T=L���"O@x���K�b|�*qiT':�����"O2,��爯��x�Q�r��`""O�m@��� n�yx�R3%Vp[7"O�hC�x ��M�>�� "O��   ��   �  w  �  �  *  P5  �@  �K  W  �b  m  �u  P|  9�  �  c�  ��  �  O�  ��  �  <�  ��  �  {�  ��  6�  ��  ��  (�  x�  ^�  ��  X � � � <' ". �5 �; B �G  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����iX���XVp���#��I�� @L*D�<�ޠ�B�"�ͷ^���1<D�<;Uc��*�"bi_OLa�'y1Oz��#�~����{���"O�@��_4#.]dᎺ)�8��"Ob���/�k2��Y��A��(zR"O\���1?��1E^�n����E"O&�2A�
��1��kI5��A[�"O��p"��kpRur�/�8�����'�!�ĞeH����d� 9���g[�l�!�Ā�iޤ<)�eϫY�f��D�	lq!�Ta�dZFÅ;;�T{�mI)�<F{ʟ&%����a���qa�(��s"Oڌ(3��Q,I��iH56�pp`"Od� 6���#� 	P�9x�C&"O��kE Z1Px8� �B��$A�"Ö��?b� �E	�7|�(��"OV�" ՞����/@�����"O4���U� ���ȁo��	�a�IU�O��̊����v	$<p���G����	�'�$`)&`*G+��K���A� 0��O4Dz���W8}�M9����
�"�Y�)Ϊ/!���T�|�&GҚ#i��ч�̑|!��vr����e�()�����*_�Q�<�'�Q>]��F<`���Qr�A	h"�G<D�X@ǋ@�^����c
M��5"�>�N>	�O'����Q�g  Q��_6��h�	�'���h�IR(b�� �N"��q*OF��e؞h��hܐ!���ӆ(�Ľ�H&�pn�/?z����
�0�m�"_;I`R�	K��d�Tˊ$�N$�-O�Mj1�p� ��J�F#}���P�0�����ɴQG�zQd�~�<�	��)�Ĺ��c^��Z�#}�<T�=�`0ȃ8(�ɗ�UO�<��*[��p�[�&P�N�^iQ�M�<���j��D�G���L0K�<9U�q D�����C����#��S�!�$_6w)�l�'�j9���ɑ�7�!�DB8N�:0� ��+
��h�4�\�&�!�����-���Ѝq|j���Ȧ!�dNT��)¦pc�$�팪b�!�dփ?�5`���$GV��8��Mhf�F{���'��%��cK���\�↙����2�'[����d��5��b'�_��	��O���¾U�r�S�`��ޕ
��R�>!�;n�r�)�g�:��鰂f\�#!�"18�5��8hY�m�D��W.!�DG�OQ�I;v.ӏJ¤bs#�6!���
,5$����V�UI2�㖂��o�!�G ��Y��C�H�i���W�A�!�d�y�]+/��k>��B��~!�$���,+�d�%*�A1��8	i!�$��d&Z��߰qX�t�	��!�d[�lQ
}�S��^�8�Q�jU��!�D'Q�(�:C��>A�%1�(�Y�!�D·���C��q��y�%ک<ڑ����)� F)�ő�<<B�2�-?�uP�"O�L1���;j��P�T)l��бi~C�I�F5&aP��e2̼x��{�@C䉥 L�Z�ʇjT�`����4�:C��;�.գ%�N�zv�ђ�3�(C�	;cDDT�*	�"9��K��57�C�6X����B���ؒ��cUbC�Ij�&�JRh�\�^���h���B�	�#WX�
uOT4(Sf�z��טU%$B�	�3���t	K1o$q
.?��B�	_�A�d�8y�T�6���_�B�I�k�੉a@�Xa:ѻ!��2ND�B�	�~��Q#��}8!�A�a��B�I�	ɖ�Kt�-D��0d�IT��B�	򒴲Q�n�i��I!l�
9��"O t3�CO�,0N�!́	-��PG"O�"1�֝6���R�l9"�|LU"O�pǬ�.��H 7���]^n��W"O4A�פÉA�, �5埶/����"O<���eh��aCY�f�2̑�"O��4�Y*���RN8n�l�""O�1��H)bt�\��a�ԆT��"OƜ��&S�}y���a˄x�\R"O�غD�	�m���3$ΚV�
�P"O��P��k$��"�F�$L�"O.=w	�'?�N��o��n�8Q��"Oj�a�*&��-:�
��0�"O����E�TU�i�R=Oߔ��"O���K*!.LṦ*�YmBy�s"O^��k�.6�FIBrOߪ2l�աc"O`5b�̢O������u�x�[�<���/1��)`k���M��A�W�<�G�wJ3cD�
���9C�G�<��^�6=jW
ߎi�vY�.�@�<Ѵ �)�j��e���ky�<�H�'e�D[�!�
G}��0�t�<���ۅ-�P�bA�������d�<�&/�9Gt`��0��(��yǤ�\�<�2�A���*�@��+/P����Z�<�b'�	Q���P�4v�zy�3m�m�<&���:��Қr�����f�<� @B��4�K��"�F�XQ,HH�<)�	�pX� ����P�<�dO�l�<q��ɡ73����I,$�4���C�d�<�����0�2��t��'+�����b�<���ϡ�������[۴���HZ�<���A�:� � �c,B:y��a�{�<�6*ւm71�iC�8^4�
x�<��%2Q"�1%�ͫ7�he�F��\�<1�d[�j���G�L0v~M�&JHC�<����?(�5�`gE�[��m;�/NY�<�'�A��zuG8y����hW\�<aEB:���q���
|���Qm�<y���;ith�@#�G�����\g�<A�!ץ;A^uC��Q�4�B$i�<��G�8n�H�I���i)�H�HL�<�f�"Y'��15F T(�t8�#�L�<�7LH�Z���S$@]�*6��X$�JF�<I�n�@y"Y�BNv��8��B�<����oc�(�af×f��s��@�<�fcן9�Dpv��2Tƹ��E��<�����a��}�D+k�P"�O@�<��$��m�tɣ@��N\�hr�XW�<q�L��P��P�K��z�ㆃS�<� �xڐ��h�%��IWdV����"Opt�˙�dy��X8��A�q"O��;�CĨy��V(Ӎq�48Y`"Oؘ�lU0K��Ma�S�~88��'"OJ�!���nD&m�G%��Q$�qBW�'�r�' ��'bb�'%��'.��'����(�0�l��\90�d��'�b�'�R�'��'��':B�'�ȂS*	�vN�|S��ǚ
��I �'���'���'���'��'���'ဌ��/0D	x��^�<z���'b��'���'Fr�'xb�'6r�'lRi�D�1I\��E(�2��iu�'K��'�r�'��'"�'�2�'E��B��KNy��`#[۞X���'@B�'���'X2�'h2�'���'+�H��	�!��9�g ?=��ep�'��'f��'>b�'���'���'ǰA�aCB%4<�(x�+bJ �Ѵ�'R�'��'u��'B�'��'AVI�C���6B��H��[��24�'���'u��'$��'���'���'� 0����)k�Ua���:���*��'#b�'B��'
b�'}��'�r�'-��Y�H���:S �_���C�'���'>��'B�'�2�'���������89�I�k�p����ǟ���ԟ��Iߟl�	ٟ`��ȟ���ş��C	˾s[*պ��PN�P}�vm۟�	���柬�I��,����M����?1"�����е�ѭLT$p1�.c�4�����E禡�6���}kfYR���	)�Tt�El4V'\�{Y���4���O��"��،G���(QD���sJ�O����THH7�;?��O4H��$����:�&e��S�Ϩ���$˘'��_�F���L�ZL@�t���`�JO,7��?@�1O��?������H7
�ر�[�Z[��Jr ���?���y�U�b>�qW�Ѧ1�w���$ȗ�D��Iv�V�9�͓�yR�Onu҉�4����גefT�u�W���r��>
�d�<9L>	Ӽi�x��y�A_���	�f�=2u��H0�OB4�'P��'(��>T�ƎJ���Q�lu�Ju��A~2�'&2�(��?�O&0��I?j�2Jܸl��p��E��Cj��	py�󧈟�� $k�h����a��p;aF�%����r�0?1��i%�O�	�=L�����0b~���f��4/��D�O����O�y��.j�<�����21�FfQ�Zǌ cD�I�U�V`�"�������4�"��O�D�O��D R�A�A�e]��G� rֆ�#)�6���JXb�'ib���'��]B�n����"Jǟ;�~�6¼>)��?)M>�|��lL�Vr���c��kX<i���L�fM��4w��	\��4�w�Of�O˓y::7��Ӣ-Q7lO9R��=S���?���?���|�/On-nړY���	%�ƙ�A�jg|��Њ��e�R����M����>y��?���^L��1�gì8ܒi�CS��]��k��M�O<x`u!U�������w$4L"��= ����� �2t��'��'}��'"�''�b	{����zOYk��=��� 1M�OV�D�OH�m�h)��Sʟ\�޴��_����weM�UM�����GP>ѺM>���?�'nڙ�ݴ���W"2�n	��ݒ4U~ �1��rd�UJ�I��?S�'��<�'�?	���?�2�
�0l��8�b�v��<9V�T��?!���Q˦ek���џ$�	���OP4;u`I.�:��T�������O>X�'�r�'ɧ�)@	@��ՁkF�)z��5ĝk� ��ݴbj��5?ͧ`���d
*��H�FM�A�C��8:�&�4}7tT"���?q���?��S�'��d�e��4~�ɉ���Ze�E�E�=1��ܟ�{�4��'#ꓨ?I�҃IKP��6m#2�P��V䄳�?��p�T�ش����<�I��'��S�/GT��"Ǖ=|��;�
Ga���Xyb�'?��'t2�'��P>����O�C���5��}�Y@�;�M�&V?�?����?	M~���cC��w �Ge��NA��:�=��e#E�'42�|������-��f7O�wC��f�d$�㈱Bh,��7O��4M��?y��;�Ĥ<���?Y��i%��y�M�
(R��)e(�u������IޟD�'��6�Џl*����O �dY�'Z|�(ŎJ�H#�X���M�.����2�O����O�O�(�p�̵S�*��3!��a~��+M�\WbB� ͢��
QO���R
ݟ\�g+�RG^��!��$wp���vo�ӟ��IΟ@�	ΟPD�d�'�:@!ҽP皱�w�Y�h��]ٕ�']�7�V5P���
���4��h
���-�Ū�m�&Z��,aG;O��D�O2��˖L�*6%?�����3J���/@�@���1m�	Q��T 	VM$��'��'c��'��'��Ǣ*a�����N@�	��_��:�4�:p���?����O�x1Yw'�&4�~��5�M K��>����?AH>�|�bI�$Q��PPƖ3nkր�b�]";��u��~~��Dd�����}�'b�,{�B&��2
L2�a�6`x\���@���P�i>	�'��7�բ=`��0@X�8Bv�β�(QQe�58��T���?��X�8��Ɵ��c|��qϊ$e����C�kn��݅d�����L���ڒf������� �����%��m�� ��!�h;Or���O@�D�OL���OB�?a�Ģ�#8֦=� @ak�@����֟,��ПHP�4zL��'�?��i�'��C��e>�h�w�A'��J"�|r�'z�O�F�&�i&��>r �x�����}�@��* ������Wbo�w�Oy�O�r�'��Z�%XLH��N�k��ȧ�%>\�(;kO�	��Mc�����B���?�,��u��1e������1?ڀ踄<O���_}}�'	�O�	�O�e�p��M�D(�Y�:�^,�E	\&�Z��1LB@X ˓�"�N�O
aIN>i�!֖`�.�肆ŉ*@���ڞ�?����?��?�|�(O�Mm�2	l�3"��@9�	(Eڰ	��������"�M���>a��M;*�j��- �A�C�]�>�`����?��k��M��O�$�E�:�O�౪�H�yP��hOh��'��I����I�����۟��	\���i�k"i%L�LC �� /�@6-�XL �$�O���7�	�OB9mz�)0�W�BJ�}"�Dʱl�4���+��D��f�)擞j<�m��<'
4H���0Z��d�lip��I�Jܠ��O��N>�*O�I�O��b	F�%����E߂ �����O �d�O����<Q��i��'[B�'{.AJ�A;�r���v\��4��Q}��'9R�|B-�,�����Y�$A�g㌯��d �r%*����Z1�
��_���*2���mJ�r*X�;B��}���d�O����O���>��[���M�|�0�Ɔ�3٪PZ�ş!�?���i�91�'	��hӢ�杢	��<Q#�a#�(換#���˟��I˟����ꦱ�u�㏞$�D�3xw����I�	q��Z�k�!��&���'���'r�'��'����AN����v�D�1q��\�P�ٴE�l��+O��D:�)�Ot<�CN�7Z[�x�`��[��]QdA}��'5��|����J�Aj(t/����Ã�V6��M@"H(\�X��@/�1 ��M�p�Iqyr.��V?�����Cb�Az�A�����'���'[�O�I)�M��J�
�?1Ƨ��7� �U$�'�ņ� ,��I-�M[�B&�>����?y��h�����˝ao����E9�1#��ћ�M+�O�H�̛��(�����Wh��ec�?%a���d��!��7m�O����OZ���OT�?���dĦC2ȳ�/��o[��CAU��d������ܴ?00�B/OF�my�	km���żhHh�!��<.��$������>�\o�Y~R�Z�z)n��U̓+b;~ k��+�����i?�K>�)O��$�O����O�liA.2�0$�e	�R7,���O���<Ⴒil�� �'!B�'哞䀣rƃ<N�Tt@MƧ8����ϟh�	z�)�sLˤC�!�4�ұKm�d�bD?��L�R�ݔ[�<U������P�`�|҅]HdH���رS�t�"
�3fR�'���'����_�\ ݴ{���Ȥ��+��D� ��,�ޙٵ���?I��d;���L}��'z	2����v\0����y���Y�УdLڦ��'�pigE��?��S�;W��~��ѭ���*�8"i}�T�'�r�'�R�'M��'�SvRR��c�ؔ�
ښ��o�yy�����h�	�$?M�Ƀ�M�;|� $ISE 	<�U A�]�	�,����?�H>�|Zs�[2�M��'�>I���0 ��
 U�S�
�'�,i�
Q�l;՞|�Z������z��B�Yr�@����XH~�٠�埬������Pyjӄ|
���O��D�O�!�� I!.dy����[�%�'$9�	���O��$>�$��`��=:VOI��*	�>[��	�vc��w`�|�Lb>E�'�'�L��i-Y�S�ע(���b��יK>��5�'�2�'#��'k�>睨Iln�itiɳl�5	ҍQ�>P��	��M�@톺�?�0���|���y��Cv�3t�W�fV�i�c ��y��'B�'� x ��iU�i��#a��?�:Tm�+`a�y��Q:`���0�E�+��'��I矀�	ş���ݟp�I2H�X�`,�E? ���M�+5�섗'�7�!h�T��?)J~R�_������<[ʶ���O�-!֘y�C_����͟ %�b>mb�%מ>H�a �MޕQ|@*0�1l��l���DP�)��e��'�'�削H�}C���R���*P�@�f�������؟�i>u�')x7m�D2\�$�p�j-R���k�5*��72��D�&���	����O@�4�X�B�M?��<+\4)P,0�\��Êe�
�98tå�� \�I~j�;r�4� �.*T�)�v�)̊$͓��?� �q�j��%Hb�\T3�@��D�O�o��"X�'Q��|Bg��u�ܜ!�i	�v�H3V�F v�'�R�����y������$d0wCHTZ&��F��NV3R/�]{w�O�O���?����?��#~|UfD�TK�h��ަx��$q��?1,Ov�o�.����	�����~�Ԅ��P�u0�Ϭɴ4*�����$�\}�'�|ʟp�Sr#�E��i�s�E�Ru<�P�$�827N@6�}�*��|Ji���$���#P"Dxbh���ş{��`s�ń��`���|�I�b>1�'��7�J F��Ҧ^��ċ<!�e�q��<�s�iU�OF��'��%�4~�L���(0vJ��O^!9"�'Wr)ײi���4n }BCܟp�S�? ��H2�@6f6���K�2,[�6Oʓ�?Q���?����?�����F���	aF��x�R��� J��m�OL"���ܟ$�Im�ܟP+����`ѣx�H�e)ު��q鎹�?�����S�'s�TL��4�y��CD>��:�H7ɶ�y4i��y��N�s"���	�G��'$�i>Y�I#J�,�c� �S�t�,�-���I���ϟ��'�H6D��z���O��āT�(��A�u�Zi����i��T�O����OR�Oޜ��ELs=�La�iӮUTl�r��ؙ�o��{dx�� �6��{a���۟<ӂ�/U��Շ[�~�T�da���0����h�I��G���'(��S�f�|1���7Fs��AG�' 6-̹0���D�O�o�I�Ӽ�dTVn�)��N�<�x@�h��<a���?���r��Sݴ��d�7>P:�O����2�L><N�<3gwm�#TY|�IIy�'���' �'��b��M+~�ao�#m���N �di�	��M FƇ�?q��?�O~b��{aL�8���5�\Y�Ҡ� 5��2�V���Iş�%�b>�ꆮ�3+��u�%t�Qk��I(�j�oZA~R�ʹ'�n������D��=�8�(�C�A��bX
73����Ov�D�O��4��lX�FE� ��"��X�!�ҼI�p ��D:[-2�dӂ�Hb�O���<�U@�&�4�kO$R˸�tHT�W��}��4��$�!J�|���O2Ғ�l���˰��0IZ�A-��ه�T�w��$�O����O���O��D1�S�T8����Y�0�rE�@�3OV���ʟD�	��M�H��|B�&j���|�f�*(�Reb# I�^ �%(��G*|g�'�������6�������	J�5�(�y��Y~�=����6PS��'���%�����'���'up�&m�UwXM�,ԗk˰�H#�'�R���4_[�l{.O��$�|���K	?��x���<��=Wb�S~)�>��?�K>�O9J���::����a��QS��D0^�0���i��i>]ˤ�O��O��2��Z&Aڠ��k�#hXҨP��O����OR��O1�
˓Oꛆ�O������Əi�a��B�_�6��',q�0�4;�O���"V���#�
8���b�����d�O:dZC�i���=p�H��f.��a���N�}ʂ�ߧ#K���ny��'�b�'�r�'��Z>}{�O�I��Bv�\�A���H��M��C�?����?�N~���x���w@j�H� �\?"x�c��l���y�'Or�|��D�B�o���?O8p���`�)E���r�;O>|p'/ۢ�~R�|�]��ן��D��FDA�Q.$"����S�	ޟH�IJy��x���H��<)�"_�u����(R�.��3������9J>���y���ş���_�	+*�ʵ��X7Bx�G
Qa�n���a	��M�F��t�_?i�� �,b��LO�*̠�DǸ^�p����?!��?9���h���d��b�6١�C�ȉ%N�:� ���Ϧ���@��������M���w���I�C�4u���0���	!�����'~R�'�r�$	������j�@-:3�);�����
�D�*���D�T�@�O,��|���?Q��?��腁�w���F�._��Ss�H;��æ��c,_ZyB�'��O����'s�z`3"��&���+8F���?�����Ş,��l�6F@:q��d�.ux�8慘!�MK�O�ԑP#ٗ�~Ҙ|�\�t��E )5��-H�/�dث5NB�l�	��	��iy��b���z7�O�$�DC��;�DQ��M	U#�@��O�nZC���I˟,�i�E��8���&��i�̥KŎ�Y.4aoI~�.+.E���'��'���E��%�a���?3&��  �<Y��?Q��?Q���?�����e!�����y?@��c卲Vr�'��}���0�:�J�D�ܦ�%�|��$G-9	t]� �]35g�T �>�I˟Ԕ'���;��i=��78x뎂+%�� �f��q��*େ1z�,��	P$�'��Iɟx��某�ɵH�(�d�>H2�Qhw��u��I�	͟��'0D7MX��b���O0��|��C��h�1D�C-pT���Yx~r�>����?�I>�Oc
ua�UG�1r�B=w�a�&�P'6�P��i����|
a覟�$��vkD"Axb��D�ł�U�ʟ �I����	��b>��'M67M�1/���a
�5<B���J:M�T�R2L�O��d�ɦa�?Q�R���	�1�h��'KB���Q�LzR�����@�Gæu�'Ӭ�s7�EܧAB����f�z��A���dΓ��D�Oj���OB�d�O��į|�Ul	�(�~�Y�LM�l�,: R"x��/�,2���'"����'�V6=��|+�aT+5Y��H"�8Im��`(�O��(���>e�7mj�����
Nc�}sԬ���Q��n�T�4"߳G���!�d�<y��?a"d��m6fT�w��� "��CÍ �?���?a���ߦ��c
ʟ���۟X��I�Q�	to�V�1�T͘G����	���z�	/;�J}�3aK�'z�\�5,P�F*�O@��En��R�@X�O~e��OTX��︵ DЛ9�|��A腗!2dX:��?���?A��h��NY����@�T�-�ƁQ%��s-��dT��*we�������M��w�V�@u��FD`5aW4X��1�'���'��O� �����@���!k�� .ZrK�R2��
D�~��+���<����?y��?A��?A�a��D	r�ۣ
�LY�d���\䦅�@�[yB�'��O?b�C� '�Q[eV�o��Աe�w�*��?���T��6+"5��E ��d�h9�4ua�&"8�剢y�tH�'��('�\�'�0�#C�^>�U95�/M��f�'3��'�����dP�r�43(�]��pw`Ѐ��e��(�gO�Z�H�
�5����d�o}R�'u�|FJi1g�4���A)�7:�̲Q(H����'��@@��?�������w,`Ÿ��
�a37wݬ���{�h�	ʟ��	��I����*��đYD�jj�pR�4�A��>�?���?I��i���ӟO��iu�T�Ox�Z����+�5 �\�4���+��&��O��4���gsӒ��J���U?s�Fi�Ã-"����d���Z��]�IKy�O`��'	rl�L�r�z�N�	WE�1' X�[��'��	��MKԪ��?����?9(����%i���´t��%x��a�B���2�O��D�OV�O��c�@�J�3zD)B��;X *�8v��H��(�'.?ͧp�r����[>6�Ajj�lm�ą-ED`�����?����?a�Ş��ݦI��#U&2#]//0L�4EG�0
8�AU�'�nbӾ�O��DF}��'9�ิ�!6G�ik�̑-ڠ��'9j�E�����֝76S�u�S�e�
IeT����6A"
��
*M�t�]yr�'��'i�'�"_>-X��"ղ� W&A,-��!;5EV��MC�%6���O�?e`���37�D�j	C���=����(�?����S�'SW!��4�y+QU�XQ��,o�z�xUł��y2��^>~�������O^����D��/��4z0�!V*��hv��O���O\�Y�v(�=�������v����O�'3�rS�KO��=e�	ߟ���f��mTЁu��7^��Y8g@�&�6�n�4�i�%�|2��O�%��I'����1\X�p#��u�����?���?Q��h��N\��� ����oE��7%�8({��$�y�U�H��`�	�M+H>��Ӽ�C��2���#�>}j$���<!���?��	�(\0�4�����$Y# �Ni�&�8tH'fY�}`��Ή�������O����O����O���ɸ0XR8�%9G%�0Ӱ�D�p�ʓu��fFE-"�'$r��$�'N|�ʁ��c���٠�\��4���>1��?�N>�|��C(�Ձca�'u�b�Sj 4��b���)���,x�T���g��O�ʓY�.��D�$V	(�#qB�H�8 ��?Q���?���|
,O��m�+V���Vz�@pa�j�ؕb�O��&�-�I��M����>)��?���Č(r���[�����'Â��N��M��O����7�z����w8�R+
=�2Ak�v�u��'�b�'���'��'B��`��ԶDG��g-J"�P�P��OL���O��o��xN��'T囖�|BBN�}�>U+�!%6\���p�
&�'�r����;zQ�曟�݃}C`�R�?(�qH�]S���PEFП���|rU���I̟���ݟ�g
�YW�q�$؏TM���ˉџT�IFy2�j�lı#��O0�d�OZ�'~��B`�U�c��J���0b�i�'��ꓐ?����S�$&@&G��#��
�7<���gN c�rW2����O��G��?��k#�$Q�$Z��q�ۿN���H$œ$�$�O��D�O���I�<V�i������
&w�x��C�\�Z,y���_m��'��7�+�	���d�O�Ps2`�*5�g�z!V!Xu�O����Md�7m>?A'�Ȅ@����xyB�Ϸt����D�3��4�`(J��yRW���I䟄��؟P�	��O�<�*�GJ�lDP���&/��a���j��(ɇ-�<A���Ou�7=�N� e�B�{���#�*A�}@f��O��d?��iȧK7�~�D۷�)a����ŵ#����GN`�\�B��=���/�$�<���?�@�Ư0�K�mЃ,�.�0ti�?�?��?����Dަ9�!�П���ΟS$ ^ 8'�M���j�b�å�p���Iȟ���]������q�N�c��=Q��2��p��=R�$�|��O0Z��,k`�u/�l�8E)�?ޘ���?����?���h���$�-�ݒ Ӹ\�f�	��^�)>��D���!Y��S̟��	&�M;��w.^��&��v+&��J�
��E�'���'�2a�E�F���ҩ�2u����Z7/�0\H��]�_w�Ab�͇h�pp'����D�'�b�'H��'���i�f-��A�&�ǥ.�ZAQ�[����4A'6q���?����?	����c*�/1�i��ɐZ��A��O~�D�O��O1�h�`F��p�\зf�5R=�2�`��=��6m�My�ΐ���������&;TlP̒�4  `��˧a|�iӌ�`@�O\�(gb<�$�*Fm�+���Z 0O��oE�����ܟ|�	�( �M�|���(�G�%]<�9#��7B�J�l�g~"������'�����4�K�D	�-�J��<	��?��?A��?و�̛�Jb0��MA�	���h��-V��'�".v�p�:�:�"�DA���'���ՁȞnIB��k�F#�t2LU^����t�i>]���R̦��'l5!
� Ru+��[H�(��P#�( E�X��7�?�D�2���<�|�i��5`��|$�Ȩ0�!&��MFxb |Ӕ��� �<���� �� (�#��+.�Ԩ@ǈ��I����O��D ��?5#����3�X��X-S�$I��3b����Ə ֦U�/O�	W6�~B�|BD�:6����@N�p�й�x�@o�n�*����h��8��B�76��7�E�D��d>���$CM}��'��	�#�u�H芁�.��X��'@��֗/��&���iݾ��ɬ<i���ls�q�I?N͊dHG��<�.O:���O����O��D�O��';Jr�Pg}������_�(��!�i�tp��'W2�'p�OU��}���RM�����'LYi3/ؔ%����Ol�O1�~�P�r���		poP��v�>}m<���m��I �	(lc0�ۗ�'�f]$�ԗ���'ށӗkľB&x�7O�P�,H���'���'�[��[�4m��/O��$��|�����6%pX��(�s��㟀y�O���Ot�O��A%Nێ �p��N�)g-�)斟��Ý$<t��l/��By���ܟD!�Ꙍ\nyX�o��a���ʵ�ݟ,��Ο\�I⟠E�$�'h�c�b��R���\�#Z7�'mv7��U�:�$�Or�mY�Ӽ��aG:6p1a�O�O1�D��<���?��K[x�{ڴ�����M��П6hՆ� �|i!T���a��� I#��<ͧ�?���?���?a�J�%E�`��T� �0��D��&��D���� ��(�	П�%?!���\xД�X�T�M�4$еNI*-R�O��d�O��O1���ۄ�2�%+��!�p�Kf�VjXt7m'?��^d��Iq�	nyBᕣ'�Pف�Q
��2� �5r�'/��'?�O��I��M�&�L�?����<6|]r���":�vE�w��?q׳im�O~��'�rQ�,�.�t���;��sڰyU��� s�Tm�j~�ԄA>��ӷ<��OH��	mv�qQO:6	t$֏��y��'�2�'�r�'M��i0���-�$�q�� 	�bВ��O��$�O� mZ�kF|�Sޟ�4��Vh����w�hГo[iE��H>���?�')nl��4��d��ƽ��ˈ5�\��Ν>c��������~�|�^�b>�I9�b=���R�o�m��	J!�"<y�i�.I���'4b�'��'��A̐$1Pe�W�Ճ;1^�!���x�Ij�)�g��a�\eYWE9.<��y ~NY�ЇD�MU�ؠ(O�����?�b�+��ݑ^�lqPB'ٛZ�V}�U,�����?����?I�Ş���æ�q1!����p�P�̳"�Q{WH%@$��ןT��4��'�����n�,�-���8gm�ԛ�O�	$����П�ZSO�ꦁ�'BlX���[�'A��h�4)����ŏjT��ϓ����O��D�Of���O����|�ጌ'E|b���H��L)��V;?��F�Ao2�'����'th7=�F��7	�	@��u:Ja�m�O0�%��Z/uO�7M`�4���H�r�Bs�-�2$Z�"y�H�d-G�4�+b��my�O\rNU�P/���A�7w���ʟK���'@r�'��	��MV�ջ��d�O�q`膡|o^�0g�<y�x1�2)8�I�����O���'�$�0K��R�ةB��"�a�����S����ɰ%�b>�۵�'�����t���kX�_�R�@$ĉ�����ݟX�IΟ���n�O��O��1Hh�0�˖Ѕ^��sC�'�7K-���d�OR$n�@�Ӽӣ��,M]��  �h�X�@��<���?���A��l�ش���Z+~,��B���.��F$�@	E�$u0�"���<�'�?����?i���?	U�
�y�eeq�Z�G� ��ĞǦ���yy�'��O�2Oſ	6֐x0�\ & (h�r/ۼ"Bꓙ?���d�
�&z��2�㝰]���3�e�#xA��-Zv�I�}�D�a�'�h�$�H�'��ũ$�I79�bq��h3R!rW�'x��'�r���T��ڴ]�8���);�$R�w��(�7Cͮ�����v�$x}b�'w��'/�!j&CA�}���S���N�������[Q��������j�Q>��]�x��T1�e����u�M�t��	՟X��ɟ���џ��Ii��Ruf� ���'M�u���An�3��?�hi�&o���ɓѦa'�l9pG�)l&@{���0H<��`�T�ʟ<�i>M�#	���'Z���s��D&O7I�5H�
�.,�I�Ae�'��)�s��ٶ'��'�vA�����3�0$YD�>ÛFg� ���<�OV�fA$K"�;e�_�;#pYz�O��'cb�'ɧ�Iޢ1���S��#0A��S��+��-a+ϡ9 �6m�Cy�Ol����c���`�M��V �HO.̾ą��FW�V��gᔅ�@���8I�MSa�ӯ.=�yF^�PR�4��'E�듮?�d�U�'8���2ft�2����T��?i��/lxh)ܴ���	�]k��y�Oq剁?�.=25ŷO�] ��y
�Ibyb�'u��'�2�'�P>uJ�ɕ�T�H<y����W�$$��ܵ�M3�Z��?1���?�L~:��w��y3+��0��9zP�E$z�|����'���|���ۆF[�60O� ��[�]K�~�ؓ/z���:O�u0�j����9�Ϟ6`��ץМUǀa�ɚ�M��9�̅+kq�ف4�T9�
H3䍇�s'�����F�b�1s-�/u����4%V�QXy��Hމ�� ��h'Uk��D��d�`i� I�~�@��ڶL���cR�@�#��i�`����^T�dȲ�ݚ3Faz�s����gL�L�f%K3)�"�����n�.j.-+��U�>��L@�lG2 � aaݯx߶Ŋ�.��^T�Bh��M�6�^�VB��%+V�7(Q�� ��?�����G-U����%)b{.�R0Ed`�$��M�
X&�n��ɑdV��K��G��v��T`X �ze�ٴ�?qL>���?�`�L6߸'���H�$�ea�U�d��9 {�M�ߴ�?I���d؏f¾��O�b�'#�t!M�2�$�&oݜJ�
�+��"O"�$�O�<@�!?��E*��L�z\�P�4+E�=���2�&�⦕�'y�1�t*w�L�$�O��$���֧5f'�l��l3e���ꡓ2$Š�M���?��'��?�N>I��d��#�V���Y.�zQ���ީ�M��픪-t�v�'b�'?�4�>�(O|q�T�UE��1*��:�I!$���xJt���OqB(I$���A��.� t�`)�
N�7-�O4�D�O���2�p}�Q���Ii?)�&\=T 
@�ߨNS�`[�JYS�8�D!sN>a��?q�p�^�{��Z����qB�'f�t=���iN�%_�H����O��Ok�W	Y}h-GA�"J(�9��ʌ3F ��$9�]&��	ޟ��gy"��8T@nѻ�n�__~�yt�T�{PJ���>�*O�d5���O
��*9R���&��Bu��wm�iA%��O����O`�a0���5�&!1o�K�~Q�3�Ц�y�A�i!����$�X�����r�D�>i0�� �� 	�H G�
HS���M}�'$b�'��	�D���������8<"Iz�X{�a�I֩bcP<lğ�'���IğH�e*F\�H��a�GО(�JMaꝧV��o���P�	iy�F�$��'�?q������x�q���X�.)Lq#�荝Mى'\R�'~ڙP"��?=����y�RB��tR��,x�`ʓ:�J����i�B�'R�OyR���,��QH����F	pn����.X女�	ӟ�`Ɍx����O�=�����
T�dEn�)ݴ�9�ųi���'a��O~����O7Q�Tf��V�pM�ׇH�S�"un�5&V0�?a��4�'� iCˏ��hQCR-�
����Jr�\�$�O��d�H=�D&�����7�D# ��z��X����!�nZݟ`&�����d�Op���O�D��#\�WWh��G�֫n�sa�Fܦ��	��
taM<�'�?�J>��I %B�Kx����TJŀq� �%�X�I@y�'v��' �	�[&I�$��> ֔x�ʇ5�2�;wG�>�ē�?���������Xf�VC��ۦ&Ѕ��i�rX�<����4��ay�O�!0غ瓀x�Z�2��B��@|�6F�5x���?������4����]�[����FOS�J� �dJ?<s\h�'{��'~�R�(;�,Z��ħ,+Q5�ͱW�X�Ӆ��TmH�i�|�\��埴��dX��&�#&��c� �J}��3 �i"V�P��4�ؔO6b�'F�\cEx�id$�4M0�Q�U�Jbμ�L<����$��\~�֝^�Qsp��chH	����?vH��?����=�?1��?i��*O�.��~̢*�;�@� g-�kc�v�'U�Ɇ��#<%>�Ha �9��KW+�2yЙK��j�<<c���O6���Ol�����S�t ЁOkܗ�d�6	����ќ�+wY��pA�'�S�OY����N��I��8k��Z�0�U2�/pӼ���O^�$ݳI��S���>Q+U�>�F��#NܳK�E"�ҡN������'Y��S�c+^���gm:���.}K�V�'�Ȑ�\��[����[qj�� вmŅL������tft�<�����O��Q3��
�L(!`��Q4Dԉe�F>6r,˓�?����'1r�O�@����,X��� Tw9Z��°i�L-k�y��'���ǟػ�jV�p��59�:`jtg�4�U1�c�����IƟ(�?�����ux�v�ħ2# h#�Ψ��=�ҏ] �ē�?�+O<�D��stD˧�?QT&��~�J�8���Ot�r�̺X�����Oz�m���&����E �n���%�j��Je���d�O�˓��Ē���'��\c��\�oR&�Lc�O�<ŀ�Ob�D�<����?�H~�Ӻۃ(����t	�`8c��YRG����a�'��*��r�N��OL�O�,�vr����LO����q��n�ޟ|��ܟ��I>���<�.���b��w�|Uy�b<YVQ	����M���/�?���?����(O�ӛw����A9G�F* ̞�1fx��O4ġ��)����5oE�)�̉HcaW�-Z@y�Á��M{���?y���<0'�x�OnR�O԰x�C�vO �ю��k��!�Ĳi�|���~��?A���?q�"K��"�� IF�Xu�2�@;���'�~��@?�4���<��������+%�8��n�<��B�x��'��������<�'J�5BУT�Ó���*��a��޸�,O&�d�O��O$�Ӻn�5qy�����+}˔ݻ��Ҧ��	Zy�'���'i�6#1z�H�O��x���v*���׼o��d�޴���O���?����?!T��<�v� �Ce딛}���j�/K1�����i�"�'D2�'���($i�)Z��z���v�[2$�<>[:0ҁ�ғ$�L}ـ�i*�V� ��Ɵ��	� �$�ҟ`��4�z�k�˜$e��ڃ�[Vi �o���	y��~U��'�?����j���v�	�֣��h����R@�=��	��@�	ԟ�ke�i�D��y�ן���s��	W(a��h�${��y��ir�<]J&��4�?����?Q�'`��i݁s�)V�ka0���D�T��a�t�c�:��O�*A��p�'Oq��dR���./:J�e'_�(��e�r�i+���5)g�
�$�O��d�����'Q�,miX��Q� �T���q𧟽[�0�4j4�̓�?�/O��?E���$<����(�\m `�A�V��<S�4�?���?��Ք��	fy��'$�DC�\ �
�d�7.��G뒛;d���'��	�Y&��)*���?��\ �H+��;�T�p�#K�p��`B#�i��vx�����O�ʓ�?�13w6A���L��`�%K�3�P�'l��ћ'Z��(�Işl�'ʑhi��Z!R	�c)�0^�`	�-SFi����$�O�ʓ�?���?a���2��܀��cψA�@J��z�Γ�?)���?)���?�+O�EZ�F�|���Ykh�p����z���5��ݦ�'d�^���П���+/��G�� �1��<'E�an��mZ�H��џ��IRy��k��'�?!��iV�8jբ�f���V���<Z�6�'�������������l�\��M�A�V��l�r���v�dxE-�馩��ٟP�'�.L(�~����?��'L�z���Y�rո�oJ]�ੳ�S����՟��I}@��ʟP����T�'@�Д ѪQ	Z�䅓d䏮+��lZZy2�ڦ#�r7��O����OV���n}Zw��=x���[e`uP&�S&P�J���4�?I��g⾵Γ�?a(O<�>����!VL��S�'� ��W%}�b(�`ʦe���P�I�?MX�Of�T�	� ř*u-\0���X������i�@U��'V��'��	�Od@ap�]�bLqj��(/9��r�o�i�I럴��%��e�r}bZ���	r?��\��n}�fI�,8rŹ7����ퟄ�ɑr���)����?��s����VA�Ě�
�@�j�X��i��-�R9���d�OTʓ�?�1h ��Y&���m��h�$�K�<�4m���%�x�X�'���'CrU�V�H�KH��XT怾g��|z���)"�����O���?�+O����O���E�U�A�痄����g���_fĜ�7Ov��O��D�O��D�<�2��E$�P�Jy`��&�^����O��O���Y�p��sy��'���'.n�I�'��X:��I �*$֮ϒ �1@�,w��D�O��d�O�˓= �+�W?�i���@L܄�0%n�WV�U�,s����<����?	�9hx���i��h!˙2�˰Id݊)��4�?����d�C@d��O���'���	*��JQDE�6-@��D(��[�~��?a���?����J~�R�\�'����C+w ����qu(Im�`y��=UP6�O�d�O��	�A}Zw6�(c�k�(q{��"�bƙ	U���ܴ�?��rTp�͓�?I.O^�>9�&NM� D�}���А!�Z��q���`����	ȟ���?�9O<A�sjb�@�&߽ب
���ư��c�i��p[�'c�'	����OL&p�솉PrP8��F�u5�nɟ��	�<����ē�?Y���~���Y�p|�2%Y�-~����,�M�I>aU�I�<�O���'��C�>"+���v@,#��O��0�4�yB�@�ǉ'#"�'"ɧ5V��r6d̑���bO@%�GN\.��dţ^'�d�<����?I����~8&YF��N#,����9~\���cMU�I�x��^�	�|�I}�t��%�
��ŋw��f��|3�?�I�H������'����s�p>�0��z�ѱc�I�M�8��5�>����?�.O�$�O��D#A�$���HAZ� P�%:��H���+�x�'���'V��ädG��'֥���=�6)3!�7�"�P�l��M����䓧?��]8�����I�2n@�W�޹:t��&�ø!�N7��O�d�<��{4�O�B�OnL��NĴ{�,��,��d.`bf�7��O^���%����<��?�f'�:kC���*FHm޹�� q��ʓ� D�ži"�'�?i��"��	f��4�r�2�DxG��0�"7M�O,�߂?����=��3� #jna���g`�f�����En�z9/�V9oZ͟$�	֟�Ӕ�ē�?!Q#<-������8��AĂ�g�&g��yr�|����O�hCp�@�2�֗��xt���	���'��N<����?��'��H�3R���ggL��ݴ��@Gz�+����'���'��{�.��G=L5�c�[#([pxI5%i����XJr<|�>!�����Ks���u�RmARjϪ*

1��oe}���rz�'*"�'6BX�ԡ0'��O�AB��ĿK�vX�gO= ��L<����?9I>���?�W�(W�1���K�~QZ���kf������O����O6ʓi���Q6�������	�tK֌�O��Şx��'��'��'^1C�'�x�P'(��u�\��2阕��%#��>Q��?����aU�'>�$�$;�hSq�
]��9w���M����䓯?��bFf ����	QwP��a���q���#��M�	ڟ��'�,�i5�I�O����U�����)A�����J]_���&������Ԙ�f���'�4�g�? ^,��֟f*R�zt$��`
Bɺ�iu剪��H�4 �����S;���I�0���Ӵ�A|0�j` \���fy�'��O�O\f�A1+�E{�ͻ �֏ol�0ߴ$~��K��i���':��O�O�	�9�j�3�IW<���۸,����'U��i�O� "�5.P�h@w�VV�J�L�֦���ڟ��	i�I�J<ͧ��'34�T�06��؛��X�Ն6�/�����'�?����~�5)�����ǔ�|��uI޷�M���n���*O���O��|rMʿi����1�{�1�o��0;@K�x�m ����O"���O��B
���(qa�x�0!�"0|C��@:]��O��D5���O��Is�x� 2��7'*Ti��b���	� ��L�ĆÇ_�)������Z՞��$D�b��?�����?���V��h�'Y����⍴H��0�҇D�n��Ѩ�O����OP���<�f-�2\�Ob��	'�J?-��y��͇�������q���:���O�D��}�O^��FcR��vP)�c��
��%Xr�i�B�'�Ic	`ܸ�����O"��D{���&��L0LDRMS8d`�|�'�r�'�2�F���Ĥ<��O�4�B�� ���q7aV�x�*���4���6���oZ���I��`�������"��O 1��x��Q=�V�S��i�2�'�$�3�'L��<a��e�1l�J�O�2	4���u�ߘ�M�3�ƍ8����'l"�'	��(�>9+OЈ1�mLQ>蔘4�
N�H���h�Ԧ=J�b�@�IIy�)�O�4	�I۝7F�8p�:��lN�)�	�����Hŀ-2�OF˓�?��'p��zb�
�~S$����(y�ёߴ�?)O����>O��՟��II�s�G"2j����ȴ�ץ�����I�f��8�O*��?�(O(��Ƽ�5č�p�0:�L@K��,T�	�G=���ȟ���(��]��';��`�4n�qYGϔ2>����q,D-Z� �����O�˓�?Y���?�fA
�(�*���=v�rmA?������O~��(��G�X,�ϧ8�6�����"[��9�tM���4oDy�'Y�Iğ|�	� �-m�HpC�0q"�q�R�� <Ș�ȕ&�����E68�Ģ���nU.����Q��H�t)�#d�h�Zh¥r��!0T*O<iaf┨\t�#�тU�TP�'�F�z��P�:��� >��x�1�֫"6�I�B�u,h���돺��m�0kS]�nɀU�K�\N=x!n۳ ��n�b�@+�ޞ-�n�j�l\a��i�ֈF�h�]��k�%@1���)�f@ʵ-ׁaS~p�T"z�P���F�8e��ő�	SYxH���W̢�K�������lZ��O�/d���i��y�l��\4m� ��Xе�$q_�#dG�����wϘ��&�� 8�z��ፇ�u��h��C3T{t��Z�0س��#87���H�G�P�f����܇��E�$i� �h��'nR�����O�aB�<J�l!�d�
#�X;"O�ik�+[�+S��C'÷r���I��HO��|��S��)���3�� �������T�!J�8M�	Ο<�I��3^wB��'#v����s��}H&l�X�&�q҄�O�ݚD/W�t�jX�wKN������ҡZU�q��.W�<-�s�
=����	f�bQf-^+/?bTR�ޟўtqr$D�*��M-4��
���A�����S�����O*�=�(O ��roڄM:����F�3�h�bc"O�ۖ�׾A�<	�S�Љu���&��@���ɰ<��ɏ�E���@Y�V�M&�!�ʍ��/ǯ b�'���'�~ �OK28�l	�cKk���۝:�����Ȇ_$�)`��:8�|���/m�Ɍ��"f�~�� sW`�4-p����9\��'�X<h��$R�zx0#hT���-bQ�'aRY�D�	R�S�db�x$�d�ݓ"Y���p��ybo��"��z�̂00��w����y�L�>�+O����H}R�'��S�>��3`��/D�Q%�J�)�x�T��O��d�O����v��%s��#�T>����N Y�������k�>)3�/�r.l�lB}�}�l$�*"��d�%%�lX��,�9�<��c��Ă�4ڱ�ց�t��>1�؄��`��W$����6O���-�O�A'dP�t�\Шt��"wҔAd�'�rO��
XNd�w��:'_��>O�@�$A�U��ş�O���E�'(��'G4l��H��W,u3t�̤%��%;w��~�b�T>#<��G�tJ�t!Q�k`!�E�>8��`����O~�8VO |��!��C��[Є��q�G�a�\��9�)��(1�)�;0"��h&�Ft��L6D����.ަIY���&�"��A�7�-Ƒ��Z:�P��ܔ1VbbM�[��I��?�UC�5w�\����?Q��?qr��x�4�dL��$V����
��/�~2Ą���>�u*G�OJ�\��M,%gfh��B�^?i�b�Ix����V�U�Ճ�h�A�2�+򭬟p�2/�O����7#��=��h�D؄��/��fG!�� �`Z���"j�|�C��D�L-���Y������4'LƦ]��ŕ"~�P�XB"��o�|Y�՟���ğ����,.�u�	���'L�I�	ןd!�o��@��\��L@B�(D�:�O��(�V��,�'\͊=+r��5
E��/9�O&a�'"mE(I��0�7L�cҜ��*���y�)̩UWе���S;L����Ԑ�y�&��L�C(�SD�@��dШ�y�"+��9`z��޴�?������U���A�dQ����#����O�$�O -�bg�O�c��'c{��[Tc�x�T�Yd�)TF��Dy�����=z�Oq���p�E\�Lw�@�� v ��d.�'\��(Wod0�s5,�!>*��)\�q�`^be��T�/���񉪗ēux�y	H5�PԢ��Eo���D�QCp�i�2�'t哪ghy�I��d���4�,�!�G�a�T˄/��v�$��E�˟��<��OlB�L3��	P���54U�E��@�C "<E���+���Q"J=���ٗ�9jJ��B���?��y���'-zY�5��
��H##@� Ƽ�' ��#F,U�]�H�AG��ɂ��DBI����L�tA�r�N"_h�@fI�N]����O� ؆�҃C�����O����OlЮ;�?ͻd���!8 %����e�$F�L��,�����:Ynx�u/��[���(@`ҫ%����=L����׌D��9�¡�
C�� �h$��$��'g\��`M8:���H �̸DeN�S�'�,����Y�LeIW�H�:��E#-�S�O�n��A�b�r2P�.�ptAs�V�1y����O^���OJ�D�:f���O��6<�D�O�4P!8p:��,\��g�'3���-O��"���qϾ0C_""la�k��p>�������;�*��-�2#Ů|����T�HC�=W��Y�a��"�Pd���/\-\C�I !2�z�E
?�v���a]mp���'Һ8��'j����O�ʧ/x.a�C)����0;���36���xV
��?����?�cm�?��y*��X�3�+XF���K];�BEp�	�BT�3E�hIR��57�*խLB�'��$���?	��?i-���"WN��P�F�
�JP��:t�vf�OD�"~ΓJ�6Ś�����r倰��p�,0�O�&��$��{��i����:6�8�Ci�RDI��M���?A.�T�q��OF���O(!Q�	��U+��	���P`DB�%���D?�|FxҨ^�=��\��E؂(Vpa��Z#�d9���)����p��8a3�����/���i ��C*����S��?yB�x){��! b����E�<Y��aBA���M7p7��v�O]�'>#=�O��]b��׌q�V�	�C�u[���'�BCڵ*4Sw�'���'$�c�~�;?�i�D��cF����K62����z�a�'R���w�ˮvo��p��^�]��,k�'�)B��)�O
}C���`�*���N�	���OՉ1n�O6�D�O�Y�p��vy� \��8"쟷a�8��)-�y�g�~��Y ����S���i��("=�O8�	�B�Q�40]I����+&52a�Q�
 .5��?���?�+�?!���$'�?Y��0�*�pd��p��QjV��3d<���Ih�ZRTJЀ^0��&�5Sp�݇�I=
�D���O	�6/G�:H�H���S("��L�"O���hDF�1�� v-#"OB)��S.����7���i!���2O��>��gş2Ǜ��'�bX>�xG�+��]���V�;�De�FL#*����Iǟt�I"L����i�S��� E���SȎ�>��% O��(O��pS�� -��@sb'WPdk���m��<����hG����71j0x�ʟ�<����$�y�:%TT�%�h[�H���0>A��xb)�=c0�!DėC�n��*�y��T�	N�8����3�\�C����y"E� ��jW%�`[�i�䣋?�y��	OZ|�B�T�UQ�zWϕ�y�2Z0��F��!Pm��2�OF6�y�G�V�dm�@[�CP�	��Y��y
� 8M #řOz~8HR�F+Z���"OX��ѪJ�y�:�ʖ'�(���Q"OT%��$��N
�"G���1��ʗ"O��׏GL2<���7l��0�"O��"�+وz�.}�)�2�ԑ��"O�T��K_�+�z���'�����$_y�<q�B�􊠃�_WZ�%�e�I>>!�D֒y�9�UBȭC���iC�S��!�d��X2RhSׄ��D�;�(��d�!��ȍW!��r�P�Em dq���]!�-_%��(���9��EјY�!򄜯s���� DǤvP *@��?_�!�� �ArX[*ƈ��1+�V�!�^{��`p�e�W$����9�!�[i�(@ƅ+Zi|�*1�	�!�d��AJ������yb`pB��M	\3!���D����BQ&�#�W!�dX�;���G��[1��s��z�!�d�N�@�_�:���P͒��!�d�'6޲�i!�3O$B�
T* 8r�!�����MݽA�=��HY�!�E�H��� O��z�ȸ+@��4�!�D� o�Dj��`�Mx��!�$P&f�p�W�φn�)�N�$!�ٕ��P��X8]��sN�%!����8�;�&*���65!��� l�f��.�� ��81!���gL�-���7�� S\�!O!���]�z4�K�	����!��aK!�$X�| �}�B!X4ADp�
�(!�D��D�`��vDSzފ�Z��ة5�!�$[w���$��s�hG�S�`�!����Ld� '�@ּ`6Ƌ�\�!�đ3Ta��ӗjްR$l��3��!�D��R�*I�	�m�(��"J��!!���o���A��s���%h�\�!�D�����K��l�t��K�!��  Kt�d���G�9xpq��>�!�$B'&�� ��G�}��z!��0|/!�dȄV�h���;r@	�F�
~!��D1t��� &W[�]�Qn�=�!��-E@B�L�<��8�� r!��]+p艅e2PAs�JE,v�!�D!!�&!y���/J����#*�)�!��#`$:h�ë�5Cj�E+�H�7o!�d��1<�(#`��-����"i�~~!򤊍s$H����K�\�E�U�!�ݳ|�����ift��E�5K�!�$YI��� �hb��;��  �!��@>�2x��?iW&�dG��!�ě�$�.�7��#,rQ�p�αF�!�DC(pq�̢d �-}�}J�.@2[�!��Rê�PjOp�؁"-�,!�ݘ ,�P2U 2�ˀ�W���>Peh��$1!�*�Hqj	6�\��
�f��}R
�b��/]�@pK�W�J�#5�ޟ
B!�$D�[ �{Rɇ^Q����ў�J��F�O�ɫb��(�q8 G�;R�|��'���1+�E�@�ʀ�JOڸt[��B0�>��O֌�(�d�+t�/ ��%9	G=�)���!D��T`Zv1Xa��،���Ea�tc���:@$����HFqO<Z�L�����D18,y�A�'0<Y����ᦹkR��#���B��S�leRpk�D2?�� ч*Y���D�b�!Gn�=`��:�� \ўP �YgL�'56�H��� �]�V���P���Af�
�9;^�"ON)� �Mv�z\"��	\ 4`���'Z�� ���g��	E�����ᓔ?�T�9��u�qy2�DE�`�ȓlP���m֮  I����(���}]f̈��K����b�d�i�,Ё���E/I'<RE��I%8Z e��i�H�V���\����G��n���O¸�_0�*	ד,7���e��l��x�g�@�t��D|��f0�O�pB+�- �p���|��`W ��
��)�"O���RǶa|ph�%>
�!����'EE�\�gOηb���
�Sn��� ��n��x�h��I��R�E &"O�q��_�w�5J"���<N�u��$0��zs!@�d�Z���'�>��f�Od� ��2g�3Gnlc|�Y�"O�)s'��A����j����2��'�|�� �;.&8�UB
S��(q���/K`�[��&�K#
�T�azBe!HD�$��^
~X T����)Ar�vMZ�����.��� �r���Q0@ɖs\�aR]�.��1*���i�B�"h"}r�ܯ�)�l;�~Zí�W�P P�� Q^�����^�<���("<<������9�NعC18�� ��3�	Q��ޒB��U9e��~BF =�j�p0F^onͩ�̇��>��ė"Y�tҗ�F1B��y���"��6�|��^�9`��&��(vO}��VQ�'�>}聥�6I�F�7m��mX0Q�����8>��Ve��%#f���N�l����w��8��[�_���� �/?�^Hx#�Q�C:�~2�f��%���ǣf� }C�h�8�M��ϖ$���z���/(�j�q�S�\c��P����+}����pKO�I�N���'� ,�0 �Em)�ĐN���ТK��O`�j��9�V*P�a8��'��C�.҂1M���+6<�q��P�����eƟGz����(ѕB���2�X	Ω���O\+���#!,��茊������	���컑��	}Q�L�g!��<y*�Mz����Z�|S�\zy,թ6�l����o�zD���<AR�h7�_��|j�L�	.p�p���"�<)sIݧv �e��
('��(*�Ó�r�|�>�ϿV����� �õN�0��L�<I0��ge֬x�D��snd5k���DC� z�}�џʭ[���67g��h���}?����<L�`H��f�u�*%Q�F�EX�TH�"�KV�q��k;ah�Q��э:�]�r�S$�?�n@95��:���%k�>Dp�c[�'锡����j5n#5 ֊r��A��D�4J�EP�G�Z7��cU1��^#���@L�Iy�8��5F(�8�1��M��~�N�q�����U,5V�2��ֵ�?�G�AJ\�Pgh�
3il\ɁFO�S�4����K�n6��S�o�����"O�Y�A�Z9d_���Ԓd�,d�c�5\$��A�y[>}���˒������0�g#^�M�ܛՋ�!��+3�O�	둁�[qb=�c�@�M���w�U( q�A�b�'���Ș�=�X� o
h�b<���P�x���c��1�ŨOW�az̈ <bՃ�#� ���sI�3 ���jL�m� IV*�$8t�J���sVj�db
 r��\$���+#�2�$���#'%J"�@!`�8��~ڶj�a���Y�&G�z~y��f�E�<I�lž>,�*R�'�-0G�ٛ$NV��W��bu|p`$��⟼G�d�HS?AR�ƙ2G�� FdQ':���+M{�<�pÕ�KHp�7O�G^���M��K7\�Z���>s�P�u�U�]�(�p��,i�@kGN�<	���"�%F +g��&�
���=�vN�!-��a��kA�r��	����(
;P٩@��Fx�(�D��*��M�T\j���E:�+�- �N9dA�=�� M��M�PBՅ6X.��ӞeNv��ԁx��!��J#El��O��aR�Ka�S��0#3��b'���\�E�@l��AW:ݛ��J馑��㐛�qO?�k'���V��{���	:��l�(�x�0��	��OǸ�{w��UDf�(��)ulHQ��#{X��d�O��0Tϖ4�p=����	�%7��г��Y�Dj"c������?��W��h���k�C36���)bd͓J�$P�*D�L�fF�B�!
������Z�'���?$P���4.��(�I�?�c��H����!uXɻ#�O��0
#�y���=
��G�T�Kxtl����5�ؠV&к1�H���O�&kq���L<AG*�cMb��ڠ<�Jט�d!�$�w�|�����a t�āl�8�aإ*�(��V�& gN�|��Xzre��zi�h+T X  �\X�'���Q#�Q�d��'K��H%JC�b� �����,�� #_����a��H�Ԁ)�NZjh<� �t@'@�4��xbqk�UE��r�+}���0ib�c ��n�`j�n���5@��&zlK�wy0v��nJ�M��Ҝ/���*��vqK��@<T������L�ZHAgʑ VU�� ��U�;�h�P��$f�cS�A>P��g��ɐ`��ʧ,t��3���
�Т?�W,��𙳞x�h̥o���Ȓ�C5.�锫�p�F]���F�LɾU�t�X�9az��[�B{�L�Q�F8�2�V�����ӏ8xE�Z�)�Q�����7[����0IA=]�Yҁ�L!��ʑ��!�(�S��zQ��n�<	�(�qO?�D �cX�x�,^�7L\M�"-��!�$N;Y��q0��f�(0@ ��qf����w�c�1.��qLJ�n��<�梃�[S���
�~mI�8OE��'O�h��ˎ.�n4��"O��Fb:,�PD�6�� 
�B��	kJic��)��Cr*� ����t��"� �!��B*&�Y�aZ�A���⦦4U�!��ݻ w����*�&2�©�`@�2:�!���5o:0Ċ�DG���QB*2X�!�d�21�<�S��Y�S���&�H�+�!�D�{����ҡ�7(;�8�\6�!�$�o���a�E)G�.M���.[!�$Ɩ!�Y���u�p���)Q�;!�$��b4YpkկZ��<p��1
�!�$�0�`���$��uǰ(�̈0!�d�F6���ꟙĶ ���ϴH�!�D׷l��(�@��������2�!��
N��17mG/P��15�B�!�d�\���i�o���*�Έ<!�$�Xk�I�ca�>8 ��y`��/�!�D b�Pą��b����*?�!�$��rY<]ÔąR�01c�C�Y@!�đ�|H� h������刾-!��^*IL�%
��D9erd�e�!45!�-me��ys��md<�G�N2`!�$�P�P�	�]��	�3m�!�D����A�6#v��`0ȝ<[�!���5�|py��J41�D�t��!��1�D,3h���v���Ę$e!�T'-B��Zf�ׇ$�h�τ�,O!�	=����;5�J�붨��s�!�䑰4�"F�( �t8��U�!򤅆6����A/H� �L=�"���!�d�)c�J�h_�]���0e�!�$;�>��E��ͼP[$h��<�!�$ɑ��5K��-��M�d�V��!�dW�Tz��ׅ�J����eӸT�!򤋞o_�m;�K�
'�,����D�Ey!�$ؕI��\�0o�+Q�%�6�Ɖ9�!�dܮY�Xq*V�RI�� ��N;W�!�8$�Nt)�b� gc�J��R��!�d��u���� ���	Ac!�ܿ���DHD�d��(�!��"&�Z5چ� ;.�Myu�U=�!��f[����Ӓ�Z �d��6�!�$_�"��L�a$H�ph��$� e�!���vTH���|��Y�Mɔ7:!��7�Y����Ф��՘e!��F� }Rek�jy���{^� D��J��M=Rp��U&X�&R.�XRI2D��"@o� #i�X�t�B��
���C.D��H��;�)� ӤB��z��(D�K����Zv��%Ï-���� %D�Ѐl�(l��tcҠΈCU� W #D���DO�=#l��	�j�P�
@# D��!�N�)�A�5mC�#e>�T�:D�� �ę�`�1Xcᦔ�d�tГ�"O��Dl���PFE̤f��)"O(�Xr�!_l$�6$5B����"O�`���Q�TG"T �DƯ ���"Opѩ��#P.���"�Y�E"O ���|����D�m��1v"O�lZ���� �ӣI�S�X�"O�)5	�:Z^�IS��v���:c"O�t���\�*K��� �����v"O�L�!��m��š���b���:�"O܍�E�g��L�2��$
�P"O���n�C�X|��NP�V�J�k$"O�m�@_#Lbz �1��9��yG"O̡'��9[�hf���Zt4"O�|9��ӤTd|�vBU�m���IS"O0�:�*���+���)nDR��"O�SgiLj�$uk����E0� �"O���&m�.��T��`��o�L�7"O  z�)K���'��"Ip� �"O�,g�D=\�h���9&#���"O�0CQ�_�h`З���7eP���"Oz�*�$	Pp�A��_�2��{"O:��u�A��Ȍ�{�JA�en��y�c��}b��C(ԇqd�5:dc>�y�I�?�`�	�ʷ~ST�ڒ�	�yB�.�PͲ��f�0�s��C��y"N�<c�Q��"�b��M[��ɤ�y���U�$���'��n�a��$�5�yb'�|�9��.`檝p��C�y�(�|*ƍ�T��4%L���CD��yBn��?��Pp��'�� [����y�C����PC*L����ZTƃ��y�ſKrp���n���4�C�ʎ�y���bh�,�1�ɹM8(Q���yb	A�H���
'�h��g��yb�ЧH�hX`	F�q�H��.��y��7g4E�7���c}l�H�����y���Tl��K�1^*��
4H��y"-L9�fT�S\�P�H��f?�yr�C����3ƪ�0 ¬�y�M_��p�kƢ@�0+�<�r����y�h<!�p1�L��33�:�y�+@�4�Zh���G�4�����y�ϛ�5D�S���H�I���۟�y�%������@�J:����!���y�B�r��y9���7.�:-x����yr�s/^XА�� \�#U��yB��&��ipU'�2l��{$��yR�(�8� ���&�!�MG��y�E��w��M{'�J��� KA$_���'�ў�p$)f�9=0�i�" _�+|t0�"O�D����FP�=R"�:E%����"O�1y0Hɷ �4��N�v�D���"OL��(�*���-۩���b"O.��p�&Y�Ɛ{4cLm���"O*�
�Y�{X8�{�Q]@pi0"OH��R��ln��#��Vr|�S"ORa�E�	Bg���t#��r9�<��"O�9֫Y�$����!6�p��"O.��%Ӽ��yzĊզ-� "O���cM�4��Y!aiήP
����"O6-�a)�*tr�I�/9h(��"O�bA��_Xza��!5)6`B"O� 1���ujX�Aa�n>*�	&"O� hX��昍+p��kg`Hs���"O��$O,aFd�Y��(*�A�"Ojp�c�	�VH`�E��/�,�)4"O���ъ8m:�QC������u"O�"�}���i7[�b�ޔ�w"OrxK��ݓ1��-��% vX��"O���D�4,�ΠI�F�(g^�B"O�)����n�X�P�EuMJT""O���$�H�ĭf�׺)E�E��"O���Π�>��Ȇ	�^! �"O(aW�U�.��b�K��5�Bs "O|ѐ�MQ<l���*�\�ޝ2D"O��z��ѥ_�T\�ъ�m_Z邰"O���3��do|�k��6J�r r"Of+w*������@N<9y��u"O̬��'G|S�aN�0���1"O�	Z5�H=?j��0���'u,��3"O>�ɡgT<�����+��Qd�T�"O�1�N�l�H���L�?Ґ�r"O���uO^>`�a��=!�Mks"OF|! J=lZE�u��J1�"Oz�x��M7b���3(B:U��9"O^=y�C��h2di�&p��ͩ7"OH�W��H�ܔSU��qjFe(�"O�jbj�OŖ� E(S�	O<�'"Ot%�!�D?B�Ɲc�L��?� R"O�ЊcbϱY�����
;3�exR"O��j��ޜ{Q��Ä�M<8\mط"Oh�B`��!d���j7�ʴ �ґ@c"O�H:� ��|��g�a��Dе"Oh��3�ʑ"�GG��5��"Oa���	".0���6��D�Xa3v"O 0��/�1���EڧW�>�%"O��q�ê#��!Ã�4vo���"OYQE�B����ᗔzU�B�"O����26���%���8�ҡ��"Od�.42��tO�
�F��b�M�r�!��K�R��Wd�KM��Zł̕B@!��z�[�"�.$<nP�v/�'*!�ȟE��H�\�nۢA��N�!�DP���	bd`S�7�j��"�;�!�Dׇ6^|���������⦢�48�!�$��t5Z��q��(Ɍ8�d���V�!�$Ƹ}��x�fˋye����!7/!��ԢD�G�a6��1�$T���ik�@��kͯ ��02�MeF\�ȓ1n4���O0h�0��b"�"}��Ň��X)#�It���$��PGvЅȓ>��x8Ԯ��@�0��ךc)��	[�'�T��f��a0�y� ��&��5�J<����iĹ[P�L1�nH�lu�e�nJL!�ė�Ef�JQ��a���R��d^!��ذ]�yJ�KQ�l���IuKA��!�dHM��0Ӓ,�$l�@����ʀ"�az��D\�w[�k��x:��6cC�}�!�ѷVgz��)Լc(�O+!��	aЦ4���N~={�FՂ�!�D�/O�<�e�Dd0~�",U&Qm!�ě6s��) �X(x%�M+!�V�HV!�Ӣ=��x���l9�(�㤋�GH!��>3��e逡d1�<�A
��A!�ŬSǒ��"�����u?!��+R����
V �f�g:!��X
���Q K��eeN�.�!�� ��v�@:6�H����� ]4�W"O�9��c��:G2ٚ�L��?��`�'"O�T��N$��APkO&O�����x"�)���V�Z����7w!fM��ӈ%LXB�[f)��	ݠQ�R��IX�jc�`S��X��x$��D��r���R���g5��?�U#E�D' �"�օ5̱I1�^ V�����|(<�`e��8�R��sn٤��h�<1P�E�4��a�/����|�<�����b�p�#�]�t���!�z�<�$vqNǄ�b��y�<��판.�$1HDC� P��L�c��s�<YgK��Ia��T�E���� H�<��'��5�&OPBX���SG�<��jZ	Z!8�.V%2H�|�o�m�<1s$ٚ"���������Zb�i�<��V-",�5e[#|��}J@i�<��aD7j4Xp`&�'����7J^h�<���a$����)�"l�m��&�O�<a,� �!�!ŎrS~��P�MU�<I�I�4\~��'�Ō1s��91�Gy�<�����j��@  I<>䪷�o�<���T\T�8u	��`�̹�w�p�<�c��?,����	4H��ljI@x�<�ч[b��C��$+�rdrE�M_�<���L�(�Z0�&'
�~L��M�f�<�T�Ə�b,�Ē�w98�I�!|�<���M�����B�OO�����w�<�qI�sj	Q
��-�qD�Bq�<A�j8wS�I�G�n2P���i�<���T��Yڀ�Ķ��u�G�F^�<�wȜ������(����4�Q�<�!�_�{<X �Ʈݗa.�(ʱ��I�<@��#&U�t*�NE)���RL�F�<a�M��H��S6���y�<�G�/n����٘�Di�m�<Yu��7!�.x宏*K&�H�f�m�<��Һ6�r��rl�������l�<�G��S�|0J �P>�XG�L�<acG�DL	`֒*f�Pa`�K�<Ѡ��${s��R压�A�8L�E�l�<C*�1�b��0l-� y�%��S�<�$n��}T�$�M6m{a�O�<�o��A��X��Ȼ���0�ˉH�<1 aE+x��H�4.��~|���B��I�<!�� �6 H��5G�t�
��MG�<af��v,�1]�}ϸy�vaOW�<����Zܠ�0m�<���
U�<�t'�e�0���&וj�|��IU�<��'�7e���۴����y�͒L�<�"�΃f�B��	D)H�Ң�n�<�Ký8�Xkb��u2�3�A\S�<�u�I�Vd��{�J�
A��E�U�<т���At��� �dP�er��U�<����r�	P��O�B��4-V�<���Yߴr�d�,�"�y��N�<!����H��ɳ��;r���L�<1���13�ڰ� ܀G�EY"�Kr�<�c-O�'^��D�<.�z�;4��o�<ѡ���o$}��8U�L#R��m�<a��[�$@��U�<�t[�`�d�<y� 	�����t-׬�����Oc�<� �4hya�@�)w"ɒ.�_�<Q��E�x](My����B���`�<� xyRG��}�$i	��8�z��"O���GE<l<�3EǱj���"OB��J��1�᠆�ђa���"O�U���� k�8jdcM/_o��"O��� ��>%>P"S"]��>e	&"O�`�u�>_v��뎼iB���f"O�����
	VČ��ai��?j�J�"O�q��iƚO��Dˁ�Т,<8��"O�r��ň�����M�)��HP"O�i���
�K�T�e���'"O�(�5c�~�@ɠ�C�aq� p�"O8ySs��8\�R�ɵ��HSH���"O��z��I�<���q��33`���"O���
��l[Δ�w�ǈ9/�j�"O8��ʞ6v"�j	�$�� "O��Ҡ�*W���T �(�"O�T�HY ?�b��Ճ�p���"Ol�X�+Ƕ�)e"O/-cx�R "O�� O�d3�q�aA�����"Ol�r�*V�.����{�v9§"Oɳ��`��c�Z���+�"O��v �?�&��2f��v dA��"O���&���˥��b��3�"O��RAG	U6\�����7F�̂"O��e��p�n��R⅞r@�8��"O@�[aߺ$�����A�3]�Z�s"O�����[�R�(]0#�0�Uz!"OV�R����L��� S����%"Oz�bb�<��p0����F�\h`"O�DkD�ъ"T
�ٰ�!�n��Q"O�髷�ߛq�>�CE��g���*O.�K�۾;te҆�/rn��	�'�P���ǔZ���6!�r>�Q	�'��i���)4�T��`͊v�V���'t��ׇ\8��TZ�I�-gY�dz�'A~��'�Ųt2u�$�܅\�4Ȑ�'N�}����kȨ�TBY>Ɯ���''\ �"�ەo�L�Z�_�e�*���'��4���M�Ӡ�QCmU3P�4��'),��i?�N`X��ī={�� �'�H�2�a^�u�x���92'�S�'�}�W�V hs�T@��*�����'Wdi�DK-`�\��J�yq�r�'u��cT���Iq�B.#Bĸ�'^�Psp��%sV!+�b�-��H�'6Լz��FrOFM�GI�8!D�
�'�d�h6�Z;D�m*���/��$�	�'t�@�5&�!����e�Py�1z�'���9��X�v���	 5����'��`�YD���9@)K A��U��'&~t��hOZm|��g@4�2eR�'�f��3���ʼ*G-�0)Uҙ��=�T���Ж!��P#���b���ȓj~�,���ŏ@��)[%A�Zk�d��PJ�-�F� j�JT�3�Αc�����v��$ꃂ���4�`D�#�q�ȓa��U�qW	�^��	��/�1���dQ�%��U:ZшߗUc&(�ȓn~=�ЇǸ#�~XA�f^�+���ȓ��Ya
O�}>�$	 �F�V�.���GnD�)�ר
O�`뗋\�p�^���w���D�3.�SG	l �����T�b��%	l;"�P
1��ȓ;�a�z	:u� J���S�? H)q�Dݡ.�4ұ���Dj~���"O40ٷ��k�ajt)�@��,�""O� ��K�1&pk)H��̩�"O��#����
�@�;��C�j�2�"O��4΁��4���M�w
$��"O��QFV�+��l�,�-b�a""Ot,"���uE�PQ�
�K�s�"Oz� �N B�r�K,<w����"O�Q�v���t���݂X_����"O|E+�l��E�8!����%]$�I!"O�qbF��b/� �7��s����"O��Xb� �$Q��̜�+�(Qi�"O��k<=�e�)��1��l�F"O����D�7I�����\w���"O�4�Ŏ�(F8��`��&i�j�"O��"��)p���	!�cШ�`"O*��ѥ��J��e�`�!	[z��v"OH����E1j$��RO@�C�a#�"O�1�"%�
�I����+��ن"O�S�C�=k>�hj1ț8% �BF"O�����ܱVQyǨͷE:0;�"O�����X�3�(�Ĩ&I�<<9!�$^;�H�7�Q(�,��%h�4 !���`G��W)Ӽr�8 �WD��P�!�$�"ܶ����B)�"Aa�@�!�d � �����P!#��uAqA>9�!��Ƴ%-�@
�	(7�&E�� /�Pyr��nv$̻��f��$gĒ�y�$�3e��x[�H�?lBHSĨ��y�$�3~���h�B��B���=�y�J�hR�a�e�ڕ���7���yb��5�L=�P'���ˆ-E+�yr��`jXU�p�0�>؃P��y���+D�X��cH� !�K�y�i؎	<�� F�ô�2x��N���y"nS!4�JL��뉲]@(j5 �2�yR	�x�\�f�[�t��5��%�y�`�L47nMj�����y2-�0G��I�*�$dozk��5�yB�
[��
�@[R&�����y�*�'ONșWMD��8����y҂K�7PaS�ѳ���xG�a�<A`��#d��Ijg�j�8�r��N�<QF�z#h}�@��X�C��UT�<�C#K&R�P���U&��ӳ
�L�<� A�Tn�pL}�eʢ�y"l��e�mr�& �І�u
���yW;x�T����D?^I����y�DŢ8��805N
�~�sk"�yE��T�@�`,_)(J4H����yb��*4��hs��9|z s˙��y�)K0sˆ�)t�X����AM%�y��I"�����U.Ib��y��X�#O̰�gx���b�]*�y�+�7�<�*��<]Jx��"�+�y� F�Y���Ņ�W�D��hͦ�y��K��!w`��Gfx����Y<�yR"�]�8��*�̋t
���y�[�!r"�$8�}�W��yB�д��˱�U�JϺ̘D�Q�y�GY
2��P�@g�%B���hAm��y��24'�!�����Ї�/����gs�m"�d�<�h�Ũ�pSB��ȓ��%	���8��Q�Z�u��S�? �IST�G�2��w[�R'��j�"O��+Bo��]ʦ`�B�p�`�S"O�a�Fn�+; (�cN�lHX2�'�ў"~"��^h��n������k��y�&��g������*I��Q%�yEAF��$;BL��c��(�&�8�y�aI(�d��Z�X6�8���>�y�`����y��Lt�)ja�֪�y2c �1��9s�A����@��B���>q�O��ZC�D�ڴ�P�!p�rph��y�d��,��x���Z� ���y�
q�*�iC�@!z�����g���y�"�)RF0m�v���Z��<�u�݀�y�(&'�A��M^�M�r��yb� ��|$h�c�1v�|��"���y�ǉ;U�,��d@�� .�#����y���,b!���98,!T��(�y�뚤�2�H���~E�x�G�&�y��>0~؃�[l�A@�K��yb唥~�n����<]���rl0�ybɎ C'h�Y��ҋ)6�t��N��y��Ȗ�n\!g�'��=��MV?�y��Q�	7~���G�I2� <�y�DLbx��\�6�V�J��?�����e�][����C��5	ӆ.T
���w"���h�
w���OM)�P�ȓz
n���X(X�`S'қr�&���M�i��ţr0��`ѝ_HD�ȓ=eXX�eI�%DR�[,"�b/D�A���N9X��/N9I�B�I�7��lyWN���t�@EJ���D(�S�OyQ�7O6V�V�_���R"O�$(C)��J�ъ@�A���Q���I�<��`ͣX�uw�S}4���e�H�<q#▕9�>r���M�a�� H�<)��&A}h=h��V:*F$�T��E�<Yf�4>.�ݰ��G�}����y�� ��z-_5I��듨�-���䓫hO 0ЗM�RY��RN? ��$!��.D�ȣ�A.]�yx��+V=���s9D��1U��""��H� P�$=TEJ�"D��0Q $j~��25��n|4ux�?D�0�6�V�ҦX��̌N�I�$�>D���0��2���y�ꞷ5�A�� D���@"��,�z��5����i?D���SaO��|���\/j�0c�8D�\�`� {�tI�HN�E$���!D�����aЧ��b���a4C>D��b&E�D{�����C�9�m<D��*$j &I��| " [��1�p�8D�`[U�:M��D>A/��c �4D���N͔Vr����QW�H0	'D��k0H�5"�5��N�	+� !�0D�dQ��{ܔ�b�b��mD,�b"-D��@�W�I��1���3`0`[r�+D����MS�X���T)ՃW |r�?D���h�!x��b�#P��}��=D�,:��N�x�`���P�#
e��9D�pQ�GL����R�΃�r���*5D����jU(��TXr�TT�D��j4D��Y���
�����-mL�ՠ��3D����a7i!T�`"��ظ��p�&D��P�BĻ;�vx����'u�-�#D���"�
�4�RvFJꖉЂ�#D�� p� g#GBF�!�K�m��R6"OX���o��7�z�1����c�:0�'��8×��'z��0˝�Y�p ��0D�p9��K�[�`����ٕK�H!��)D�xH�IµLw��o˧l����g5D�d{s�Ԋf�$YX�	�%4@1�1D�XA�!D
M<|��g��s����=D�xsr�_�/���էN?KQ@��%D��Hf��,f�R�X�h^ξ"�o0D��aB��"�5BuТ1.ԍb�F<D�H�$	6	dё �$u�M�wI8D�xh@	�2�p9����q��e1�e"D��2��έ+���AtF��J�Pً��#D���v
�nf��5T�Z%
-�4D��p��J>"�h�L�
k截v�5D���I�&�ع�S�ըO۪�1ҏ0D��qe��D릙A�S�o��;�B9D��U�_��ˠ	�IGR�y2��O�C�I�UPD���@46�L��A�5^B�I�4�ƌ��5X� h��8�*B�Ɋ1|�zW��<TP\�`'"ٰ1��B�	�=;�, !���V��U�K�0��B�	6(Jl��.�M�d4"�t�C��쐃r�c`�Sf@T9jC�I���:��6��!(Ŏ�VC䉰r�e���cP�a�2S��B�p����+ϗ+2Ny�c�K9B�>[ �V@�N�҉�E!1g��C䉳WjF�bӢ1y����b�vu�C�I3mԾ�!�XdV��{/�B�ɬiX�cW I����[+�^B��0X鰨�Lz4���X��B�I�E@*����,i�8Mw��'�C�	�w�T��,�r�V�@$�НP�C�	.-�jxZ�U���Ɛ�C�rC���T��40n,{�R|��C�1CU�p+%.� Poh�2eNR�
ubC��(�P!�1cxp����2�(�/O����B�>���ٖ���S�EH�!�$�6w*�"oY�C�T�0Ϟ+L�!�dݏZ�.U@�,SJ�\�kR�Y��!�$ϫP����0��D�1�:x�!��G�o$d\ff.�����\ @�!��&C�0L�O�/BwнKw/ٞL;��2O�	Xc@�X�XŠ��`� )�W"Oj���GI��~�YbD�0D�	��"O*�ʃZ�6H`�!�D+c�>��"O"��,��d���d�X�]�4���"O�x���K�]|}yr/Ю#���IS"O<E"���P7ָs}4��D"OD�Z�"�.�847.֫j^A�"O�[��9M]��p��9�ֈ�A"O�yv�	&r<9F,�q�Jأ�'�!��#y�C�	DH��	����K\!��Yzh �aN�N߼��u�ީ0R!�DG�O��q��C�0"��e8���uG!�DE0Bh�u��șzV�H��3E!�D
�����G='������Q�&@!���o���3�:8�'KYEP!�Dɧ|V�����	;Ҙ8z�� G!��R�\�ZCj��m�x��/V�5!��FA����G�C�.���.�!��1hE��e�'-����7"Կ-�!�ċǪ+�K�A�|���R|�T���G~
� ����
�*a��PB�"\%^�3t�'�!��3���#�!��� ��JU��)�'
����a��`�% ����	�'��D��B_1CJ��`$�(~b�%Q�'�n�K��8�,�*Y	E`�,�'�����e*�t����:�4�{�'�6���-w�0���*N�I�'y�@�@�C���9��-�$#��QJ
�'��薊V�n����#�="�
�1�'�$�deX�\�|�{v.�?QIZDb
�'�!X�%ԐmjF	� kM̞��	�'�h�� C-Y��Zp#ќ\\^\�'�@��)�+8��B���_��8��'�$����MN�!��dݦQ�dP����)�V ˃�o��)�Oغ:�N�S$�'��	�4P�� ���o�*��=9e�ʓ�hOQ>�{v-g}�{���,v+!C�����O��"��SVt�)�C&R2I�r��-H�B�ɴrH�U)����YY�Up�ȕY@B�0ю9� � ��U#��U�t2B�	�: ��3l�,z��{��S�F����+�	�:�e���ɯJ�Lq���r9Ԣ=i�$}:�%�]���X�,!��m�ȓe��F��)2��$Z�^qʔ�'�ў�|�ŉ�.Ln�U!��=f)&��Р�n�<�Ra�#�`H�D �``8��Ņ�D�<��A�r�r�Iܱ��$iqG�}�<1��<hU&͚p⒄�zQJ�y���Γm���"�LK�������:����IB̓9*LQ*��+o���f[�D����332Q�f�<�t���F�E�'7��'?ɧ(�����,D*CaH�AV�\�yMQf"OƑj�"A�8�r�@�ċ_n�� "O
���C'A����-��<��}�"O��c�DK*bJ�@5�b�p���<�Va�;t,({'$�(W���	�Bx���'H�P�w��K�����;Z�I���:������0��E(�g�3eM��-�yB�Z#.E�S�o�2<���
��!�$��"E�IK�#�6d�����D�!�R���K!B͗G�����`�2}�!��,B�T��lN�\��9�Tj�%F�!�"3N����	1
�T���/o�!���z��v��S�PI��7k!�d�C���D�[X��%(ŕ�!�>#},4,RJ}1�\�`�!��3Lވ;ecX;O�X8�&A4�!�d�%�n����E�u���p�eQ��!�$\/�ʼ�E�Q�f��Px�C��!�S�l.��1��P�2�U��`~!�D�-H��3�ӦC����w	�4c!�$��H؝��N'=�R��7(�=0R!�d��Ow�x�@���zd���g�!��Oh�hɅ�2-��%`i!�Z�EF,=� �|�3��!\!��M���2���=���`�9_,!�Z�S���am	� �`�vOK�5 !��%�3К �Z�G�g !�$
�&���5W4�H
aK�k�!�āu����_��zVE��!��#:^�H�l�\CN��!$ȴ.�!�DK<�V"��SCJqA̒D!�d�	bqɲ��	@�:��&�̿%!�C7���r�&Ƀm�ű�.ӕ!�!�� @�slJ-Z�2΀P�J�"O�܂��ƧS�b�5�H!��"O��$eЅ?��p8���W���r"ON8�r�VS�A�G�"*�Ѐ�T"ON�� �N�S�b[ե^���"O�ձ  _!���BM wP&�1p"O�Y��ba�B!�l�ф@�4!�DқR�" c��.g�l������OZ���-9�P�	K��R5B���!�S� O:��@�I�r�,Q�3��9B�!�����*��_���(�Jp!�d��u�X��%�L/�ԸyV��^!�d?}v)�R��(���q ��!�R|t�X�u�2mbS`�.�	m��\����@
�H�-��j����F-D�8p�W�-�����®0av��v.(D�`S��@ܔ1kF(�m�#U'D���d�{H���$��wK\|Iri&D���f�Ң]�*��.:gy��!)&D��d�_9���)W��!���AD�#D���S#שs���Q���6�~	��!D���a��*�4!)��+��{$E$D��i�)�9T��p�$n����O(�=E�h�00s&���ȜH�v�6� G�!�ɕ3CJ=��f]�M�.tu X�!�(h�j!K�h��c���Ec�A6!�$�.�B��Aa��
e�� [9X�!���2}�@�aTg�?Yx.���*��!�d�:h����Ӂ!wd�R�)/C�!�D�����s��N��\�T+P,d����dqr#AX�f���A� +hkRB!D�L{��;<u �˓5��U��E=D�D����p��s%���!a��:D���ڷm��Ec��΁MZz1�q�7D������I2<跭��;:�	s"�<�
�sV<A$��m�jt�3) 'JF)�ȓus<�	�`^�.R�Q���p^�ȓea���5��pD>�qfIݵ�J���f��F�yO���G�D���P�ȓY��J��w�l���*0Ot��w���$�D3:� @��Qv�ԅȓ6��\���������2�L0�ȓ��=��QF� �R(�xt����<�Ʃ
%l�D�6��E2L�FϒN��O� tǉY|N��r�X�\��"�#D�x��FN<�v����ثl|���?D��p$E�,e�l�a�c�;`�Qk�"D��zE*��I��G��3�	�9�!�d+rd���$ �})�P���H��IX��(����������$���J���I~��I��
�|�����C&Y��b3D����U8w�jL����/��	��/D���pY�<Zp<�R.]#!����� 0D�<r�Olq�P9�`� K	8�d3D��°ʛ�Y7�}�DB̝A��\ڂ!,D��Xb(�R��,!�m�S��L��*D���B6Q����`���\��<�G�:��V���ꅦյ@,�#�	� j`�+D�P@�È�jB������
��Y�3D�P�A���WD�qږ�\=<��r�(<D�Љ���r\�\�@����G�6D���`Ֆ}��B����5�O:D�xiD�	4=: Xpk�1��ٻ�.7D�tqp�_�un�Y)����P�@���'D�� |\q6MZ
{��-�*U*
���3�"OX��� �%�����RpJ	�C"O�
%KYy�T��v�Z�oQ��AQ"O �+��R.�|��U�A�fc����"O���h�  2�`c�gF+jQĈ�"O`M��苬C�F�H�бh�6�rԓ|��)�9Y�ahR��5S�9���H
�rB䉽�j�Pa�	i�I��']�n⟜��ɟtDv,[���r���C4��!F�C�	#yHh]!���AllkQ���ܐC�?�V��@j�UC0�ц�U�H�rC䉢D3�u!r
��cM� �H�\^C�I�}=��:7�C�W�!B!E!��O�=�}��E�T�q�h�:\��6]W�<	�bF<�΍�ՌֶW%>�9��TI�<�C��! ��zp
�3I�j-��\o�<�C��)�ʱ���!���󅅄U�<� �9��%�K��@c.�� X�<1��J>���x�R��Y�"�Mo�<A���y�Q�W͓w�캥�ex�`Fx2$�>����F�^:���d��yↀ[ �����sD� 5�D�yR,��n~F�h��8I�]���:�yR@�}~<�v��6FZ��hac�ybW��9Ҩ��:tR��03�yLÂa��qF+K�0���'E͗�y"C�7�x}��∱�Y�q�7���O�⟢|R����W�(�ȗ�R�d����{�<�d� �N�q�ɒ�lo�!���A�<q`jRC�}X��[�А��X�<%a��X>(� I�sB�%�c��{�<)�.�4 R`Y2�Y dպ1:Ad�R�<�D�}H��.xe^��Ni�<q��+>����@<@��C��c�<y�KI�yJ�c������a��S�<��/M�[_���(��i���K�<QF���^{�Tr�� ?'f�����G�<��a�H����U�R�`��%��H�<��d՜.�dE�7�
B��9�0��_�<�g.�;V4!w��; �|!0�U�<�6�T	lY����Y�m��p�iV�<�LbC��BjM%� �"o�M�<!��Ώ w8�q�	F�-b�{��`�<QĂR�z 0��d%ݾtI���r�<ׇU�Ef<AN�;E�cw�Dx�<'��q^�x��^>x�<��s�<i�D/;ʱ�2�<k��<p��p�<i ���ƭ�2��Q�l��G&�Bh<�eɫ&+��`A܃s8��fJ#�y�)��r�%g`�!r>ΌR�k��yb� u���b�	L:|eI��X!�y"9"�Ð�,?�$��L1�yRa�RH⳩G&iJ�c�o�0�yʆ^�p�a��#M�I���y�DD��e�0��'QMf�t	�y�)�4v���BQ�U(�Ы�Ų�yΈ)h(��[S�J�"��@J���y"LH�G��Y �*�>!�v@�B���y�eK&����`�ʴ��#�Z��y�䓯=��tj�)S�aQ�F��y��ժf��U���B�u�(�@NF��y"�Z���)Y�}�~���ܽ��=q-On�� by�M5&�6*l�|AC� ��B��1{Sjp13a�a���:D`s�B�)� �0�q'�mY��²/g�L��"OR1d�S�2g����"��h0"O��`.L:�x
p,ç;�,��"O"��ц�l{�9��YKk�u�"O�d�`�w�F��U�ܠqM:-�'=�ā�w�&K���4���I��Y~!��P�H�* "P�]���as�"��!�D�7tt^��̆�2��tQ��ף&!�d��f���p�N�,����!�d�[^4 ���y�@����К&!�L�9N �"�6��
"�N�[�!�$қLN��eh�\$�h"Wl:!�DL!�>@��N1>?d���� ��)�Uc~�k��U�aL~陑�W'T� �'O@1g$Q�z�*���c�=TD*���'��r�
�1öE��NԧKND��'���z�!&rD�` ��E5d��'�l�Cn^h��9��Ӯ=�$ ��'7�{�-[�J߆R�I62c�}�'�>=�6`t�BP��\	6̌��
�'�a	���b��x�Đ�'���2�'d�C#�ߏWc���ǀ'!���'����Ak�,<�;��"�x�2�'���[�GW�q�U��.?����'�x�[��_-^�
�%�w��A���yB� I��1`O_	�e��M5�y��)A�ne�s�ѾXy��<�y��L�<YJ̰��4l���9#�[�y��6��X�o�`ArZs�J��y�ߑ2eT���R�J�����&�yR�̦i{Vs�P7J�M��,�0�y�ͪ�\AH3���Q���ѱ�G	�yBFú�q���*M�rL�s����$(�Ƙ'$��+�#��� A	 6踚�'��	�G�#F��)  d.o5X��'�� 2��U���Pz��	m�$���'��OU�6��Y*B�ٙR>�a��'D��b��������6CX���'�x�ao�vh��0f�_�HP6�q���d�3��i�a�3"_��f
L�|��	۟|D{��4
Ѧ>����� âK%F��y�^�d��Q�r���*&����P��yr/J>qw�M e/�x��E3��Q��y��Ə~��	�������5�����y"h� =�Eg
�n��mⵤ��y"��J��}�T2��A���\��y�×�@��CD�ץ7��A�#!N6�yn��#j�*6+��?"~� ��  �y�K�2�p��ˋ-��QA�,�p�<�R�W"7AT�Rp�)Znn�Cs+�P�<�J^�L'��!��t���#QT�<q���Hidp�mV�Y�xw��S�<1�^C��P�2�R�+)෭�N�<qu)��q�<0"�F�4q�Vx��FxR,Q(:���d�)�0�R��"�yB�I�-��,�ț�O=N�`Wk���y2��6
R���@T<��W6�y2�	����,��b�D�����y����"���g�6/(za#F��y��F�)�|���$C4Q:r��<�y�JЋl�Dy�g-ݳ~YD�:g����4�S�O�����IV�^��
��	%��Z	�'��� �תb	4�IN��=��T��'@V�p�N��������;�:�{��� �lI�N��L�-�5�S�]بJ�"Ol����Ӆ,���Rdb�1bp"OL9�U�G�Xg8��B�p�ȼ�"O�p��mRgT���AP�@��Ի5"O����(d>����5�6���"O��xМ �X(�`FR�CH<�pQ"O�$��;e��l1�k?�Ȼ�"O6�pC
c���ZS-F�3L�S�"O �"V$�:���J9hI�"O�,�"C�/LΘYPɘ�M-���"OLЫ%	�>�B��Q'�,﨩a"Oh��ľk02�isŎ'.�ܕa�"OH�HL�C�=��d��|�K�"O@82�* H������z�)q"O��a���%ߘ�X�I���
��g"O���wk�(]�������.�ҰA"O�1*1��p��Q3�+
=TB�B�"O�(�7�YKl|q#�E�VI�Iҥ"O轱ՄG�Q2�h�tˊ�zG~�Y��'@�'��O�����3�b��3��?K6!�>�(�6E�Ysp�(�텱 {!�Dɤ2����8U��S��"!���"0[���j�$GJl �-�!���� [���]2�Y� �[n�!�G�?J�թWi�w%�%���^"X�џ<E�4*ѧ5���s��wĠ����x�A7���V>Z���0��aO!�d�T��1C�,<�6���K�=>!�D�Bz,��!k�(~�v�hRu"!�D�Y1D��'	Z�gj��I��)
!��q)�,G�Jd.���C6(�!�S3�T�H�8D1�f�.n�!��$o��4	JM!�$C�k�!�$T3Fd�)e!��m�~�SN6[�!��nF�����h�������Nq!��D���t/�HZ��nK\GB�I�8���v���l=�K�F�0C�I�R�*�*E�� �4��펑]�C�	�3��@��	rjiC����2o C�I�D�&��V����e3֭��-��C䉰;=� C��>N��*�-�7��C��?��,���#N6�#���x۸C�ɬW�m��*�_��\�d�A)Zd�C�ɨ6~�Ո�� `�^�qeGݩW��C䉢N6� ���v���rV �q$LC�	�@ՠ̙V��2��$+��B���.�X�Q��ω$����A9xq�H������%A� 5+s�Ր(����|n �EAtI���qv����L�ٰFѣBHNLk!�[�����/��"���{)v,C烐�bc�Y�ȓ&�XS3(Gk�̰Z�	�l��ԇ�81�i�1��*mV�9��K ������K��^�����n��n��(�s'0D� ���C�sTDk �9(�Z��1n.D�죥B�-�T%x#o])$J�|�'#:D��H�.�7/�4;��'δ�R�K8D���$� Z�cP���P���&c4D��ceNڼl��Ѓ��:�p���e5D��y1�0���2�D��:A�3D��:�$���`��T�H7+���Å$�O�ʓ��S�Obp�G�¥e>��A%i^y�"OF��ѠM]V�p4�M-a�$q�"OE��Z�|
���}�Ԫs"O� (9�@jF<f�P�:T��\Ά�SA"O�Ͳ3�O'}F<����9G�&A��"OT@ۤĀ6=�h�M��O��a0F"O I�e^�Pc������-����FQ�\��Ii���QC�M	:h@�alƔ6�NB�'~ƭ���k�N�	��n6B�ɗQ�(b��m�HwJ�c�"B�ɲ���2pI$awn}@G���TB�&87�p�R)
�wN�˖��>*�fC�I-�X�I�����iXW�*zB�	�R�B���
�	��@�d�ݛrB��C(D��'Ӗ�HI�E_|�XB�$z�1���1#�ɡ0JX�a,B�ɻ?v�ɠ��V�4��y���[=�B��:Tl�L���_�@}�=��aY6t� B��
`-�iJ7�9f��9�'O>�JB�	��|@�a�=jq���7b�q�0B�$�!2RKS�	�qKY�쭘 "O�Ix�ƳGA ��l��/��e4"O���Gc�~yR�3D��K2fu�0"O�M�A��#�� �Td��8��b"O�a�C�1C�\��-�M����"O�x!�c²�NlJ����i	�"O:�9��T0$Q�c
Ppʾ2�	~�O���j'�Ӽ5��9�
OI׶��
�'}^�J2m�P�`���/U�>��
�'i��{�h�&ݔ�eB2^����'��Y�ra�XH�aQ?W)�Q"�'���Za*�Q��h$D�(S�����'	b��A�*q#
�����z	�'ʂh�Qo�)�,%ʱ�~��iA��D!ړ(�-{F�J�N��Ih�T�r�=��'�4u���c�yq*r&���'?
`��{<�4��gG�d�!	�'�@Y�또s��q�o��x��'��EC��/hx��*�!�+�d���'�,	S�L�9uo�����ā�'�
qC��8> �8s��)CO>)+O
�O���yrjV?�tlHF�2N<�Pr� ́�y2��S;z!e8D�:��ɱ�y�#\�������e0� ��G:�yr��4K=���\	���W��y���#�D��D�H5qL�}r�a�y2!A��\�J�	�c�<c�������?��I�6cX�؁LZ�N�N�Ġ�V��'�ў�>u��'�._~ �����%e�$yЄ<D�8��Њe�|3�a��A� a�8D���3E $w�=��C��
h�P�P�8D���V$�_8H����'۲��6D��P�i^�.r|)��S��\�҈6D��TeS�28�ÀFN�h�c 1D�rg^����\2/d|���.D�pD
T���ի�Gu4Hqa?D��s'��!���h�j�_�&\�"F=D���&��t�֢̟[��-��<D��c��THt���M"���`�:D�\j!͋~^�$�aaLO��P�K8D��!HPNT�L���5#Z`����2D�3SBW0)s�m+1*��F&$�0d�OΣ=E����0B��yQ ���c���0G)Q8!�D�J�A$$��V�`��J
!�dB�r�F 	ҦL7&�1	�eS�!����D  � ΋$�t�'B�0!�1T��i��ɢFՈXY�'�3!�� F1ّK�'J�̫���mKt��"O�xY�KGrd�!�L� ��XX�"O�q�󦙓&:���#&D�~���"O���%�V���I2D�^�T��"On��$̞�⭘�oލRT�hӄ"O�8�#�L���3�I�B휤�"O�u#��^/t����L=G.�$"Ol���	icF�2��"���R"ODX³.h&)C�K͇I�`���"O֝b��W��pi:]��MC�"OTЛUO>b\(��h�/SW�9��"O:HPsA�;g&(J�œCU�]Sq"O��+��,N���qT'ژIL�@T"Oz�
F�#p$��F�>P3��3�"O2DJ�E�S���$��R �|��"O0�P��%7��Y�fH�b'�v�<�s*ŗ>��qqG��D�ɶ�p�<�r�
�(J!��(�m��$Kk�<��a�8�`�� M�s&�h�<IC��>L�x$����8̣��L�<)"��8Z�!H!��� �qb�H�<�q�E�.��S
�>�H�xS�z�<1!�=}����A�:bk�P�S`�<т�d�P�C��>A��=`���Y�<������)w�F8I��x nY�<�a
�<h�:L��ʴF>D��E�X�<Y@�PVAB��d�[X�X3�Q�<)à�zx^�qAj��C�@(��
U�<�G�0:��J��۫Ժ�TF@O�<�R�[�B4v��=
a�����v�<���� �t�*��ȅz"�a��p�<9�+�KlF��� U��֭j�<a�L�,Cu���S��L� $b�\d�<ga�:��ԍ`&p�yc�f�<A�`�	^h
QeR��Hp�l c�<�Bg@J�4�:w�ȅ77|�q��Eb�<���S�-ص�&:Ir��%�y�<�$�����0"I
�
�a�Au�<�Gb��u��'�4X6�15��w�<)G�ͥWVZ,)�B��`�Y@�C}�<!!�ʍyEbE	s M�D�Pi9�%�t�<�잺3ظ��E��R��I��.�v�<�1 ��~E�|���C1�d�[�<���;rX61Z ,��8�|=��%I\�<�cˀ �L�J2'Qf����ì�T�<��X�Z�$����2FN�<���I���[P��k5�(���[L�<i�Ύ$�j1���	�
ap��HG�<����*�x���� �Ȉ�&a�{�<y��K5#�B	j�'�nL~��3�E`�<a�k	N��W�?3���� (�Z�<�T�)(D=3BٻN �(Ig��|�<���ކ��� ����e�`@�<)��?h��Q�oW�2���@y�<����"@�>�3��>7����l�~�<Q�K��h3ٸG�8>{�s�H��<�Q�3�,��B���8I��U�x�<1��A
54�q�󤝻��f��[�<1�e0uŸt����V]���2�FX�<	��Vn��S�!$v��QCLT�<���A����ՠQ:�����z�<��OM���`�ߙ&� ��N�<�fξGEz��6��]�	�6SL�<���	#K� �)T�J}��s�N]a�<� ����^RC�99u�G�w�@�C�"O9�� ��I��j�mXY�T\�"O�,����T3ʅ
����"O�PI��fSF��w��P
�"OL����ՆizZ�"�EGu�I�"ODiѣ���k�9�3�:GU���W"O�0�D
͏g�غ��t��@�"O����WPa���׊rǬY@1"O4	K���K�^3��ѵ5ɈܑA"O�͡��	={p��d��=��\Qf"OpU�tmV=s?2uz��nVQ��"O4���؉1�u�E����*c"O8P�-�T�}:�D�
�&Qq�"O������$!s$�����"O6��%<��5*gl��z�)�"OY�a�bێQ�^	e�=X�"On�i���9|xs�H-l@� �"O���Ӎ��x���K4��;,_�8q"OTL��敐H?��E��a��2s"Oʹ��g+��E��"��`��ܺ�"O�Րd�ġk�ș�����c����@"Ov��(��U�B�	E@�(���"Oh-��M�0c'i����"O�5ʕ���j%Y `'íC�T��"O��(��2à�h��'.�Y�"O�)�
���]��b$^>�t �"OH��A�\@C�: ,Z�	�"O��h�)�%>�"��ޯ{�A��"OBa"	J�z�͙-C� �"O�)���j�%c��C*0:�*u"O �#�[�}�9qaR+Wz�є"O�S�lX7j�BL�F %]���˗"Ozx�uZ15���BU�w�H��"O��_&>�p��FQ�$ߐ`�"O��)rlOq�8$`a`�V��y�A"O�!0pl���6ْ�-��-R�"O���7�M3��ঌ�#A\�Æ"Ol����fk�,�K�O�`�v"O�a�?M���!��@�g�� �"OH�j掤��Հv���a�lQ�r"O���5G6p� )��;R >̂"O8X���3j���J�tXy"7"O���'��I�����-l��`�"O<�K����ʲ��7Ơ�v"O|0!ƅ�� b T��R�"O��	u⇎XBU+Ů!ؖ`�"O�Q��/ÒR
R�: lB�$vN��"O�qpGj�0#tl��LŞD���"OJ����\�}�ڵ�M��)3�"O����&IVĬ��J_�CD|R�"O�	�ĈE�*��e	�&���$"OX��tO��"�~��]4W#r$#q"O��HD�'�~��"�ؚ#D3�"O �H�`P�:����5^a�"O8s��-J���A0j�6SE"O�q����C?�-��$ǵ�4��"O�����cb���i'�x�W"O(Uh�@���fk	%^����"Oz���D,	i���B*Ō|����"O�P�#�UX�Ԣ1�S�f��h��"Olz�Iҩ ���th�[��h�"O����\�S���7��o��z�"O��[�+]��8P���!���5"O�� �>y�JD�mE#�Ip�"O� t�����SM���O�_��2"O|%���HK��0k�	+Ͱ&"O����ҕx%�U��ߣA*б"O����ӊeu�8�ʏ:%:���"O�]��߹ +D��I�v2���"O64(E�ӣ"-��O(
�~)k�"O@�9t��: [`����Nٖ�"O��1̒���m��$��ic"OB���`��={��Q��0m�.�q"OX�C�E�r~������1�P� �"O"L!w`�p���kf�~����g"O,�&��RHB������"O L��>M�!b@,O)$��2�"O44	i�.͘ ����MؽYG"ORܸ6�˞	&�yF#��]�:X G"Ozݺ"kM�}�$R4�K�.��E*P"OX���Tc�аD�J5�x\0�"O6i#�.я4�
��֯g�>��"O.Q��[� ���>0�`d�R"O�=�6�ռ5I�X��
���"O�M����'+�ԉ��V��*Du"O~is���=���Q��1r��*b"O��5��"s�qbH�;��`"O`��V�Ǩn`(!�;`�<�g"O*�+�c >0S6��E��� ���f"O �`��� O>�`���#PE��"O�)(���*4�h�fC�3r2v!"O�Y�j��������'tt�� "O�yCU윏p��Xa��O�,|����"O��J3l��x� �&Jt]��"Op�׈����hԪF��@�У"Oޱ�sB]����8T�j�9r�"O�� �N�u�jlZ	_X��5"ON5��Nyq=z��X�Nm:�"OT�*����w��C�Ɩ&�^�`"O6�q#
?_%�;�ûzt�$�u"O�A@u&ˣ�$I��׃7�V��G"O��Q�����KR�	�|V(��"O��چ X�AB�]�^��!"Ob6f�_*�"�+ݛvUН:g�'D��MHd:h��v�ǋ5̙�'�%D��n�,'.�jӥǝ8����'D�؂T*ת)�܌���b�D����7D�̛%�\�`8����ID�rv�"�L"D�h*7ؒ)-�52��h��˄a"D��KdZ��Z5� �ܔup����>D�,�cA�~��	
�;ۚIa�h>D���b��g���烌�H���yS�:D�p0�×�ht��
v�J�+��(c�L4D�H����l�'	$��,�E3D�@�.�0!ym�Y،$(V�>D��d�d�� r'�ˊ`�� x�a=D�\����fmP<"�nK'[-|hq N/D�$��#R]!���.\�H�@:� �ɀS2��W�
�R��4Z4��C�ɬ=Ơd��ي��QQ�A��v#?y�,�'�h��B� <���A��H�ȓ7�\�s���X�a����Eu�'bў"}Z#�%���"��1ɼ��� �h�<��Ĵ#PH��G7a��� h�<i1+Q(6
5Z�nX�-cp1PT�e�<���X�sP��C���|T�d�q�e�<�����e$���o�x�x�"�|�<I釚�4�����g����aQw�<� ���g'�.�@h��_rx2Т�]�PF{��),�R9 g@0t�����ƳK�!��@�/�(
6��n����j��h�!�[�:��Ӵ
K6A`ⴸt*ǎg�!��ћ2��Z�'��+,���(C6O�!�ć�a��:2H�C?�T���[�!��ěs�p@jR ��{��ߟy�!�E�Q���s�ۊ�5!!��.8!��@�gn2�i���Ij�����<!�"�~�*g*� �`qQ\��'Pa|���7��xs�-��u�d�C� ��y2
V)k2`�Fɜj����3���y2K��7Q��&C�cU���aS-�y�-��S6�Q -|`�ђ����y���;i��ڷ�H!Z7F� rlɩ�y�)\j��q�2O�Rja��NJ�y�$	�$� 3`�%:��� ���HO2�=�ON�X��04�}���_6�0�'$})�M�	|��HaE[��l�ANL�<9�#̀VhppS��e.�jRi�KX�P����5$���OL�n�nE��IO�H,���>Q��U(aD���ưR����
W,�',��'�I��O�Ĥ �ԪR�\t� KX�@j�(:
�'�T@�WC�X��8�i��^A��0����X������y� ��E�~��e�M�*�����,�2�p?��O�(	2�A.TdT�`f̖r�&��"O�`1C��XP�u��eҽlF����'��a+��YF��_:��n_.�N	�O���d�'Ĵ8��������$	CE�y�቎Ejl(�cO0i��zVbɖp�.C�	,;������l����nG�)vHB�	�
l=P�'d�d!�O��:B�	V����@^8�1K�aɆ,� "?I��)��@t�5�p��+`�Ԉ*7�A���E{ʟ�(��S�Xd�T�?k(��� _��F{��)S(`M�p��Gqv���E/
��ay�E�*�qOj����y����5��0�v����$|O��C���r�h��c�p��"O����,�N,��u��������"O����-v�4T�3����!�6�i?��E�)nZk�(m�̋�Y}��=X�ٚz�hC��1Yæ���!˾p�R%�g�[s�bC�ɇ6�R�+7�>U�N�P�X�Ɣ���.}⏔���m�:z��qP�dO��y⇙'�8��ѽB iFN7���򤔻���O����� �����sL˿f�q�'�Yr��V�x�(-�4j["���J�4l>���3�~FxR��:�R|�$,ۮJ.� �c���Oz�E��@�JĀp���U����/�b�,��p?V�8��cdc�7[�8�VHX}��7�S�D�|�@��872�5JSVg��kY+�HO����).��|�A��0�FA#aKߗ9�<����Oq�2��<��J^�b@�,Y�l��|c
h�UaCK����>�ʟ�Tlr��p/��;~��#��C�<��o29��u��#�dy؈3�z��0�'KL�ڐ��4o�m�J�y�x5j�'3�+2��,�N���! %���'�PW�� 8�J|JIۋO��y��'t�As�D�3t\x�4읊LX 	�'sў"~R�CZ�2H@s�$��s�
$�c�c�<���	tJ�X�4��M
�M�b�<���ȜxV��7g��e���I_�<4$�"��aڕ뎞\�V1AHI]ܓ�hO�Od���Ί�k��)ycC�J�v��O�O0��� D���>N"��9�Ȝ�B����Q��SX�t1� ��2�"�rD΅-�l`v�8�O�OP��eA��05X!&ˣ!5��Z�"O`�2�9ZNb5"�D*c�0e�x���_�Km��	�d�@A����d	O!�DG���� -�Y��y��M��9L!���9�4�����"e�|(�E��_Q�p��ɚO�"TyR����=�""�8�f�Є�I,
��l�$>bq*��W){�rB�Ij��i��W�Hd9���fB�ɚ�
q��I"W,���������$7�S�O�t�n�F:.<�oZX�i��"O"X!Tm��t�X�%��4{�� "O��i���N8��gL�bT:�*v"O4�g�>������s:dx�w"Oz��!/�R�8Y��V� ۣ�$]<���D�	;R֘I���)G�@y��@ E_��oӸ%��M΋;?���f'��,lHrS�HD{���Ҡ`��lW����$�/>�=�ȓ>��=��h\�#l|1�&Շz�x��ȓ-��i�'ƪ|ڴ�Ч&��\����o�y^���͹jI��(��ĭl���ȓ�>��V�1J:�y �W'� �ȓ�
aa5�	\4aP'�Y&t�zцȓ\r<90n^,'��) Dg@�\���>	����D�c ���nL��R��F���y��B𰴊e�Ҧ"F �ӑe�/�y���.��8	�a��l����V�$��>��Oh�n;+P80�ҫ�n#p�e"OUr�IN*ba�mJ�
ǎ8��2C�u���?���wRF=�N� :ؤR#b�9}�M��'� ���e�4t�f,h�D�@�۴⑞"~nZ�l�V(���N;5QD,�'�1C�	�)�%�&�Y�lt`�uG�,��	:�MC�1�`٫�f)m�(I+3�ӆ���'�x��)�� B�A!A�Y>�� s�_�(B��&n�=A��[�]�)�#��_��7=��I s�T��~&��ƈ*]�1�E ���.<Oң=��F�+S*�H�F�,/P�I6�p}��'��\��".`(��eH4��Q�
�'�PB��]����T�J
�'

[q*�2��e�E���J�'2"�<`���$�t����!Iq�<�S��ؐE�T+�Yf�,7Ȅi�<��#�%e A񭌒&�`�`!G�K�<�G,P"��f �/r��ìLF�<�#
� p���Gc	�˜ap�=D�TC&��(/�aT�$�R��9D��9&��N{d��qvPT���:D�z��6Y�$��ǮG�6p���:D�T2g?i�ГЅ��D`rC6j7D��Ç�,$E���(�'$~��e8D��a���-JM��'�@9!TΩ���2D�����ϊo2@���^7Y���9v�1D�@A�� 2l�lD�p� de!+0D�H�eB3�b����[?�BA`�,D� �A�öU��q�aM� u9Ґ�#=D�6$�l5�T�s� ?$h����O;D����+,/^,��Q.ۼ3� 8D���sh��x��]�!�3��=��+D�H(V�O�)�19�Gf�:�'D���" 'z�8�%��K���#N&D�ܘ� 
�/kl�pf�G�UJ�� #D�d�C�T�L�hR���g�$���"D�� ���>R�¦��(j��Qc"O8=�0k�������s?�"OF���h��B''ޔa  ��B"O�ݫ���:*	��)W�.hܔ)�"O���FL�*BL��8��@�S�n�I�"O���2��(G�l���p��`�G"O��O�ۦ�2#H^�3��]�P"O�	�̱%�zL� ���%̶ňU"O S����lB���VGODaJ��E"O�tk`�.U��#�\�e��"O��6��+5f9;YHDaGN_*b!�$@�n��h&���W�2Yqb͇�g!�DɏWQ0��o��|{�˅1,�!�䖤.�ERЩ��@�ke�!C�!�T86ňT�����Bm
�!��?V���g��>ko�����<t	!�dTl��9�N��pg���-�8{�!�ӍG�i�ˀ,TO"@!����}�!�B�B�y�9Jd��+f'�!!�D�7>扺��(4QN,(�`ٛ`�!�<V?��р�U�n^T��F���i:!�$R9-�l�:NU*<[w�02!�Ď/	\2��:4�2�̑�E0�$ĢT�6��Q�R�4��"�#O���F'U+3H�����7��}�'L"D�,Z F��\�2���) \F���l&D�Ĺf��bQ��� bV�h�g;D�H��%Jml0���oT6��`b-D�\g�ޡg�`��@l�
kL�̣��-D�ly�>?#d�yV�wg*�(B�*D�$�&�@�,��D[Q��[:�(�F?D�H��'�1RcV���L�>e����!D�(�Rd�N�"�a��cHp�<�`�T�@���(­Z�4T��O�p�<!��r�>���Ӎ4}r��t�<IG���c"4m 1�
	Z��s�nOH�<�g�5Ȭ]�1O�l<�����F�<y�/�6aƴ�@KI�^�Hl��A�<!�5Y�{�f��uC�hJY�<�5'V8����hM:��D�AfZ�<�!�X E\L��/��Uv��D7D���D�B�\9�1��A>1��a�E4D�`����;Ҋ�G/KI���� �>D���Ơ�<���2���1y"�jfM8D�� ⅊�B�2 �$cǡ,'�D�-9D��c%�5^Hz��ӕ3@43M(D�D�cӜV��9��2�x8PJ)D�к�I53?���R#�:@�X$"R�)D�L"�� E�PŘP.ݭo+��#D�����+V@����)/����4!D���"��j/\ +g�ɸ�����!D�$�D�^>c�薬���F?D�8;w	�"2��-)��/*r��rǋ D�d�� �8j&<4��F_6\j�H<D��zm�9HNU[G�a�Z�4k1D���SB�+Y���(��1# ���//D�P*����n�hgEB<H�"�1D��"'W#8�	9EGݽpG�1�4�:D���dM,s�HU��/�^4��vM"D�� e�Ν~.�i*�CGB^j�:u�<D��I�h�9)F��#�Z�v�"u�$D��d�#�l�de׮(�p�e#D��`��
�]�����4�qh!D� *1O�{x ˴�G/ $�S�!D����G	V@r3�}���kV+>D�� Dp!�Ȭǎ��CC�=Plqp�"O� q����}����&]��x7"OL CT��3#���n�;c�\�"OL�k5�ܕ�DlB� W�(�P"O�� 'F0n�`���X�EI@=�"O\8���M�a�@�^JAX�"O$Tqt�\g�]�ץ�, ,8L�"O"`�Mŵ# İ�0��yp�/�y�&\��<��Ϡ޼��e�7�yb�ץ	��H��8�b�J��y��OI�}Q�	E�9>�K���y"bȮŊQ��&(��bӧ��y��ݲ)�"|S�m�+.a�d�3@߈�yBH�5T���!(��49�&���y���[S.5Rt�L/_�,D��"�&�y<X�ִ�2�	�{ְc��y���	R��3%��1z	�a�E)�yH(��(a�Y�X�Z}�D��y�lJ�:!x� ��Ҥ�Xe���@��>��C��'���Թs���
�N��`�Y��� kS!��X�9tF�K�@��k���4�T�EZQ��I�E<;pB�G���O���}S�	0Q)�
�y�ό3g�	7@U�r�~������|&��sP��O?�I�q��,�rϞ5������Z�y�&C�I�ik>�cፊ e�qb�7�2��9ظ ��&4��z2��<^{&�ӳL�U�QB�A��0>!�h�	h�#�$�^���j#��C�x��3�͏y���ȓ|:tHȓ�Cf0@`S�l�BGx�힉g�j�����_�O"�=�SeK)j'`��@��P����'�4��j�p�@�I
l�
���/g�� ��I��	!Tӧ����Y�t�Z��AΓ ��p5�Mi����٣u�2�����	2�i0�	� ��}�l�@���c��
��H<RAG<H	b�4�l�
ml��.VM!#�g^|��SE]x)�B�� x6�C�,y��P'��p���(�����:����Etx�!���7(x�m�^�µI2D�O,ij�"W�-ܸѥ��&A�	�d�&���7L��2n�$Y(b�aW^.u]*i��N� Ȍ��bw������|��5ۂO���.�Ac�:�>��'(_�,�$��*2>�1�#풚���ς;�(5ۡc^ӦU�;7[��I��׹J��]┏A�V�B���	>�V�2���ge��k5�3E����ĉDp&��pe��ꥇ�!F��X!xh�C	�rg���gY#@��d�L~�%�C�EjU P�T��S�ʺ�(O�������y
���V�@ș�/ʻ���B�5��s��?O��s	ʣC! 1k��A?��Փ� �>��j,�Q������ J�K������7M +� i� �B#���qL߿x��,��� ��<}��4�"M��>udUaӎ�('��3ʞ8������W0�Ɯb
�!ޜ,3�J�;~�`�U)�6%�>dC"-ȱV��d�#%_��E¯B4#،k%�M<u�`�5)��#�*L�;=Jx��۪�.��sI��f����	??�d;�n	8Mv��ve��q"̨��O���rt�jP�p[wa\�(H�
^*AK<@�&�I�t:��� �C�S��Z��'oN=t<�+�.9�4!�?�eG�$!\�(e��
~�H��֌Xz�yR�OB���t�ʦN9:Q�G�J)N�ȨI���K��6�'(�"D	�	�1��3�p��	��X����]I�VuP�J9�U+2򤰁��H�\m  �9���>	�WE�tt�|�@� ��ASGBυ�r�)�+6#�@��YtX���&�A(�$�ȳK��-#R�˂ɔl'�j��C�:�J��"�'�H����0����Ś/&V��'��D�d�?3J��;�@0�l�ߓB:�@��O�O��6��0j��B�ĂN�$�)��Գ��F,6H ��
�4w\!���>Q��4&�<5DI�3�]1q��D����'���"�'͆}b�F���+�nY�V�iH��C�͊9P	�J�����q��'���	I�uRF.O���� SkN8\ވ�D�1}�s���E�7��Z�:^?����K�& Ψ1���0?	�″c�@��6�/S׾�ʐ���<16��>hv��:�yZw��/,���E4?ygc��V}�]R��p�t�w8�xC��S�:��d�,�D8h"��6��ɡ�W�U��'n�=h㣃.h�����SD0���f2Q���8�K�!�d�#$1�	��eB��8Dn�+o��4JJ>1d�ߪm����'Z`�LO 44
�z��ˣP��s�'<D�CQ� �2�l8: ��;�6�#��;'T��)� �����sP�y��T�|�<�8�"O|��SC�I��uS�Z4;x�=�0"O8 �!�<v�ԙ�N�4e`*���"O�U;��Ҋ Hy���ʗ	�%�%O��ӫ_�C�:Tp�P�qϪh���1��1��sfa�`�a_x0C0�R9��I�41�q�%@F�	'tX��S�P�R�Z�Ɵ�B䉒NyRxZ�	G�d�$M�B֖Q�(ʓ��=�tZ_@)���3�'oLɈ��l&2H�$T+lM����3�XX
�S"�Zl�ԭF��@8sE%#>��E�I�bPҐ��r�3�����=z�@�X$��5,��-+���DE;!^�˦M�~IҊ�-QN��b�ĳo�����O�#�z��D�./��ւ�j5��!h�6�ў��g��d¢���[�t}Lz���|2�e��u�\�����u����o�<ck�4#��q�۸h*�ӕ�	�&Ă3:�l['B�'z���TF��H�k̓iP4�p��()�6nW�K�!�DJV�4i�瀨#4#�,h>�d��M �B@��1F���Vӟ����P�>&��1ǜ�	������|�>Fz$CT�+�ҕA�O1/֝y�Q���\�a�� !����=I!�6=��8%�7���qd�y�'EL���58��x�"�1Թ�!�D9�R'���}�DP�����[���ѢEp�<AcnZ�'D�s�M^�U�4�xSH�/4䬩+��U>2��9e��1�p�z3�;���[4fEą�M��@N
�y2A7K�
��d#̎���M�H�\�N��8G^�Qb�	�K7�<��O�1�r�	�n<TM���T�\��p>1 �SvK�|8R�Za~^�!gֈ|,32�_�FQ��p&gTw/p�p���q���2#�K;{%~|1�O�5U'ԥȑ#.�;�
S)˺x-lTm@n�^�{�C������+T��3q�R�#6­c��X�<���']�^���)�5P�r@���e��뗪s0Y'��\���w�Ͷ�H�k,؛D8�5"Rj\
pgP$ ̛N�!��Cz��!�C��"�h�eF+z����G�=�i
�Ҋe]v���]>�DxrMۛI i��/܍R~�����?�e�75=
L����V������
N�lB�j �*|��C�N�!�p>�$�A%�|��FQr��X��^Z�'d�2�EC�6� ��ď�>��� 
@R, &b��6nH� ��lF!�T�$��H����.]�$�/֮L��	�Z�xyҌ�Z�4���`���A&��Mn�!@��P�^$�C�L�"�Z;Tm+��O�c�2E�T�!}B�E%��i�}&���qONH�`��s�X��h3@�<4��9q(�$t��H�Œ8푦� ��L�Q�'K��;i{<�a�� \�?��y��'���ⶦM�{G�<Zr�,?h��'[F����	\����a�% �4I�'�,�;���1��m�p��H*�%��'������W�%:�i�SP^��'��	{Ǯ�j�[O�9��I�'��r�%!v2u)��+�'��8��`�@��V�M�m��X�	�'���u��z�l�bG͔r�(	��'^��/Ub(@��H�(>� �#�'��=���� ?l����+����'���+�#LhK�*��E�#�����'��J �P���tR��<+���@�')`d�R�<#Q���&�\�"
�'wv�G-��0����ˌ�\R�'?@]P� ��4�ӭ�7} �`�'�l���a� `T)�b «h!	��'���H�G�#X�v�����P���'e�p�t��n�zI{�#ȴU��A@�'H�0��ȍ�W����A�Q�BĲ���'*sd�^62Z��9qHL�d]��'hՋů�FH���G��R���'��D�I�Qr��`�*�����'Ƅ����[� �ndZS,ĳ
����� �����#<\p��@�u8���"OZI��nb����:7N��&"O}7珿���31�,A�u)W"O�庄h�YL���Q�"�*�"O�ę&F�%���P�@5�$��$"O`�Wd�!$�P���t��.�!�$J(3�6��1�L:u�Փ��O�f>!�D��l�ro۾:�Y��ˏ:=$!�$K"Q���O�;��GlƿN&!�d�Q����e��/r� -����!�<zF��c˚7����gMزtx!�:m1�i�5o�r��=��]�~!�,&����WY��}Q���`!�$Ȫ4ռ�`��Z?8Z��;�LPo!�$�:`

	�ŌG�\8mp��%>A!�So�,�[���:J4�Qʊ�E�!�DEi�m��B0z'�%"ND�!�@�o������8���Sb��$x!�d�6pn��Ye�:�v����pT!����� ��և�"5=.!I5g̓RT!�J�o�!�&�B�MJ�	�0_!��B(L�%j�BP�l� '�$TO!�Θ`5�H����W��]@H˘ �!�H�b�84)S)~�%ch�r���b�<��F�=�Fx�v&�v�9`�	F_�<I5 j���3�X=欜�Ө�U�<q��=�~��e�κU�m�&��V�<i���M 	� L��c��#!�Pi�<��S���AT�W>1��WD�'�!���
f��:�����I�����!�$��}u"�R��E�a T�"�a �Bj!��ȑ�(����٤~�0X��U�^R!��ʐ�P��,�:����P��M�!�D�V���狑Cu`D����t�!�P)�p�K�#ŧLiP�R�R<D!�D	�g�X��KR 5�s�E�|!�d�?�����ꎜOj��@IQ/|!�D�7��ٱf�ED^p�A(�E!�$�_�¬fƜ�"���F�n�!�DS�������!� !���з:�!�dL3}����\ah�`v�Ѫ!��Ķ	$>$���U�a���ƍJo!�0`0!�7lX!S~��Gf�0zS!�d�)���o�r8F�ce�Ӳy�!�$�]����Ҷ?@�E*��1�!��;tѬ�@��իn\1研�6�!�$ǹ7���w�	%g�TLZ����b�!��Z�p{g�)7�Y0m���!���8=�´q�Q'�I�e픰M�!��(:$-�4�6 �R��3!��E�j�hc�	�l�xx��<4�!�D�3*���rg�0�B��攫�!�dQ3Z+h �MՃ_��D"uD�(�!�dM�v�^U2gO��M�
����Y�:�!���<v>�y'�>�v0�#"�-�!�Y/
^"X8F	U/i.����ߍ.B!�$_lK=#$�,�F�����n!�ĀHK*�"��A)T����ԋ��g!��?}�iHGoO?C�rMY�K'!�DO8����L�-E�,Yq_)@�!�I�37��!cΏ� `�}�t䂶x�!�D�z�L����,niժ�j�"G!��S�h����ɼw�iC��j>!�dÂ 찤��'F(Lx��Z�FU�)!�� ��s�I�%pV�!6��RSj��#"O�m{��=Om��5#WiH�8�C"O�h	Ջ���mGB[:,I��I"Op�X6�uyL�J�̡ E���'�����H�ݪ�Reh_��Q�'��:�+96Pl��.�7Gd���'6���U��L�ҩɵ!B8�(%r�'�~�4EA�a"��E��b)^���'*�L�ү�4I����X�[��%y�'fiz4j�wi�l�1�2f��M`
�'(�3�N�5-V�#6(Y(T��s
�'<���֊��\ ba�jzԠl[
�'/~Y��l�.LW��a�E�2|ZN)	
�'����ȝB��Q�-�<ga�1��'�l��Ԅ̋!���Q�!N�Y#�L9�'�i�� V	x���:��[�MH�'-�dZv��	[�*�b$+Ůl�B=��'@�X�s�Z>-`E�f���$��'�0��3GJ�Z��yv��x�.�K�'�� �˟w����(�t���C�'D8�:ǀ�Iz0�ktIY�E

�'�⠃v
�	J���ɣW#�r1	�'��ͫDB�/87x2�H�H|���t-���O�pa�K�I0�0B&<d�C"O�� �5aR<k�Cۣp��IT��S��u�O� �qc ��cak�q�
���'�H%��J��/|`��:�n��T��;���ۡ��w��s��&�:�H!�D5`]�(���-D��bf�L K�6P0��Bx���v���i��>�	��'Z2��d����+'�Z�BC"��`Ќ<z��A�.�Rp*t�M)�Zm!�8:Th����\�<1� ��=���
"5׬]���A�'r�k�. 3t|��E�D̂!b�,��� 2`�{�D�<�y2U�� :�e�Kˬ񨲆P0q�Z髷.	�6]LT�O?�ɴ>< @V��j0���I�r���$Z�?8�`��ԄJ�R��Dӝ$�z�� j�G^JE�ThT+D&�i��x�P�W(�H�<����\�v�9�.4��F�J�'̼���c� �z�)�d�qZ��ǌ�%�A�͘9�D�cw�:�s��d@G���<���S�L@�I�r�P�# ��)���w�ʌ��!?8�Qj�R	�'@z8h@��0�88ڦO������a�G\��Z��lX���	�f�
Ȉ���!��8���~��*���*�z������gᚫd���2�� ��4�A ���Mc�w}h)�E��n�� C��,AF)I�Uܸ!���\FrU����h/�!���=�M(Ḑ<� �&b��>�����cQF�t�sO�k(�9�3�+�I��Q倀Y�*��:�h :VB۵Xۺ�<��m��T96��<�pj�ڷ[߾�ӣd���92���#�Ғ}ߐ 99J�c�P.8"9�wM�|Fy�.Q�hn�a2A���0L�$���H�q�F�% �kc�N1n�x������'i�n��d��k]�9�.�%�U�#�՜`�ؔ:�E�u��(��?�O�eb�cJ�5�������(��A�Y�7�0X ���M���p�C�L�}"K 4���`	��2ܻ�4�|��(�>J��E�4��ja@�� �'��5�fFU* `����.&b��6BC�m��M�`%�i�&�ZBF[h(.Tæ��Z�1Ȇ�ү%e�!���4o��Oe,���H� f�y�!�<%e�Y�u��L>(�zqұ)��B�ڶ��|@�ԃB�v>M��E�Y��x(ƚ�oQ�:��ULV��ݴ��L����@����O-!�E�D��}�1��?l^��S*gLBt�Μ����Ӷ�λ=�91�)��R��+2��p�v<;2�\�,�f[�S��A8��G2!1*����ג��?F�T�sE���@˄k�81�d�T��TQ���I��:�I<C�X��E���	��}���0<�2a���C46��dSLP t��S�M�P�LV����F�4�X����p�/I-p�j(�D�Nׄ��O�c?M�p�l���r�# �R�2��$]̲���&|؎��H*���#�T�E�
G6�ȉ�>��k��t�>�O.�i.���^�7�wꐑ����e��	��o�D%�禕Av�$W�)S���Hw>�p���;;,pe�\��a~�"Z�O�)�m��9q��K��6�y�$� �Yo2�i��ƈ�<v�-�'�@��3�K!_���
J�lp��(�z���r�L��M�5/_��sa�O�Y
2,��K,}�V�y�xh���X>� ^�gH\.E��pF	)�~i�E"O�����X$:�b�e�#v�z�b C����v�r�Jp��x�D�c�vM��F��l%��RH��xb��'M�|m��A����}�f*Y�u�4��f؟H���	9�9��DV'x��(D�H��G�^���s	�j&����'D�(�L��R�D!g���I�(��I(D���&Y-mk�hJA��FҤ��E*O��L�!�&��s�Pu�a�P��y"���Zr<�#gU��&�
�*^�y���Q鮘�
^���2d>�y�߃%�a�K>�"�/�y���JRԑKT� �R�ċٴ�y��0s�1�j�-�L)h��8�y�D"Ѡ��N�7.C��GZ:�yBLظ*�
�Z�扚TƶU�2I ��y�
R����
Q��<�y[��Y��hO|��tb�!�H���Z7��7]��s���:H��3"O2���X������	�:|����i����S�Y:\ɧ���&#�4�`��� ��g����Ί�yr�ųj�B��f�\�z�J
�~��5p�&�҆�b�� �'M*c�0]���"I��P�"�O y�� � ��Y,ÚA�1A��W�8��q#d��%�yb��i��M���N�KM0�	M�(O��8�(�o��Y���N"��h�@a�8;\�{��{	��'��-�r��ec\Mr«�
QZ��橝#-���;^`XbJ�"~�	Y���CЏ�tے]�6�҈�4B�h�yp�FϟSbP	��*U�{���	�7}�rC
�$T�az����E����J�<�l�%�\7�p>Q�%��v�� .��p���*z9�<���
Oi�C�	�qn\{�F$���@%F�e�v�<Q�̗!v`DS�#&§5!�|��e�Ei����\�7�
Y�� Y����!v�ڈ���ܓ;8��o`3���n[�)��ѡ�'��p��{����&vHң�?D� Zc��b��ıE��[�q1�<3��1T��dJ�Ǻɧ֜J�a	 ��.�!�D�4�8��1�^�c
��Ԃь@�!�D���|��/���$������!�D� /V�9��7�XIzҬ�C�!�DA�:�~Y�҅�66�} ���=&!��>��\�3ȕ v�b���'�-l%!�D�+f�̳0B�.[�`� ��7s!�$$U�Z̀pN.|��\HK\'7U!�Y%�l�s��`�TG^!�dQ�E=����c�Uj�L04��3bY!�� �v&�9 )ԑ%jH��KL!��Ã=� �X��� IJd%��I�C�!���"*ry��d_�o��\��G�2�!�Ă�*���Q�‫E����`��K�!�d�[�(�c& �>k��S gQ��!�_'TT�*0%�E:H���l!�dW[���0r����3!�D�:)ve�fe�r#"����R!��<f��J��DJ� ㊙ZF!�$8?�����ǃ�4�=bqiA�yM!��ש*�0E����+6���*.L�!��3*�z�s��
O�`Q�&i��j�!�Dܓm�X!�Gfʿm���Q.L6T!�H�"ttu�t�k�N�[�-�/Ge!��ƌ,Ø}b$i%����+�)X�!�ă d�P�v����j�)�/d,!�䜥L �S���!>�dep����,!�D�Ζ��A�X%{�����6}!��9)uFt㦅J�xQjtAB����!�� �}��c��B!w���L5j]�"Ob]!�m��{��U�N�	*��Y�"O�}c�"�;{v����7?s���S"O���)�>|�e!�lF	��""O�᫡�T�N�>!�RkBl�z�b"O��9�.�?m��YJ�m�p���S"Oza� ��: �����`�X9�""O(��DE��Ԍ#f-��w"O6��U� bY�T�Jɸ0�1�P"OH�s�ǓC�J-�ȗ��t�;"O��p&J1D������A:M��ڧ"Ox�P�bޠI��yP�ΥzB��+�"Obچ�_�@��$s�iHiB���"O��F�^$*虒�J�+d�ar"O�8�
� �졑VJ@,;���b"O@��@�RG.AAR)� \��(�"O�p2Th�$���cÆƎ;Є��f"OR4k���*��u[5��ո�R�"O.��I��0��pn	�t��q�"O`��e�?7 >	��\le��"O~iEJH�
AB��tM3@��hG"O�My�I��|�����#z�,��"O��H���9M�P� �P|`�"Oj���$Gal0�[u��~.B��5"O�@���#F�dM� K� N��r�"OVye�U(�y�!
2��c"O°yw�ԏE�h�0�TEP�"Oȝ2�#K�O=$$�Gi��A���S�"O
y���(�Iw�O� E`��d"O8���@��5e���T(�z6T%�e"O֐�s��D5<��r�Χ(Q��<O�T8�#��-x�@�aѦX�ȬɃ�I >C��k�H�A(��8�bC�ɛS3�� %)$> 
�pQ��:8bC�I�g}�]���������+�N<C�I�T0�0��0vv�r�l�92VC䉤ꦴ�g'ԎGd�B�V5q<JC�I�s�q�j���Qb��6\Yp�O�Uj��!�)�1{X��[��_��U��`A8;l��~Dp�z���)�-/��1؁gI�;�P��ÎI�E��*[y�O>�Br��(�M�f��K�l��g#�@	�����h�<i�'�nD
5�Ou
��*W3<��(I�����xD�@��~Be	ڢ��>9�˧<��e*�$_8xh$*�� (R�+��'N�����""a�ڑ="N�?�qb  ��Ppq��"�,i�c(��R���M��*�"����M�F�O�z�S�^�Q/>�b���,@زĈǹe��1��ì�M��%�[�����O
`�E�Y�����Tk��ض A�[�h����`���C�&�	�0|��Iŷ
y�����-W_:��� E�m�Vxϓo�j�z�ӿ9R���?�}���6��A��5���T,�Cy&]�lG�8��o1<a����y$���X�����y�gx��I<�2��B�SV�H�Ӥ��}�T�#2�	HA�-�$�ѸM��O����ӲP�&L`��V@��g��~�v(EN�D��Z��.��M׀�+�n�Z�($�&xAt�O~��AM�$>c��A4E�?`���&)ys�h>D�H)E�)j�����;o7��v)0D��
�GF�4Ȳd9eG�#��	 O)D�(���
}�B��s۫]�Ze�Rd(D��Y�(���!�s<95H'D��ï�6:A䠓��E4k� ��#D�$��M�~��"��c����`"D�̭<\v�9��#&�H�I3떄�yA��f��%,%Cp��2%��yr�X���Ae�&^�m*����y��p�z�as��68uq�ٶ�yRf�"{ܩs�o�����h��'�y� C&D�=P�	��������y
� 87�P�9ꤓ�մ(�`+�"O@A��j��r�8�B�.U�Mk�"O\�$��:��2�K�NI�#$"OLq����g�bY)D�?HG��8�"O6��v`L-I�����6�ջ�"Oj��΁8?�բ���}�@I��y�!Bޤh����R<�}S�c���y��x��(�!�x�
`�g�yb᛽T���r�� %t�&N^
�yB�Q�_^ ��J��"�|MhѧS��y�\�o}���U�/J�L���y�-�R��`Z�<(p��w��yң�8a���z��D�+���q"��yҎN�(�FΚq�YC'�ݶ�y���7���F}�d#'�ԍ�y�G�^Pư�S�CA(�D���yrJ�
V.����
�2k~>�uF���y҈ �]*г��(Rz����V4�yB�P�EKd��$#I&�<
�M��y��A� U"�a��C�r���H�DN��y2g�]��#��(a��I ���6�y2��_ J�HOK�R��5+Q`��y2�`r���阸L���V��	�yB�(]{���dZ,q�F������y2BA8򰤲sF�n�l`5"� �y� �v8X��m�:R8���ǳ�yb�	��ᙖ&/	d5 ���yR��PQ8���Ό�2�Hِp)���yr˂�4��5�fa<'���Ҍ���y��O�x�Sag/$��� rKK��y��B>�Qc"�O�-��Q��-�ybh]�4ȸ �tg��{34���o���y���M��I���2MJ!$�8�y�ʫq�ƉC��NE8taiD��yRNK[��e�
u!]X��ٲ�y�����x�N��p�X,8%��&�y�(��kvp�*Ɇgb�$Y�+B��y��ӊAb%*�n�-���0�ω�y�Y�@
�E��(I<-/����O�yL�'b�����p���#���y�;�y16cI�`��������y��
|	$0�`I�6G�X�W��9�y���.MQ5Zj�FU�
ǥ���yb��T���`gV��y1I��y��q�R="V	[����)�y"mH�`�p�@ͮ�ȴC��D�y.R<tnА�*�2Ĉ։�9�yBi�I��HH�� �n�@�B��yBd�+JR�<�% S ��D#�����yB��jer�(nא���&�%�yrL�:9�~�c��&��ѨVV��y"��-��
��$m}腪*B�y���9*-�E{�҆fm"�5cK��y�C�`����Lذ��%]��y��\�w��q�Փwo��p7�6�yb- ]�^�6-��aD*(X'ŕ�yn^��1��@�"V�p�(0 ]9�y�g��ICK������ ���y���)��Q�:
i�y�gDC�y"��z���"�n4ɘ��C0�yr���G��ј�ぞ�MS�EN��y�D�R��1��&�+t�\|����y��B<�hZ�.�s֊�FHA��y�+KVš"��3l�`
��.�y
� ���E���CA����.?�@ A�"On%�����uՒ8Xd��<s�ޥQB"Oh�@�lY�z��`N;K. �Ф"O|4��!9�jX�sn�y� ��Q"O��xG�T����r̀7:�S�"O��Z���s#a+|1V���"O�ѨB!��B��[������"Or��e���T���6+����&"O����Z,Tؐ&��EwT��"Oȑ�Ń�4=M\��N��}�^9aV"O*�*��$l�D��uz)r"O��Ť�>:��!5�W�Ol޸2�"O4c4fD��$LC%=h�� &"On�ЩR�7`-V�=U�y# "O�p��ۃRw��KU�L}����B"OꌑŃ�F��# ���5C""O�S��	�D�a*\_넍�"O�;0a�9 -�͛"#@�.H�7"O�A���-c������	w)<��"O�i4��*p��UX��lG4�҇"O�̹Al;p8�B�Q�u4\�Y�"O�I� ��)Wfd93�S-  �"O8��L�O�2LF`�;x���)�"O�|�GGGJTp�ˆe��i�"O�ZF��1Py�xZ�*�/t��"O@�r/̾?<��`jF�}j�!S"O0��aN�<N��
�N�Dsl"O4�q1��0$[�<Y�Ρμu2�"OP��q�@� �B��W皬�DY�"O�}�E�FS�IƸQ�fE�C"Op���*1Qκx:B��-d4�"O��q�I"��@K�Lϡ$�P���"O����H�H�`%g��J�8re"Of=x�AF�$9�Ez�c���@	)�"O¥[��Ɛ �0%e$݋U�V1jW"O��:��j�x�!���:xZ���"O���2DՋc��x�A�><t�x 2"OZ� #%ύPk��)����v�6��P"Oi�(X�"�Ћ`J�  ���*O�@�Q�,$�iHt�y��}�
�'���lE(/�B�Uj�T�
�'"q�F��{̨��,W�u�x��
�'�B�x��<l��hr ��ef��
�']��s�����К�'V��
�'悵(�Y��$�3��%R��!�	�'�	h���Dz42èZ�H�ʑ�'�}����J�s#��)ZV�
�'d�dC'
Z�q���B�J�)vЅ1�'��]��Ĳ%*��ʵJ-R���'y@@��iB ���	q�k�'$҅:�%�=v�N�q2��:
�'n�@y�eI1�й�W��8i���
�'�fͩ���i��LC7	�9��,i
�'d��"P�G�s���+G�9|UT�+�'�Z��⣞�2�<i�Q�^�r���
�'wZ�S��F-_[��X@��,��B�'t-��� P5�B�D&fJ8�(�'�5�a�0X,@�Ы�XA����'e�1�&�׀���I�T���I�'�fM�q¨w5h91VdF�Z�j�'���[(Nϔ�+W��H:�((=D�t����?�4�T嗩&���O:D���D�F%ִ�sKS�&�h��f6D�� �/��HeE.#���-3D�� 2�y�D�) �X� !�S D�*�ye"O������P���T
�b�teA""O*��%�{�dA�H��H��I��"O��f���|�BHD#��)�d"O�a�"jF�rP��Aա�*��2"O�h��K�A��B#� ���"O��pdD��`4�7X�L�0�4"O��ꏱ`焄Ѡ`_# R�(c�"O��:cU��(�#���e�&���"O�d�g��t
���6��?��@�"O�$�3�� i��8j#(T�Y攰�"Ov���k�|��p��N��$
"OP�5��# hm�Fh�/��%"O�EsC ��~+�Ũv��$g��`"O|m�'��?q��А�R4f�,Q"O�𡰄�yVp"6h]	S��h�"O MC�jD����ƈ����&"O��;��vsΜ��V,} �i�"O2(�$@A	+�1��Az���"O�%`1l(����V �m�����"Od�8X���0���@�h٫4"O|��͔=g��8���O1aK"O�lIJZ
-���w��p��&"O���T��tv�	b�b�FFEK�"Oޱ��
��P�툵��" "OD�����,�����4T��T��"O@{"��6�.ɢ��~,-��"Ot}[��ت<�����$j.�`"O���5��Gh� #֢Y�c�+"_�<����Oe��h�oB�uA��q��[�<ф�H&l ���D�M;W�,�p��@M�<1�*k�&�r�j5ID��(�cGK�<�a�+�n=��
1�ӗ���<���x�4�:�۳u�*�s�I�g�<9@�F�V�`Q1�-�~�;��Q{�<�j@46/Z Q`��L���u�<Id�T�]�r=�C!�4=�x��G�z�<a���>/�I�U�#}��Q��z�<!�K�a
�Q[G��
J~��%y�<����E��%c������O�<iŇ5{(��0!ţ)f�aX�BA|�<���+}���7 
�)�`��&J]�<�#j�3h ;�!�rfި�Sg�S�<�"�,/R��Ì�I�N��4I�<)Β���P�1�C9"���2,�F�<�p��$ٺ��S?/z��BB�<QEEϫw]�uۂmG)"f�%��~�<�n�"/��ܐaA��*��8�u�{�<遌_���2��O���j�@z�<�ׁŝJ��A�K�o��:c$y�<QŇ�O�^�h��CP��F�|�<�'��D����`�8+�ēQ�<!U$q���إ�Љ
hRT��j�u�<��= )p��>p����v'_u�<S��(O��@�U��<CI�$��JPq�<�Ē,z�u��	\"@N��qw�<�bk#PR8�if��q�F�����q�<�VJ�	"�=:�j�=s��yH�U�<)6�Ǆ%	 �WD�:7���2�^H�<��o��;���:@�Ёh�d�c3��B�<�gE^   ��   �  B  �  �  �)  25  �@  �K  �V  b  �m  �x  q  �  S�  ��  �  )�  k�  ��  �  W�  ��  0�  ��  ��  \�  ��  -�  q�  ��  ��  O �	 z � 8# �+ q5 �< �B &I hO nP  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e�'��O��P�]�۴$G��d�q%"O����bN�#K��X	0�O�#�yԮ���v+T�4z��s�����yR"?�EP���2.�R	��%z�=E��\Ȭ i��3Qlh׮�	.���<
�<����$�`�(��@�ȓ|�<��TL
!��qC!o2䭄ȓ~��s�X�\]��9�E���F�<I��^�C�}�R��-�h�J�L}�<�A0ho��+��ݐ%�]bUC�^�<���ɸ{�Z\y���6a.�Qe�Oq�<1t
���A�G��J5�-�3�o�<q��w����EQ�*@�p�S�<Qa�,��ms��Q$i�QzREY�<9�����A�Ђ8�3��R�<nM7w�jǁ\ۦ5#�E�N�<yt�g�zQ�EcKU�Z����q�<sK
 1rT�h�$��B�O�l�<!$�x�Z���U�����M�<�V�h1�\� .jV�S �G�<i��8�V�+s"[,hn��UaE�<��_�P�S��$t`�(;���J�<a�C*!�$�r4�KZt��҃�Q�<eب)����.��{3�����P�<A��]D"A�Di;c��%�ЩCM�<�B�<.�j�D�g���RbaDL�<��!İ<0��i�H�k�x�$�Q�<	�mO�
a2�*kC���[3n�H�<q�M&eP�(Q��^� ��%&͛]�<Aԇgގ�Ƞ��$~�$���s�<!�H�E��q�4�
,g�<	�c�q�<#Դ
���(d*�E�VD�9�!��6x<y�&F�(9&P��G�!�D�;(G�̨#`H�4�=�� �!�� 
%���J�]���"����"��,�u"O�$(�%)-�+�GT�=x�!Zr"O�EK�/**Y��W��!	�"O
��G�M�x�ؓ�I�#����"OԠ����$q��Ç
J�ʉ9�"OP���a�)a4������$U��"ON����m��� �0�,X��"O���+���s���X�)�w"O8�+��f�D��@%�* D�U�A"O��aR#k0�Պ�&28R(�'"O�E� cO5=�v���oϢn�@��"O�́��2S�pmX&�
&<�x|�"OR���A5L`#GD�4�8�"O<hJc$ϱ4 �p�!`��3"OLIE�%q�D\�/ � ����t"O:4Y�_�6f8�F�۞�`��D"Oxd�����p��!B�eN8,>���"O�@,ƋS��lb"'�y� �b�"O��aM� �r��4���M�F�C�"O�a���&P;��y �?�H�@"O�=�#$�/�J���/��"O� *G7Z{�����1EGl��"O�̈��HS:\,��!3NF@��"Oμ`��y�%�`a]�N6A"Oj���lW!+@ �p�9���"O�j"	O����:�M�&
�i��"OD\����4%Hv�a��K���H&"O��zC���L5ȩ*�,l�"O�$���]�}Q�|ɴ�Ul�> a "O��a��O#D��)�,O�v�"1� "OЁP���
DS�z�l��+� c"O�!��@�8��t��o�Ti�"O��8��$}ܶЁ-^�3�dyc"OTT�a&���d���"Z8y�Za��"O`���
�M�,4 'ĩ;���p"O���bG�F��%D�7^�M�"O��b`a�l�P�B�?*Y6`�"OxL�C��.�$4T��oA2q�t"O����a\������.$��"O4�* @d�����TE�ƨ�%*O�Q�O��t�4/ke>���'~�P���!3m�d��f&k,0�	�'3�M��@�s��(���Ǒ`9��b�'��5r��l3Kg��Z]z�z�'v���o�2t\��Ӂ�0A}�-��' ڼ�E��?t�����1S�@�
�'��X2F����FтV&��
�'�\�Ж���Kl>�(�CЗUք!K�'s����i��'(l�	RcJ��S	�'T�օT�Bt�,�ْ�)ƚ�yªR2?�d���W*�Fm�WͶ�yB Ò\��9��Ɂ)������yB'�7C�r@ϓ�8������y�,O�E�"u�B�3o���E��$�y@�`6A�a��4�����I��y�	ΐT�:�J�kY)cf1�%��=�y�.Q>H$��+�ꄾ�,��O���yb�j#Ԥ)���y
Z4��&�4�ybM*G���Q:l���9g�Y3�yb锴x; 4h�)�a�lŀ6HN9�y2A[�5��<�D��Qk!�3�yR���[�����L�T�����y"�R�N��Q�F��G#���dZ��yr>h�c��_W�j���V�y
� ���^�)AT�BP�M}�萗"O���&�ӱv�c@�k�p��"O��d�!Xb�c�� ��Ȋ�"O���M�U��\F���"OLu���/P�l	�����3��ak2�'���'-��'��'��'���'�vA*"	�;?��xU��<Z���:��'�"�'n�'~��')2�'�2�'���@JA����i�e�{�0@��'���'b�'v��'���'���'�ȸӢ�X4t�L��&%h���R��'u��'t��'�'b��'�2�'{@0,M�f�3�f���$ꍱ�?!���?!��?����?����?����?Q��"~����N"96D5�T��0�?��?I��?����?	��?���?qf-�JΔ���K��Dxd�,�?Q���?a��?����?���?Y��?!�c.!�1���_��\��d�1�?!��?����?����?y���?���?QaBD�)�R�a�HV=%c���u�ݞ�?a���?����?A���?���?����?��3gS����gR���j�kM��?����?q��?��?���?9���?���O{���do�;#0MZB��#�?��?Y��?����?y��?	��?q���&b��h*�/X�m�&!)$]�?���?��?Y��?����?y��?�ƍ�8t��q�P��(�`I"�?����?1��?���?��A��'_R�ڗ�LL��$z~�Kc�J߬��?�)O1�����M�`a�d��Xku"��o�^(���H,#����'rH7m*�i>����c���H���Rj(ے���&��x��/?��nZW~"5�҄��v�I�|��a�V��<�R-��
�3{L1OP�$�<���)ŏGk"\�b�҃n�`](�Tc0lZ�33nc���j0��y7�V'S	D`���?�Z�(򌕣.3��'���>�|�R�@�MK�'K`R ��q	�$����"
l2�'.��	�(� �i>)�	�N�\a��m��XO�� ���
e|�IVyғ|�&y�4q1��e8��Pq*1��D�vj� 5���X�O<��O��|b����m+j� c ��q�>�bu�|~��'���c�!��O�����!3�.٫e�
���N"��i�$�/B��Iwy�����d =�p�"�B�X%�ĺǦ�Yq����4��ĕŦ%�?ͧWb��p3&/5^	S5�G�N��X��?Q���?Q����M��Of��7��&�8?��xƇۗsx���D�MJ<�Op��|:���?���?��E5��z!@Z��Ӑ��!���.O
qn�K���������l����8�L��s�c�X�fNl�bOD����O��b>mc��ޣNV�(��L�T^R��F�T�B���^y��
�V���3�'��ɳX	x<Z��E%La�Tf��Ψ�	����I����i>��'�D7�
�:f���5D�P`�W�\�`�k���[_D������?)�]����˟��G��y�	)j$\�v��6��ܸ�$ߦ��'Q����?MBÞ���w���cL)&��Ш7'хx�b���'Gb�'k��'���'��l#���
h�KP)�:�Ԁg�O>��O%mZ�lt��T��|��*1M�X3�)�;ƌ����+e�'F����� N8_��&���A�I�8�Pȣ猇�,��d�݉I�@���'�x�&�������'��'߰q�0*��V���т��d,pI���'��]�t0ܴy6�A���?!����	ʀKݮQJ���[F^��6k޹-��I��d�O ��;��?�C�$�[��Q��ל{T@}H�E[<Ty�b���%V��|b��O��K>QƄ�x�T��JӉ@R������?-�M#���?�Ş��d�ܦ�SbH�.W�p����Z�nc H���p�I��l�ݴ��'6h듐?�c�+���4`s�l��DC!1�<���O4X�iӰ�Ӻ�D�����D�<9�-��/F�|�`昚H�t)��X�<�*O �$�Ov���O��$�O�ʧy*��b�v���,�9�|TF�ipD�S��'Y��'��O[�I~���R+�����C�x��� uG�����M�H>�|aT��MK�'�<p�Ί,��)���&o~��'����O]b?qK>�/O�	�O�tApIIO>�`�g��j8�����O���O���<��iW�E�#�'�B�'�XL
 .Pq^,���׃�.���$JE}"�'�B�|��	;_vఖ/Z�&�(A����d�j�l>ø�����MH������'�L�3��A�č4u^��6�'���'_��'�>9�ɼ5����LZ&�S�Dͦ�P��	��M�7JȀ�?��/i���4�:���
h�Y ©Ao��A�19O\�D�O�D
2l�7�#?Y�Ñ�zQt�钢!߂)�A�	�(a�U`O�r�p]J>�-O�I�O4���O\�d�O��ֈ��mq�P�p��58��)ғ-�<Q��i�P��$�'4��'X�O5��M��`�&!7C(H�x��]����?A���tNO)C��u1��M r�a��¾8�����92�I�
��xK��']��%�h�'ܲP���1����5��9+����']��'�����dQ�X�޴,0ր���<�vɩu�Ȓ����i��g�f����	E�f������O�g����eC�n� �(��6����M�O,hhъ����P�2�I��� �p
զ]�|GJ�hq/�lK.͑P:O���O �D�OH�$�O��?�a@-�H�R�j |�r��ޟ��I��q�4dpvP�O/7�/�� Lh��E�CN��QW��1O|��<ӅY�M��O� p�&�!{��Ʃ�bAL�'�v����j���O�ʓ�?����?q�>F���o�H'��aպ�8��?)*O�oڡc=��	П���q�� ��cN�y4�rU����d	V}R�'b�|ʟHI�ѫD�w�bՉ&�F��ֱ�w��46�<]8&U�m�i>1� �'��$����Y4p�}�T���e���YUޟ������Пb>��'QF7�C/��@a� �
3𲵚�剡
�d�H��Ob�$��!�?��Z�H��f�-��C@9'��-���)N[9�I򟄣e�^����uwF@<&����{y�ЖT#��i#��(6?��c�CE�yR���	۟���ݟ�Iڟ��O9�*�ɉ�Hua­v��i��`f�HMhP��Oj�d�O~���D���ݦ|=V����0!!TbV�M�g�Zm�	��'�b>���o�Ȧ��P�(���K�3<9`���/C��0��8K����<'���'�B�'ZV��� HRช��@,}j�'���'��P�h�ݴ`��A���?���� O1eg<M�v䅋I���ƘO��d
�O��D�O.�O�d�u�C+Y�d�U�\�j�,�ۖ��,���&H�p)��3擣H���ܟ�1�ڴX��-[®?�x�����t�I㟸�	ٟ,F�$�'��U@(��H2
����=<�8c��'�6�M�5�����OX�oZm�Ӽ��Ӈ0RLqQmޢ��M�� ��<��?	�)>�aٴ���'|p8P�O޽JU��iLlQу"H#.����|�R��ߟT��ş��Iȟ`r�f������ �Z
y�[��qyr�d�"U�1@�O����Oz����䚢l�d� �y�δ
G! �]�� �'�r�'ɧ�O����,ɄBQC�+ؕ(��q��*�^ޒd��OR�c"!��?�0i(�7?)g�:
���NM�\e��:��ן��ٟ4�����SSy��pӬ�cC�O���ЯS�^:���+�M���Ov\o�a�K���ɟ��Iӟ$UER��|�Ȗ�	p���b���.�m�j~r�ūjFYE���w�t�B��0!\9A���1Z�����'���';b�'���'�4�wL��~�Lx��Zp���J�l�ON�D�O��mZ�}����,��4��M�j`��(z��(�&ϼ6�N��L>���?ͧgq�e��4��d��:��R�e]J�2D ��3'�^��!�+�~�|R^�D���������Cb�j Y���?q�2 ��m����Iay���O*Ģ#�'�2�'	�S.y��ɐs�ȇ
���Q�b�	���Y�	ٟ��	L�)�-�� �����.D9���_�i�`NM��M{\���sn�$1��O� &�"�ȞHx�	@�G�/��D�O����O���<y�i��-X�\�`v�@���:�\AQ�-eh�'��6�4�I����O�|��̅�v�Z��/>W�T:��O���^�O��6m8?��>�^�b�';W
�s0��u�ɔ�@�iЅj��T�����O.���O����O(��|"!҃7C4ɓ�;f��#��ʭZ/�v�G�yV��'��)E��ݝ3mpPz2JW�g��P�D��{d��	U�ŞB̼+�4�y�%�$\|�D��7zDHBD_�y��WJ
L��%t�'�I$���B�� OM!CiYP�b�~����՟��I����'fV6T>�
���O���O�n�R�k��=�l̐th�8���©O�d0�	:�|��a�}�$���D�����|�XIz�@!i-��H~2���O����O؀P���=�.��7�әj�ڭ���?���?����h�6���4D:�ِ�I�TDfR�W�4���Ӧ!
s	]ʟD�ɮ�Mۉ�we�]����~����U��C��y��'mR�'�}{�i��	�W�b�)�O��਀-��S��I;�!��r����-NN��Ey�Od��'%��'
JT-b#��d�!E6�څ&��2��ɽ�MSc����?���?iN~��9w�kMA�s�ĭ����@K���VW�����$&�b>���ΐ �����E�$�DA:Ux�!lV~�`�V�������$�,84`"��/�(8�*܆�����O����O��4�`ʓ��`�g����5�]�wd�	t1r�ڥ&N2�yӞ�xh�O"�D�O(��6v��D,�7��ur��s�&����jӠ��nE��m��,�>�ݙ ���@lIcj`�s�_�QA��I�@�	����	ܟP��^��[�����#K�B N��5�^8	U�5���?A�Cݛ�,E'��d�'(D6m1��.5��@b4(�M�\YZ'k<���O��d�O�I� ��7�&?�;�v�#B�;`�A�I����9D�ջ�?Qf�4��<!��?����?�B�
6"����/��M�Z౥����?������զHn�ܟ����ԖO��Q(��7\���O�*1�<lj�O`��'�"�'(ɧ��K�_�dAЋ9垽{Ve�%���n�d��7-�ay�O=�5��� nrBH�
V����.�$!����?���?�Ş��ԦyN�^
 ��5�D�lJw��_�fm��ޟИش��'�"��?�SH�tl��ir*�`KT��GG�?Q��.KR�Q�4��d�b����O��)� *���'F�p�4���Ցa���4On��?i���?)���?������K�Z�,��Ǩ=pv�Qw�O Bެl���e����IV�SH���{v��S��Ȱ͑%#�ك�ŉ�?1����ŞC���ٴ�y�"(�a�wLsڬ���%�y��~�P��I�o��'��I��l���m�b9���S�Oy�H(%�&��|�I�p�I̟Ж'��7� �
\d��?���߃�4%����������'����?�������Ya+jAcW
ͮYS8��'Wl�����}����i��~R�'BlD0�`��v1*-bA ��`�'R"�'L��'�>�ɓo�N�j׭ǘ
u����3t���I��MF	���?y�qݛ��4��pi�͠Œ��\#!�6݉">O���O���U�[�\6m ?	�HB�Gv��I�%k�<��%��-_f>�Jva�9[�U�N>y.O���O<���OL���O@D0q&֬QEΨp�G�t+���*�<�B�i@|R��'��'m�O �F�"�>�{��ġ="�Y�`�0S�`��?i����Ş]�T��aI���+�AB�P���$'�>�dr+OF!����?Y��$�D�<!	EdA����	Y��t@��?a��?���?�'��d�������Kb�˥&�{���mFVh�V���ܘ�4��'�b��?���?#��!&�9���ANV\�`��{D�|*�4��䃵3>�Z��Lfޒ����!z��3��?%��Ցu�D*8��Oj���O��O���)�ӼVJb�`����<u��С y����ɟ��	��M��ǡ?��ɀ�McO>1�ʓ�TG�I`@��i�t���?�䓹?���|�1��MS�O뎘4����%K��LON*F��c�p˓O�O�؃N>�+O����O����ONy��'�87�9� 聊vf�t"G��Od�$�<I2�i��y��'�2�'s�,+�q��C�E.��sүϔ_1
�r���̟H�	v�)��C[*��)�h�{xꝡ��{;��`]*�������P��LSu�|r%	�?��%6N�O�P�i��A���'��'��d[���۴w�T����)rt�aiƶ%#��[6g��?���J�����e}��'�ȵ�$���ء#��l�,��v�'�"��'ЛƔ������l��ɼ���L��?q�rńƆi���\yr�'[��'2��'�rU>U�E�D.E^ms��]���1)�MqF�"�?���?�L~���#>��w�$�jc��U����Ԏ�A��}��'Qr�|��$l@O��F1OtA[_@�貍G��D(b �,�N�4�`���$�Of��|��,$�eq� Q=Z2\�1A��(Nz�$����?����?�-O��lo�ΰ�����	f��dH�T�ԐT�R3;��?�Q�d�	˟�$��b�FJ�4A�޻(.�E��'4?���<2|�=*��NM�'4}���O��?��i�tI�c���2��\S��]��?����?����?y��I�O�����/|Jz��c�"'!�
�O�nZ�&|N������Yٴ���yWd[:W�<P�$�hl�*@�@�	ǟp�i�m�6bS�m�N~"�ƫ^���8W3h�0bM<%�r�{�G
�M��!�|�W��Sܟ��	ʟ�I؟�+�����1�b�.Z�t RDZuyңmӴ(#�K�O����O�����u�1�3��B�CR,ڒe�
��'R��i�� ��}�� ���&�ܓ��ǀ��ʓLn�4 R��O |sI>*OT��!��1�m�5#;h�~����O���O�$�O�	�<�%�ii"}��'ܚ@��T|L=�j�&�C��'/N7)������Oh���OfD�𢅶[ix(*��˧2��AYP��i46�??��G1>��7�S��u��됚`� �j�f�$�<L �j{��������	֟��	ȟX�rb'�hH���Oɪ �i�2���OR�o+p�����Pܴ��q�H�M1HDH$Z1`ˆ��O>Y���?�'N�]Bݴ����H��'S�L|���T�v�6E�GǮ~��ŧ������O����O.���fuC�C�U1�\rn��%����ؔ'w�6ɠt�����O8��|�kO�~�,҂B������Çi~rO�>����?�I>�OjIq�@D�&�@-�u��.���1�W�r%�p�i'�i>Uå�O̓O�Ĳ���8 ����.Jr�钧d�O����O����O1��ʓ3����q�r��3O�8+�\\��h޾�l��'�"�e��<r�O���׼K�QȒ�Ƥ+s�us4&�z*����O��ٷA{���z�!I��O�jM���I#n��P$��#)�8tY�'����D�	韘�����b���5@A�!q�H�;C^vR�ߑ1(�6-�O�d�O��D"�	�O��oz�ը�
G
=�������\+���Iퟤ�I|�)�S���lZ�<��';t�ܘ@c�Y�ȉc���<I�̅	<g��Iq�	_yB�'#&ТUE0�
͑A#T4b�pK���?A���?�)O0�m>_����Ο�I�I�x��+�K�MS��(!��T�?q T����`�o�"���� �"�14���*�z��'@v�J��1Oi���g��d�������'���S�oǞ�t@sG�B;�а��'�B�'���'��>����iT��!�W 9i����D��-R����M������?���Cћv�4�$��c�b�p E�'-N�`� 9O�d�<�t.A��MS�O�}b����"�� lE$r�(��W'5T�0Y��/��<����?9��?���?1dKҟPF��w�šW�܀�;��Y�����Fퟌ�I�'?��IG��c��B�*-_���b�O����O��O1�`����T�]��`�E#
�F��U҆���aP27�FDy"��&��������l�3��F��ED�0���D�O����O��4�V���Fl�	TD���5]�¡9�n��Cд��sJ��B��f|����O ��<����c1�X�d ]-ʹ��i��1ܮ���4��D��Zn��A��0�x����.�'i2v���f�Fr�����	/&��D�O����O���O���7��->����	�:���	�'0>��	�P�	=�M#�G�T�n��O2��u)ʆ���3�7sׂ���#���O��4�>�ed���}�]�Ƃ��A.��2���	P���b�\�c-��������4���O��\5}����&�O
kj�*�.	6P���O`�F�FMU�r`b�'>2R>9S6垶/eڙK���e��-!f#?Y�Z����K�S�DmǗvlF�h��ކ90��!X��v�iWb��2��y8�W�擋,g��\L�I�z�Ty� BE�����k�7GD����d�I��|�)�Siyly���2]�8����=@<��������O��o�H�v�����4r���k��A�a�D�7 Z��@ß`�	�аloa~��-h�d��}�O˖j)����P'��X�%Ζ�<�.O��D�O��d�OL�D�OJ˧A���RS�ǟ]�|�3�5>�����i������'{�'��Oym��.f:� {t�G�`�JSI�#�"���O>�O1����$(kӢ�#�fS���HثV��ah<�I1�@��Q�'?�I$�ܖ����'6�]�$�P�S�"���eB�$�q9P�'y��'erP� �ݴ�u0���?���R9�$k�7z�"h�c�O�)z����>���?�K>��EP3�6��#�%1�mɦ�Sc~�G
"[�@йi1��@�'��#G�B_��{HWr34d  		Z�M+��?���h��N�z{2[6��gtq3�aS�k����T���Yeƌ�`���MC��w,�DkK�<_�t¡�R0�q��'���'��N��Ui�f����0�m��A_8 7h�)��؀(��Cf�|�X�\�I��������IԟȚ,��D�٤�%΀ �Ua�y�t��\���O����OҒ����O����+U"��K��C�>����?�M>�|zq'�#E*�e�E
 Wc$8#4��p��Eb޴��I�qunȫ��Of�O�˓�v��m��fլ%C$�%^���k���?����?1��|�.O �m��o�֥��l�6Q�#ϒjeXE�v�M0]�Ɓ�	=�Mk��E�>����?�;#w`��C>I���lH0���1޶�Mk�O\�P1Gj����|��OE���S�(%�T��(@�xRoѽ�y�'NB�'�B�'�����D �B&�� 3�c�N����O��������	t>��	�M�I>��I�*"��q��M���Шtɛ��䓳?���|��	�
�M��O�dr@�C7�0��!U8���B�(-(p��P�O ��|����?Y��O8�14-n��L��b��0R��?y/O&�n��#�q����x�	J�4�ʹ�~ct͈A�&Q�!�����D�Z}"�'3�O��7�Ҙ24lZ;=��@I���8	�>Tx�*͚B���s�Fy�Og���,jQ�'d\���C+�P$�U��:R||�1�'���'�����O��I�M�U,�S"|���)$%* B���/��T��?Aw�iN�O���'�2F��;ذ��F�7GP8�ɜ���'�6�cѰib�i݅����?��]�TI�B�~v�)I��D�2nЙ�����'���'�'��'��z�Ra�q
�$�p��b�$N9��Q�42K�%���?����䧌?���y���3�ݚ���	L��a aD�)t�2��	ɈF6�o���"���Og*��D��<'0z#s�|�|��N�R��b�IZy��'�"&���]�aHAC��ʅ�[%w*b�'���'s��%�MSgG�!�?����?���T ��L9����i�)	5����'"��?9����'Lq��Ǳv
,��"��O(���'� |Yd�I�"�P�ya��t����y��'0�x� gަ��iVLפl�:��'?��'�2�'}�>��	=S[��dFT�x���§27���ɂ�M��X��?���,����4��PX��h�	�1ET�r��Y3<O����OL��~�^6�0?!镜5{��)�Ѻ	C9M�ܠ�o�>b���JH>�-O���O���O*�$�O��Z�Ё\ei�Yk� �<��i?2Is��'	��'�L���i�C!��"��f���AaH}��'��|��4G>i/�@�%�T�N(��Q�@R	C��X�f�6��ā��½��h,�O�˓!�����I�~�(\����p�X���?����?Q��|-Od�l��su.�ətub|�e���PtS���B���ɿ�M��"e�>���?!��G%�ySb�-u��)��/$Ti,����޻�M�OT�a�fӉ�JrK4�i��ę�!�^�#�D�!�Ã�@\y�6O��D�O���Oj���O��?��J5$��yc"�Z�<ţ��_ٟH�I埀[ܴ\�<�ϧ�?�!�i��'��w�
%?��([(w���y�'a��c]z�m�Q~ �� ����'	�� {�k)Eڅ['Iښ�?���&�$�<���?)��?�Ə�v�ӵ�k�ժA���y���O*˓^,�H�@c2�'�X>�a�U�S�!����9N�Z�!�)?)u]���I֟�%��?��B���+�����R-�^��Ê!Yz�58� �l~�O�����Y��'���
����uɖ��D%��`#F�B�'�'w��OH�I��M#���
�^�C�މ��e'��R�����?��i��O`H�'�҇K52X����T���30�J "���'F����i��i���֫��?)3�X�8����	AL|Hq态& � $#g�(�'�'`�'1��'�Ӷ5����U�X4���5N�8� B]զ���������	ğ|'?��I,�Mϻ}�,a���U���b	 2�|���?�H>�|�q���M[�'�.e3&�8q�>�؆�]1�]��'p.�G�ɟ���|"X��⟴[�×(n�4�`6[�S�rM���럄��؟H�ItyM|Ӝ�"�ͺ<��n��k��))�B�+�`�*��컎�ϱ>i��?9M>�GR�u�a�!jJ�Cq�\ȷ�e~�CT�naN��j�	 H�OtJ��	 �a]�QS�i��"�\��1:��?q9��'��'8r�ǟ$
�-3L b�h���cn�n����3���'�?��Û��4�$I�u(��/�&�
�(W0UH�T�v3O��d�Ob�Ė'={�7m"?��<T��S
;�8��j��+���2!���:�$�������'��'�2�'08�2�nT���F�f�j�W���ٴ5%z�+��?����O��ܣ��̕96�OVB$��!�>���?�J>�|Rj�XZ�h�bK�8�^0YA�9W�H���4��D(�H:�'��'�剈U��U��_,C�F�w,�������I⟨�i>��'��6M�&�@�$��L8��"����H9�p����?Q�\�H�	���I�G-���#B��[��1���*����3����',�(���?��}:�;I�H$��퟽(�j�(JD8ϓ�?����?���?�����O1�MqW,Cnhq��=q�nl*F�'�"�'٢7�f��I�O��lZw�	p��i`�AD�{>���`ݱR�%������#B�>o�u~�$}��e���V�Pq��O�'E��U�t�\w?YL>/O���O��d�O�a�@R�a��2�g�6B~���G�Ov���<QƽiR0MY��'�r�'�哳WJ��Y�GS�eG���Wa��6o��@�����	_�)��D�3Cd�G�R�Y�:ղ���`�b@e�]d>�������T
%�|"�*�~=z�$�"8\f�"�H�k��'��'���DQ���ߴF̫���eP<(��������<�?Q�y���$�^}r�'(��d��������ٚ7~�����'NG�0lᛶ��<Ae�"%o��~���&2-BH���ޒ7���4Ϥ���'n��'6B�'z��'�哳�ab�폟~Xh���ט'{
���4�$�����?y����'�?qִ�y�눊�x�S6Ό'X�T���דi���'�ɧ�Oq6@�T�iG�/8Y��lV�+4�)�%K��ē�C�B����W�|�ON��|���k!|%�C���[$�,r��N�Ak��9���?9��?�.Ohlڃ/�����(�I%�޴�'�\S��D��T(I&̨�?a Y���I�L&�l���^H4ĸ8Jڂ�t��Q�8?aqH��6O<M�e����'>M2���?�4a=ܴ-�CȀ(�Ѕ���ԅ�?���?y��?)��)�OF��$�Y(<��NR,�q��O�}nڇ3:�A��ş8��4���y����@~�@c�/n�D��fň��y��'�B�'��$rV�i��5Q��	9r�O��rq�ƃi`b��D*@�H����[i�	ky�O��'���'��]/'�D��1SS,��D�\/W��I%�Ms�$�?!���?1M~*��Kh`����w�ƈSF�;?$���T�<����%�b>9���;B�YE �|-�"SH�Yc��"T.)?E������]�����$ $ꊌ���*5H�Ļ���;KA<�d�O����Oz�4��ʓ2ϛ֤R8 I������(�Ev�(I�i��Ch��H�O��$�O ��?SLe#N�<
��u�&�юo�͉�&���F;
�[�/��Ј�L~������î�EGT�1�f-��xϓ�?���?y���?a���O����D��a��ȗ�K<�����'��'
�6G��I�O�oB�I<f�,XF��"Ct$	��F����'���I��S�A���l�k~�Y-����+_��� q� �YV@ RH�^?AM>!,O���O����O�\Cu��bJ�ٹR� a���f��O��D�<1S�i��3R�'�B�'V�S�0JE�\�t�ޥ(�
Z�(�����Iןd�	b�)jS�N���9�Ȍ_�(k�%V6�tX�`��Ms�O����~�|� �c�$%��kϬ;��wea�-��0۴���AI\6����V��1J���;�*Z����ݦI�?�VW���I�O��h����h5���ּ�	Ɵ� �`�ۦ��'&�"�&Fn�*Ot��낪L�	!7��fN�i?O"ʓ��=I�+�'��;C�Q�E$���j�6L��fg�>c��'M������]��A�ǋ��d�b �~�	̟�$�b>���b�ئ��S�? �TA���K:aA�"9�Рa�:OX�aV����?��)$�$�<)O�d��e܅K�28��<W��QIS�'�R6-M��8�d�O���O� _�hP0��2��f�/��⟸c�O���O6�O�L��8`��R7�T�dZYؗ��k�D�x���N�E���Qܟ iY|-�m��m|)�@1D�`ؗoŪr~�Q�j��Q�\���şp��4g�iY/Oj�o�f�Ӽ+��M���� �Q�"����E�<���?9��ƙش���8X=B�Ol0KF��dL^���բ-� a�S�|b[��D2-Νj��yX�#�s�R�qU�������a�6�U��H�����"W�K:�8�Qt%D�:���ş$�� ��M�)�ӀaJ��Q�ҩ��i)f�d�\-ؓ�η��'>��s�!���T`�|�Q���ը�$$���9�d�/��m;�.�OB�mڠ}���ɒq�q�#U+;/���e�ݥ?;��I/�M[���>����?I��r��Ⱥ��2�9�3D�E���H>�M��O�{b$^$�����t�w=R��q�K?f�h�p
by�`��'����<U	3���(�Eiؾ!���@��4f�X	�Oc7�2�M� �x��Z�D 
��C$3KԒO����O�:1>n6�-?IS%��($H���Ą�`
�h��"�2}���R�� &��'�b�'�"�'�V!���&��d)���4�����'��]� B�4.�P���?Y����lN�i�� o�d]�1�>��I�����O(��''�>x���X>.���T@�8? �\z�*�<��*���4��K�F�0�O��s�#"�${6`	u�T���"�Ol�D�On�$�O1�6˓3כ댤9U�(¡�.al���Ń
U0T��'r�v�㟨��Oj��S�!	��A��31�@�F�[��ʓ&y6�4��$�_�ؘ��i�(��P���N�<"l\X��R�W�y���D�O��D�O
�$�O���|�@Ő�B��)?h��8c2�L�j��]�S�2�'G����'�b���C7�X�U瞣*{z(�E���(��9��?�J>�|B6J7�M˟'�U�#c�C�V���jA�Hz�Lc�'3��;DIM?�K>�,O���O�X�d뒹E�^�"��F~�9�bF�O����O��Ļ<���i"H!�W�'���' Е�a\�Jk�=�񇛽	���(��
[}�'+r�|�N�aJ+Uc���)�p(ϼ����0:.��Ypf}��c>m���O���o�LMH��ۡ���
����O�$�O��$>ڧ�?�a��f������ ���x �/�?��iL|��'�n�����M`�(�"V96}*֠�5�*��������I���'���h���kz��si�����*��Q�ID�<Y�9$�X�����'�B�'���'�hm*PN[ 8ր]�gΈu�ʆY����4W,��(O���:�i�Otx��\�j�@(�D�P4��a�G}��'���|��T(ӵ3�*!���p�!j���j�I�iq�ʓQ�=�F+��D$�`�'{X(3#N�:��8rK���Π��'���'����\���ܴl;~��#��1Ec���j��Th��q��i�6�F�|�O�h꓊?i��?��G';d2xX�׉�B�S�L* ؎���4��d]3U�F���O��O���]$������.!'� ��y��'"�'6��'���)P�+f.0q�BN����4͔*���?��fD�&�V�����'�F68�$�1k�D�9���*A�
��j+ц�O
�d�O�I�%8B�6�'?�;F��\(w��U��HJUI�1*3��DkL�?e�%���<y��?����?	�ꓨ~Xj\PE
�g� m��[2�?������񦁀�n�������̗OlЕ�-L�U0�|XJ�Q���'��j�>���?�N>�O3�mz��"'=� 33[�^�Q)�]�G?�����0y��i>�X��'���&��,��Pp��X�"���P[hU֟���Ɵ0���b>y�'J�7�ҿa7�Hl�8�b� S��(����d��O��dTϦ�%��S�����O� �_J+�/YL�;7�Ҵ5���'~t��is�ɿ�%�L����[� &-S"q���v&ݴ/��)1��p�L�'���'Z�'c�'��D��yA��0��=��jk��x��4s��:.Op��-���OTQoz�	Z�!�.,�x���@W�?�H�����l��L�)�.ɺn�<�fKϧ<j�D@p�զ
�N�����<��F@�T�	d�	Gy�'�2@O6//Nf�U�PIJ�B�\5Q��'t��'�剎�M#PM	��?��?�6�:S�
pB�"!P���� �䓐?Y�P���	�$��C�J�%N�ʐKs-�8������-?1��Q%�y"gB>��-��$C��?�T��&|6��g�;��5r��޸�?��?����?�����O����	�\���r�ϝ%\�D�b��O�PmZ:����ӟ�1ٴ���y��V�?� �0��N; e� ɗ˞��y��'��'"��i��i逐�ս������_D��#7��c&a�D ԡ{7��O,��|
��?���?��1��i���?l�c���;R��1�)OPl	7Kܙ�	̟��ID�S̟\���Th ㊵��15M�.��d�Ol�9�󩉺�� � �f�)!��	����
��<I�`�kR�	�=Dx�!�T��v�%8 �l����pq�ˆ#��И�G�3^�:8!h�r�R��!	�n,M%*Є��IA䫘5"�xp�"A�)j�����o�N����@0,Pat�
E�l	[��Њ�㟼R��6nx�b���6����e�$����a�o��
��ҽ>B6幱�R��*"�X6I5�Z�ˡ6#��t�ʿ�d�r�$P�OT��dĻD�k��U,}�b�慅�n�>����Wd\�뵮Å`Jp(
�nP�%X-� H�f�ސ���	�\���1Gھ-M��q�42�J�1���i��`*�@�-���g�i��	ɟ�%�L�Iɟ�H�l�>	��(�,YX���g�)¡�O}b�'��'��G=᨟
���L�NX*t�E�|O�]8`ǈj�l��0$�����xS`�I�x�O��H�l�s���h�ِZ,�8�iR�'l�ɽ�tk������On�)��+���H�$~<��m�6�B�%�|���dK��0����/qp;P!X�e���(�+1�M�*O�L��f���Iן�I�?�(�Ok�Q��X�xp��.W�^�a�,ΰuJ�F�'B�W: 	�OZ�>	��햚l�h�!`���xJ�{�T�p����U�	ǟ����?q��O2ʓu�
|h��L�?X�����5�ֵ��i���@G��%��tp�m�'�\��-����W���M����?���3iY�V[�X�'�B�O�퐠��1���!��M{(Y����FZZ��O�d�O�d�H�Y�R�����` ��n��@�SfS���<�������K���g���L冐i�
Ǉa��c|`;O>����?�����D����%i�'�"n�ܘ��>^&E��˅R}2P�H�IC���L�I�T����4C`J"fc�M#0�0�Qq�؟d���H�'���� `>QX�瞴b�,�#	x�<h( O}��ʓ�?iN>Q��?���T�~�b]�`������G�6=#p��5��$�O��$�O�˓0�~D3�X?M�	�`!,x��g��	�	��Q�F6$ڴ�?�H>A��?G@Y�¸'�.�����~w��6M$=��ai�4�?����U-c,��O|�'����*l��T).!r�'a�eTO0�d�Oa1�<�	G�s@Gjƚ��冁-�T��F Φ�'�\(�Ol�����O�����p�է5�L�Q:���Hɏ\�|a�5�M��M��?Y"O̱��'<q�&$�G�Βd:h�!h����M�Ms�n��9�v�'���'N�4M�>�-O��	����sԤ���χ�w���H熎�ISì�u����Our@ĳN2Ψ"I��`�ɺ����7-�O&�d�O�`Py�i>��IA?9qlө!��H�UE'@��-p�Z����	Z�	���9O���O��D�)AY��I��<R��q��WD���l����j�nZ����|����Ӻ�VΝ�;�6�c���/ĦIIq��A������'���'��_��HdL�?�BS"&��1�
�0bG��6��K<���?9K>�)O��ݠ���+�&{�wd��aB��"��i!�V��I�IZy2�ÌY�0��uۆM��"Č:V��2���*���?����䓗�4�"��l0c�n��U�`7��:��>����?����ب㪍%>�ې�Z7����'nT�$�:i˶�\mZџ�%�ܗ����'��'4iղ�Ŏ�2�����3z!�mZ�h�	Sy�C�	4jl��D��k�W� ��j\�z!
ԑ�%%
�'���̟��|�s�֝�^K���¤A��`��H�P���	��9�Iٟ<�I̟`��cyZwny�B�	B����@�7`��Ua۴�?I(OF����)�Ƀ2�d�ʱfH/���f1M��*[��'�"�'n��P���X!i��B9��ȓr
K�f���XW]�4B�!�S�O�\D�adN83��z&KF�5M����z����Ol��7`6�S�Ĝ>	�ܧy�
ѹ���t��T{�l�(!�p��4�'l�������t.[(C��ӓJ_B_�6�'Q�}CU�x��� �,�6��:�0�`��T��b[������<8�<1���d�O�Ѐ���bL�2QO[��6�P��KL���?Y����'��O��1S�C�#�X�"NB� j���i�����O���OF�Ĩ<�&d�<��Z�� �`K��;�D�97���16��ğ��	y��Dy�OM��Q9O*Z�1!�Mr��aI�^OP��<Y�yEά�(���F�'�T<�b��XX������\`l�Z���?Q+Opq�!�x�]$qH4j���	Z���mڴ�MS���?1)O@q�.�R���D�s���å��T�9ƍW��%��'2�<���?	N~�Ӻ��J� ���P�F*2����J}��' �(Z�'���'��OQ�i�-�7f��+�ڜzc���e�Nah�c���D�<��T���'y����o�h"�"���MpnlZ�+y��gӺ���OL�����S�D��#<�ZQnB=Rz9C�G�����Gx���~��:E우P���JU'̀Ƅn���4���Z���pyʟ��'��Iѽd��FN2#�>"O5={�OA2�'.rJ�V�
�`q��n�hh�fb����7�O�-����M�i>�	]�i�i��dA�|H�(jW�?m|��A8�$�O���?��?9*O2Q��kV�M�|�᥆�c,����җi��%�\����`%�X��u� 
(�"()�"�
���M��d�ix�W�����\�	^y2m�)Axj�ӈ+�d��
A�$�����@ZX�7��<)����O^���OV�t:OXD܆(a:�����#?d軷�K����	韤����x�'�؉��i�~���d��5� �@�=D�K�������UyB�'y��'�� �'���OtM(P��MN8��D�<f"��ձiR�'��3%�$����R���O���B�`)��ծR�����儹L�r��'�r�'&�ꎠ�y��'��NRg��;�,���r����٦��'�X���`�4���O.�D��
ԧu(S-|��5�ѐ_�� :�#&�M���?���<�L>����
9��4a��Q+��`D�#�MkS��_����'q��'E�t��>�+OH�	#��bq,D�a%(}�֎ߡ.z6�\�so��O����O炜C�p�#%B�s�:��w�օpOB6��OR���On+�H}"R�X�	i?!��7�8%;��h����^Ħ�$�P�%b��?a����$Lǚ���R̔� 3�MQ�2�MS�,8��$P� �'9RX��i��@`��#n�Ls����^�*��>�'G��<�-OX���O��D�<�6�Y&7q�ɘ��;h��BrhH�i�a�$W�l�'�RX�h�Iҟ��	|r�1f��8�.P��l7�I�s�s���'Tb�'j"V���A��.���l�
5��}�䪓Q��A�C���M)OV��<��?Q��|���ۣ,@�F)�E��kڦ2h)9�Bզ�	���	蟌�'�1���~Z�!��tD�I><�w�J�FK���M�����OF���O2��3O|�$�����^��9�,�(5��#�s�����O�˓���Z?�	͟��S2TqB�bf=Gt�Ѩ���J�dm�>����?��nϐ ���9O��SG䭋7L���0� �ح��6ͨ<A�G�.ƛ��5��� �S�����<@�S(�5�MxѦ�	�<-	�i{��'Ѹ���'d�W���}���y$n)	�h�T>E� �V֦���D��M���?������T��'�h�u��>�u �0=�t�SFkӴ��32O���?�����'�~�r�P�}���(��y�5�at����O���(j�Ё�'�Iџ���)ꄴ��%F�{�:��c�)�nen�Q�	J�F�)"��?��!m�� ��9;ӌ
���#�$𡂲i�ЇC������Oʓ�?�1�ȍp �bq��b a���l�|P�Hh����՟t�	ʟ,�	Jy�+#���2��{���)I֐�;2��>�+On��<���?��c�J�i�ِ9h�L� ^Ҡ[�a��<�)Or�d�O��ħ<A� F�!�	_�a��9 Rşd���;��f��\���	my��'A��'���ۛ'�vH���')P� �UX�@�Q�u�����O����O��&���Z?1�i�Q�!O�� �P��ρb����t�&��<a���?���
#�u�>�d�.ٲ�*xu6���c榕��� �'j�J��~��?��̖�ZU��S��(s0b'LXgR���	ٟ�	
\�IO�Ix��&[L��y�ǚ����A�Β�a�'�� �w�m�F��O����޵էu�(^z
�%� ���BT��MC��?�g@�<����'*v%���%k�֡KÉO�87�A���ql��\�	ß��S�����<ibh�lr�9k@�KL�֘��@�=~�����y��'P�v���?a'gY��H�sW*�P���@E��N{��'��'3�9U�>q/O��Į�����JE�y��
,���9�n�r���O���Ԅe��?e�I�|�I�>���i�XX6u3&+K���Pڴ�?�p.����	Cy��'6�Iß֘��>!H�'_�I����!��\ܰ�u�V�Γ���O��D�O$�rȼ��E�[�Sm��#CQ@���'���]y"�']��ݟ����h�_:v�@!����A.(��F�S�P�I�����ɟP��� �'VT����t>���D�TOĜʅ���IG �f@t�`ʓ�?�*Ob���OP��"X��	3G���b��&H��ѫ��Z��`ꓩ?����?�-OD�ɍ~���'��B�� #�Y���G���A1�nӀ�D�<9��?	��QD���'@�$��P� ��u�-Ԯ�a&�{қ��'�RP��z%dP���'�?���X��鳍Ⱥ�ǫZK��`��x�'7��|��|�ҟP�R/O��>���V>����iC�	9�x��ٴ:z�Sϟ������KfJXYcC�ZO�qy )a˛��'j�R��|B[>	��RL�Y+���<�����o"qG�pn��U��m��4�?��?1��qV�'er��v�"��-�@zX��¥��".7���X��d/��|�'
"-�9HI�@�cD�w�DT��/�W#�6-�O��D�O�Q �j�^��埌��r?!����ۮ�8t�ǀp�A�rm�צ�&�prGN�(�ħ�?���?����6*͚���/Fa��/��
B�V�'��L�v�(�I��&�֘�Sv���N n;�L#4C�'*:N�xP]������O��$�OjʓF��a1h	8� �ŀ��j�.�ZHTj��OT��8���OV�%&{��b � �|>P���OT�rN�g3Oʓ�?���?(O��r���|J�D	�.c������:0�a��H\x�	ǟ'���Iǟ4�W����0�7iH�?θm��R�-*�@�fן����O>���O�ʓ%N0D������l�t�Y��Q8$L�:��:Ql"6��O<�O����O���'6OZҧ� l�KD"Uz���4!F>r�64Q��i���'��	'Fb�y�M|��2��xI�m��Ɏ�{X�u�!	�87ˉ'�b�'0�h4�'�'o�)3fh�@�U& k�ϙ7'��\��q$X�M�rR?��	�?�[�Od�)gk54�)��7�M �i���';��i��'�'$q��9����V3��r�lU(c)�8���i�p�i2f�
���Ov����$���	�&��m���j� X��
��[ٴjB��Fx��I�OZ\
t�P;:D�"3�[����+& ������x�Ƀx�$��}��'���~i�X�
Xk@�rB	��T��Ɵ|��ۤ/�����$�O:�S�G���g�C(O��M�DoL�7��O�\`�)O~쓛?AK>�1%rݩ$囊��e��*����'~&�������O����O�˓Lb̩1�_�{��Z���6���C���f��O"��;���O ��G����GQ�tE�|îºW&Y�u�d�O����O˓��X�S9�� B��"�RQKG��?1s�rX��	j�'���şX��Jږ\�p� ��P��|*"i -��$�O����Oj�V]l�R%����E74���S�FF'e4rP���'Q|7M>ړ��d�Oh�'p�������V9r!��(UW��ܴ�?���?��#�S���?��y�'|6�z	^7	 �D�0#�-.�J@���x��']�	47D"<�;c�*}ZC&�	
�~,�&�[�v��meyB@˨Yn7��O<��O��T`}Zc֜��V���5�EcA�;��M<q��hOP�'����/�,z9���a�*�t�ݴ$�dJ���?i��y����$�|B'�*Q��qmc<�ȑ�i�����0�&#<�|���Q����o�n��l:�G�%�I"1�i���`2!ɦ<�.OT�Ĥ�h�NѴ"�����&�~\"Gd�?�Ov�%>Q�IϟH�	;E@��'V���'-��_9��ڴ�?��W�������'�"�>�c���:��TycL�U����Ʉ[��Z�	ӟ��IПx��ɟ��uN�	\������t����TI�."d���ޟ��	�l�II�I�h�u�JD��)֑#���aӜz�.�l�6w����?�������O���%�Z����<j��L��B�<e*t �M�&T6��OP���OԒOR���<Y��ʦE����W��0J�KT�4��>����?����D^-F��D$>��@�M-a@�$j�GP�7؜1����"�M������?�����>iHjD
���/ˈt�ഀ��i���'剡Cj��XJ|������<4Q�Pn�;"̰郂e�h�'E�'m4����?��%ƈJ4��+o�X���H�jӺ�2�\�RP�i��'�?a�'yV��3�DqITf�T	�q�Ȭo�6��O,�䍘�0�}Ұ�^<wH��1wo� h���G��˦y"�	ǟ�I�����?9����ėO���W�\�%��MD5#�hk���>�`kH���O3�Nh@y��~+ ���.��6�O��D�O��`�`I@}�?��O��xKM�qtR��f�
<m�ƨ��z�'�'_��'V���	.�p����Z�b��hB� 6-t��D��O��@���'��'�p�d�)���95�J. ��=	p�=�*#��0O\h;���B�\��\&����݉`��!�!���VnMk�dH����h/L�Q�h`���5dJ�Sp*ۢn�H�JT�\x��q+ȻSN.�F뉟rE��:RIF���[$f�`���ɗ���)�L�Z�.í����턅F-(��NI�?�J��ʈ�a<�iD�	[7`�p5/���H��D�L� Q���	]��#��8#?�@`g��iQ�l9�I
=���Pç�=�`�C�ǅw��*&��:I|���O���4U�,��E$	ʂ4@�F�M�O�\��V�.1˄��t�Z�^�s���G*m��<ѧ�Ӧ�Xd��O_��
9o�(��O��| ,���J�Q�4��j�OL�:��4q��0��Mu�B� ,�jR�	L���
v�'<ٔMa��~�Ax��0�O�$����!$fv���KS�y�����n������ �MC��?!)�D�h�	�ON���O´p��R� tR���"Zb�MIE'N� ��mQ���>u���ö�͟ʧ���?�t�Dccp���jƍB&6�9��G�N��y��J�X�&�w��t���'2�"��'�X����͒�
1[���)[��'��)��1�$�P~��
`�w
8U��@�!��ٺ���!D/����R%�H�g������4�����=���(n	�l؄�Jf����O�� _�!���O����O��d�����?QrM�!lp2q���\�u=.�rOF��/��!��V�W����g�'��xsw�ۙ'� �
�IHI	�)��.�O!�폰 �HT���*����D�sڪ�5�B-T�X�LH�]M��׬92��'vў��']DX�Ϝ�f�����Zo�IJ
�'SvcSi�i"<���M�p����8��|�����ҕ#&��n�'UT�P(u"!�P �8*���'W"�'�R�X��r�'��*|R]���f�)�%�6��X"���'#{���p �j؞X�'C��+9�x[�oH�0I�p��f*Z�P%D,�
ۓi�A�	ğ�  Db�F@f�xR��B�t��]�'�$���O~�iU��~��̃+_7��(ڕ"OdlIR��Z�x<�dI�5k^���7O�lZϟ�'���	�L�~b����i�#�8�ڶ��_k�-��/ÃO�F��v�O��D�O4�
	 Y�b����Q�h��|����Q�b)���4��X�H�'��<��� �AӰᱶ ��'��⢋�S��j#��nx�Dy��ǎ�?���iNtc?�ֆ�;��TF%Q�!����w�e���	ex��Ӥ��gy \�w�P*�DM�&(�Ot�&��¡�$�|�����i�;}2[�ԇ�	#(B6e����Q>ΐ��εa�C�ɺP��ͣ4�֖zp��`����C�I[���%�9��t��h�5Y�C�)��۲C�p5��EOà@�C䉭>#4��A�: j8�
B�N}�C�i#��kf*��3=��05C�yfd��(}��;��S�BY
���~����-ǐ4!�!S�D^�#��@3]A��8�za��P�u3��Qi�$�ȓ*4�ĽSUN�<$~
��ȓj�h(ۥ%F6[��0I���vw�i�ȓ<������o�֩r���I��Ņȓ�8�A�C�T��}��#X1�%�ȓ+��Y��W�|���ڱf��ȓ	���E�h�<��Ǐ*,:�y��~�x}rA)��Ne�}r��1K(���hԀ�8�� gj^�y���*R����]kD�Ca��}o��ナ'3�݄�s���q�N�(T�F���҉
;D��ȓa�еH�i��E�$�SC�P�2x�����m�Q� .Z$z�� <|^���w*����T�%��tX��?*Ɛ�ȓj��`iѭҐos:�Ӕ��r�hH��S:�ਦ��/:W�����*ʍ��g��y����~l���c@n�ȓ�$��F����e��Ly���o�Լ��L�sn{#gN�90^��ȓq��4��16c�	[�O�����ȓ`�l�-�&���qͅ='$R���D1�� ΁#���J�Qd�m�ȓ-¦}*�!��r��N�<�~h��X?br�&(qn�a���.L���ȓ;̆���>QV��"�Ч>LZ��ȓ"[�ͨB�U&OU,8�)]$_w��ȓk�"����<�䂑e��E���ȓX�8v��qax�J��KN�p�ȓa��z����<��L�����v$Ɇh�*��0�VB�\�RC��J�\�rE��-b��!R��)pFC�ɭru�����X"v!�uP�g��HoC�I�?�}ؐ	��f��)8�>B�I�q�ސ`�[�N�h��HV� �X��[���#��(XxE�A���|V(�8��?\Oz0��(>�Xm5���@텬`ʊ;���-!�FXb�*Pl�Mg�j�'� �qOj��.�)�)�GG �) ��9}5��k@�X!���l����8m/y1t��լ��?!6�;�gy��Y*Q6��C��ܚ�h���y�kjG���b�S�01r0�K�&����/�O0��"#��ȴк7��A �'���꣗xR"PU��X0��	ze29�g���yb�E9\B������t��ē�����'�4�*���djҁn�ԡ�fiP5e��9�+޻�y�ɒ����@х_\�p���W=�y2�	/5d���N;M�~�a7iE��y
� ����h��>2��iA�Z�&e� "O�#�ȥ�x����>,FH�xU"O|�����+�r��Q�K-��"O�ȱ�CЀ*��|SҤƶ���a"O��c��R����aN;��I �"OVm�AO�9j��S#�"w���%"O���ӡ̆\�\�Ar�s^��"O  �ǎ�7j�Q���2hf���6"O��U��)\�Aa�/DAb=�5"O�ћ�L�	f��RS)�BP��s"O��z�.�=�ج;5.\/3(�-��"O�h@M�#d�؋�b��Đ�"O����`�34L��7�B�i�X�Q4"O�<Z�0]��-�b)��Qƌx�R�	�
�dٳ�yrhL��2ff(r0�T�"+��̃�'�`��K2�G�ǘ/�T�8*O`�@.��Yl������Z�i���_e��:ޑ�y�+�;b�1ʄ1U�:x�q�@�N� b�bG'0�'�֝���'��@N?�� 6��	�d���Gt� [�'�h���l�{t�� �*wH��cî	�N�O>��c¬��<�(��E΁A@�|*X�c��Tk̓x"H�!�'Lj����D�LUA�V/6��?E����@�^���xb��6M�5�C�د~�d0�Q��=2,lQԬI}<�ܨWDX�X�a�O�
����W�&��' q�Q�ao8p�3n�|���|mp��0>�F�YZ�i+��
��uЁzV�[Ƃ��Y���I'��'Q��BM<)�[9̪��e����0��_�'1�4�Ǥ�!ҖA�$B.JN�+�;g����i�"j�����2m���'xY*aL�47pĪ1*B�ZZht��'�(���+F��
��F�ۼM<,�2���Oɾ=���7,f���ӔX(���'��|�BB�]��%r夅�zڀ%��Cۧ?�$U�q3OZ���H���Ӗ.��O���ԍֶ����M�L�S�'�
�,�3=���:�^B�R=A���#�=�G�M�c��d"�$�34|�`��I�{��3tm��VI8�(G�>S�"?�p̈�+�|�H�IWR����ݦi�k�O� �L*�&���˝Fh<��3Y�������&���١�I_y�&BO��=P6n�f�8h��D��M�R �-'���'��|�F�0��f�<ɗ٨GK�p�d`[(d�1�uC�<ɐ�x�L'oF6�oZ&3n��+�8x1�!�"��/�@�86���P,䠚Z�� ��(�Ot�J��˦C�������O�0=a��C�ȅ����Ph���3f�p!:��L;����	4y�Xs���	z* ��j�XR�lcG22�������StTT��&61�!�"�Q9,�LhJ�F�@r@��A��f1\��4���#�¤kT� 9U��3D��x1j0�$T�&U^�W�[Ժ��_ ¥iP�?u�;~�lTC�jܷ��љcNS-��i�ȓ\bu��)��m
L�r��B��M�!�X�"	٤Č<wخ����Ժ#�͒��6(3'����	�.C�R�섻7��xN���V���9���N��d` hU
W�@]���۵ukؔ�p�N6fV�r��x�\Y��]�N��x&�~�B0	��Cr��җkQ	�O�,)�T2_<Ԅc���vd��'ǂR|�%��gL)0��f�@�qnY�T�����V��}��az9�)�5rA>�c ��>�`�0���P�Y!�@�|��9���� L��J'�-0�KW�8p~�Ro�u�<�#,��R��\ӤBŨ-�|�eK��xB�(���'ibĬ۰�ߎ;v�ͧ2ML}�"Nܚ��?�����N2�<L�Rڵe[���	�J>��)�/ ��x�F�Q������2pX�����a�����},N)��UOx�����E/l=кD�E�(1�ө9�f���5͘�>�=�s�4hP`��Cy���U%f֐zR�6+#��;�+0��x��;�y��D��썺�cȻI;��7o�5^(�����Ƙ������!^��x�����w�%���8UHH Ir��cn��'�2�:�¹)3��ģG<DZ�� #��sQ��ڰ�תj|��@R�]����ډM�~��|riI�{�����À&H@�Q����0>�F
�2Ĭe��(э�Mi�%�,�wf�?�P Vfߗq6\���B�1�&��ӓ7��3�bY0C�@	B'���.��-Ey�dĢo�~�0�nA #p�@#���n	�SrX���F6o���2�g�S��B�I�l?�Q{Ā2c�Έ��\=G���	�G��)0����[��q��(���/�1c�q
�OU��H� "O� �=;�ϯi�`I�$�UU~=��ȓ�~CRyW���������$J�pB��)wXl%s������M���7V�Z��dGm����P�� ,`|a����~�Ԗ��āȑoY��!F�L���O �AW�Z]8;�%8����p=h�BEU>T�rЮJI��C�?�v�����)�Rp��Fë�.�Iy�}�t#*�4����2�J\;���r���"C��{�)#�"O$�e
N4b�� D��I�.|y��PB}�:��I�r�����I% ����&(��~=���l��H��$WR� �h�c�Vd�((��'�Z]�@�V��F�h	�'RD�pC�A�\R��q�	5q���
�'g&]8�ɒ[X<%:a��Wt�	�'��@p�j� (��D1�� ;�iP	�'��q���Y�S� c��	2r�����'�:zSC@9w��٪���+d6���'0�88v]��@90g�b|qh�'�pl␭8u1�\	D�!T��5�	�'��R�K�D�L�J�Hz&z5�	�'V�@��$��;	8Ac��4l�ʨ[	�'e<1�%ES�x��\��h_g���H���м:�pc��3}R�Z	X�CF˰-dj��%��4�p?���Tktx�)�青-��u��O�>#�4�jT]����Z�J?�1�L�	�-֜�!Ď�/n�Q�8��&Z� ���?�K.�n��ņ��X��(R���@��㟔G��'2<�ǧ��(�զ�4j�]��'�T�@�iĪ���h����%
��M<Z��0�Ɉy0 ��'�pɛD�'H��I&l��*y��Q�Z�z�d5}rd�7��c�}���$�	{��9�
�
Uʪt��m=e��~�O��r4̱N�=D%�YM�ђ W1��'�4$����~�)R�:'��1o�� r�1'Ws�'�2%������O�2�3�)[�Q��QO݆�ء�(R;��'��>�ɐN�|���"��BR��baW�I���I�YT5�bf1�)�'y��Ј�"7����"<�@��	�l$�q���e�a���>,�X����*��'uH�����ا��O�\+�GP'�)��U�-r|�c�'W�����5�قE��\�g,ܷC��}r�Q�@��O�'NR����CMu� �#DdH�'��E~B��b�����@�pI�T�btBx��>5 ����s� ��ìU��H�/��m���gn/D��1��[�x�f@�������Se2D��脮J�T�4����w�����/D���7	�8fҠđ3bT�`d�l#�n D�4̉�&�p��ߥ
Qްy$�W|�<)¥_1\'���!mU�#�<�A'��u�<�U,:71+TE&As��C�I�y�8��T�p`��2�
�F֖C�Ɋ
\Ƙ[e�"��0t��73�C䉩	Y�ѻ�Ç�[�^� ��19X�C�	6X���ŏ�1f�8%��D�.0��C䉞}ԔY6ʕTc�Ӓ��}�8C�	�<)d����$�:�MJ�4>�C�I�
: ��$ɷM�jI
A+g��C�	�J<Ƀ#!X� ��Ql�C䉷@]�劕
01\P�䂃!:؀C�I�$y�	BSA�*3%p	`��̕]FVC�	g���$�ҔF�L��b�M�+�TC�ɘj�*����8Fްx�%��IWzC�Il_���l�06!��ڇ��A�C䉩U鞤�R�H5j}�T���]�C�	0>����O
�P-L��0FlǰC�	;B� �� ,�)4q���Sc�IO�C��iN ������DЀakJ�o��C䉅t�����V�`����@șX(�C��4\d8@K�B�mH�BΉ[{DB�)�  �)F�H&<�q�7���(2Pq�#"Oh<	�M:`�ځP�O	%)L��$"O.��s��F� ����*4/T�B"O�8��I�\�Q�9+\� �"ON	���L�b�8����c-q�"OЭ��eG56�\�����"'�d-��"O� ٱA��W% ������t�q"O}�f�OC��5�]��z+4"O��[��>Z��!C�Z�7:L\Yf"O(Tr�s�za��L�<]i�"O\4SP��1Q�pqWBX_\�
"O����C��>���P��SP�R�"O�HA�Y��~�J�K�=KL�+6"O~a(� 9pRtC%��~8J�p�"O4���e�⑓vkέ!�]ځ"O��w�\?o�U;�݇�\�x "O�=㱅ݦy5�H����(T��0`"O�UŅOo� ��>���x7"O��Q�dZ*��8Z���T|�ѳ�"Oh���-x����F�7_�84"O���ޭ0u�Ykr�R&7�YXf"O
�8 F#`k���"�@��"O��wĀ)H��%PDb�$�,��"ON��u�F�!T����cE�S#D=y�"O&��#�[�z�fM�`M�%~�(�"O
�3%fZt��Y`/�.@�	&"O\9�1$A�v�xs.��$X�"O��ٗm��9����Ġ[,��"O���+<�Mj�̐�O�t+4"O���8"CV��Ď�<_���4"O��7CJ�a��@E$P�c^�h;�"O��i�FI\���9c�KB$A�f"O�9��.��L�ɨƫ�[*a�2"O��˃d-_�F�ëY�KL<��"O����
*=}�8C�J�!#P��v"OV)P�g�.�������Q���"Oe��P�DGZq�#
�@�Dh�c"O�%1!NǕ
4(��5���t"O�u��/E�a4�pU��&S�hH�v"OĨ���7,���a�9g�~�˖"O.��g"@�Iq�LB�"%�2��$"OBH2�dȣ�u &��4~��I"Ot��bQ��0i��H.N7�'T�P�vO�>&��P2�S�U8��*O���c�
@!��:��6�ҙ�'����Ķ��Y���H�.L\��
�'T6���AH�d�lTˆ�GpaQ
�'� i��E�%r� ���-��~)r�'/<�Q�O�GZ�B�cG�1ݲ�)�'�J�i�+W/&���#���-�����'P2���I�|�3�--����'؝а�:
b�yctR�#�Px��'�M`��#Y�w�L8,�(}�N>I�2�a���	=h��yf�	�m�(L���pHR�ᙲ]nL��m�x�y��zV@-�@��j4�R)	�X��ȓ&`��V�U�(7*�aGnϗf�d�ȓOlb�BC��M��	�nG�L��y��E7ĸ�ai�4�t������T�B}�ȓj�b1H��� )�n_2s\,l���XaF ���kCmV�%��ȓ��!
��~aՋ�	�t��=�ȓ)�h8�e,�nn Z�CC�]v>�����u;wGB�={�hRQ�[g^�Շ�S�? �� ��1����a�I3/B5ڄ"O��i���U�|MB�	h�B�J�"O���ƞ�W�Z�Y�+��(��p�"O@�Ia�̻%=`u3�A�T��Ջ4"O\hY���2T����)@�lN�)yE"O��)�K^�TL�M��gҔKb�Tq�"OF(�%	>���"�X: Dn�+B"O����FٮBkX$Z�,� N蔠b"O��iš_�8����p�)E�و�"O�]	���i����P�b����0"O����#M�"�N�����^>�U��"O�f���f�j0z��">0��x�"O(���	;~�(��*�Ƅ�"O�a!��2���E
yF!��"O��13����㮛�`_��G"O����O��ѐo�?x�<�"O��4eةK���'��Kp�L�"OŻ/ٻ.��ձ�e�:R<�2"OV��e@y����EX�s�* �"OQ����T��I��[��V�y��'�Q�h�8�zT$ň&�F��N&D��;�B-`�B�j�4�#�#D���mʻ&�4M��c�4$$�!�� D�X��D=L���)�N<=Ն���K<D��2F �o�Xyp��K3pK����:D�����D�Z�1 1&���N&D����H��D��"V[|�إ�"D�d���<� �@S	8[l٢��#D�,��ɸ`�0����$k |f�!D��1��Y�``��:�Y�?D�0 ֆң&e��0&�˩v�0P�l<D��1�J[�&�< %	�l ƭ���9D���3&�,%2bu�qc:K�@K��)D����B	8Lv*��Q�h�,5D�,ʰ��3~�bMբEI� �G2D�"�%C^Җ��@�H�ZX;�C2D����
�8k���1��!|���+D�\Їgܾ'���	�/X����$c(D�\"��5J�0t�L*
J�x{�� D���T�^$�ِF�cE��i3�*D�$yV���%�xL�o� 6e����&'D�l�s�Kjl`��S��8KƔ���*%D�����V�Y�-E*~Z٪��>D�ص̏f^$5l�.�^�T/D�@j5eH�MH��P��]�J�Z�� D����*�vE&P��F %�����.=D��(�E�-8dGF�+�I��;D�t�c�77xE���@�(7��SPB9D�D���<��С�'��(=+��:D�X��F!��,��(ə�DJ*7D�İ�����²BSw�LЇ#D�쓱C���^'!WCF��$� D��P DP9�=�ԅm���s��?D�0�4�,m��S�Nl�~���;D����\,Z��:�=(v����:D�,q嫏	m�� aMF!�r��-D�0�R#�cv u�b��8rԂ���)'D�p�J��e� %*�-�5C�D����%lO���AmB� �T��[�6�ˢ�-D�t�d� D@6��D�e�8EO D�x�@D6r��!�i�<P�Q��#�O������$�&��3����ik�	�ȓ(T�{�jB����tj�-�^��H���B��l0� 0Ɓ�+��u��S�? ����NQ�:q�=�&"C�J��Aq��'����{��w�J$?*���-D� �W�,'hQ�0�Ԩf�Ґ Ǫ'D�̛@�-�|C&ћ���p��$D�8ʀ-�#4J�J`!�Z�j0W�>D�� �W�]G"X���X��@��=D��k�cǷ=:��Fb O���3�1D����J�&�R5���18��e<D�\�i�h(>�9��ܲ �1%�8D��{3	μ ��@��)"��:�7D�� �Ņ��l]!�,�F����3D�ʶ���H@��pZ�P�1D�� f��;���M�(	�x�%0D����ir��p Z!SQ�A��3D�,#���3���c��k�na
��.D�`7��=���ae�Z�M[���ň6D��97E��X�y5j̉sVdM�"*D��5K��BN�h%E(NZ`��4D�2T�S�L�ep�G])Y�8yB�1D��!������skU�P��e"D�|p�T�S�B�%�!�B{�?D�ظF��.U���r�x9��2D���Wѩ!9��hd7��p��/D�$�@�̢y����Ԩ�DkP\E,D��#"صI%l�x��JDA-D���/ �^/
	��XD�0�`��8D�P�D��5�2ᱴA�?|�¬��d5D�x�n��^�����K"�X��l1D��A40�"�E��xk��F%D�p��lQ>	O�Ə{�H,�6Ɠ�y�%͵ �HU�B�ۧ��Ǭ)�y�ɑ�7L��tb
#L��Ճ1�y2��#�^U��הE|"�<�y��0�Ba���P�l�
�J���yB��XF`�c�eƢe���q�:�y �T���ן-L���,�y�&�+ O���`+Q-P�bM�q���y�"R�E��ʕ���@���{�M�y�iΨRd��&i:$�nmK`V��y�ֿz-�ܡ�X�{�G޲�y�픅
'V%�Q� ��  a�%�y��¸ I��d� &�7o��yb× 4N5����"Z�x$�� Έ�Py2�E���Qu.Q�i�C�Q�<�R,�nmbcj^�!RHyv��c�<A1�*5��V&�#
��3"A^�<9����|$)fU�5W�!b�Y�<�T��N%t��B��6�ҏ�N�<����?�TaI���)W
D=��DQ�<�GBaz�a���V�0�f8v�ZJ�<a�D˥\Iۖ$�DAn�P�aAC�<Q3	.���5�v �R JH�<9�+_Re���$�!s�&x��n�<�!dȉh4�TdF#�bs��k�<i�m�1�I8e���R�xe򖄓@�<�v�%�,���#�����~�<��!zlm#� ~�n�x"�}�<�T�_�1� ���$�ŋ�Q�<��
���`CQ<p4��A�GL�<3���O�0dfE�L~�ɫ2��|�<� 3�,-�C��t���a�<� �α)�R4�m�z�q����]�<!׫�&,&�XB�=5���'�Y�<��,G��0⥋�
ar�7ɕ��y
� z����l[���aB�8G�Z4��"O��bJFFbU�/I�8N&x�g"ON���O��3���1P�J���f"Or��"#$�H�l:�H9u"O$�-	4>M�Q��
X4*�f�;�"OT@p��!��q�
*]L��B�"O�tx$�]�/r�b��O�
#�<��"O��g�'�<Q��&]ijJ(��"O8���A�jtq1oDK�,Ju"O਒�.:mb8`� ���1��٘�"O�!�#Ej��C�ES"����"O$1Q�,WZ��׃��QvZ��3"O�ř�(Ǻ"h�M0q�ķC��a�""Ot�� �23v�"a�N�i�(���"O�l��M�.�6a�G�ڡP��[�"O�Ш��ŷYֈ�2$�{cN�D"O�$�������É�)y���"O�!�dkO�)�������)hV��e"Ot��v�	j���Eem��Iۇ"O�8QC�E 	�eP��ܜZ[~�u"O���֧]� BV(~HT0sC"O��h"�2��؋��ư5D��;�"O��qj�82mJA���>z��"O��z�է1�(!C�aױs�@A�"O��;r	�
z�h�V"ӔG���"OP`��m�X�*�S'a ���"Or�2ub��HЪƃp.�� %"O���,M|�=�G.�/P��)�"OjH{d'��v�z�	AHӌw�%j�"OzQ$��A>~��p(�|�fmr�"O��:���$]�*XN��j���!�"O�c�;{9V���-_�e��i�"O����ɍ�_t�]�%���OH�ag"Of��Ǒ$ƶ]��eJ�SEZz0"O��1��&@vT�����>s�xH˧"O�E9�/��J�r�k��΁[� ��"O"�j!'Q�
"<c@��@���i�"O�Y�bM�nʩ�R��?Q?��hb"OU���_��+5�D�I\A3"O0\���Y�l�+V���%N��B"Ox�C�n����X�́pf|��"O��#�A�|U�q,ςg]��[�"O̴pr�D�X����$")pX�"O� +��+#�t=P���`?p(�"O^h����(a(�h��
K8�hr�"O�a����'cu�D� ���:E����"ODa;����3d ���T
O'.��A"O����B�4c��6�('$��2'"O\%�� Q@��	1"��Q"O����f�n�Jj��<\x!"O@��j�>���.Јl����Q"O�����3qrDhP���r-�d"Oj�zDX�%�J��&�͙f���2B"Obi1`O�H��K�I%%�� #"O�H����Z���Ti�4��!�"O���$D��Y ��[�Q��P�A"Oh��K�~���Sfܔ�~e��"O��b0`A(kz��@t$Ēn�=�$"Oh�`����z���L�Rn�ٲ*O������q�\��� #Q0My�'˪Y+S�ϋA-J؊f	
n��i �'P�d9Eᄢ�������mn��;�'O��9����L�
!*��g�L��	�'���:f�!^ʼq�NŅz�aq	��� �(���/���h��Y��X�*Oڨ��hF8a��+��	cH)�']b��Z�B�H��g��tRh9!
�'F��PPK�̌��7B=A 6 ��'9̅��ٳZ	(��w�D7JII�'A0�("��7H��0����7�b�s�'��#�	V���рWCC/,�d3�'���)��zF��v&˯x�dQ�'��+��A>X��D)�"��>�j��
�'���Ƅ�MöDܝ.�EKa"O�E�e�:wږ��"#%z��"O���%��X�Z�u�� 7"O>	��c�O%�#gԥ��YB"O���gȬ{������eU��`�"O��a&`ƣA�	�a��Y.���"O��§;���aT获m��� "OV�D�>���R�D�� ��$ B"Op��F��9*	rё�����6"O�A8@*O'/m��jD-ɊBZ��p"O*�D��@���1���=v �)�"O���C��B�:�TEB�ec��"O��`���V��9��Jj�x�"OсQ ˾UC%� 0��"O*��9q�]��ŉ���j�"O�$yD/W6{(M�c˟>�*��w"O����/B,���A!A�x�"O2H%d>���rV�;��$�"Oz�@���&n��
ġ6�4��"OX����ɑ���%H3({����"OfA��K-x5>�Ն5`	4�"O�A�V.2+�XcD���Q�P��"O�����Q�*oؼ���S� �~5Q0"O���%��IAtQ�&N�Mo��i�"O�T3#)H�o Zi���?hp $"O�y3-ܸ

��#B BIvp["O���5GQ���l���Ŧ4=P���"O����n�?g
����!�� :Blr"O\\�p���fe��G�0�+�"O^,p�_�B��c�?��!"Ob�SlL����xW��f+.�I�"O��0HB�@�K�Z�4�N�3"O����]�p"�ԃw"O=׀�D`�����R�̜a�"OrC鈼d�DY{B:6�`�k0"Op��A�*,vVQk�jW�zf0�"O@��B�Z=]�zU���2E��H�5"ONiU%^3'��]af�B&����"OR	ks"��8����Ei�p���"O&i6fH;g��Wg�1q�0X�"O�T��8r�m���f���"O�H��U�'CH��Goe^XXC�"O�0���p�����V�o#���A"O4M�S͉� ��U��Avf���B"O�expa�I�����g�"c"O�(C�͞�@b��2��6AL4��u"OrL��U'-׺a��OHl%�Q"O��ʷ�L�&"~m���Z�|>hV"OJ��R��	/;�@:A����'"O�3���?4���/�����"Ob�àOMߔ9��g
0�X��y"��e@I*^= ��0f��y"�U�5`�
���(dZ�IwD�y�N�;1l����IH�6�bi�5����yBiY �K�d�YTH@';a�Q��S�? \}�2�8DR����IuB	{�"O��1h�,@;^�A��L5^��Ȩ�"Oc�;@�,�B3ǌ2N�2X��"OT=;Q��l
&Y��O����F"O�d��%��,���d� �p�"Oz��`��
,jz��������ɧ"O���`N�u�LE��!�7��p��"O�e�НiƄ[U�	1d��ȋ�"Oּ���?=�*�B^� �&D '"O����z���A7�P�~��$Ӄ"O�3eĝ�hib'��z'>�jf"O�)�󅋦B�>�SR�ŨoT��"O��#E��j(U�u	G(p�T�i�"O��b0Z�C�t�R��,�.���"O ���?Qh�1$(�.ڄ�3�"O�  0b�G-�M��c��(c"O��#�IG���$ T$�)�� �"O,�p�uq�(�u���A��̹"O���4;�4U�f#(8�R���"OH(��%V�wj��኷h��`"Oؔ��b�a���z0ձ���Xc"Ox�1GX��H�AT��4�AH�"OT�8ģK'm�<�0�J+.�F� "O���Sb�':$@Tk�D˛F�MB7"OxM��BJ�t�����!��X�z��"O�-
��|�N���@V:L���g"OzXh�/h%����`�(|���˵"O4t*֡�cۂ��g�М"w���0"O�d
��"�R�ƙnG8,�"O��S��;a�1���3G8��ZA"O����O�T��(�'
�8Y#x1U"O�YRܒ�PX��5? �Ÿ�"Ot�s�J�Eޔ��I�/#���"O� kƍ�$�^�!�o�P�E�b�'��IB~�
n�����,
���g�X��y��'cUe����G�Ķ�y��9Y�ҝ�r�ɴP������.�y���!�Ҹ3�DЅ �8Q�d�1�y"�� ��h0 �/v�t8��/§�y�e�
�����kF�vll�����y芦m�T���/%�n,��@�:�y���ehĂ��Y.8WKA�y��0_F�c� ���$1Ri՟�y"� v�I���nga��nE<�y��6V>�I��";^�DLh�eI��y�)܌_�FE�2��Y�,��M5�y�m�J)J%Z��Q)2�&��*� ��Vd��z��xivj�"CNP�	t��������H�<D|;s�˰h���I��/D� `��׈7�>�J6'��P��(K�-D��3���6B�C�ɂ8h����,D��q�A)\�ؑ�hI;z=����*D��v 0ZR�z*Ǽr��[u�)D��%A�]��]�%�Q?ybf�J#�<A-OX���^�re�l%��X���3��':�!�H8�ܫ!�  �:ڤAE�H�!�$�Tg����Z�ޭ�e!]+,�!�D	�c�~ ��	�$8���?�!�ДY��b&� #�)4o��7�!�Dā~(�أ!kOY�����0�!��Ȁ"
TlC��ը(�(��k�;&�!�d/O�JA�0d]
T��K!ʐB��OJ��j6ʡ!Ɇ�_掼8�ɉq%!��{LqQፘ��x�%��J�!�� �m2�d	*n1����� 9��	7"O2��eKW�+�ř�
@��bŹ"O���qa��L���*���Z��p�"O4 b�IMH�Ȑ�D�m���"O��cč�hS�!c����L�zX��"O���Ф��k}�ia�#��@�Qh�"O��¨P�q��͛ �g�}�a"Of���,F;��x(�)�J�d�"�"O��B�@�;X��`�q�S(����"O����Ja���P�fЪ�!���)�!��&c�]P���
�Μ�HՒ)�!�$Ö/?�4Hg-G�`��ŉ3�<z�O���E*	[��A��*�jɩ�X&S�!�$s�f�d��!���Fk��!�d��W�8DPj�4 �����ꋱex!�dΧ$�2�3�bÒv��ze�ɪR>!���t�q�b��
z�8��f<&���>
�B��������@��y�.�H)<�ʆ
L���b�G�y�ˇB�J �.4��PH�D(�y��Y�xT�j�ag8tæ@/�y��͔{�l�w�7Hό<zV��yhgUb}��+mf��HU)��y��S���p�p��!Xe�J�y��	$��NWmqF�wd��yr��(�!B��Мc��%���S�y��-^�v���k8,��q1gⓏ�y��[�������8�<��&��yb�q�Ȁ�䋅��eb�ك�y2��"hlع6�ק	�
}�\��y�Еjk6��N<����y�H�?���ӍI.x-�"�D��y�"�8:��b2N	#q�
/��?	������(���)��%۷�O�R���f�����L]H�;c�A�h��Ѕȓup���� `�l� ��M�ه�Z��H@0��>���"�H�:Ǫ	�ȓB6�R�`ӱr�߬V��*
�'����5@������CA&=b��(�Il~/��������n�
H�o�7�y��5�>��gbÖ0�1BĘ��yh�"Md���䙴%p�t[��,�y2F]��,�A�*#y�P�����y��C�C:B��Ō�`�i��yj��`K�uB��ԔW5��`���&�y",K	�۱FP�E���"��yRH��H��t+B&&ݮ�����y/�)s��%CZ����ۣ���yba �L���x������R*L+�y1��wo���3��H/�y�d��~���kߟ
�����6�y��ʹLj9�F��4_-�←��yB�R4a�@��H�=V�9�����?9��$8�f��qI�ց6t�� ��#���'V9�f��4s��:���%�H�'�����T*Q/^�L�rM��'���HT�y=J��YN��dgFa�<����O�r�����rI4�z���`�<Q.ӯn�P�1ᇁV�L����Y�<d��(q�/��kZ�{4,�T�<�g̅ ^��t�C�75Ҙ���S�<A��,Ҫ�p �N�}���'e�W�<���M��E�b'��K@E�G�<�a�ٲg���q�9��#��E�<� N��L�_G"	jA�.m����"O�e�Q!K��Y���YM�i��"Oi�6�]e��93g���4<�{���%�S�	@>[�,�*B�&w\K�QR�Ia���b��ުKv�I&h�@
�ꡡ,D��`E^[6��ɏ��5g,D�@ҡ�K2/�h�kG�����3��.D�4��Zx=��+�͘�p�1KTe7D� Y�A�c>��@K���DA��7D���F�7a�����O�,kt\�4²<)�u��,�BO��,@.�ʅ	R�~�,9�?a���~�G#A����kU�~�&���bZj�<�曦#�����9sh���HB�<�5K�#qI�����&%Ι���B�<!$�I,��E	5�E�>��-1A���<ҋ��C0�Ά{��Q�	K~�<��#*2I�PDK9��CQ̊v�<)�AO+N��������afh�W�o�h�?�}Ra�6E­��ƥZupP҇k�<y�Db���6��2 ��D�;�y��8 &�4ؠ.~�&�9+� �y�ω7r�p�ֿ}�|��F���y���w��!�o�'{_�����y�.Xv2@y(c�Ř'��`���y�K��&3zq�gDS7j� �8�y"�Z�XCb�^�
�
@(���y��J&@~�:��T����l�"�y���n���˵-Y	lEh�����?Y�'�!��n]G�f���!�8�H��'�z�B�D]Bȹg��5>�=2�'1^U�ҁV�dz>�n�%���'�^%��,k�j%�fC�s6���'��!㠒+j_e����^����'�1�e�I01Sd��V��QM�!{	�'e I�vIZ���%�'.�At�tZ	�'�d�H+d~���G qWd�!���?�Qn�ػ���;�F4�C@�Ht��ȓ����	��8��mcPk��J�`!�ȓwC�JԂ�tN�Y�u�_ ^��D��R��!"�ڃu�,#���=�>���I��Ӥ���>G��(���;^�5�֯$ܪ�:֮]5J�E{R�OGn�[�l�)���#)�]���
�'�����>g6ؘs 䊸\n@<
�'V�غB��C,����R7T�������3ʄ1��n�2!��̜j^�'�R�|�Z>�'���"�Q��6��BQ���
�'C�4s��S4v.����d��p[	�'L�p��"-�����LF����' �myG�y����GMV#8� Q��'2�xk�Ɵ�R��I闇̕:6%h�'G�X�4|�j�X6K�o�XWL=D�0`��΂F#��Eɚ56��sd=|Oj��#?I�'I�n״QЇf$�P9	�D�t�<�g�e�D�
 �!�%�@�	o�<����.i��|2�BQ�]�:����m�<�W�ϋ[RD1R�M� [�νj'�hy��d�O�#|GC�5[:X���O(F<�*�P�<��V�^�6���ʙ�0���J�a�<Q@�4�p��Dgɮu��]Í�X�<qU-�i����b�%\���W�<yD��,% ����PFj���&�W�<���#,�y����u����aC]�<�DO'm~�)���K4)�Dir	\�<� ~�3��<p#���;g�Y!A"O�P�cMǜ(vD�v	ĎP�'1�	�G�b\��� 2�D�1QC�7XK8B�	w�8:�.��S},��b#Ʃ8 B�I.l�"E;ա�%ig �#я	���C�	�N�f�.���8���_���`�;D��禇�J�4��sj�1 @l��F&��~����[�4�I��ڙ�Ĉr!���B�I�c�81�+!�i#l�^I�C�>�DH�3@�5\���Ir!��| �C���Ur�^")��ש�&e�C�I�@x��F'R�>5�����pg~C�ia�k�a9��
7�Lx �)D���ˑ#c�x�D�T�E`s�1��0|��W�l��|�T��+v:���Fߟ���Ic���ƥ�:�RI(vB�.Vc�]�ȓ9Zm`S]j$hUQ�EDY/`Ї�bu ���](���w\�H*�ȓB~A�P�n�,�Q`K�t
ڨ��,i��8���t,(ҧJ��ȓ��Âg��H'��%F�5�Ƶ�ȓ��`s�6��P�^[����'(a~� G/e�D��>�$��g���y��۳&-tx2%�Q:gН��+���y�=WX~	���>pV0�q��;�y�	:��٨Wa�7�α�F��;�y�5V]��"FJ��<��u��CՃ�y҉$Y���@g��%��!�!�E�yB�ƞcb.8x���	���RT�B!�yBC)o�d0VA���|x%�1�y�H�6g�M�揊��ИB���y2�ު)�Hq+"C0K3��`�9�y��K�N�
Q��쟯u�`c��y�KF��2eW�x��õn�,�y�K�#��爉�P�e��j�<�y�(�'v��e뀕hr�ԤÌ�y�X�J�/ڄ.����Gֹ�y�B93T��Õ��"#S��1��yb�@�� �l#���AHʪ�y�w�%���5n�|B4���y��Ä� ��,�^��C�� ��>	�O�x�'�I�3��:!�w:fث$"O�h*���rhر�N"X*5�a"O�L(���XH��0���<Qp�v"O� �����O�@m��M��?��"O$�*�N33��J��K���P*�"OJMr�J�:��TKV�S���K�"Oڹ�g�!vF`��'KKn�
���"O�IY�e[�I�� ?=�y����#LO��Q�!�;� ���JU��Rukv"Ot��V�X�g�2�3F)�&K)ʌZ�"O�	k6�+e��`���/h�d "O�L8�EC)B��6hBY��i0"O�H�䋯E�>��M�9�4b"O�������1h@CT
~�0ܪ��'���+v�D�p�NC�C�$zG'1���=qç�hA1!Ɠ9����JһS6���0�$�"��<����-ž��ȓ&�h,(���j���)un�3_AT��ȓp2��#΁�uoѱ�)ϗV����ȓ�ؙ�׮�,�Z��b�i��0�ȓp7�$+�&�.A�`���ϋ�q�<��i��թƮN?}&dP`��!vE���i�>��g���b���M�}ܞ}��S�? ��H�EP�DXR9��j�6	�z,��"O�MK�l_�m�T͸�o�+ ؖ!�p"O�M�Մ[�v� �����':�Q�"O��fZt��(�c�69��)iF"O½qdO���hL��V�P�"O��HQk
6$OЉ��7�� @�V�<���9q4Pi/�0O1�xx��;H;
B�I0v)��U~���ԠW=oB�I�D�����Ԙ^=J�k��-Ig�C�Iee*�9Dl�0f���K�j�.B�I|���fC7J�&D�ǺM7LC�	�G+<�g�V�^M��*�أe�pB�	^�
�c�ų�d�i�l�$+SbB�9o5J��j�~l���ȫfNLB�	,�h�ңL��_F��8��A&B�I��h�i�ͅ'?�ʅQpEƺ[�C�	�uL�`������ܢw�� z��C�<���㘻���E�@ �C�8'�Nmi �����/�:v>�C�	�E��H�C?���@�Ć@����$&Kf&q�؉K��h��	tp>���b����Ȓ�
8�0ꃈ9k�ͅ��J����U�&&�HaV'��8��(��U��,��Z(վ��%�
��@��?l��x��ԘOmzܨ�wĄ�ȓ���ԀG9{zDa�G���@%&8�ȓ���3D�\7�m�t��5㞀��\��HO�D���A4��?7��ȓ/;HD�BD�<{N<eq��L^��ȓzӴes�F�a��*5��E�Q�ȓ`0�!GƄ9x=�R ĩxl��ȓE��(���65������4��a��z�6E�&��ni�����a�hY�ȓ-j�hs2���S���(p��$�	U���4-ϩ~_2%i�H�d"�mz�e#D�H�#CA�D��	pR��`��-0�j$D��a�(Zp�0��^�^��p�d!D�x���b< ���b\<؊�x��4D�8��B[	z�j�r�.��9�^�T(D������.P�:��L��D�j�o$D��*���2�Dh@�a�6�ضA-D����2�� 
A.&U
�!�&D�Њ��ͼMb$�$��4�b�/D��Y�J+Ruԁ1�Z-uz@���.D��g/цz+���� ��űr�.D�@���o,҉	�
I&$�81.D����R�9b��$��H@�9�O�I�8 .$K��ݺ4<H����2ش��0?I�*Ӆ1��WnًX��-���]u�<�D#�%9�
�z%��Ƥ*���p�<y�f��5& y��#K���1&�w�<���~���#PM<R8И�U �v�<�l�Y�¥	�#L�l�(Uq �v�<q2D�7I�Ls���m|֐)�J�X�<�V�T�sU���C��ig.0��ML�<�Ӂ <��ѣ*U)60�)�Q+WD�<�3.C�F���0!���j�Z� �hNY�<qGKF�AxH�d�2@�|-���U�<�FmR�j8���&(:eQ�u�4 P�<Q��A<�xB�Ց�D�5D�K�<�WC�<7lp�ը�*g�)��a�R������i���2Z>xق��:��	�<��'�`�f��&[�`]T����b�<�O��1�����M�fѺ�h�/�G�<� tJ��Orah !��Ή"(*�"�"O��r ��-3^t����&y�&D1�"O$�QlP�R蝓)G$0p�̂�"O��٦*�l���f�C�7^ܸiW"O*0
ǭE�r�,�b�?[􎐊!"O�l�5��?a<BYg�t�4L �P� ��ɐEF�ᲄ�?�ؘ�G"��!=.C�I�,,����*s��E��J��H�JC�ɸ8L&���&�k�R怚;S�C�=pl �#b݅�ڰ����I��C䉇/�1js�M�M���bܕg�C�I�N� 8�����a�ԡp�Z��C�ɑE ݙ��ԉ)�X��K,@pC�I;
f<�J�_�90�)dF�iW4C䉎Wҙ6%��O�5xP@L '�C��:��!���2? �B���;CJ�C��,e��(�����P���V��C��9&�Vs�E�/���2�BC���C�Ix6������10ԝ�T'_#;lH��F{J?19V �C$$̠ �Z-���!2D�t�K�(%P�L(�iD�v+�xA��=T�$�`�Z���j��\�$��R"O��K%N��`�(�ʅ�����"O�pU�ʠ ���aC�vrz�J�"O6�:$�|Ϯ�s`F�h��G"O2Xq�Ä�ZE� ��C �R��'iў"~�Q�� �P]KS����Q d�$�y��?26$��E)d:�(��"��y�M�:��U�G�]��X��)�y`|#��DOZV]�&
6�y"��.R��K�F P� 8�v���y���B8X�M 01=����Y�yR`FX3�qel -��k5��!�yb��B;�����|-�ء�Gʢ�y� ��C�LB�@�q������y��v�Y��.Q7uX�0�����y�E?�B�K�g�
�d��-���yr	�\m�����,+=�
Q�A�y9p^�)`!˾N�Ɲ��ƀ#�y��S�C�8kƥ&J66 ��g���x��C���X���F��ݸ���6�!��8Ux ��)�u72m��8i{ў��'�>��$�U2"b4H�'D�
� 1�F�.D�P'@��)�����,�C� D��zg�7|���4��R���R�9D�iwA� #+lDS���)4�H�g);D���R(ZE��`G)���ր9D� �C�*2�r003�
�KƱY&�$D��C"b� @�3E��B�1:�h$D�$r�N��Q3R�#N �OkZ	Ȑ`5D��Z�BH�p�p%-_2[�8-�e�3D�,�GK��n^I��AJ6P�8�;�D/D��:T�Y{����C���#%K.D�k�h]w�f����7C������O��=E����	WC�݀gG��ĠВ�]�[M!�䊁<"���T%��ސ��\5&�!򤃅TR���͸\$e8FK\�!�ě�{j6��'N�;����� ;P�!�$V�@؎���!�4':l�֥��!�!� |_l���'�QV�A��7�!��ͧ7 �)�"ζ_8([v��/,�!�䋟s��\���D9E0�	� ����!��|̸���F< A[�ʕ�|!��&�U���K)%�Pñ�P�|!�� �D	ĮV:�����B��)kv�q"O��Yi�(p�`=WÃ�Q�6"O�5P�n
�1���h	/YB�=:�"O�1��l�m3��+�ǉ_/.�e�	}�O!uI�㝖3�����"����'���蠬�4cxލ1�i�� �� ��'������΄�0�iaW�k�t�'�j�񐄒(;�۠��	�Np
�'�N�:��LJ�^�3f ��`�	
�'�HhWρ�
$�0', (�\,���d�O.�O��S�f�"�Ss�� 	a�IC�P��Ox�O��=��!7*��&b�7 �\0����:�y�@7MԆeq��&:p#4!��yb�܎,�噶�֖NO��# ��y⨉>q����E	R���K��/�y����	�@�!��ϥL����qC��yB��#}W�Z6&�L�.�ADm��y2!����餎Ⱥ9�X���J��䓲0>�Ǔ���NΝ_�<SՋNZ�<A��7��m����bT.͊�gGY��d�<!���
w�L9�\!��"��U�/̬B�	�d�2Q�|MV�xW�׀V�vB䉛7sP�:���*ȲW▧#�:B�	 &��E1�"�t�������>���)N�����A,W�ࢧLҦ!Y6���9�b`�-@$M��H!dH�Z:Їȓ	Иȷ��lv@|`����e�ʙ��`�'b��",�0|�8@���VB���'*p��Gi�W^|̀�/�H���'\DB���M�+aG�%��b*;D����kƗu#�1��Ҩ]�*墒,:����T��"��%�%r
2rz�7i�<����S�
$�P��N\�k�Ƅ�Ɓ�Sg�B�ɴq$�Ӕ��F��p2����<�*B�	;N��i��٣Nvz,���ڔP3 B�I\�H(�F��D��7��+6��C�	�=�\�&	YiDu[��XѲC�2m|�m�X��҂F�XGf����<D�����#�v�C��ɱ(��e,:D�I�l��WX��(ȡEml��
3D�,���t��U��:o�����<a����6�
��^�	'^�#'��0anFC�I#r���9$���Q�	5�C�	�%��XP�ɹs9j���A7�C��*Pl �$��Be�x�⛨dH,B�	+[`��k�6}��I���*=�h�$7ړ��Oz�E�ɖQe���.J��Uu"O�8���Љ ڀ���O b�Ԁ��"Ot� �XL����@ ��P "O 4�Q#�v(qAB@ �K����#"OXm���hbPۇ�)^����"O$��E�Ϳ>~44���!4��D�C"O��r4L�2B\d��؂msPe��"O�R��u������� �mj�"O���snĕ2l��eL� ��0Ւ|B�	d̓cHd�0�̚ ���C�K>
�fI��:���ę� j���k��<�ȓ�lt��G�/B�=�D�����s�2LS�)8,��E��"�r�<|���|�H�� !�n��f 0L� �ȓHĶl �'#��ܰ��$`u�9�ȓ~�H���
	㶭���w��̇ȓ�,�`RƑ��P��.C/%a��?�ӓ�.m����=w���� �;r!�u��S�? ����\GE�V�U�ʤ[C"O��N�`�R�8�j�\݌�
b"O�42�i�&^�BБ�� q�؉����O��d?�'p�z��V�'rlJu���HFp���IX~��C�Q��$����8�:������9�S�O�Mٲ��MJ4x�!�ڪN�Ĝ�
�'9�L���X*i�`�XQ��<b����'2j��霝T�x)���-�6���'!����_-6�x�	��"9� �@�'�0���T�A~z��o
�7_�e��r�)�$A0r���P��-4��r!���y�ɀ�_�P�9�
** Q3�]:��D4���'��#�(�)���	�#�ThR̃3"O��	���2�MY�"�\O�M��"O�{ӏ��T,��Q᜵k9���"O��c��	h]J�#�/Є7�qbV"O���#κI�2Ċ��ж,��������O�d+�( ���d^�vN!ɵ.�d��фȓ�:L(F�$;��9�BYYфȓx�m��>%���h��V�?\�ɄȓkF��a�~��΂N3��$BK�<)5Ȍ:G�`���'bR)⡁I�<!�;*Ͳ�[��P �tM���P�<)s䝼rH�9�e_�!� ��O
M�<IV�׽��-�� 6�|��l�H�<��ʘa:$�U�*�ɒn�E�<q�IRfp�d"b�T�v�D� ���wyB�'R�p�#�
T6��	��(��k�'G�@XЧ�%X�ar�Q�h���1�'vNH�E
�k�ll���˳b<M	�'@��en
6Y.\H V%1��"�'��35MFGrnܪ�a��x�D��'������҇m�^	�d��H�|�����̆)�~�*`�ňH{�;S�*�!�d�>|ıy�΋�)�� ��n�!��cP�M�W/�H��2!��BEF50�ǎM��8a�ƍ9�!��hn��y#�͙
��i��2�!�>�֬�#�F,D�z��FV,{�!�D��jPT��g��w��i#�*�!���Wݤ�xaԝT�4��ĬУS�!�ĉ�,ms)��,(��j��R�!���Q+v�}F�i�)"�!��>}�1!',�eI��e�!�d<m�̄��瞿^@�JJ!���ޤSc�[����j�>oN�O��$��6�ֱ �._�^L*�3��c?!���	^:2$ȲQ	h^�3�����Iiy2�'�����O6�0=��!�<���'�8U�""ގ���A�_y��yr�'���b�+I(�8���
(N b�'�t�*�S&��뇬ֻ�p��
�'1v�s�kĆH��,�G��U��{
��y(��O��c���[�}�-B��y,[�fE�Ls�e���ŉ�C���y�˖&nF�<����D�X�B� �yr �4"O���^{5��S
�y���]��9�+D.|���ѥǬ�y�#�c	�Qy�* �eA��K�H��y��ў$���I#n\\$4����8�y�˟7 ;����*[�N��������yb�	<g�@��L�������y�i�ϜD+�fC$JOR��S@���yB��Aؒ53bFXU�,鸧���y
� ړ���x)s)W	�vs�"O@q�.̨d�X�኎]�`��&"O��q�D2l��d H�x�|p�u�g>}��@	�&�i�&�̋-�����<9�q0�
��e����%�W�~>H@��;�e�2C�e��X�2��8d�Ć�Z,LѷjZ#w�����/����q<���b@f� ���̯�p`�ȓ���y�K�P�i�$B�/~i�E�ȓi�4��f�]�N��6�D�&�هȓW�`r��C!B�X�'�W�`�VT�'�ў�|�
B�מl�`��"Tn!Z��U�<qp-�:/��1P�_�F�6�yb%L�<�ǔ���eh4���#��w͞F�<G��}�B��3d.a�
���E�I�<��K�T�J�s�ʀ2{a<�4�A�<9� �:Y���۠�@/d�mj�'�{�<��+Ə|��\@�+M��4pS�w���0=	�ѡq�b��P�1�P�3��q�<�f��&1��t����G��Pk�o�k�<�b%�~��)�(�\hiG�B�<i%ԥN^�Es�Ɯb�x{�CT~�<�qK��H{��h�����,3B`�<ٳ)�8�4��d�HͲ�:R@N[���hO�|Ǵ-*��^�D�3�(<E�u%�8E{��T�)fnؘ��)�������ρ��y"%ܫ覨�D*�,&�!
r��5�y҇S��0�D��S?�H���=�y� �1!8M�q�L,]nY��W��y2n;j  �z���_��x��jN9�y��R�cǲI�bܻV.������hO@��	C&"u��1���(��� ����O�!򤎚�t���Z�N|�%{Ѯ�o�!�߿jh��cd)V�9�hP�n�!P�!��B�#7\�a'	��Mlq�b�$�!�"1��D�QR
m9�aA�!�$D��9���O.@dS Qw!���8�x�*_1��$��i!���%�|� WB�v!�U�__!�D(Ml�F�'�<�`/KpE!�� �Q���B�L�-ez�R���/1!��Ϲ\��Xw/�96~���f�#g!!��9a�"US3���p�J0Y�!�DB����Ս�:)���悔�M!�� �jp��D��,��ሙt�!��2U�J`�g����JL���C4�!��?	F�qb둌/�����M��C�!�ċ�����l]�j���"� F�!��h
9rѮV.�����N܎a�!�P-D�90��\�q���Em��7�!򄕊
-ؕ"�gJ�{��p�b�V<�!�$�d�@��A��Q��ө�!�$�	A�hD�0�-P}�%�c��n!򤄵'?�}âh5����Ǝ�w�!�d��|΀�A�F�E����� �`!�$C=Xl���2���s��Ҫ]�!�$�@2`��	R&��lb,��|�!�d[?)]�3�\�_�h���Ӂ1�!��1u��:cۺ-ʃ`0N̕��/.�Q� �G<z>�:�(�)���*V4�QiL+C���3�G�tH��ȓh�D)y�� $�k��[�R�D�ȓǌ�s0䓢�����aX�Qq:B�	�l����R�
�WF-y�§TW�C�)� ~�(��� �N���փk�^��#"O��3S!+����o�;Y2��"O $�H�}`�<	� M� �$(""O@�B�@�A/�Q�#o�d (b "OXX�Р���� "��/��b"O\� �Ȝc��I�Ai#��th�"O�H��H��kTftYD猾�N	��"O�y��)�)Y�N5B�
�[�� v"O\$S���+<�jP��%�2c�x�#"O �Q��C�g0�|c���@��̰�"O���VM4?fLӒd�3p�JY�%"OTt����2n�����BL�1#"OaX�c�!M��IR�6lc0�H!"O��8�������͋ZLFԚ"O>�y�ˁ�=� �/�QKH`s�"O�}sVj��Hc��XS-b:Դ��"OR賵͈c��)s��	�PA"O������h䀥���g����"Ol��.���D)Bȓ1�<3�"Orx��*T1�L���� 5��`�V"OQ��N۫;@�"s��;�
%�D"O�I�w��+td�	�@M�	�l�d"O`	�(���u��	�!�X�d"Ot�cU$�� 2՘q�ֺxk<�Q"O΍H3�_�<��Ǝ�*P��u"O���w�7T�k'T.m�`<z�"O.�k� �+D\Ҩ���2J��<0"O,#ä� ]�L"�&��3p�a�D"O���3
H�\��e�?��I�"O<�d ݔv.���B�%)
�e-�!�D]�6C���f�F(�c�"E�!�DP4B}"�Z��"(���&r�!�ڵ?�t��aĠ+\2��^ ?�!��T)
ұ���25F�C��l!��<�X�b���'VA�magjԔ|+!��D�x� �04�d�T��H!�/T[�e�"�I�{��k�Ƌ�!�䙮'�5c�L.1j�!!)T�Z!�D�1at� �S��� �'߃)<!�Yo��c�УN��	P��A�U6!�Dӻ>����C�],�$s��Ѽ{!���&.Ff���Ћ"��{�E)>�!�$�x���"	��a�M#�!�$33�K ��%9�b��b���ux!�d�S��@�_9 ��Y� '�':�!�D��F�,(�ćڳ.��p1G�4I�!�$>-�,��wkH�D~��gg#!�d��������0���Q'�N7!�d�Y�6UY�/��(�(����m!�N� ��3��lPS�e�4�!��ʩRC(��i�)kj�h��?Z�!�u���w&R� Sz%��\��!�ȗ-b��J"��%#B�	2�ޘ:�!�$ �d\ճf!�n-<�r"��-B !�V0i�Z�Q�E$r�RDtF9y!�ڤ8�q{P뚾c��ڠ"]�.!�dؔHb�L�! [�$�Y�Ӧ4�!�XW	�4�M�"� �#��hK!򄒲]��tu�)v�veң��4.!򤒥n��`�W�Mh���a8!��4����r��6��4���&-!�d�#h��s�M�� 8F�7J�!���oĺ�`�*͝J�Ѐ��e��0�!�P�&�Rɝ�F��LJ�dʹg�!�� A���_'N���pQ��/Dh�{�"O���,�?}2�sTL�W?ƹ�g"O�*R�ɓ-�2Ѳk�1
��"O6�h#nO�@��A�Jʹ-=��U"O|� 0�I(:*�������v"O��KP)�L����hC|r!��"O�TWޠ��pnL6\�Е�'"Oxx��L�}BR�ʕM�mel�1"O�([5�S�-�H@G�˛3��Q��"OE��bJ�c�(d1�]�^؝"O"�v��Vf�� *<[2��'"O��P��)�x�x�(�b��"O��� �:%e��Ɯ�N�`��"OB�d�*������?Mo����"O��bghחI�Ҽ�T��'jV�{t"O*�1�L_�U� �,,(���e"O\���oU��1�%��A��m��"O�x�.S�e}���m�3$|F�y�"O��Q�H�\;�`s�b��z?�j�"O�uC��տ|��y���216^�q"O���a��vt��+�˭`/@�"OT����8}��u�����B"O2��T��11�ᓱFǡZ�����"ORQc�eM����eǼVE�w"O�%� �ѡ[A"`ٷ�C�?��p�"O��`��֛�Jк0�	�W��uH�"O�B� Ѡ
cdK��A
N�"���"O�@ir+$��eE[ Itt!��"Od)���I$`�� ��YuZN���"O�ɨ1��-�������j�0"O����i	0 
� ��ǭgՒ��"O$\r�c==�q���^�:p�"Op��!Y�(V,���=T�x`PB"O|�CdP~	Bq:P�ڳB�h}�"On�X�Z�U;Z�O�S|�L3T"O�<��>�2��w�0J{~i�%"O�A���6,��OAi��%"Ob0�(l�|�򌐾/��l�s"O:E۲B�Lf�٦L��L�ĘSt"O�E`��'LBys֪I���"OR��$�T!K��P"�X�I|\�(B"O�|br��&�Ub�W�_�H��"O����K�v�h,��
�>N�k�"O6q�Ȏ'�0�{i��L�\I�"O�!!��p;�����j�����"O8y8��� ��P��K�O l\y�"OF9��͆._L��F�ݳj+8|�"O�����6~�D�3r�Ձ�D��"OJw���{?ha�QNߜ�� Jb"O�h���~��]c4�G����"O���k߆%���qn��z�d��"O�]y#�ӥ"T��:r�Y�M�}� "O����Pfh��WD�3n΁�A"Oj�t�B�E��z�K�;S�x�a"OZz1�
�a!���d���zd��V"O��Cq�f\�hҢ��N#��ѳ"O� �W��9inJmz1�E�,xau"O��� )[?8����,f�Q�"O�����5|t(J1�XA��)��"O��hP���
E��� /^ hɴ�� "O�� ��_)}VH��@炅:�Tpr"O��"��8�� �2L̸k�X�pW"O��qAF�z�hH��kB� �r��b"OF��BeėOa����~hz}Aw"O� �ɰ ��s3n H���!4|uxa"O��Q���+�2H��#�`+�C��!lO&p#@H>�@�����
��5"OR	
��_;|Y�`�
K�bȫ"OZ�	�e�7|˼�8� 2�<��"O��Sf�#B�D-Y�c�$g��l{b"O^A�� ��N��v���"O:!��͓]©
�i�H�:�kr"O�u0w$	����H&	Ǝ}���#"OJ���0 
�ڇ.�rزܸS
Oj6�]��Ph*�̉Č�5!�Ė�WPN�)Eo
���'��:�����k�KϢ,z���Ov�U�`��"�d�ȓQ��܉#F餈���7q߈��'H��(�)ʧ_iv���E�]u,��ٴ �\p��C ��83ʇP�$I@��-O�*�Gy��' dU��tر��Q
O`���'pBy&�.#U�U��/�fn��7O��A��q����x#�� #"O�䳧nC"x�H1�a��.H����P"O� u @�N��T�ghH':�h)0 "O��P�K%����E	F�Zp��"OZ�K$ �:v�ֹ�3�܀|��I�u"O�u���ه/*񰍄?�J��"O��c�HG�OX�E�$-�,Ey�u�P"O�t���K���8��дbK}
�"O��!cF[�w�N ��P�e+���"O�㢃�)Y��P�dO	2t��"O������~
�UB&)�XV��"O���2X(���W�aR(����"4�t���F�bW�1�'$ؾzD��I�"D���Ӂ	6l�`�H�o�H��ؘ !D��zAQ�g�l�rt�>e�li��f>D�|1Wg�j�5Z���T��IxR<D�  NN���X!��ޑj+�-qs�%?!	�]�>��w	�	 �u��&Қ`x���>�˓�M��Ō 1}�� ����e���ƌR?i���l��Y�A����O'knB�c�"O U`B	$G^��"��vV���3"Oy��L�Fޒm�K�����#R��G{��鏠p1�m� �ճ]��B'Y���I�<	�}���ʋ%{
hF�*]�`���Q�H��I�eGx����w����$ޙ+d����*�0���>Oz���5P��h����Y�"OP����
�0K��9��1JĿiʡ�$�L:�S�˒|��q  ����y"D�+
����a�
s
�
��'���'�1Oq� �Z��!�P�#�
����CW�D�O&ʓ1�>i��J-3J
 �jS�<
�`��B[��yȆ�g �i�KV�&d�%3P��
q�������%��O4� Ť =���7Ċ� � ���"O�)��E�K���xfM�C޾��D_��oZ�g1Q���>�+��W:ʭ�`'Ǎ2?�1#rNoX�4�O����(0��@ԋ`�V� ���a�A2�MB%��'�ɪv�؅�d֬�,d�$�ѫ0�C�I>�za�tAصB������<�7m5��:\O���S˪���B@<.x�h.��'�ў����W���Mj�ũSA�>Ĕ���"O�t�_3}(�I��!r���iPT�ĕ'�2�(�3��a"��Dn\��H��h\!!�0��k�矶\��s���:Se�'��O=LOT�c6G��4Kv�-z�\@�O<y�ÏY��n� H�$�$`��n�K�<��UZ)"�D� DV�*��B�'S���"�g�? ��8���No��35I\*,�9��"O�l�a�Ķ�<��ڬ!��Y�@�|�0�S�'+(>�:�,��\ФP+�i�;�nh�ȓ$�.)��ꈵAܔ�G�N�>��=�>�ד'�r͐�f�$�{����y4"��ȓ}��M�S�ڀ�xY+SI'C�t0�'F0��/�9��P.�H:����{�)��J��PTJuÓ,?��=�W�L2	�!�$GU����n��.���(���!��R(��������E�r�3�̋�!�Z�c�ZXuK�3qtЈ(�#���Dx��'��H{�.� ohL��l�)��+�'����V��/?�����Q���
�'O�=�5��0��8s��T�c=*	�
�'�xxIC�D
]��5Y�i��P	"
�'#:� #냠H�T��8s���'M> ����?\����	�p P�"Ú0|�����*�d�+C�܁���zG�����ݍ<�!��z u‭[�;=>�Qs]�!�!��o�8!����`�P(�&�;B�!�[V���f�F�|!҂@г:y!��J�E�Kc�#ⴣ0oT�pg!���,[�=ٴDҁ. ��Ѭ}:�'V�6�'vL�!j�`�~(XPr�4��	�'ۛV@�R�����wlp%HV�)�yR�My��8���C#w]�H��/��x�lӱYd$���37�@��	.k!�*DZ9��
�Ɛ��w������m��(�:�r��E3^� Q6&�K�*aI�"O�ʂ�
�j4(�"���-JU"O⤳�� �g��BG�x�; "OB�"#��{�9�U���`���aD"O�آtK��9�f� ��6	4��م"Of%�.��=����"�V ~�ބsb"O��u)�1P%j�
��B=@~��$"O��X�c��'����4C˺4D��H74��ZPF��Cc�r�AD�bۖY�D+�$�S�',]��� ޚ#�y��ش@��0�ȓ{���w.عp'�8�5�J�gB�5&�,�'��x���-�d���*|\xX��F���?�'�����#]�$�y�v�_,/=쀛�'�n�/V�X�����Iݿ8��ᨍ�$7��]�I��"k�(��kH�^��9��e�?(�!�_����ⴍ�2z�b���E�I��'���z���)�'9Ԁq��
#��'B-�!�Yn��I�$d��PհĀL��	_y�)�mM��h8#P�LFXY�L,��O^@���OΈ
�'�w%�=F��J
0����;O���㍣a�� /P�wu�Pbp�'�'[J9�*�?&=�V&L�+��19���xR)�E.&��զ�(sz���r�����y��)�Tȹ�eIF���b�������<�Zu8�Hۡ�2�l}� ��&�!�Dү*��́�o��t�`Љ	�S[a~R\���i�3 ��ɓ�	�#b��Q�c�)��p<�� Na.1���.W���pqJP�'7�?+��M�c�쁢(<L�*D�<b6&��JH@�Ҟ�]��C����t���iω9"��$���L� J��D(Y!��q���:5�.:[.�)F�y0��$�������b#�����i�!	�F���l��
�Y���ZNڤ@�!\�E�ȓl����#��|���ٶ���'���G|"�ӑ
E��T &�����%�9H" B�)� ���6=,=������4>O��=E��D�$�v쳶�4l<� K���y")S:Ԡ
A��
a7F��e;�y�@�.M ���GH�g�B	ӥ�yr��8��:g��Y�n����\�yӓs'd�r�e��OK�!!�*�y"�A?ct�`��B(�|7$�*�y�_��� ��I�����y�#��Ēd��I8��$��y�H�	a����^�j�:����y�@�Y���3	ͮ�TI��:�y��Ky���L. YCd��y�iߨp�yJŭ�0�d��'j�7�y��C.�ʶd7����N�-�ybo *��)���>:h�ʡʛ��yrgƄ*��|˵��L���� 
K�y��x������<4P�d�pf��y2��c!�`��!�8wR����y�.��q3�/:����bȽ�y�GU�K���T+\�*���2"��yR�ȶj��x�`Ӧ /:9���)�y��m�� ѓBU�Ј-���1�y2$��S�B��Lq4lK��y"��;�~�����&�����-Z��y�&�=�lb1��?`]��̆�y҉��@n0z���5�YBP(ú�yR�
,MN|XRdd
9 ʮ�s���y��1X���j�)��"����t�D��y"C�,�L [&W6�X��W	8�y�3�D|{�J���=�r���y��B(�$��f+V�1�X!D���Py��R>����1*\]�'.�J�<�H9�jLr�6�d�֤�F�<�#Z1��ˣmG�QڤH���|�<�u���O̠�2�8�6� �y�<A�b�0��){�ѳuv���b�t�<	U@\-. D�D�/�"B��<�⃧MK@Ūq أ%��eq���n�'������P�@,�Վ�8V4�:�'~��T�� $(sE�K�>�` 
�'��dk�o�����#��A�6쩂	�'�����eڼH�$�D(/=8�[�'�r�q��?TX4	������9�'�FQ�6��:Yx�L�d�S��PX�'kf�2��Ǡ?{~L9t,���<��'o�a�Lu
D��P�S�f-8E��'�x�l�ec������S��}a�',0���%A�bfɘ���+��'��\ 1����BI�@-ӤQ�!��	x+�iKr��&�P�0k@:�!�䞭C�L���H��;S
Q�~�!�$)�XP�d
U��Q[��Z�#�!���&�LC&GǓU�(��Y�|�!�d��XZ&�c��3T������$W�!�D��%�̤�rK��{)h���e�!�d�:5N���� �07��9�2K\8J!�䘰	�	�i
#Zj����X>!�$<Q��liBcS�r&�-�b�	�5!��*-Q�����UJ9�R��!�S�K�"�yрM*Je<=뵧�c�!�d��ZZ�=���֬s@NA�����!�
)���!� 1o� `�C+�!�$]���8X�k��T,� A^�!�L��FPI'j��)�0�"�4'D!�͢�&�
�`X�0��@r毚q?!�� ���fҷ*���6d\H�:�"O,�˒��B���E�\�"'���"O��#�3I.��[�c��J�a�v�<���ˊV'45�0�!eȵk@K�n�<�P�C=}��hK�OA�,W�o�<� ��|�±��@B�j�*��C�<�T ��Υ`5牻!U�r�GH<�=���
����Y��\��9���+�O�PC�l	�)Gɓ2��!!R�����'��It�ʩO��'X�H��J<K�R�)Ԏ6%�r Y�'�^�����E���:ԯV&��(��OH�,OBqYH�"|��J��L%apK�d P��O]�<�C�
�n
n��g�S�1�"@Rw�C?��'a]�����Ϙ'����H8�\i�jE"�x�8�'��X���4��m���=���r�A΂u��`��\v���z0��g�D0�Al)6}�U�'O�,��dyf\iH��3�nŴ\8(��ƬΗg�=R�!D�D8 -KE��E���*7�4WC5?���H|Yv�Qr�&}���Q�t�ĥ�=&����2Qb!�]�s�(����V$2Gb}�5oX�M1�*O��҄+�3�vb>c� �Mϖx�4y��EÉK���"�!�(1���9��������C� ����QhH��
H;��~���6d�q�Mz���h#h^*�0<���ӌ^g��[o&}"��00\�v�N�i�^����y��1I�V]rK���5�䪁���'>aS�iՃ��)§B���􎓚f�F84�q�H0��8rUx��<�8es��1����3�|©��3����}&��S�G#j,9`�.�<���
p")$���1��KK�	�p�Q�H@��I@�!�@���'T��3uf� %�����n�`�Ă�'Ɣ�� .��BdK�3hm����'�ba)A�I�Ya��	3gߧ7+�m�	�'j2��ؒ?�u�-��(�l��	�'l����3�b�
w'�&ebA��'N��X�B�#%kZx!W/3$_XL������Z q����6i��|{H�3��Y�ݚ`c!��ƀU�<�D$6`����G�G,¨��NAp��|���Q��`K&�ː:��1�!�,��C䉳%p��KXr�v�{�� �:�_� ���c]�&v:��$Q���l��|#�(j��D"Ta}�䑈@4�,c@�A�Oi��x�3�ൣ�bC-ѥ�(4�x��� ���yD�Q�C����W/$ғ{$2́��Q<��6�щB������v$�a͟�ΠPH�N%O�u�"O�쩄E���A��'���ys�i�ڼ8W!7-y�� �ճ<j$X�C�s��Iѧ�fd���,��#D�Lh�._�}xH�KQ���|P	!LAE��������Сk���'=!�$zVA�/���H��DDmN�:\h���Q��u)TLZ�2 �!!�n7�0Z�lb<��嬃��`��c�,��)G�|ܽzq"0[vT���~�v���]�e�(�EgӘ�cp/R�69��o��?��\��!۲�ywJ@�&��=��g	�:�Ҥ1tHU�y��_�Gsv<J�#Ȥ ��1#%�l���[D'F 4�D0��2] �&-�Frr,b��%��s���ywHg�> ���R8"�)��MU'�{b`�A��(aP}�(|�@�[����)�x怱� !
��}x�κ��i�G.�&`�����[�DW|S|��cI$ֆ��+"�I�Z�nmb�=��@S�J:�	�EJv/��*���D���-��l�2P����#�W'�l��VF?�O4��"�*mF��"N�5L�&��q+�Đ���2/�h����:�6������uw��9�>��Ď��[th_#IW����|_�@��j�_�<�6��8*l4�¢�!yR��F/̙jq���B�G�. >-���"k�ܔ��;��"i�ր�]� ��-�@���j��ABНRe ��ə#�I�Fэ����#�i�"@�Q���5. kp@5� ��59��l��d9���b�2.�,{�&�::U�O��b��K>)z���S5`P0IN|
�/�)0N�FX�n�t���o�S�<��ŀ05���8F Ί+����*��?[ kc�`찀R-L�[�lG��'f<����]�z�C`���d��,k	��� ���!���%�A'v��|��!�O2�	@�٬]�`J�
�l�?i�k?"Kvع���:f4����/�f�4�!F=�>-��a�j��-� �è�+��-ԡ��H;���t a�M��{vD��=�ɝQB��P�O�g ��eF���OM6�Ѡ_"HO����I��H���	�'�����O.Y�
�Kc	�0�h�XV@�L���(��2\��ӭ�(�剎w$��A�\F��פ� 2�(C��9K$�0vLT<��(���Xl��t�A�a�H�{q�	�H���xх�y�'�Z��@ǎy}�E�P�Qd����	�>�$A �H�A��� �G6&�(+0m({��U�X)'2��2�ͳ�a"�P:c������
S����䏝Ҙ�5AN<~X!{4�ٲ:���T2��'I��<`�@ٜ<T����m�)��%��O���SӅX�:��$�EPd�����O��0V�����H�wVy���{�'"���H��v���OB�Y`¬Z81�Ɠtc����ՌC
xJ�l�'�zE�U恻_%L���$�$�DQ��(֖[`"?9`�K+>���{eL }W���VBx��c%��y]��� Wl���q���d�+� �']@�@��E�H�`�'���aO�oM�@*����h�:H>!�A���|�Z �I<�` �v��1(�V%�v��x�*�b5
˔51�"Oz�s2O�+�D��H��N�U�åF�"�N�:�/E�����$9[��5��O2Q �6-��JcHèM��x�O޵Z��%t�PYa���	
�~�*!/ث�|y
�l� ���/,���F���F t���̷���YF����<��������-�^��Ĭ��>$v�"�kE�#b�bJ�&< ����*�:���N�~�z}&��%�,�<	+E�&���L�x%���7�S�H�F<��F'0�X�yF�M�0D�B�I"	~*�Dˁ�+@t�A�V�2	0����E��R�u_h�8��!�g~2/)��p���]qN�8���:�y��D�'xF���i_d6Ԁ��lI�V�L�[�ǔ8;���q�Iʔ��dX�Г��Fi��lA�"N4;7�z��$4_��Cm�cmJ���?k�~DЍ����w$U�;|�'��Wdm����$_�~�[�q,�XGi4�IG:�]:U�L&	�zy�ş�&L�	l(Z��ȸ�� vb�& � 9��`������KJ����
�m�T)�P-N�MΤY�Ą*>�$Ӧ�
��6�O	��eGg�ԭ��y�!V�VPH�ED��Q.���#�7�y��R�A:��%�Κc�<� ��
�*��I�XG�a&��	����R�RG�1D�\ 0�P�����6kr� �ጡx/�X&"�Oൈ' �`~��f�F�6��9�T`L��|��O�3u�b8Q����?���A�h�ki&�au�p3!��'�d�g�6D$Gx�!�	f��0�vtG�x��ϙ�ZfL�h��ţ2��2/L*y#��]&_f�� �߾)&���đ`k�x��ҍ�8@��i��}]1�FN�~t*�P���]��u��Oi�d��gӎ�2H��O�NLr7�Hb��=��< �	�2h�a~��4j`ޔ���Y�y�b<ԇ�8M�Ӱ@
3����g�ƱEs`��3$��[���?It��;I����0�y�o/x��y7GSZ��H�v��?�hO�������Co���־.X�m�G,��R�W�%�n�)�++D6�Yꀂ�+pd)b��O@�jcX$/Ơ2' �b�'��A�$G�H�\��tcȆt�h�ڴh���s)��l6m]��4r���w,�"E�ҏ"��� `�8y#�K,2�3M�+�MK�
6F�x񤢓Qx�p�"�aJ.p#�ɱaYv�;��K6.X�q&� 2ʆ,c��8A���0%��!�$X0,���5Ot��daÍ|�C(A8�&�U�'r�Q��*��6�&d����"f�bfP)�b�9����;(~9�Q!�)l ��R�t��Y��)TJ�Y`ġ��',z=i��� WRD�x�BD�^����� ����	A��*�Ms���]�����6��<z�@^�A��ı��9H�b�B��"T��r���hE�ՙF�">��1}�U+Ea�l���}�؀��FA�I�̴z�m׼�S@G͹�h�$��,Y1m��c©۪�8qQ�R�V=K�F-�O�-1a�Hl�� k�P�(�Ը�se�Ď���(�3k���m��'E~��93�gj前f֞�8�͝tl�x 5�%l��DL�/,DĈ�lZ3��W���?j�����"t 8�O�ܠ��\EO�XP��Sm�:���܉�h0��Q!,�=����2��(8���W %���^�T$��	��}7r��q 0}lN�`b?OD�q�%�4kP5�ua���aA8O�E��Aճݸ�h������ܞP,<	��ϭn`�s�$C�=~��)��3�Oܤ����Y ܒ��J X��Ѧ�'j��ce@C�$�\�V�asj��1T�Hp��C�0�!�؎/�Ze��16���l@"bW!�� 0����_�)62i��h$-�L�r"Ot�9��C~�!l@a�"O���UjH#pa��I�"^,�;�"O��ZW@��|eJ�"�/:��piw"Oؔa��L�,N�T����-�p�B"O�W�lx*f��e��B�f�<Y�a�,&�;�Լ.�`]�N�\�<�ū
,�	a��8
H���a�P�<���ϓ
���۸+�nm��N�<�t!��ˡQ�����$E�<ɵ�ƿ3Ј�"S�E�;P����@�<AQi͎S��"� ��F�YP�K~�<� ��gg�y���;o�T��CV�<��&܈jզ���ҽ,u���A�Q�<���PO0Ɉ�K� {`1�b�D�<y��i�R��2�XPe95b�D�<QI!�Z�qk&����]�<���4iԐ����}��d�Y�<y�+A?/�yh��A�����D�~�<���I�a��lQ��RT�����<��,	.6?<�c�Ҭu�,����C�<��&D�r�����c�0$�V�w�<9�a�`Eۄ��2��`�OAX�<�J$vGv铒E˘v�	Kg�|�<Y!�[$���&�+�^�b��`�<���T�g�B](dХ5zn�Hv��w�<�7G������!�Fi��� t�<�����>�(aDZ� p`�@���h�<��
�WDR	�F��"}vEp���<i��:����d�\�va`M�m�<��I���5���A�Iή�96��v�<y�]+UV�H�B^�?��82cd�<�"ˊ�[�BL���ܨ�ޑq�c\`�<	2J �B�t��c@�V�eᤥC]�<!�
�/�-ۇ����Ӣ�^�<��Ȳu�fLRQBݭ$�^R�g�q�<!U����q��[+u3h�2ˋe�<Y��X�q�D��g)R3ktܰ����[�<�E�J�&"R����,eDV��C�^�<���+��p�O�(l�Z���D@�<��C��<|'O�*Td�"bB�A�<	����)����[�qt�Y���}�<� �����Y��ģ! D���#y�<	5MR�6C��1����#%���2'Jl�<p��lyN0�q��j�x=h���W�<14%��{�A�Q@�(-L��;v#�F�<YQ"Έ6D�P���MT��rˍC�<����p�M8č�� ��0�O�k�<)%V_�$\�s��(�4�xE* d�<Q��	Y���*h�xm�W&�y�<��aɝX$l b�O [�X�y���b�<��E.˶E�Ј[�TJ0��c�< ފd���!H5�>�v��P�<)%�U�5�b�q�mR?6ȜI���k�<Q��S�\ɘ"F��W�IH�e�<Qb�3^�.�"&����)`˓o�<)�B�$v�S%+�3:��Y��k�<�� �h� 
G֫l�����f�<��E�&F��mSVg��y��ł�R^�<��w��]r���9M�qil�w�<��K�:ڀ���]L��a��r�<��`�>gP��D��m� D�q�<ѕ��<^@�ئ=�6U`"�t�<�`�F"A5,MR�A�K�|a����<�  �I��B��0��/�@f6a��"OT�ڣ���E�S �/_^�= �"O�x�6˃j*$�s%F@J@��"OL��:��a@���_=��`"O�ز��z>�� �j��"�\�P�"O�x���K?½Jw��JE����"O@���ŽM�sѐ)I��@�"O��r'�W0�ʔ�4���L>�
"ON���Y�/Wj}ī�EK�-��"Ol�8E&�D��������L���"O�I�!c��e��@A�C�0�V�6O~���b_&\�6`b�φ��`x�&�)�m��M*���!Ƌw�|ձ5fZ#��	�+�����X�-��`
��2�؈����(RHB䉝W�D)c#瓓]�������uk"�'��Y#A�z��ҧ�h�S��ȟ6��9C�c�3{61	�"O\��i�rB�4$H��[i�x������	63����)0�3�	'n�N �A�D�� R ��<�C���l�Z��t�^�A��lB�@	���a��*L���1��'k�	�$�\9I��i�N-=bI!�(��Y("��vϔ�'�\�k'�L0,��a+�G�C^�#
�'c�}+���:�*�!a F:L�H8�OjA0�B�r��H�"|b��Q$| zq(6�@"7`�06�\R�<Yp�I�r���; �Y�fX	iѯO2��'ƬBB^���Ϙ'�*4�qgS?:�����nJN�@a	�'� (���a�R�+RL�
�6}�u�	%q�Jƍx����e��`:Y+6iӨGQ(1�1�7O(�0S�۳L�J-�J�$��
�:9���a��=!��,�9D�Ժ�����^�S�B�%@QbX{�2?чB#H��ܘ�d7}��)S<vO%CQE �iL��
�a�!�ď*-ǜq�țE,j�.[���&�(z�.��Y�q��'�4�����%5$�@��8^��'���%LqC�p�d΅�o�<�[P`�9`_���I�@�6���Xw;�|��f�$I�B�I�BE�p{���o��b���+ojB�?V�l`S䌋:<K���R��� �hC�a~��'����ǝ�-��C�	�F Py��	�9X.�Y81ƇB�C�ɮ/D��I$Ć"L���.۽=�b#>����3���|b����rL���պ}b(s��R�<�w�
:`�}35�D�	7l������Q�T�%�"~B'gӷ2#�%+B�B0G�}�%B��y�c֍v&�܉�ц�T�cB�Ӭ���Δj�8�������<)��,d&LCC@1=L�i�m
yX��9��Zw�Y�"�ܕ|q��*�C�?R?�up�
�'@��d�*���1��6R�4 �U�������D�L��X�i�0(�u�Y�t�7G��˳��M�~�h����y2���q�<!�s�D�sH<D����Mca.%BzV�0&N�h�i��撛�h�k�
�#����0`��M�Nd
�`�9�!�d�=X��v�ޛsyh<���:�j��� i�YWG1,���S0Y?A�����<�Љfl��m{v]JR�\e�a}������@D 5� i��7� ��u΍�'��}QD�Q
�"HL0�O��2A��A�d��A�ɜxI�U��LH*��Y����ę��i=��S<o�7mǠ#�A&I��K�cө�XX`��-y�-I@%�T�<y �ZI �iK��\�qat+�)�������Q��}��ៗA��*pIڛI"�AE��6^�eI$�A鼋!b�.R��E	CI7d�j09��Yk��tS�h�`���Q��_��(� G���iV�ߕ`��d@E�v
zd�1	�e��Uv��'X��8� �V�'U0P6�XY%�4Y��!�R�$C�S �Hx ,ѳ"�^ )��#:C>�S�
��x��q�4m�h��c��-�qQf��q>`�Ɖ�8Ta|rH�	�y��a���}�Pm������� j���I]5�r8�g�� �W5	zP
��4L�睶R�(�'ȏ�{�(�9����2�C�	�fex#H�%Y'�<�GCL0O��[�!4�le��� ?�(�4���'>�8�d`��b} �B�yNp�1�ՙ!!̐��:|O^�!�B�
�Mz�dC��X-c'�ŵ	�l�0d��\J��;P)���'����ʙ{��� t�����^�R�U�8�H���d�j�`�B�E�?z96�@"e����' w\%�'#]����4�f��ȓ8Y���	c�r4S��ܰ% �Q��e�ٔ�	�臲��K`]e��~��;Z��Qi�]�)bL�y�����y��T�-��9B7�Y�.C�(� ��{�̞�v&��b��#�TAX��	2A���TCG�|�Xu�3G��~k����N���Y�P h�XP��G#�ha ƃ��TĲ�(�%�x`���|�b���p��g�'��Or�q�J�)�9���%C�~&���>�r�	@G�yRǨH:�ʐ	���b���ҭ�~򩖇I�4��eKLO��S�D_�-q1k�a{|$��K�d"C�2�ȥ!���w���h�(� ��'��0�+�)MV�	���O���6G���mr� �Sg(����'�&�!��۟*m�mu�	)vB�[r��\Y�����Pa��_�}��I�սlF�I o����O���� 	�A�D���!4�)ޚXaX]07C�%��y�ҿ4!���e�6.B5D���!��c(��7s�	�f�^�z�D�S�O�(1n_5"<�	Q�X.����'Kz�����n�vt b���~#�}���7?� d�$.�X�B���}����[�V�a ������C7��?!�!�]����`�uR4�ѬCjϒH "A�H���'qh�:�n^/`���X�	�џ����Ѹjh������ϗ}.�؇�U�ca�$'���y�`57Tpx8���+}0�	ѫ��Đ�dt��YP`Ц��)�'��	�G#O `*�)�phF\�^t��1��{�� /�Б��'-�K>�5K]�/��|�<C�@�+R��1�Ɨ�Z-bm��MF_(<)q`�+c*�k1�#1,60xo��k0�Ġ�"��[ HX�NQ*��⩌�HRڸq��4D��&��L���ȓf�U['6D����.HJ�K�>DX��`�.D��H4�Q��r��#��@Ð�ɔk.D�lⶫ�7,�~p�ẁC�8D���S2\u,��p��,l[�����6D��%�_�b�ze1���~>}���9�>�:Pi��'w^(�@K�9cxQY"�^�*���xb���1�i�+���^�ɢ[b�yEØ����ɼ��ݹ�����(�Y%��*���,�Iı����-P��V�����v�d���1��IS��˧�y�-
� ͈C�X������jW�u*�Γ9P�ZѨ�?�x�Џ��O*��$C�*��T��t"���B�)��|L#	Ϣh���J��n��!hK�$-���S� �R-�`��q(���#	D4W�>�*�ɤJ�f}�񢏞{��a����~#<1�`�.K����Vc�9�D��A�?��$iگ9���Bw�K+��=�G�Q�c� ��k٫v�a�	��4��Y���O�^����B2K��q��$y��@%2l�$0���5��q�pG�"[�ϧ�y��ȭ~����5S��f��0?9"�R!%Dl�3��*?4�iK!N+siN�`M�!f���#��BF���^-��@�N�*qkD�B����<1ЦX8O�|��c��&��r��[�'n���Β ��ɬ�Dpi�f�`zXc���"�b�Be�_��;� �"$���'�������?@Ihb�)ړV��v�Z�
�a�-L���$�r��9 �7�<d�ݴ: a�$��ss���-a�E���S����j� 6$������!��s�z}�%��-n�Jx`�'�u��	I�[�F��n-k%(t+�������+U���ժ"�7������^�xX���?�Γ�.�ř����VGؙ�|%��	01.�*4 �;��9��ׯl�b(�'�\<����#-trݚ�m�~{�x�G%���'���Y"��MA� ��!]��k��ݖ �AvG]$�ў��V���@��i�����s_
�
�@J ?��)���7�ұ��-N�$����B~r���@�{�'���{c�ĭT{��:�酛n��X[�4sj���U�N4^"2�D�iny��:�'X_�4�w�D6j�9�v A1:"���UE� xDp�	�?:��%��8��}��'�_Iv�`��8^�0ܻS�X5|u�@띧�i�W˲�����oy2KI;� ����-(��l��֗��>���,,h1A@�P 5% x9͚}�`<S��[���'���8Fܵ*!JF��L����mbU�O�w�x����hO13q�4z�Z#|J	>]�<=���x�G�G�[�ޝ)sꉾ��I������L<��� ?���LɯY	��2�@��<���π@Ȗ➢}� B Q�
љ[ �L�Pi�={M���f�����'v|L)sg��*t,��a���R]�
ӓ8\�j"}�
�8�� �eI<2�L[��y/��Q+���ʥ0]Rty����y2�V&[�$�C�%��Q*r�Y&�yb�C���b�-_;^&�F���y�(�V���مD7îx��G��yh	���Q(�-��;���g�yR��|T����@��l$��Z�CH��y2��e�U#���!X3�d�ƌ��yRK �c�x�H��W�ZW8�VbŔ�yJ����d�.�5����y�a�� x���̆�z���7Q9�y�iF'n�x�J��C���G���y�F�������U��LDS�5�y�l�iψEb`Þ�K,0Q�� �yB*��UH��đ�(eB���y"�O�YʀJ���3v6=��#J��y���A��̄��B����yr�M�	��y�m�{������y�c��w��E�4qv���@Z
�y��Ґn�b��!ѡZ�n��J��yR,�c�P�K��G� Ξ�����y��U�r�%��(��o�(��$�/�y���4��
���P��m�3`]&�y�ӚU�lpc$D,W`yARP;�y�ψ^�,%PB�P�F*
 �ʨ�y�,�d�&�����-�����&ˠ�y��E9A��1f��s�0�+���y2���W%�a��k�>n�.5!�L=�y2��:Ze�ܠ`I�f4J�
�GԬ�y���)��)���x�� ���y��k�ȁf��4|�8xḘ�y�����r�k��q,ܜcB�$�y�{�JjéG,jn��Q`��yҩ
 5z�ЁY�p<r����V��y�o�*|��d�K'E�~0`W��yR���t���EK\G�j����I��yr�ן����Ý�J��V�?�yRmؙb�-�-�	v�R��G�3�y�fM�hF���ĸkz��J�G �y�g�bh=��UJ���r�䑹�yrmF�PrykRM\0L����$G���y��?yz��Aܧ4Ţ-����y�P�;�a��ϊ:5Y>�"gA�y�إ	�+cR=,}���$��O�i��۴�>�i�*A�X���"O�Y�ƥ�-a���P��]:9/��"O�Q��Ά�q�D�g�k�� �"OD�5ϛ�9�$���f��8VE{3"O:)�����=&�h�2�F��"Oذ���P F�>��\6ʝِ"OHx��R���5Q�-�	{�u�7"O�QW�	37&�:F��*t�����G٦�9�3?���X麣R�?�zq藩Q�t��W�O�hPr�o��lW��z1��D�Fy��)��.�ijvE]�e��!���#km�"!�&fV�Q�ʽ<��S?||�C�H�7��-�G�M�F�����g�T��x+O���T�l�a
&,��Hs�_#[����bmH")�dj���O�1��	ɻ+ׄ �
�'�$eYt��:�!`�Y7��'�r�HQ�C�xd�ecM��� /o�Ќ��B�"ZE���2�'����WQXYT�6sS��S�O�8`�LƔ/�p�PM&u0lh�6�C�P�fH�"/����d�u>¨ò@�]��\�9�^���E0!�8(�O��`��K�'��Sr�p��6�d6�F�f�<�O�`&�f�>����9@Ʉ��t�I�r���%�ށ8��d�p�1��'�qA��0lTAr()=������� �+`@��8������}�@�`u"OzX�D֬A��d���$��"O����!���L�j��u"OfTS'nH+Bu����J�����"O؝�5�PB1r i��^�K�<%j"O:EC T�3vU)a엻3��Q�"OHhP0��@��-�V"�_m�ak�"O��;$h/7l΄Zs"�	, �;"O�=�s�9/<��go�i����"O�0@��]�e��� �٦b�@�"O2��
�x=ڭ�G�-�̒�"Oh-3B'�,/��h�D-T�HҙiU"O�S��cB��so�]� �a"O6@҇/̋p諱,[8 :�	G"OL!@��*�x%A��,x���"O�E��*<�v��X���Ç"O�ap�7-!�iQ��I�w�H�S"O�۰�D�U1���~����"O��R`��o����!C1	z�=+�"O��!�T�l���UWp\��"OH�� #�bT���6Q\�� �"O�`[�$kڦ�xA���
C����yo�=������e
���Q�X*�yC�X�N�)2.Fx3����y����gl�Dge/|�L[#j��y"D�$�����JX�%���C���y���5���Ӣ�E���RӍ�.�y�	נ"}0���Z�n���3�L�y�.݄��+�a��5#^I��-���yr�R������f�*��hI�H��yRn�Ne ����U�a�2�yr� .?$e�D�@�{� ̲� O�y�e=��Y1EJ8+f*l���W��y��ީn(L`C�twL��h,�y��	%��"��Y�oSԁxu�D��y�I��Wa�₣{)�p���� �y2F�O���K�mO<@Jd�$�y�-H<N����2l�"��v(M��y�6}����+[����`�4�yB�$.����$��NΆaI���y�$��O��aș[�44W���y�HL@��wXY��1Ղ:�y���:\2J [�'� Q�p�A5&̸�y"�!9fD��ٲt����i���y�m]�"h|�����].��z�#��y��E)�m���֜XA�}�u�X�y���_�Ȓ��
f���[���yҀ��jT���1�S�\�duj�P�yR�Q[ &Ub��W'X�T�n��y��9�� ��H�*�Ŵ�yB�E|�z�a���!A
�L�@��(�y���>Ko"l���[�6en����4�y���oӄ��$�).a�xb�M��yB�B&�:�z��+τ�B��T��y��U�yc�-R�0(�h#�פ�y�� x�fJdԭ�"��U��y�녉	G�`dgB���IP��L��y��ij2\[%-L����+����yb�ӅAP�!C�%��]�A��y�-��d���s�#��x��&�y"i�8E��~��){r���y�E��m#�ȱ3�M�rͮcB A3�y���/"�n%t
��bdh������ybjh�p�ई�60�p��%Y��y
� *@� /ΧF1�jE��i<q�"O�¤� K�	*�耘[LM�#"O�����>8���qg�
UEd(3�"O
���ܦ3�jEy�%֬}=�Pc"O�<���X���� �b���$"O��w��=D�(��2i,�"Oʜ:C�ƣK��X��I�3���"O��B�,�>�LI	�XT �;�"O숰UטzD�8r���B<�U��"OR#���0�FQ%f�t,�l�b"O���`�|y�;�$�}��!S�"O��` �'BeP(��3�H�#"O��IҾw0��M�E\0
�"O�I:7m�&=������\&�N��a"O���h��YyTM�3�E&��P�"O4�2��>2�I�̖�b����"O6�⋜h'Ҙ�#n�;Z<��"O�t)��6j�鸓,�b'��V"O$���;��9�v˘5?���"O��C&�B@��i��{����"OX�jP�T�,e �X�&R��8���"O4aе
�0ܨ ��8q|RI�"O,��Sϋ�q��	��BcZ�"ON� p�%ir���Ƈ���T�"O�� h8zA�<��EK.A�T"O2��v"�~$>�Q���/�t�;�"OPe�#�Dv`��jD�~֔�@q"O�����N+IR`��bB���"O4�E*W�P�T��Q��#����$"O�Q�;xp!��/�:R��*2"O�!�&�X�Z6�u��͉�@��"O$�y§�Iq���C���R�g"Ob�K�#��Of
�� �6��Y"O�T�4��5Z�+c�:w��*E"O$�c�!ǥ&���JsD��i\x���"O��t�	'[�00�zL���"Oް���ס�t	�q��M(z�y�"O�xUC�	����j�m%���"O�t�t�͛�J��C
M9)�U��"Oly�q�:��͹�	�s#���T"On`�eKA�[�����ԀW4�ї"O�렀��p�r�I7�B:��#�"OP���@��e!A"�-�P|�g"O�Ƀǜa�!j�Nh{�"O�|��"� �̺@�9n�H�sV"O�� ��c�j�H�o� T��D"O�ŉ��?h��(�/L464�}H�"O�ؓ�N�$gV��e�+#*���c"O q 0A�+GŔ���dGd�6�<D���o��V[���g![�)d�L˅a;D�� p6kgj��\@��L@E�9D�4pF�L�}�\��-Ů]���qI-D��`S�W��8����Ĭ=x��V�,D�PZg�M�T�H��O8K���+��-D�����	�(! �	�Y��}{�)*D���AO����� J*|�V���d=D�<8�� �*�t�� �}�(b�:D��' �>u~aHp���I�����j-D���&N�)]������;5��Xj� 'D�p���
��lBN�/&����&�%D��3�!���'+L�t�,��%D���)B<FPX�@*�0�����?D�1��
�B�*��X i~�d��;D����EM=AY�F"�>@��|Sr�:D�� H5�A�<(����i
D�D"O�(G� 4��*R�o���"P"O�� S#i�)_�O�8`�"O�B�O�,z5ܩ
��1
�@
�"O��y��'Q�̄�`H�<h���#"O`)`��խ-\3�# �B��q"O�dy�hń^t�%� A7,�laB�"Ox�[B�"iq�h�!$
����E"O�A5I��y���
�b
�S�����"O@���$_x����`;9��z�"OD0�@a�j���)`o+��r"O�A��,׷}3H\2���kJ���"O��0�N�g����f�� :��"OB�S���0��$B�e�k0��A"O@�#/�3��U(�n��y'qY"O�ғhW!i�"ѳ�A�As���"Ot����٨yx"alN���"O�)�:)NQ�˒	ZRb�(�"O$.�p�	 *�]D�"f���!���,X����J�������!�d���a���c�6�u��;r!��?k&�:��'	�(��u/{d!�\_ ��6'S�v�$q�G�,R!�R9`�����$�����E�P@!�$J�{*(��-'c�>U��A��#R!��f�V�%CI��b�0!�Z;[y�a+���:m��8Q���!����x$i+`a<��E�!b�!�'=��iAQ,n
T�wEExA!���!:p1���#[d mJQO"!�d�@����`�
*\�\s��	�Py"j��F�)b��*`HLs ��yB�s�v�Tj2(�p��� S�y"��.fD0�u.����&�D-�y�.G�d��������}~PXG��,�ybI
~3�x��+8��	B����y�'�+�p%��)2n<�/�y2����2�A/lz!��]��y��q)\HS�")�R�nB��y��E�0��❂	<��*C��	�y�-�+#Č��@�2 �써B˜��y"��q����Bu��Qr�:�y��S��t+rhW����Q���ybeޛiW&�Q����H Uт�;�y"�K�f�m�u	/� F'�yJ��hLX��h[�K�LQ��y�^�o��q����a��]�y�h۩:x|�ie���b��g`\��y�cÿ_����n�~JuG�o�<A0I+
�M���Q�p�3��\�<!#��v�z� C��;cJ����W�<I$�4�����Ș8:>���.S�<��*ZV�<��Z@��bģRR�<�D�a,����K%b�&Ir���P�<�1��
j ٵ���sRA�J�L�<ɕ�&l�Z��ƙ .�llhQ�GG�<12�ӑt"�x���R�"��F�<�#�g���(��0����F�<�P .}	^�[��V�jo2�z%��D�<)c�"���ƌ�*b���:7�\�<ap	��j����گ.C��R/GX�<i���#O�8D@��'%�	K��~�<�f�ٌ,U �)`霣
���*W��A�<��O�K��p�V�;k�j��4B{�<� 4�T�[�zZ��W�]����"O4��WL�uL=��ɔ�A��u�"O�t3��ٷ+�L�i�g�/yX�QA"O֙Xd�W?e� �%�Kqh��"O$Y�e�;e��u�H	Tî���"O(�� 쎑�J�r2�ۛ*��e��"O���&b�u�q�ԉ:�Fu���B�<9�)7;'X8��˂��D�&��<��ݬ^�|�1,��Zl��ӵ��{�<����BMHu��P5@]>	�"l�ȓ� � @�?�   �  Q  �  +  �*  _6  �A  tM  Y  �d  p  �{  Ɔ  �  P�  �  �  b�  ��  ��  >�  ��  ��  ��  t�  ��  :�  ��  ��  �  \ � � � y �% / �8 �> �G nO �V �\ :c ;i  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�|��'����F��a��������yҁ�0��(�A��>@j���S(E��y�M�-o~�C�X#?i&�s�*�0<A����	)���̖7����vW+^!�b,Q���ؐ4l������Py� z�ЩW+�5�)Bc��y" ��g[�䋷�ݘ3OΤ���y�G��@���ף�8Yj�� ���.�y�/A�yz�97O3H�vyh�{#!��J�:x���� ����RN!���8 ��]K��ʙ�2'�<c!���`L*�*V�q������ �P&!�D>�dY�Z�T�DH22��!��!�U# C]�Q׈Ł����!�d�4���{��J���7�I:\�!�d��x.��)�J��W��<[7��]N!�D�r5�	Sv�)~�@H	r�W?!��q5R�B��\�b��
�N��A!�D�+"�@*a&�&7^({�m@.�Ia��(�n$�,Q�+�����xqԠ
�"O��G+�Cΰ%�Ek�
j���"O���[�Ȉ�#��'�`cGB���yB��B:�8��|\nt ���)��d9�O�RRGq��H��D?( 0P�'"��(@4���B�ҶiW8yX��w�NC�	87WX�`�jE��
���(��?q��)�&�b�@ś��%M�cb|���� L���Ȃ/:����#6\@I'6O̢=E�t��,JL�t�� >!��2┇�y�2^��03�1bQ��%���y�,�o��Q��	�zH��������y��bat�ɇ)I�s��9c�����hO��R�h�b� ?Xz������0�"O����oL�P0��s�@��P�� ��Lw�����R5��Ыc./���e���x���N��U@�Ɗb�������Ḧ́��J؟�y��(v��C��8]f�T�f'<Op#<�4�GP/�d�0�,GŠ}�WAI��� rJ�9� B��0�&L�)�bl�Ia�����Xؗ���p�	��o�0��j-5D��"���_XB���.��[���#���fh<u�E	n�ڽ���	#�4�� �h���<17�I�0�Ҙ���g?�$-$�M��K_i� �<��)!f�q����=)����ܒ$��x2��;��)(��ӭ�y��_�xD@A�
h~��(!���y��)�v���睑
?*-����bV�8�ȓE�m;s#�4>��S�'�C7�9�'&�=��w�܋t$]�|��ěg��e8���N~�A��<��*��t�\ңΑ;�y��F:5��2�	7i@�Yc���y�F^�o�0�맡��RpSs��y��Nm�Y��e�2M��k�	���yGx���G�j&�0&�;j�LQ�u�0D��qc@@"��b�%Om����1`�>i�����(E��&~ MY��F{
^0���r̳4�@��<q#������ȓMkx)����; ְ�%$_�1Kv|�ȓVB�p�U����q�#1x�E�ȓW�4y���;� @�� V#�y�ȓ<�D���
/^!Æ�@�8�ޱ��m鮬0 �� �<��p���u �E��!��qg��)@I��Y�66���ȓW�P�!�끅V�l!V��++(L(�ȓX��,Q�B�$_�	�s������ȓ��1zw�Q�5EX8wI80�����j~Y��.�K?�� k:LK�݇ȓT�R�ņ1
bAb��ƫ4�`��(��)���9r� ʗ'�*|�<��oQ��XQ$�*Ì�F�K�aBf���M�ب	�!��O� �1a
	05�8H�ȓ
鶬��+ؖ:�ЅѷJ�/�&L��ZF��5 %IJ8A1`֔d�N��j�Y!�Ԟ!�*�05/�i%`��ȓx	�xk���60w����Hh��ȓ}��J5f��2�!׮�Sk���ȓ��EѲ�A1"��R)=4�0��J�^��gB��<Y��ҕ�޻u��ȇȓz2-X`�+��TzqJ��Fv�5�ȓ*��������>)��3��5��Ѕ���&��@���H-6h��ȓR����� &s�����O��쑅ȓq�fNE�t3��i�R|�e_W�<)Q�V�+xs֏��j�����{�<I6
ͺ_�Ĉ]�>����WGN�<)�����c�!��H� �p&f�<��#�&�|�pb��#7���FΆZ�<QB/I��Zu��&u��� �VV�<����1�>Y�f�	2$�M���T�<�r�E#/�Ҍ�F�~ Ћ��S�<�Ə'M�`�1e@�mq�%�R��T�<�  ���K'P��xC�QRPqR�"O�q��L��(Y�sA�2B�m9�"O.��&������2!��6憱kr*OnP�уu�R�b��^�[�>͙�'�t��"z̰�вfɲUG�U����?���?q���?����?)���?���mfƐ8�撞v��H�O�%\���8��?���?���?����?I��?i�+��8��c�^?�`mN-]�:is��?	��?���
ߴ�?Q���?���?1�@�CQ���	F�V�j�)���?���?Y��?q���?Q��?9���?�D�^ʝ٧��&��
3! �j�$�O,�$�O|��O>�d�O$���Ol�����U(d&J�#�h�"�/R����O����O��D�O����OD���O|�����-�U� ���P�*�V�d�O��d�O���O<���O����OB��j�`j��U�E_|��s�h�d����\�	��Iϟ�	�Iӟ��	{���d�YO,�e�B�֡V�^E�	П���؟��ş�����	ן0�	�&��HB!$�'�r��p�G1]�W�����X�I���	���П@�	���Ϳl���vꐾ*�I��@�ܟp����0�I��	��t��Ɵ����dP!�H��&.)D�Qa��^П������Iԟ��ߟ����x��ҟСE��I��e�a��Hy�$%�ʟ��i�7m�O6���O����O@n�����I�RI�M	�	C`�Ӗ�.l�,e#-O$�d�<�|�'�6펯D]�=�3K4o�D}��J�=?�N8AǕ�,Zڴ�����'g���mYv�Y�I+:��X8`�cN��'M��k�ij�	�|���O�B<�(*��s�n$�efH�6��<�����0ڧ����$&�-���G���"��JҾi�$ḍyB�����q�:4�#T3a%@���J�-�I�`ϓ����N���6-a�l@Ӫ���Zܣ���21�����`��̓�#������'����b�m�uR�lŮwY����'���r��6�M{E��J̓��"#iT�O�6����>f��,�R.�>!���?y�'��Iz� �J�@N���h�'��f����?�Я�%�^=�|����O\=��Mʐ��]�a��y��T�oN��+)O���?E��'c~99b*�;X�xe��&�sQjD�'��6�����MS��O��t����Jj:�0�
A)=� h��'J��'�"ͽ!������Χ��č֒W2$	ХE�	R�T0bØ+�(%�P�����'�b�'H��'��h�(ŐF�����Y��F-��R��s�4)��8��?!���O3�$�7K� ��c��ʲ�`|��>	յi��6�L�)�S=�8O�6~zl;N�"}.L���h�+��`���c��5�'�ľ/�6���+��M&�˓Q���q��.Jes5��E
@����?����?��|�(O��l�ԁ��-J�t���$�vu��
�)����	.�M��ɾ>��ip�6��妍�)͸5z����K��nʜE���\� H|o�D~"��rw.X�S]���Ϻ�;`h�樐�V��L� �]�p��ϓ�?I���?I���?����O�9�E!إI�t����ׁǚz�2�'�b�t��5x@?�"�d��Q$��zf'�k��P����(2��1������/S��d���ىz�6-#?1��E�H���v����?8�%`7!l����i��˓�VX������	�H�&	K�#�L9Q4�خ���3��ޟ���Yy�iӀ�����O����O�˧uJ�å�J9�4$k3/ƐÀ�'/p�U�fi�f�&��B�.Ḇ�ޮ-�f�⦎�>ef�0��5�2�+s�m~x��!��'3hM��yǋ�;yK�Ib���
� �Yq��"�'}��'���]���ݴ(N�I)�&��#�4�{����	9�iJ�g��?1�E��&�d�b}��o�F	�&�� 7>ip�0��\�b��ش�,�{۴���D ><a(�����2e�P�MS#X��`���2�h8[�4���O���O@���O"�d�|��	<�,���H�q�-�A,Ԅ
ʛ�ɓ<^�R�'8���D�'�7=�H�2���0���OԚ2}$x��ԦU9ڴI����O��B!�i5�D=
��鸒숫? \ڔ�ۻ!��ߎɤ���Jy��~:�6U������j�$�\���0���oG�t�	ߟD�IEyi`�P�N�O(�$�Oj"'Έ"�Z�I�j�2�F����6������ ݦ�K�4Pa�'�A�(;Y�2��9yN���	h����,#��4�$��(��ZG�[��?�Ԩ�O�t[�ˇ~zi	T�1B�`q9��O���O��$�O��}
�C���Ae�	=>��
�-��x�Q��vl��	T��'�"7�<�i�݈
]�%<�ݫ��T���ST�n�$Rڴ��&ng���֧n�J�p;����H��\�n�8Nm���"�bx�)d ��$�̦�����'s�'�r�'��<��'C-��-8%B	$��hAwZ����=�f�	����b�韀��ɠ}��ث��8�	4'B�D��ɞ�M���i��O1�T�;�G�/:kz�PC��C�P�$��5a���c����M�j	B�Oy����˓@F�5 f�U�$T���&?^�R��?a��?Q��|z*Olmn��!�j��9��J��T#��kaA��<*j��ɥ�M3��+�>��iJ�6��Ħ�@��ٱ0�*���=�U
@� &�n�<a��I��A���ej$�O?1)V��� �)$�N�HZr�ؒdX*n[���:O����O����O��D�O<�?��e �� �tIT�J6&�:����^ڟT�	ԟ|2�4(����'�?�ӹi��'^Ě��8�@ ���Z�MdR�Ct�%����j��|��ɕ��M��O��3�>����$sS:���I�u����:O�!@�fT�$�	��������#�j��կ�:5��8i$a����Icy"�x��-�Š�O���O�ʧ�� �h�Xi��":%�$��'���e֛�	rӌ4&��'obB�`��w\ Rdc��t(�I�&&T:�Jť��d�غCq��O  Y,O�>;��� �hy���W�Y���#�'���'_����Ow�	0�M�d���<��M@#I
���Z�H	�s�������?0�iN�OR�''7�ãY�����f3L#p�q��	1��1nZ��M�e���M3�O���Ħ׳�Z���<�3�ũ-�\��@��dܸ���'?��U�$�	̟\��ğ����X�OdFl�P%w��G���j��c�"m�Jh����O����O��?����KFI�0���c8vp�B�Č$����sӾ�$�b>a��hM¦�ϓm6�ӤN� t����*��CP(�ϓI�T`q��O��p.O<�o�Jy��'�BZ�U���zQ��}����nvs2�'���'���;�M󐡍��?Y��?!�h^�P����NK=/��"``̳��'-$�0���}Ӹ�&�lBQnݲ3��5��ښ(�8�� g!?I`+�5/�@�Ꮁ����3r-�O���l2B!"'+d����Rgԧw0�̺��?9���?��h���d�$/:�E ���!
��7W�<�d�㦡���U��p��.�M���wv��7W�p他��&�02���<qq�iWT7MCɦ�;3�ϦM�'J0#�J�?���x�h�B���fTɀ�]�/�I��M+.O"���O�d�O\���OJ�"e�M? ��cp��qv�	�C�<�a�iy����'�'x�O�FD�w�QAb�X��$�@�DBl��?�4$ɧ�B��e���X���Y�4F%QF(y�d���=���*OV��Q�?9�ʢ<1e�i�剚~�4x#����M�$�d�!E���	�h��ɟ��i>E�'j�7mZ<-���{VRY��)�(w6 ����f���Ц��?!eU�l#�4 c�ki�ȥ�b�̅���9&'M�Z-T8�ϛ@P6M*?q���>}*���ǧ�������BK����Ř0����ʽ`|��ϓ�?)���?!��?�����O ��SV�P�M}h����^5Θ�F�'B�'�x7� k���M�O>O�1oR��wEQ%&_�a&̰���?	��|���S>�M��O뎗ff����f�Sh�D˸XE4v����'��'���'���'S@	�$%�,���U�u���Sbӟ(�Ivy"/g�A2�)�O��$�Ov�'4L�L���ԅ����0x��',��?A����I�*cPP���dzM�6�̙<5b��%(b�9����-W�o�I�x�H����/g�8ܺG�z�j�����I�<�)�hy�cw� )
sa4=�iK��E�!X���	������O�l�C�=�	�d� ���f@0�/])t����R���c�4m 8���4����+ ���������B�H?d�|�24��P�q`Du��'�'���'���'c��`]�!���8�Ms�.�P�4&�� ���?a����'�?I ��y�Δ&|�y4�L���T2�霤m�H7�Ϧ�:K<�|²�˭�M��'�a���&l]�A�c��� ��'y�MʦGZ��ؐ�|�W���I͟@�!l$&�Ճ�C�*s��ݟ��I��H�	`yB�`�̑�%�O��O4��E�:[�-;����!Ft8e	"�I������J޴/��'"�� G`���2�I[5���j�O��u,�'D�q�-�� �?	j�O.l[�k��.|��;0ĭ���O����O��D�Oh�}��]��P�!m��-!�XA��ʲW=���>���Cć+K��'�67m/�i�)
V�T(P��H<j*��U�g���4%�6�fӠ���{���z7�P�ԋ�����a���\D��*f�_�k���#�������O��O��D�O��$��e�K�[�bP0r���BHp�`Q���۴��Z*O&��4���O`գ��C����r���$��*Sx}��wӌ!l���ŞݰA�(����E�.�,�pJK/b�\�K*O2�� ƨ�?	� ���<��(�)������n�� �����?y���?)��?ͧ��$U���� ��ş��U�"uMhu0��(6T"3�ϟ��ߴ��'���!�V�l�x�nI��)Ƹr�ma�˂������3�֟���SO�K����k���9��G��6�ı��&ۚ�&xp�d���Iş0��ɟ����,�:�!I�-��L�Bb� ���C��9�?���?9��i��2�O^2f��O���$��f��k�3d�Ht8�Np���M#Ʊ���B̴xf����f�	ui4l �"�א��Z	���p�' �I%�̔'S"�'#��'/��ie.��7�T����XgZ�aP�'�BZ�X�ݴVo,����?	����-k��� 7S??t8��΅/
b�I�������ݴ#9���	��4`��%�Z����f�Ұ<�Vi;B��1(��E���bWB��]�~U�8�����t3�D���ה���	ɟ������)�S{yb�v�ZȻuB�f�PӕO�*�B�(�аi�&�$�O�l�h�<�I)�M �R����oA<���R恙s���q��c4(k���W�:������π ���U�6>..t��$gg����6OB˓�?Y��?���?����Ɉ�_&��3�\5W��1֎Q y[@m�e����՟ ��S�S՟�������i��H$��+c㗏E.�y���^{���d���$�b>9��/�Ҧ!�\w����C�2xbrꑉy��̓:� ����O ��O>�(O���Oz������(H.�b1�d�޾"(��OH���O��>A2*��?���?���:k؞��4��:&��Ũ�a\��'�{ٛ�Krӈ�&�, �ūA���7!
�Ʃ��N+?�/�9�X��-�e�'3�V���%�?��ќr�K�W��Q��gRKZ����<���4�IR�OdR�����t���4|yX��rE��=�rg��t��O�O���]Ȧ��?ͻv��(�GJ�8@�Ód��C/t���?q�48H����U��v���A��ɤ=�$D�����̀>��c�����$�ė��T�'*�'m�'�"mB�#�n�����ٖ*�`�ЄY�<ٴX�~P�,Od�1�I�O!B��$
b��-�;|@D8�e�g}�}�ҽo����ŞQhƉ #�X-ttp���R�?��h����A�'|�Q�a�����|�Q�${�CA�m(���K6�n��M����	�,�Iʟ�GyroӲ��5C�O`��kT8�0�C$T� ��@×K�O�o�G��W��	�Do���M+��\�"fB���u�t�kb*��OC@$�ش��ĉ�E��(�'��O`��Z�@}oʕ\樼IGH��D�O�$�O\���OV��?��#|VHp@F	4���T�����-��şd����MS���|���|�֘|rAB�Y��	ا��g�I���� z�'����T@�jW�6���ݐYu�q:�Kܻ���`wDX=C�tIZ�ǜg?�N>�+O����Op�d�Oų�MW���A0F���?��(Щ�O�d�<Դi����'�B�'��S.g�=1u�0m�Fu����*0�O�9�'���'Lɧ��<E�t@��ٽU��!��+L��#����!A 7Sny�O�v���h��	�bɊ>5\m����b� 	���?a��?!�S�'��S����!��g�d�	R�G7��x����&� �	ߟ��ٴ��'�\��?���7�4�����+����_��?Y���dHش�������?ї'Q  ���H<�@�$	�I2�'�Iɟ���ğ��	�\��R�ԉ�8ʲ]�/��zk�@�ь6͒�s����O��2���OD�mzޕ�'�ϹDX
��G�̌r��Y�
B韜��X�)�#�<lZ�<�㛺#�L=S�˕�w� ��S�H�<!B	�30�X��L�IYy2�'����|ui8�jG�xɒe*�O�@�r�'���'��ɂ�Mk�$��?����?�V��fw~$sL����ېJH��'2z��?���I��F
��:�pT[SO��b�
!�'v�Y�֢ϱn��Vl/�	��~"�'�ܸ�	�i���@��E)aTp�1��'���'8�'��>a�ɢT6���5H�a c�c�T���M�2eYt~"�w����)7g怃�E�	N�]���M<�	��M3�i\�7MI�)<�7�7?ٲ�\%� �	�]�n�طc
�DIqk"FT��M>)O��OH���OL���O.i�6�˴/�ĝ��LM!.]%��<qնiތ0x�'�r�'���y�n��cc4�Q'� Z���x�]%d������i� �'�b>����Ш朴󰦋�R�*(�&��+�n0?U�<Z^��� ����dB3 ��ҳ�� �:�K�..$ʌ���O���O��4����Fl���y"�U3a�2Q���Fv ��o��y��q�J�ˬO�9lZ��M��i5����F�"z�x�c�؎uR�yKe�_؛���T1��lb�d�������b_�	m��ă�j�8 �?O����O
��O����O��?-�B�J����RbLEP���	p���	�`Q�4&����'��6-+���&<hڍ �^�'�p\��'�"�>i&��ܴ{��O�:��U�i?�ɤM,�XS��ʎ�R�����'W�x��nտ�R*{��~y�O���'�2$�Y�$�C�L�^���p�Ai�'���
�M��+�,�?��?Y+���r���48��qJ �x{3��б�O8o���Mk5�xʟh�)$a
#?�<��B�/�lLB�FF�F����ճ����|b��O<��H>Y���~\���T$ȻP ���g��?���?	��?�|b/ONoZ'����0JQ�[���I�OM1WW�t��Ο��ɑ�M#��&�>�3�i�@���o�k�DK�K�,T���=����o�x k�j�0�_~��q�d�2T�*O:|ÄB�+-�vղ�,4uJ�I��4O���?���?Q��?������օVO}2�e�7�H��M�umZ�Mɼ@��� ��n��蟔����#��I��I"��-o��;���b�&E|�L=%�b>����Ӧ�� h r�D�b	�=��Ǐ�oq���!�X�נ�O�ؒL>1/O&�$�O�a ���CZ2	QԪ^���" ���'���'�I�MS���?���?�WB^�z�����$i:������'4��j��e|Ӡ�$��1%�o����`
]R ��<?��U:N��9Y��[
��]���$Z��?9M�
.-��q@6�
������?����?Y��?q��9�:���J�kJp�2�C�$-{�&�O2�n�UI^��	����4���y���[���s'��"4V����yr�{Ӯm��MS��*�M��O`��d�Jt� �L��W,�@��B�^ mjU� �d�<!���?I��?!���?���8Q�J��A�~Y*)i�����ͦ5sQnIʟ,�����`Gj�d%� �B�N�Nx�U��b���t�	n�)>�2�rG2�.,�xy1�Nc�d �'�tـd�Q?	L>�-O��b���JC�D�!S S{�g��Of�d�O��D�O�)�<ɴ�i�.I:W�'T���O��$�`13 �Τ<j ��q�'߼72��=��D�O��4�,�ѵ�Ԛ���������U�ʔ7Mk���I<L6d��۟0�����c�Zx�@��10��;�H�=A�v8̓�?Y��?y��?�����O_�K��E���)W��r�R����'���'?|7���mU��O�oZN�I�N� $� J��L���j�BV�3f29%����ԟT�I��=m��<��O� 0����=4�Y���T,��A��[���'�d�<���?��?a��$I���p�Aɭw�6�?�����A��l����������Oj~0*"��r72�7��%K�O<4�'���'1ɧ���'-P��.q��d:2�(�6ju6B5�i�����a���$�L�P)��I��4�͐a^zd:�����	���	�b>I�'��6�M*u�j�b�c@A���	s�dx�d��O������?IQ�H��96���B`��DATU2#d�::���������M����u�fPDC�i�<)��-!yN�:��$,���(�m_�<!*O��D�O�d�OB���O�˧wA�e30��=�&�	���0�����i�����W���Iz�П Y���;�P���)�M��}��q�V�A�F�pӎy'�b>����Ц�̓7��"h:$���7�E(
�.�ϓ#�F�IsB�OT��J>Q+O��d�O�p���]vI �#��y1���OD���O��d�<q��i������'���'�R92�m^.O��jO9>8�U���$Bx}�'~�(n���K�y{�$Š<>�i���@�,.�'||����G
=ZXr��tg�ȟ\r��'�Rո��9h��2u��-.���x�'�R�'��'��>M�	(uzB4" � (�i��(HzlT��I3�M��X��?���D���4�,�5ύ=o� ��a"?%�lEq�3O���O��o�ye~�m�O~��K��$�ӯyϰ�X�S-�q��� �3s�	�|�^���ڟ�I��矘YGg��;d8��CK�0N�p���_y"�r�bAQ�<���'�?Y����[\���˧��i���B0A��I����I���Ş?Y�h��Cʔ=Rѳ��G;M�l��fmO/A9�x�'���3�ߟH�|�\�|�t�K�K��p��ΰ�5ń� E���'"�'U�O�剷�M����"�?!P��� �" �ڜC2�1 �n��?!��i�O�p�'3��i�7�O~偁4:�8/	%-�LՀ����Iϟ|�@Y����7?�����CE�[;[.\�6�׋tTRE���Z�<���^�Z�l�#�&l�P���i�qJ��?Y��)���B���ɍ�Y%��K��3����7�M�9�	��c=�ēnr�&�n��ŰO��6m4?�����|TY�OEڠ�`߶S0	Æ��OJ�HJ>�.O����O
�D�O���t$�8e	 ���T:'�vQ��	�O�D�<��i�D�3��' ��'��S�1| �H��X� i��O�`���5��I��M�iJ�O�� ����CƽbFք���.��R��;~T�(��T{y�O@����S��'�X|�t�6�$M \K��Y���'���'�2���O��	#�M�ԇ��o_�A��(p�0��h�8Qx=����?�i��O�)�'�rdM������&K�6��v���'R�'��AI��i�i�M���Nf�(O�9QC-	��m������廗1O��?���?���?���򉄱�Ɯ��DS!qW��Єl�Ox�0n�
��d�'���Ob�Sܟ����!�i�b���ڕ:5����GA�6�vӼM'���?A�S3aO֑o�<��#O
�%��E~��b��<Ѥ NQjL�dŮ����4���dЌx~��D헤$�!+�/YM�l���O��O��i��&�����'�2���83�4���ى��!�WDZ�FZ�O��'��6-��yRN<e��b A#1gǶ4���r"�o~bΣmFh8�#D��ON@�I9�B�h���#Z7i�ȩZB0&��'cr�'r"�ܟ��2`وB�	kӬ��AT�AK��Eɟ�9�4Q�����?�io�O��P+#�@P��8x ��1D�։��D�O�7M_ݦ��������'��� �j��?	�f�3+:8�c�H�y�%��B�vj�'z�i>��I꟠�I��I�Yd��â��6�(�V�R��y�'��6M.+�d���O~��3���O�,(g�_��n�q�G/|@�e��Gy��'���J/����L�R��e�r	��LS(���!>.��uNY��$C�M}hq��,�,�OnʓPE�XQ��=��9��(S.�����?����?���|�/O�o�	����;��ܠDO߳`P�EC.z�Ҽ���Ms����>9�ix�7�ʦ�c�����:���揝o�h3`M�!�~mt~�̀5�Љ��l�'����"�N=��UV4�hcK�<!���?���?!���?1���H1�p�r�#H�(.�y��B��&���'0��uӰ���4����Bզ�%��� �ʀuh�*m^ �z3����%؛&�m��	R/a�6�??	3�Z�? :�Z����O��Y`��1\��T�P��?YD�:���<ͧ�?����?�`���+
P\��KGi���r�!]��?1���D Ԧ��1�X�������4�O�B(I������`OA#A��A�O�ŕ'�"�iF�O��N��{�O�.���ZÎ(��%{�oؼ�2���*&?ͧt!l�dW�����0��#85X�d�R������?���?��Ş��Ċ���Wd�<���/��]���O*-u� ��O��$�Ц��?�wU���۴Z���h�"��^1vubg[�rI�8��i%V6m�u�r6�;?���#R5b��9����˴L�K��o�=ୂ2�y�\������	���֟��O2#4L�+[�l���I���;jK�7mt��$�O���!�	�O�1oz��+�JX.T�Y�&�qƄ�$ھ�?Q�4�ɧ�9 ��4�y����l���� L�"<�!NU�y�ˆH ��ɖ��'%�i>E��`v�)��/O�,��D�p�b���ʟ��ȟ\�'f��\�K'�'"2����hyE�׵7W~�#�	K��O`�'mB�'T�'�8�YM�:0|�1�H��H����O� �`�U�=��6m�c��(y���O���f�;P|��d	S��y7d�Ox�d�O���Ob�}R�X��С*�I�񨧮I�Iu���8��6ҩ�"�'��7�.�i޹jr�T�G�r9	�.��I�vbh��h�4c���d�%�P o���~%f}[���Ƒ�F�30��ܙ�@{`@�����4���$�O����O�ͼ9�b=0�ݝc��0���)t#��Q=�Ɗ�d�2�'���'L�����D���;���	a?LqJ�B�>���?�I>�|��B�	�V��$� G�6q:D+G?� �4'Y�	!Zg ��O �O�3�1��3�(�f�R�w�f���?���?���|B+O�1o��s܈��	l�@�z��Bp��J5Aݮ>d�����MC�r�>���i;6����vM�� i�@'z���W��n����IЦ���?Qw���m����>�������#YD�p��`����D�t���O����O��$�O~��0��!oƪY� ��0h*�=��I9� �I�<�	0�M�cGS�|��uě6�|r.��!h�-c�ʎb��ۖ �.��O�$mZ2�M�'"���Qٴ��$\-B��9���V��r�P��>]	�d��?�`"��<����?��?Y�@�G�haW��:�r�:��ݑ�?�����d]��]��uy��'��Sf�r�X�㓦[��X�������Y?�� �MK׼i>�O�S�nj��H���6'TY+�E,���&Ϗ�Jqi��Fy�O��ɉ3W�'Ô�����mADH�CD�1M�����'���'���O��#�M��`�-�,(g�A
Z�* �̻+
�����?�a�i�O0�'76�2A�8��Ci��S�\�W���|�0%o��M[C�+�M��O0��S	�3��We�<�� ��?粬XR��2j�J0QD��<�+O��$�OP��O����O �'4������X��jC"ގ�#��i$>\���'���'b�O��Fy�󎂛9���2
�v�P� b��3��m�"�M�r�x��$-�=%���3OJ�F(yʌ���q�L�[�4O<P����9�?i�j-�Ĩ<Q��?��#�P��<CD���wn���7�A��?����?�����DW�uH'��nyR�'���+��Z�$�:T�R.��M0��$[~y��'�֠2�;������� Pi�����X������䳴ω�?�b>���'+�����w���jFBD�me�H���?82��	�p��៸��@�O�@	�J9�	S̔�"d,�T�4#��r�J�@��O��d�צ��?�;i�{��Y=D̪�w��V^R�̓78���y���o��V�80n�B~��4����Sc�N�5!d���O�%�(l���|�_��؟H���@����D�%�~}3���0!��T���D]y2�a�Fq+f��O���O������X>�8�$��*�䑒��{޵�'a6M��q�O<�'��'|�<�W/S��	A���>`)��B�?�1�'|8�_ǟdb@�|�_�<�æѧn�R<�D˚�8�qK�֟�����I����by�$l�������OԬ�@lS p��[�kT��:\o�O|Ul@��K�ɐ�M�W�ic�7�I�V���3��-q����ҏ�`�D�t�g���d��d�R���d�>9��-S�`�rC��u������q��I��x����	ݟ$��{��qi4�
$�	��Lz��LD3�����?�����F@,��D�'Z7m �dٿkb!��ϓZy�ఀB�%���'�@�	��|�ӖpMl�<��d����i�$_7��Cw!A�>��5��&_!w����ϼ����4�X���O|�Ĝ�5��9�0�06O�d	'��?{����O�ʓ0��l�h�b�'A�R>)��-֟u��$�&%!�� {�.,?�\�8�I���QO>�O�,X��b4��ԊV'���Q���304���.��4�LhP��Z�Oh��U�
n�A�#KA'#2*M 1��Of�d�O��d�O1���<���m_�J>5QǃG^�
q��Ԗ[9�����'>�(r�f㟀*�O���}5X�P��
C/К�,$�6�'�
7M�Q�6�|�`�ɩBI��f�OdR����c��n��V�
	-�����D�O���OR���O&��|��	�`&���K:7z�@��	�L����B����'����'�6=�B�pC�q�9#�M@�k�H5��!�ʟ oZ����?��S�?�C�*ͦQ�S�? ��p��3,���;�K,HF�"1O�=��=�?��@$�$�<�'�?I���G�2u�G"D�`�$�ه���?a��?�������;�A��p�	� P��4�rqZ6�Z�r����A��hu�	��M㕼i��O��s@̀
z���a�w�b(q�����gCC�pX��S��@�rQ⤞ӟlJ��Ç"u��I%jU�+��q �g������ɟ|�	՟�F���'�"8�p�_�
p���_��P�e�'�x6풁Y�����O�l�v�ӼS��� 'V,3aE�7h�0�RSA��<q&�i��6MZ��5J�ʦ9�'�rA8�$��?�Tȕ�/�PbrG؛eU ��U'b��'Q�I��	՟P�Iǟ0Γ2L�Djvg�s>�ѡ���j��'SX7�@�2���D�O:��#�	�O�yg@�Qhhx���WT��stU}B�c��}mZ���ŞF�X��h��������{ӎ#?�R��,O�J�I��?1U*:���<YP�X/N!��	U/� {��4"�D��?���?����?ͧ���_�%b�� ���l���p�* � �Js�@��i�4��'P��(�mmӖ�nڼx*9�����qB��2 �P�YQ��r &���'KfeQmA�?U*���t�wm����F�Q1h�BL_�/tp�؜'��'���'Kr�'�eBP�I4�m8�+�RZXQC!�O��D�O��l�kG�Sӟ�{ش��]�±��Yu�ZQ�T-�N� ��x҅zӺlz>��ed�˦e�'�d�k3�_2"-����(T�mb��.u���	1Y��'��	�������	�2c���hR�]�D|J�AĽVf���˟Ж'��6�q|V�$�O$�D�|��kG�L2N�3��ͮ ���`�'VD~��<����M�4�|*�8�%F�/<�����C���,��=bX��gg�xD���|�1��O��H> �F�3��cl����q�I��?y��?y��?�|�*O�`mڕD��0'��Jޑx�³xB���⟼�	��Ms��������M���
`ј��A��4������X2�6	zӨ0�!�u�V���F���S�����fy����Lu)�-�<"���'ޗ�y2Z�0�I˟������Iן��O�d�HI24L�h_@�T�E`��ـ��O
���O2���$�ۦ�]�?蠁q�[�:L�pC��<X[���M�D�|J~*W	��M{�'|b���g�
�`p@�*.���'{�����Pɟ�Bp�|�P���	˟T:1ʍ�|��I�����n�Q����(�I�X�Iaybhv�:��t@�O ���O4��B.T�Odp���O�&0m:��v-"�	��$æ�p�4��'��2Ȗw�q�r��$.6�"�O����=Rcnmr�,8�	ν�?Y��O"�᥋��6�
d�=.o@�ҥ�O����O��D�O�}���P����3F�(uj�aQ-4�i���M<N��'��7�!�i�{���#YE�t�e�Ӌ)�`<�������劣�ڴ9��d��4����m0�x��'*d�p��Ǚ�.����V3�#�e&�Ķ<ͧ�?Q���?����?q�r�Խ����G�)r��[��
ݟ81���<A���䧙?��F�]s��H�ee�ir���Iןl�)��S�",��!U.T�@G���p��8l�0u�B��9R���p�aBfe�OʱAH>I.Oę
p�ɮ[r�Y��ɉ]zPD��O����O����O�<QѶiD@�y�'.<���@�D��y��c�0G��I��'�$6�4��$����Φ��޴���J��%I��G�u*�i���Sd�黑�iQ��0�N��Oq�\�N͕l*YB\�ޚ�rc�֞3���O����O>�$�Oz�d?��{�(�3�E�D�b���4>Uvl�I����	��MS�$��|��&��֜|��4P0�@�Dc�JQ��.f�O����O�i��K6�(?ic��"وH�U�#S(�}�A�K	s�胲m�O�8:M>�*O�i�O��$�O0(����u؊�q��O74��d�O.�$�<QV�iS��CE�'��'�哃iN1�,J�Bs:�J�(ېh�F�F���蟸�	����|��V�R���x&�-��^.em��j�;�qc��a~��Or(��0C]�'�8A�tfG*4�ҤZ$�J\�z��'Ar�'IR���On�I �M#d��p�n00������b�6B�t��?I��i]�O@p�'$�헍$�ղ�a�m�ta��1a{�Nx�z8�ce���t��YP�n䟮�Ob,�@�V�h![SCڊG��mX�'��	͟���џ��I럤�Ih�ԅ (��L��2<�X����
Y\7G�Vۄ���O�d+��	�M�;-If����[�U:��@�*��	��ұ�i�Z6mN�)�8Qh>(oZ�<YSe
8܈q���Z떝h���<��C��M���	�䓛�4���'8���'���]⢆I�����O���O��J��vi�n���'Z�G�9fCҐ���-^�8(�+ϵAw�O$��'�6�禙�H<���U�3�4`zs�++��X���G~��̩V�n���#�>i��O�f��I=i�"�T	5�Ys�N�C��h��̘\��'��'�R����khػf�|,H�ϓ��2�,����:ܴ9͢�a���?Q��i��O�n�|���Z��Õea\��l�0sj�dB����4V��o�12A����� �(c��d�ڢ`�����	(5ք��V%��'���'���'�r�';R�'��I"�ɇ�Z�1����_��	�M[`���?I���?�J~B�3����#��=��pa`�W#;@��z�^���4$�Fg(��Iݱe� ��X�ߓ[V~e��7[n�͢GiN2�b�K�|�Qv��O���O>q.O]��	j��ܰ�ݍV:]`���O6�D�O��d�O�ɥ<�Էi{(i��'��%S�ȓ���0Cj��
�2�1��'�7m#�I ���X����شG��f�2C|���.�|�g(K�3+����iu�	�,U�S�OOp�&?�����FX�S-�'yޮX�'ǀ�A+�����	�	�0�	l��e��()@�5��H�uۨ����'��'s6�͈O����O0�l�]��.:dX���--��p�!J����&����֟�Ӣ{��Dl`~Zw
X�(�PD��!Y��[�'
���1���<a���?���?���+�t�P$G��p�T[���0�?i�������aJSCA��	��0�O��a�=G�Z��)	�s꜅j�O���'���'}ɧ�i[�OG�}X"��5�����'S�>����wĀ�Q�7�my�O�����
�=�c�#a��Kف}���y���?����?��Ş������������]�HL�x�N���m�IџD+ܴ��'�"��?�+�'y�a@Oĸ<��� ���?i� T��޴����@a8�?q�'���i�&�n�(���ox�'j�	���I���	�����P�d�դ`Z��E�c����CK&%*�7-A^����Op�D,���O08mz�y�a,"2N 	��K�]��i���ן ��R�)�Ӽ=�T�lZ�<!.��)�l�
��ɞ>�ԙ��M��<��
۩����n�Cy��'���3����*��׌)�"�'��'���M���I�?����?��&�i|t(5��9HM��������'�x��?)����5��MA��&����*Yǎ=�'Op���B�R`�&D$��Ć�~��'z�1��K�'�x�bE��39�����'+��'d��'H�>��ɪ/m:E��aؕ*�x+��
�2��	��M{�����?��AK���4��ꡆ�.���`+T�m��6�O"�l�R�l�:8��n�i~���lr
%�S
5�:�P��1+�^U�$�c�B�;�|"T�����h�	՟��I�x��@U�A7lp*��`�6��Lyr�`��Z�d�<	����'�?I�O.7
aJ@-��|	�]p��I"�M�T�i)�O1���JD��N��D1C3s�hb���XV�@D���фoQ#$U�cy�i�4���	�� 
�3�W���'���'�O��I��M�#b��?�PD٠7��;e�
9F���scӎ�?Qҽi��O�$�'R�6Kͦ}8ڴƥ��1�d�PA�#k҆����C5/��5l�s~B*�^���x�'ǿv&Y'ld�I$�4���ࢍO�<���?����?��?I��$	EYꢌ:S%�`��y�
&:���'Y�v�\-�V7����OϦM'��X�<7$c�$�$#�U�'���ēiD�V`�� �=R"6�8?ٱ��,YDxP�+R�}&�x��$��!��O
��O>*O�i�O����O��jL�B|J�3�O tc8��dd�O��$�<�V�i� �'��'�哲c4�u�P��
�q��k�O�h�H�	��MST�i.O��,{�D}x@.B4|��W���Ѳ'hT�3*�I#��9?�'ofD��3��)��#C�_�4q�ӏ�0ZK� ��?����?��S�'���C��tn#���2v��/�\�A�䔖/��!J�6�d�W}��kӶ�D٪)L]zꊲX����B`�S�4-��P��4��Ę�Y:�'��S4�9���		�P�a����+D��	cy��'�B�'�R�'{2^>]��@N� jte�d/ΈB(�8!!��&�M/1Lv��ɟ��u�s��������ɔjd>aIw/S�!�v�(5���{��F�l���'�b>I��MŦ��H�Dذ�m��?�ȄGG܌hK�ϓX�>̂���O�̀N>�*O��O:-�q��#~H���.^��x��+�O���O��ĩ<���i�]y�'L�'�
��ת�l2�#'��ha��D�U}��r�dnZ&��jF�թ�i����e�ZF$����������}��Kc�3��!}��S���P�U���A�.S)jv�����۟@��՟ �I˟xE���''`�H�&��*7@�1��l}f����'$�6m9%#���M��w��U���WZXc0Ϥ4D�!P�'�J6��˦!�۴ܞ� �4���I�chҠ�'H43׊�%"tjs�M�:T����$���<�'�?q���?y��?A�%]%l<b�S����Hf�-q��O�����ئ��wJI����	���&?��I�*E�(��
]�&)f�:� E�p@�O*=m���M���x��D#[1 d����*<@�0c�R�{t�����
�;Ƙ����#���O�˓4�riA2lݟt�(l�A$�{Юx���?���?I��|"+O�8lZ0'����@�"���2��x��9Zޚ�����Mk�2.�>!״il7���3g�W�`l�{�^' �D	��"�$zZ�o�^~r ��L�����E�'���cD9K'�!hQ"ۻ]��{Dā�<����?)���?!���?���d����T0��$(^���ֳlr�'2¦|��H��?] �4���|�,��+�@�
2���K���'�"������X�v��h���-^kFe���˸V��[��!>�\���'\��'�������'���'�|D�2�,
N�1/[�XԘ	It�'t�R�`2ܴo��h�+O���|b�?3A,��hP�b|2 �
d~��<��Ms3�|*�� �q�f�M�#zzAb��2V�����6�Zو&`$*��i>ݒ��'@��'���SA�-�r�02Y�?�.��J�����@��ǟb>ɗ'ox6� 
_����$��ŢpB($�x��)�O����Ħ��?�rP�p�ݴ|�"�d��Mᎁ��	��|l"��i�h6M+(�V7�7?�DCڎA��� �T���&	%�'@6^��lW+�y�^���I����I�$��Ɵ`�O���@߬s~���":,���Kb�6���O����O擟��d���]0l�b��uh�#��`H3
E)\/����4����(��Ѿ^:6�b�l P̻k�^H�A�	�@�x�xSGw���v�œ����X�	Sy"�'[�']�I���!�x���#2��'�2�'��I��MC����?��?�W�ZX���.�	%�\������'q>ʓ�?�4!�'�f�kP��5yׄi��F�0
`!��O�	sW×�\If��󉔪�?A�Z�j��Z)8`��É�m8�����	-�2�'|r�'^����аo�6�L���	n�(y���H<9�4#��=����?a�iH�O�.�U���BrÊ*t��9 ���^�$��Cݴu��E�
k����c@�K-���W�iq�A��)�P �TJ�_��$�,�����'���'!"�'Ť|�c�	|�/9�r�mT��ݦ����Ɵt�I̟H$?q�I/.�ɇ@2T&|h#��:�6PR/O4��mӴ�%���R�b��6MYr��S��"
��v��/P�asD�� �s� �]���N�Gy�F�8���ƃ4�.��*��0>�Եiݴ�q��'��y���A[qX���"�>�y�W�'~66�.�ɕ��d�O�7������l��2j\�Oؚp��;�`(S���mq~���E*��ӛ_�O07�Q )h�vK�#a�� ���1�y��'�l���F<�]!�o��U�'���'�7-G"=����M�M>��Y�*2ٻU�""ը1H���.~��'Į7-E���0b)lZQ~�O�1x�*�r �:��̛P�Ny<T�.R蟔#`�|b^�\�?!(ƏR^MB���!�����f�'lf6��>X>��$�O����|��A�1��j���"Z�֜z憚X~Bj�>y�i\6-b�)��i�"Y\\h
*D�X �a*�cBH��(R��ָ�H��/O�	Z"�?	A6���_�~���-��<N��͜�[����Oh��O���<�B�i��؂���$L�����1^�L1BbMH�h���'�27�?������
Ц�xg��A�x�(�"��a)�}���Ǩ�M�i�x���i�	@�zq5�O&�M�'���A�߳|�ɔi)t))+�B:�mK!�� t�9V���d�J��e�ڹ
&@��Κu��)�V��,�#ڔ*��J���P������)I$��I�i��H_D$�t�ޭF�$(���=ғ:��L��*zN�IJ֍E.m���"Ӌ�uܸ�B'���n�pT���!(��H�� nf���W�B q��mbR��5]DmX�>n��k=Qɔ�0�ك�F���`��asT�����48>pA�h3M��Qp���	[-ޘ��@/q��hT��?:��[6� Eڮ�nZ�$��۟|�Ӈ����<�b
>IΈ�X��>����-	���� ��O"�?��I+g;�� ��V�<!��ED�f�<�ݴ�?����?�Q�C��Iuy��'���,<�F(pc��Nh��w�ٴ/ѱO�(�i+���O���O�4��½X����V`��2A0��a�ԦU�I�[�,i�Ot��?AK>�1V�̨H��Y�k��S珐6G�Vi�'�i՗|b�'4��'��~8��!���u��E;���o0Lp�X�����<�����?��8'|,��nW2�:�Ӓ#�(z04(:�dж���?����?)+OX�����|¥���h���U 2<�`� Ԧ!�',ғ|��'-rCޏI�dKq����!� &3(�p�!E�WD�I����ޟ��'i�q��h�~R��q���Q�J	�R�G�<P��"�ik�|R�'j�i��RqO4Ԡ����<�!1��+p9��G�iQ�'%��&)Chp⨟B�$�O���ʇg�����*&�8k󧄆��D'�@�	ɟL����d'� ��y{�< eJԇY��W�P�D�r�n�Yybj�.B[<7��O��d�O��iRg}Zc��52KF ���I{����4�?��>c8}���)Ǳ/�1�!dߝ?\�pѷ��i�vc٢F��6�O����O���P}�_��适�M9D�ŢKt��,A!X��MsW���'G����&6�\)b0�G	j��1$[8Ye@hl�䟰�	�������$�<���~�]>.բ	��Ӌ�i���8��'qr`i`�|��'8b�'����
:����_q_���3,q�����4��?�4����&�$���ҙ4G�qЖ�@�ϹV�|�'����ԟL�'���'O"U�d��@vE�soʣM�̽�G [�����-���O���?��<ID�D���eQ�*��$�V���������$�O����O"�4%�+w;���;�JO��@%�˗����	^���ϟ��p��Oy�$:;��bU p+\퉵��v�R���u$&OX�d�<Q��Y$���+�|����-�@h�1#�4�ʽ2��)*��nZX��?+O4@�őx�1��e�S΃^�Q�ĉ���M������O�-����|����?���K��۶[�*�b��Q8Ha�&&�$�OJ˓$�DxZw�f��Ђ��o@ X�4�S�D� �4����0W/ܕnZ��i�O.�ɀi~
� �I���Ȣ!�&���; C~!cD�i���蟰��)�ħ���ݲ�]4m�N����-g�=#t�tӘ��
�E��ٟ��	�?�:M<�'>�H:�F�:	�y˶$^��H����iD��'�"�|ʟ��O2����^sو�.��q�\*�Üݦ��I�L�I�cH|8�K<ͧ�?i�'����qU�l�l���-ЛX_ȹ��4�?H>]?�?��'���D�ZQβu��@�`h:���4�?	�6��e��D��-�hX'%����a�sٯt��%�8g3?���?1����D�SB�C%������ �,�uY�!Y��ޟ0��򟘔'z�؟�X�7o��W����a��$:���1Ƶi�BX���	��T�'8��ד8��)����Y��+���t$EG���'�r���O,ʓ:��4mE+H�R�))%� �V�� K�O��d�<Q�Q�D-�.���d�:jd�R�F.rW�0��*ŀ%_�Am�|��?�/Of��x�=]���7E�=�������M����?!*O:���CC�̟��s��3"�\� ��Ff�v
�u�&c�Bʓ�?Y��?a�����<��:��us�(��5�ؠ!I۶P��lZ{y2�L�Iu�7C@�4�'��i;?q�$~}Ad�X�R�S�����'�r�'�����g�s�6�����/��4䠁)�MkqK��F8���'�r�'��Tf'�4�:��R>@�Fѱ,bx�9@l��M����Io�)��?����;m;���ޕU��Q��֤G����'��'p���tg�>�(O"����|:��L77k� �+��$��샷�>Q+O�49������P�	���;�W���dW�D�!�8�M��Y"���Z���'��\���i�u��c�@����q�N�3 b���o�z��<��O|�D�O`�d�ORʓi����3+��e�꼺��\�m|$uJ(D�E���_y��'��ߟh�I��憕& $�2/΂���q���ͪ�ICy2�'OR�'剤-8r�Ot�y� <v֨��O^�?��3�4��d�O�ʓ�?���?���<�¡�'_ը��E�49�4�$��'����'���'��T�$0� ����OzU�0�/Go攑���G�dA��(����	Xy2�' r�'g��c�'��C������T"�P��ߗx�tnܟ\�	dy�n6W�b�'�?����"�Ph��񵪝�����$ɰcp�����I���ADkh���	NyBܟ$e ��ؑ=��̃��
�R��ði�I�]��ݴ�?I��?I�'J��i�Q��l���,�KvM��"�Ψ�IzӐ�d�OJ���	uܧ�R}a���]Wh�ic���,|m� TW:U�޴�?!���?���6���Sy"�K�&�P�R�h×h��\c
�#�P7�؏=e�D3�2��,BQfǸ1�lk#��C�f�e���M���?y��I:1Y��i�R�'E"�'�Zw�����D:xsZCra�(e�f���4�?Y/O�7�g���?���?i%eW�~<����(�e<꽂aB�����'Vz}�7�>9(On��<1��#�87��I��Ν <��Mҡ��r} ӭ�y2_�D�	ƟT��|y���c&���fv �:�G:N�ʡ0�>A(O��D�<I���?��[v�1i����X����Ѓ1�ָP',��<�-O��D�Ol�����B@�|���\�,dB��6��7�㤠립�'a�Q���	ȟ��	�+
:�d%���&�48(H�
h�+G
`nҟ �	��	Ay͜�L|�'�?��5�H(C�	f*��B�;>�l�|�'��'�*Ͷ�y�Q>1�p�6%��;Ra�<l�B��aL�<�M{��?�/OD\Hg
FR���'���OȔ�:� ��7� �� ����E�>	��?	�9���Γ��9O��5>��-z�ݴ}P�x�@ݖB�6�<�G����f�'��'
�t@�>��@��%�$g�!J�4����!�6�l�����ɘx��Ig�^�''-��Y��
$A{����X�aj�l%"�����4�?i��?��'.��Iqy�'��-d��A�� �m��t� ��M	J7M�7*��Oʓ��O�$�R�r����A�cټ���
	v6��OT���O ��"�N�	�����y?!qAS�D�.�r�N� I�Ck�Ǧu&�(s�Ø�ħ�?A��?��MQ8P$+2���kݩ%̍�5�f�'mV���#�d�O��'���&�"�N$e���(�O��-i�^��顢ɟ,�'a��'�P���#��ucx�ҕ#[q���`$�!9DD���xr�'�r�|b�'��ѱbT�0B�aZh�Ef-!�xZV�|�'2�'�	�m���#�O��)��G�@:b����bI<����䓓?���rj��'�f�uBȚ0�&a��DT�����O��D�O����<�I�$t�OiDm�Co�uꉑV�H��mCd�s�*��#���O(�DY��5}BdIh��jd���1�J�	���
�M��?�(O�p#���t�Sڟ<�Sh~ |x#$2>��ĥ�0	�<H<����?I�)�<qN>q�O� Z��Ű|�vaذ��ABxYش��ę�/]�l����I�O��I�J~b��?>
Q�Gڋ5bH�;pƟ:�M+���?�JS�?qO>q��T�}{�	��X73TVa�Ga���M���"dB��'Y��'��#(�ɲ}Zޡ��"������D�v���:޴�6@z���䓔�O�bc�X���@�i�>v4��h�>G_7��O6���O`�s��b쓨?�� Z�k�#P�&���T��1/���C��iK�'��s���	�O��D�O��x�%�V�f}���2�2u�t*��u�� �`�iM<���?!K>�1 �M��K͖v4(ʱi1~���'�ȑ���'A�����̟ �'̽P��2w���:"�� P�t� �.͞5fc�8��@����<�	xd>�"�-2'#�����E�S��-�����$�'�R�'��O}���6�~>���'��p��u�c� �($�>Y��?9L>Q���?�
�.�?���ԋ'��u%�1U��/X�]�I�0��Ꟁ�':<�2&$0��ŉ2h�9�aΝ<al�e+GO�QmZ���'�,�	��B��c���Ol���!��ڵ���<���i�2�'��	�95�miK|����S�#$���)Epa�u�� �h.�'�R�'��ِ��'��'��i�u,BȰ +D�6SxAլ��i&���'B��H�2�'�B1O�d�'�Zc���"4�D�K�5�'܍R=�Y�۴�?���3,@xB�EA�S�L\���& ����TjR�~���m��
T���4�?����?���g���d�$�T�o�p������0
C��Ax 7�F,
����Sx�Iܟ4�q��9!w$�����/fu��g�3�M3���� �r�'$�	֟8��~䠥�� � ����U�����DZ�S�T&>u�I��I�T��q���3C��:�A�D�*Ձ۴�y2A��?���8p����&��q$�A 2�l�	U7�)I�դ��$�]&UA֒��������RyiݯC5�m�C68%�ܺ0)�6q�p%3�ϼ>����?���?�r�gx4�@`��.l4��텝�F��s�|��'���'��'�t��ޟ:�a�D�aZр�� =�`(���i4��'{��|��'z�������4B�� ADIHG��D��ɵDE���'r�'|"�'f"�I_��'gBȩ��$�o�+�hYI�٤n!�7-�OO@��O��Х��Tv�'$x����!��EҤ!^�Q
R�`ݴ�?y����J� ��'>����?9�7n�)������N�9�bƇ�M��o�$��8��i�h3(�0?&���iņ6��!ߴ�?��B�ج(���?���y�����L1x���<h���0.X��\��Ĳi��'V&�G����Oni`���<'&�pۘj�ƴ�4Y��qr�i"�'���O�hOX�d�t���V�"�&�ǮW��@m�2x"<E���'�f�#v#(VgЉ	E�^(_f~p��f����O���,�r��>y��~��n���c��*ϔPa����'[(��y"�'��'�� �D�]%�ĉ�o�)#�)�b����U�z��$���	�P$��X'4aH-9v�ȌshT��6��:
�zq���<	���?����$�)j��٥��6�=��b��cYɓ�F]��?�M>����?�E&�%R̮aɠ��&j�[�b)nݒ��<Y��?����dH�_�hxϧV��ƭY�6j��K�l�	~G~]�'���'�'���'G<���OtmA��W7[��A�J�k����Q���I۟��	Oy�t߮��q�#��!	TG*�2T`Vēbg ���IF�����AX�c�Xk�V0t�����Hs�����xӺ�$�O� Ĥ�Ks����'�����8�Ġ�A�Iz�#Ʈ�z��O����O�EQU�~�A=
��p,����rOЦe�'ъ���K`Ӏ�O���OE�4�����a������(i�<nZ�����#<���Ď�� ۼ����.R;y�R�Џ�M�!��7x�&�'���'��o/�ɷ �i;�'˥^�v3F�+�9�ߴP�րDx����O� s�ϐw�}�g�==lY�K����I������"�tɨO<����?�'��=�e���+����%r�}��6Θ'�b�'��xa����5��Y9p�Ķ-f�7��O��B�f�<a�^?��	j�	��T���ؐ0����%ɉu"��O��ؘ'K��'��V�4�TIW V�P$+S�
@x�-2� Y�v%{M<q��?I����<iE-�,1�e"��'�B��g�	�aH2��<	���?������# iV,ͧ7V�k��M:
0թT��#j��'h��'-BS������%�~Z�g�v2 ��� �/,f����J}��'32�'g�	�d�@ꭟ��D����I���+TT�Ւ���9g#vn��|�'-��'�B�_6�y�R>7m��~�~}�C�Ԇxˈ�(B��3Dt�v�'(_�d	RhM��	�O��$���=���H�J#H�~��r��V}2�'K��'%(�'��s�L����"����C�VD9 嗮)2J�n�Wy��L�)r7��O����O����n}Zw~2-�t�] S��%�)�Z{JA��4�?��j��̓�?A.O��>͘u��+��S�E�X銆nyӺ��QB��1��쟤�I�?�y�Or�f]���'��O�����?!��B��i<L[�'��'��b���v!HUF\�q9��	_dQ�!�|���D�O���!E:t��'��ퟤ�{���e��T���`�)it=o��|�' ��R�����O��D�O���Rh�1�����L;���Y�N��	�n�	��O�ʓ�?�(O���ƄP�����! ��;�$R�Z��@�g���	ʟ<�I؟��IMy�S�u�\��Ő�7��U��Ř�"�l�Qǎ�>),O���<!��?��l?� B�ZEkE�A��Y��9x��cCU�<!��?I��?�����C=Q��̧6Ai��b_�rб	�(�."��(m�by��'�����	��U`x��ػm�R@R9%�r���0���?1��?�.Or���Q�t�'��a0-�! �"��©G�o��,��Ak�d���<	��?���
 ���?��'Qv%H��g;�h��h�*p`\ij�☜y-�9��>7�>)5�.�P9���	R� ��L�O�<@˜�(�xT��S��|�$�� ��1)���
B�H5�O�T!*|�������T�[�B�����!Ũ�������/u"@"�#��oY��hV��^� (��K?LI�HYU�V�P�XK%��5AJ��cT&��Cթ���J�p����D�&�֠�奌�w��8QS��*)���a��y&8�(�mA��@��nԌ�?���?��+���)*Ӿp��V�Z-�6倨(�R@'� �e���8b>�O`���@������8d�p� �
iB�Ha� �A�* q��'ޞ�0X�5�*y�wY={����'���'�ѳW�������OV�#p��2JuA�Cұp�8`���74��	E���w�PU��� ����!v%#?Q��)�/O��7�4"��s�G�15�͑d��8�(��&b�O��$�O����ԺS���?I�O�<L��"ё9 ��n��Ht���;CΝ�����d��'Mp#n��c�D����~�^�(��]��z�Ae�E6K�=�d�'�|��(�K>��UbF�J�`d��8�?)���hO㟄������C�"dU�t�t�LB�ɀG�\	#ĂExX���EA�~+�c�lx�4�?�(O�!2��c���'nIS�!!<��4�ݝO��� 7�'U��H�b�'#��:'XDو�i�i�>A!�d}Ӑ�SC`K�a��� t��>�����'-XA+���-u� SԪJ7���OҨ<Lx8K�mH�sk��b���Ɏf	����O�L�! �ߦ;k&�
f�K?�\�<9ߓ3��dSѣHFH,҇��@�^��L@�FA@�<���m�5$a��ȏ�'�[����aգ�M����?a/�R����O:��5-S�Pw@d���'|�&(�b��O����<�4q���9�ˮO�D���B�KÂÂ'+/@"���i���a2HD`+^1)Q�T�O�.� �GM�^��e��3Ps��H��� ��O�b��?QS�C�$��q�dᑪT�-�4 =D�[��^j�������:���CM-O��Dz�j!38�4F�w
6�a^�O�T7-�Od���O�2�Ѫ9<p�$�O��$�O���y�,��E��a9bQ��p�!�6�3lp�$k�%�$-�0a4-7�3���^��$���k"��S��)O� �$�e����U�������|��8i��A�?�L�pE�K>	�1OB�p���Ϙ'��d�Tl�	�Ҝi��٧f�v<���hd�NU c�A�wT+<��1�'9�"=E����^#*�e)ԙ#[�A��f��C�P3W`�"Q���'42�'%(���P�	�|�P�R�3U�x@�FdLdzV��,�DxAĬ2fa}�����J�jc��]������,2��Ka��4 3X���^�i���A�,!C|�ӱ�@C�����'�Z7mϦ9�Iy��')�O�9�ʉ�~��H����fQ4��"O�e:v/T�!P*T�*G/i:��ڇ�ĝP}2T���l[��M����?�A��Fq����	��f��aݖ�?���9�i��?	�O6P��!��!�&����fp��aG�P�!q�G0
,L�O^O8�\`DB	�)��Qe�%O����� h��Q�̋&>~��)�� <0�x2�T2�?�N>���?���E�$��s�.OD�<��#I@���G����Hxp�[B<A3�i���(��,�J�(�ʨe^��x�y��fZ�7��O��d�|r!ك�?���RcT���7��
� ���A���?1�w�����̠X[����d3*�"�'\$��Z��8����3v���O��ɴ%� (Fn�:r�J?n%�#}b��/6VA�G�4I
ڽ��#\[��1h��'��O��O=@���M'E`�����'e��*�yb�'{�y�������2a�c��P� F�
�0<10�	�4��P����|��΀ |�pY��4�?I���?�1�S98�����?1��?�;��58��Z5����� K�L���3�hei�'�� �W������q�BɰQ�mt���#gb�!h�)П+Kl���'\p�S%�J�g�Q�X JM�� �d��Gϫ� -�<��G���>�O|��&�0n�!q�G��k��(7"O�8#0H&X�P�ɿht�	 ��\Z���ӕ@(>|�Wj�AGٰ�G�;x�C�	�:���8Ī�2Bհ��G���C�I��MHbM�m��-�5���{��C�I")?48��X�3]~�R���͜C�)� Dd��&A�Ťm�iF�J%j�I�"O�cdmЯRP����ǟ�:��Y�"On�[�F�F���I�mж�J�� "O������c,����<d����5"O�tbŕ8��ha�לf���(#"O��0�J�BLҥӦ��u���i�"O
�B�خ5� ����x��"O�9yUO�6E����
�T�<y�"O�2TNƚj���)�U$p��L�F"ON�3��](5\L�s�i�9nu��"ODE�f�e&�)"H�>��X�"O�;�&��f��UpP���.|RQ"O֡��A�!��l!����3"OB��ADک5ֆa#�Z>Xp�"O�q3rM��3�(�R�2j�!&"O��XN.fTH�Tf�bV|M�"O�5�TɊ�w�ԼA�O]�7�=:�"O��EIO��H�F虰`P�J�"O��oV��zì�:5� �g���y�(Ϭ}Ͱ%r�@�)Q���y �/~.x8��˯�>��2�y��D9K���4@8���VMć�yª����%��K�0þi�uD�3�y�l��7��uy�瓐%� ����л�yɔ�]���G�. Dxe���y��E�U��� �L�������̸�y�k�E��h�H^,� �6僅�yƃ
 ��)�e�z/Z����ĩ�ya�<b���% �\��ѩͣ�y�	DlN�'��q�
��Fϣ�yEĽ'�dȘ�oM�YT��G�y��B	@5�m��`�Mo�A��U�0=�O��3ϰ�9E��`��K�F�e�N�E"�2scR8�y�nV��PP��Q�O:�s���'G*�Y�s�v���$�'KA�| !*d�x����L����s�d�����LP���L"�pGJ�"vNp�Z�@��!&�g~"o�<d�pXxu�J�w�]�B�Ѕ�yr��7m����K�G !�����]�v�X,{d��:� 1lO��qV-̙?U�ӗ��rx@��'o�ɋ�@;, ��o�J̛��ݾ}�x EF �j�j&"O���kQ�ꈠuEۭt�F�z3�Dگp�V�:��>%���E��`[�\�𭳗 Ӂ#ux�ۑ�ؔ�y�'��-v��m��0�\�$s���=���5��E��O���$m�($� /��6%&�+D"O�Al��U�!; ��% <-�+�
̆I����|}��	%�=��	ݎAH����ݿO����d�"���
T�ޥ|w8�lZ�CI�x+M�I�(-+���22�C��jӶ=���ȃU���Y
3@�c��XX7H���m�!�H����d/Ǚf��UR�gX7!�r�� "O���J�sfڥA��,>�b�)��,+C�dx�\X}�kL3���IG��ʆbǩ!����A�-#C�ɻ������W
2D '��r�P�;�/.Z�n��p B��=9`�.	׸��� ?TP\��^[���0�(,��T�����M�T�E醡��a��Bt��s�]N�<�l��h$␻��]�9r��J�Y�4y򅅈
��Y��R>�SB�D�{*�Yk���e�p81F��C�<y�bV�Ph��*��x�C�'� 8b,�'9~�s@9���I+;���P�,D�p���oX �B�[�W��l�G�	5m�����(�g?����s�D1I�,��7
p7-\"�yljV�h��@�Z��e�!���?��E�$�p��@DX�ԋ�1U�f�#�ߌ��d��;:�qp�O�t�P`�G���Fj@ -��"OK�*p~����1[~}Qԍ����'��1ذ�B����� �!:�Uvq�a#c�3*z�{V"O:�I!���zgZ5�Gҙdg@usE����:I�y��(�7&�-c�$5�N3t0��X�-D����E���^x@�K��NL��ԃ�O)� ���|R��t�����
QXza#��	���=Q�4V��0���AZ4(�St�b"�����ćȓgz:���@!%V����D_&�%�?�c˅�@��TD����&�Zd��/�H�r�0�B;��'Nu(��2�'t/��٣�J�_J=J@g�l�R�wBș92�b��E��'���"�])p�,y���Rr4�#v(Ь)J1O4�a� !�'�yG�1,��4�E|��!a�`ء�?1���NJ��	�$L����L�)׸i����k+�K�,��D$i%��)��L��DRL��}�'��0ۖ�3߈uB��6L�1)
�`�j�(C��l�P�6vܘH�2'�(�#v�¥IU�iaÅ�$a ��dٝgd��	��I3g�P�(D3_��O�(fkа�y(��X��M�6*A�&>�IƁJx�����'���%�;x��ĉ6"��R)_K[MY��$4�Hc�J`����M��E�z�	�˙��OA�n?]Y�����Q�L�<pBF�()!�D71��}Y���1&�:�bwN��Dpwe̵1G
9�6g�]B��O��]w� �ɦ,|�ू��	ވ��CK�>����*[6����'�|qڥ���.������S~� !
��xi��)Q��Y��I�pt���^�|�m��&.[2��$��KG�;�ϝ~���R]6d�+��eO����(�@ �ԩCN�G}r��T���|�2&� �,��f�c��r�'E�-k",��>O�H2"�	7�RE�6.� ��O����?��]AC-R�R��W�:E"�
�'_�p�c�B�S�O�>�Y��|]B���	mh�Y��䃾Q*�S-e��҂����a��xU�O��A��i4�d*cM��20L���'�x���#H�6��i��4�`�#jݲ]�ؐQ6C^_|�]�F�vx6�ɡ9%�����/�a�T�=���	eb��N�.=�������x�d�[D�ӄ�Z1	���\)f�����ˁ'lq�������I��ʧz�xx��L$&	��A��?xK���?��oH��Ѱ�G�����qE
G��pnH<dx��k�f�\��U��(�����<���Z���i)��@���E�D��b�o�ld�bI`w<<\'�`��h����
V���UlȓQ���t�S����b�A̱E�=�m\��:��TW?#=Q�bد�~a�'D-zjf����ܺ�4tuR��'fWL�';b�ր�UCn 31��G���vT��N0�ӁS��Px`"�|�'��x���
����f抴 6�R0�ߕy�ԙ��`��ok��|YwM�(PB(����jL�P�\>��.^$SJ0$т&Q�/�$��M'}"L�W�I�`��:�����JD�OXt���/�U*9B��N?ޱRٴW�����Z�tЫ����?7mG!f!���`�ds� ψ/�$sD$��&��qVD8��L>���Q�/��tz $HL}���`p�y��	 $PH@Q'�'G���Qѭ��^�1q����j���8���֙���b�M��.��@� �OI��1!��w�X��	�XG,	��O��pVe�,δ�1��Ƃp���+��i0�L���d�'�̙�fkѯ��O_Ԉ��Ѡ��5��;i<[K<ɑjWs��D@�| -ʉ��#=�:���V'x���(�-�u^���`����ـxh��z�"~nZ��p
4Ⴘ,5�4 �L�ܒ�I��E�1��DN
�D&� .h���7	�j�C��'��	��O��|�t��~Fz�G�7��[ElS� �FљD�C���ɤx	x���	�D:E
�O�w� �M��t֔�,��C�Z`��ɟ!`[�y��I	H"�s���
O��\Iv�R�L����ʝ?������m��>Ʈ%��	��٥�t�I�㛼.~���ѬZ%lW��(���� 3��bᓵ�j�-ƼV�v��G�J�2�f7�N�^��Ě���z(QUn�+�����5�C�+��ب�"W�C�<���?8��F��&b�z,O��}��Ji�����6LhݫRGb����q "aӄ ּ(q,��ϓ2Zr��8�6�Sæ$���@�i�v6mͦ@�Jaڐ�A�3�Dz�H�)&vт_cʬ,���8V|�Y���4��]"��ڂ���ޚ��O�ư�G�Oe��B���?�m�������7�(��A�G_�'��uȲ�V�\��᛻(�z����?-����N�c�/6��7j̒a���F{Bq�d�и;#���L��6�D�E1�� �B�T���%�Mç��F7�BV�Σjrݡ��}�'�����YgnȲ�hNm�8;�4�~r�.?�Vq���sC����6g�O���6cE��mχd.��
#�?/�V��'�џ�H��-k3򁘢`��tY|�����''���9лi�m1�&��R�pF}��u�z���9�I 3�+%R�Ч�p�"?ٶH���'�H�J/:��%i�֚\M��l�a�'�$���zG�5Uc]�f��Ap�O� qST�A�HYB4�2'J��Y�,����I��Oz�C��)�8�TB���+��92�	��ԧ4�d@��լ�Mc6O!�2����S�L(���1&oyR��V�~�����*�8{��Y��C :��˓$"|�0��G>l�h١ѦO??h�H�ҩ��,HҠ̔���c�ЧD������<���\�oɺ�x%/���(\�wL w<d ��ٷ"�B8hƆڕ<G�r�K6�hM�#�i�d��/B���Qu��`�.���#����x�x��v �|�7�*�1R8T �=
�M�*�V�=Y��c�i+�̓ ��C\�=��㯄�_�,d!�'pD��1+�0����Y���oߜ ��)%�GK�H=	DK̐Y�Xcw��]hd� ���D��<I0�ΰ`�Yas���e���syb+O&�J�{�ڇTE����i��D��ɣ0��)�C,;D%���3+��<��&]�[T��h ���' ʈ��8
��4�A̨F��x��`�\�������(��Ph���D-O�^�ADy2���6�LՄ�I69�����Mj��,�48�jd�W�9��y���ݞon��F�ƀU��,bÍ
v���d+X�T��DeߗN��r�FA�H���1���,=H��:��'�"�PV� 
?3�!�6� 3>ܩ{'B��*�X9�V I	a'j]�Bd�Y�'ӈM:�F�,)��pr�P�RB��E~��z�ڬ27��(O0@0(���I��a�h@pm|!GI�fF�\`�ub����\6���2j֕A���S�(�?�!�aKʏi#f��_�atT,���{��QOc���BO�2;�L�c�o8|O�mi��o����O�6bd��˶v�p�<i��4��˓�J8N+��97܎���O��ɗ	b8��qa��qm@!�VBј  aC<S�<��*���	0"���se�2�	����	P��2a�ʹ{�
�z����d\�"��(���3��A��O(J,�8���;'~�I��-�]��	#�ƒ�S2��1f���J�21���o����3	R0J��<Q���A٠� ʠ;&H�%^�@��%�Z�&@�'�E�r�z�A+WW7R�|��t'h�`n&D��jDcަBj*����۶/��,cЪы��l(�����M�''
��7��~�q`o���ηb�x��厓A��psm�uF!��ޗ"&v4h��(iap����G)5�$�@9O�ВV*	�|�V�["Hf*��)�p��>QTƚ�6q|Y�s��0�0��i������'����l��)N((gE[>K+��b�9<��������屰�ПX���C�ʚ��=Qw�[�1���b/��)���zuC
B~R�N
Q�zta��4Dj�}�7�Ŀ�?Q��FR�nh �k�u2���X�teq��48`��3n>D�p��6U�\�ɒ��.���ï7)A�`Q���lYl�Ѐ$�tt�Q�N~҄$�p|��ݲ�������|�zyz�ON��C�I�S���`�I�9���Nw��zo��ا���D��s��ɥǎ�Ll4�2�=1�!�G�w�䬩��t�EH��Jvy!�d]5X��� J�CT�I��"�5Ik!�[R�tD����f���)�.�B��"t&����ǟ�t?P�ا�Ώ�lB�	<n�~�h����@^,���*�u�4B��<=΁;&� 1T�8���B䉬K4���Q/'$ڝZVaB��B���B�|�ʙ���;-A"O֕`�V�v�n��+ֺ0�"O�i�@3[��墰K&0�t�"OJp8�����v�;�)އ\Kx�"O���Ћ4ֈr�VZ3X�;"O��� �
�H���FT%��q"O8\+�iЎ^|@�Pp��6 �ؼ��"O�L`�h�Y2�h�L+%�X���"O�}kK�  �9��O*I}8�C�"O�q��D0l4L)��H?;|�5�"O|�{eFl�Ȁs�T�*k����"O��:���B� ��[:�4�r�"O�ኵH��JۺeR��tb�*�y�K���@����%3��u!CN�+�yJ����9���}��hqҨ���yb���d���$��%�Lۑ��y�J�(B�H�д�X/T�
�f(��y�%�Td8��/\�{���:#��%�y�%�l�lAS�*ׂ	-�x�ρ��yD��4#�e�eo�2F(���X��y
� ����9:���g>{�(���"O����K�@��4S��W�e5�pB"O���&��n!J�#c���"O��!6N�
�*�K�@�$H$ �g"O2����q�,�8 �R9�:t��"O�\[���$v.�mX$O���b�"O乫Wg��q��yK�*K���å"OR�pd�� �� �s(IR"O���.�
�\���HO�~��s�"O`����|�R��B'¿i���"O�й �c=$��&]�8�s�"O��[K�-l������J3:��"O:�;¥Fjc&��D��'*�:�"Oܴ��M�`A訪��[��p"O��unS����G���6"O$ �j�: 7�Ձ#5H�F�"Ox�u�Œ9�,�H� �
�ts!�$��.�ł��-5$Bűg]�=K!�ә}�(��&�
��+�Ń9m�!�$$�>$�b� ]�ظ*7�FG�!�Ė@��H���&"�)��$�f�!���O벌�s� $�4x�Sd��!�Kq�CDӉ/�T)��6�!�D�G�(����N\h���&�!�&q7�p����;;Q	9pϿ �!��{��� ��xllL�G�\�8z!��K���ؔ�Eq�� )�N#3]!�_.�d�e�'��eȓĊ�]=!��ɛj����T��B����cێZQ!�D�>=���pnſ��Q �b�:xd!�Ĕ�G&lg��D��ໃ`D�OP!�$;Xi��2b�%1���`i¬0V!�dQ�
�<��oX�h`��;ӈ>u!�$I2��T� �$Q�͈ (]�eu!��֍{�pX��L-<F��B�	z�!���*K�P�.K�t���	�O��>�!�d���h��OR�Z��a�M��!��S��eP�")M��E�0 �!�D̀���q%��vNi�,�h!�E�y���9�!��i7�0f�NXa!�$�0Q���g�Ʈs ��%F[�f{!�D׏[zڬ��$�65������sc!�$^#z4��$�@��u��,(E!�_!�镋F�>��10��B��!�$^�k�r8�d�T�
�0�/3H�!�dBRf�%"�O�1{�L�2��8.q!�D��8���!DH�O�xP"n��,g!򄒣i�zđ0,Y��J4A.��7.!�$��6�2 ��? �`�ٗ_�HʱO�=%>	��І`R�|1W�Ҳ~tE .;D���&�DR��ps��  �lI��(8D��9�&��B�0d��<i\Bɐ��0D�@	���':��`��1�"I��d2D��q��T%�@��P�%����1D�@!�j��[�|̡s� rɾ����$D�,���ߏ`jdx�q%��~�~D�F"D�#c�!�2��/ӘE|�(�"D�����U9K��#⏐C�~ ���?D��C#��'�Q��#	�:Shh�h?D�T�B�՝T�ad+�^�J� D<D��8�
�6�7�S�D��=��-=D���n[?�B()�ASN��qL'D�؃"^5��*���"ӆ����"D���@�ʙ-��dZ���=l�j *� .D�� \V	�)Z#�XsR,޹A8��	t"O������
���pѫ֊����"OL�"P��9"6���x�$5"O��"6��l�4!y0�_<'�D�"O��Q���I��ЂG�p���Kr"Oz0*ԥR�TM�x��O�*4-Pf"O���×�,�<A���X�K�JzR"O
iѨک}lP�7F\?~g�!��"O�q�%3G���A�)H����d"O�5YaM�'�b� ��"�e��"Ot@�Rc^)B7�Q)6nܾv.x� q"O�l�!��-M�˧́$o?Xs�"O�b+��Xs,��+=r��""OԌ�0 ��vl� ��͈�-0pʁ"OjH{fC�
�$Ph�L�>�� �t"O*1�#%�1�vȋ6솯�u��"O�jfE��s��K��7E�Z��"O"��(C�G8:��� O�0�Y�"O�qP�
W�QI�՘�`W�R�E"O�H�@�%!v��A�Ƶ@��4�@"O�%h���Z� Gę>��D�$"O8���d��P���3�&�b"Oh��C�I�����$�P>���"O<��J�;����)S!/�̐u"O���ޯQ�`���5$�ٰ�"O��7Yi&q����c�r�"O.]A 푋z-X��i�&|:y��"OJe@����! JSf��`"O�ta�cȰv>�|b�� 3�1��"Ot�q���+g�eRr�O�{{n="OЕZ�J�?n�&�_{^�0�"O��`WN��4K�՚���jH*1 "O2�F��9�rb���!Cl��"O�87*M�b��e�%��i6֥�"OT�0� #���W�^�kU$�XP"Ot0ɣ×�3z6X���ٱH����"ORir���=5}nH�.S�lY�"O|s�n�!^=	�m�l.ū�
O�7�M�#��Ʃ�*+��� �@�<�!���"T��Y� ϭYנ��3�ڂT�!��Q<!���u�IҘ[�.G�Y��'dў�>�"7�1Z{.5z�*�&L�	B5�5D�8҆�M�w>>l����}T�@x��'6�ayҤ���85:���=��ʓ��yR,�<a�n��`E�=O������y���L�H��D�;-�0(��
�yҁ���fH����6&�J���C:�yb��X;b�au�4"�&(��-��y�Ɂ;UBh��ޘH�������y���o��=9`� m	~)�%OG3�yRED*Ǽ�Y�+iasd���y"�	&1�|p(F\xX���a��yB�ҸC��=xb��a�������yrǉ;�l����a�<�f��y2.ϱ��<Q���b ���[�y��;Y�Z,�+E(0l�
�y��+c&Q����yFe���E��yRÞ�s��`��j �I���I_��y�װD��y�2hN����3Qϙ�yRf	-Y��e�U$up
�Ѫ���y���4�$�XH3P�P<Ptz�'��H���}�UJ�lJ�Ds�Ј�'��Uq��Ґar�Y�,Q=kF��
�'{��%A��8]6�S��Z�9�n�y
��� l�C
�g�Hꕁ��r��X'"O8�#�J��5���Ɠqx"�"O�l�]7%�8ʲ�I9Tk�dQ�"O^��d{�mb��ߙa�b���"O-��※-�*�6��-4Ɩ��"Of�Hp(]�Fp�����)2�"O��K"lb�*w�E�eI��:V"O����� 4L�R��`F�e
�x��'r�-0��D���f��#�k�'�L0�%T�LU��{��ޖ^`�R�'x�iҳ�)Y fl���P9�ܣ�'���0��Q<�x��c�"�F$S�'b���)6(�Cd�M�3�
�ۥ�c�<q� ���Z�y�̏�:8��M^c�<a�!�t�|��F9�.��{؞L�=)�$O�3g*�G��$PeD���N�<q�/F�	(��'A����%JK�<��n��3���H%d��H)F�WO�<��D�pc��N<�vԨ`�O�<I2��]��-\�7~���-�L�<y7#ӫ
߄��'��=9��iq�DOQ�<A��ʉr��Xp �8p̀��M��t�'�Pѱ!��"1����A���s�����B،Sv�H�M'��#R-
O>Ԇ�A�̢�(�M��2'�*���ȓ6 �i�*(nE�#Y�^�D{��'�R�걃�l3��:1l�F��Is	�' jT��TOF��#%ո>��E��'��H�&A�,.꜃���'/�����'����w�ڣ������#�)��'Jq*"�	�%G�)��
1總��'�V S�IK+�|����[3x8T���'a�E#���wDd��ǰ�:� ��'۲��2#�806q"�'.�N8��'�. �cƆ/_�����(O6|��'l4	�4,6jր��A۵5r<Z�'���#^�Z��-R%�*�R�'J*�*WBؒ�Ɲ�W P�R)�4B�'8�m8��ה]�<lصśJ3��
�'¼����ХMXn�N6P��%
�'g�U���A�|պi����6y���B	�'��P�q��"���4ʈ u ��	�'
�*��<]�u�G���1�
�'=�I��ڶL�j������Lu*�'��1�D��5uP��Ã�{*�c�'3�a���h�ܱ��	>6�QP�'όԛ���c��4b�%�"4�X��'V|d��#̋j�n�7#�]�� �'����$�蔹
�ͅ[�
X��'�t� ���O�A�6,��S����'�>���h\� q����B�Kbp���'�uhr��#\�)����%@A���'��}� a46��j��B%fv�3�'� ��2e\g�����N�b�
�'6�U+�i�r��p*ἐ�iъ�y�TX����׬A:X|T�����y�E�� ^Q�t��Oٮ� U'��y� ��V&�)���܂7�h0��J��yc $S$���a�,&�l�T���y�$�[P>�:u&���@�bJ� �y��R-6L���S�Ϧx�5A��Pyr�Ĉf���k5��AdDaP�e�<��m�6*� ��!�*M7�8���[�<9�-H48�t�P-�6�\��`CEW�<� aR���].�i2'Gؔu� �"O��c���Z�Jq`V+XKj`�V"O�x�sk #*!�iU��QA���"OL<a�/ü0$Wn�(�@�"O���H);d�K�=l�l3"Od����]�6�R�BՊ3�!�"O��s��-)n�k'�7"��՛1"O�IbWě	`z��p�Ӎ%gZ��s"O��1��M�f@FLKr�fÜq*2"O�Թ��^s�X"d ]��H	�'�.���D-xz�Q�
�<3v�
�'ۚ��L{|��J�)ʺ4d��2�'���f�Ϧk�N�#�.���a
�'[�`���"�z�jg�V/�\*	�'~�Бe%uk8��e&ڊN�n��'�r�2�aK�T�QH��y"F܇ȓy�k�.��Z��L�Ո^�F�.t�ȓ~S�LQ��C*l,p񙵌Z?;kb��ȓ���͚ؖsq�)�U"M�c]^ن�wj��ٌ
�"�	aBEpѸ�B�'D�@�$ز7�@�u�X�aj�a�'�αZ2j�52c,��J�SZT�1�'����Ƙ'`�J�c�(՗����	�'$v����0�޹�&d���	�'<� 15O-�^����Q��'�VC���±�
��r%R
�'����
8y���Ic�"$�	�'G�("$+��#����K����	�'n�1�0OD����զ�w���'�.l;�Հz��#�Y�s/���'Gd�@��\����0e�g�r$��'� �Lk-B�
�E�)G ��'<�i��q�n�ض)� �$���'��I�f�V{����T,N��Q	�'��[�k�]�2�+��EH�^� 	�'��<����
���v@;2|Y�	�'��S�ڰNޔ��/:���a�'�nh�P�M3�S�:f�#�';4��TL[-z�Y2q��5I�2���'��1ä�&v�������Gʞ�Q	�'��ѕo�:>��7���?� m!	�'Bh�w�܆@�R�"��K�9ɞ���'�<P��5'@�4(L�[�0K�'4l�R`��$rXP�:�H;P�A�
�'x4`���
1�%֋KZ6h��' b�i�.T�!�&��Ç�k���y�'ݞX��$�,N��̪sc�V9����'��Q9��,<��5)��F���'����u�ɌE��fL�uo, �'��}�g+��R$E��ޖl ny��'�效�/�wάŉ4���b6�(�'�Z�R��B}�A	��
5
u\UR�'rp����X�X lQ��P��*<*�'��t���F��y�.�s&Z�j�'�$��cD�/l~��48��	�'N̽�!I��*�K�E�(<p�A�'�Ј{�E�FЙ:��;j��'�
������ɀwHݲM��'�z��G�����I],,h,Õ�1D��*.�j����ОT���);D�X���6-���� �� 5��i��,D���M�=l�2�X��"��=y�,(D���w���v�����)�����*4D�h�4J�>Ϩ���I�uR`����$D�� �\�Sˑ�V�������6���@�"Oxͱv@��#`}��1)��-�q"O�����?�����/{�F��"O&4�D>�|�a���/�̉J�"O�Rb��.�a�S'BG�1�3"O ��M]�n�^�R`F�:��at"O�����P�f�����$J3��c�"O� �`lׇ!5�C�8 ��T"O\�{f�?*��*r!��q0�IQ"O��W��`���w�ąX �9�"O��G�	(�����/A&���"O�<	�I�j�Z]�W�;<�n��"OXPpE�FN�ܝ+�%���:�S�"O����ל;�H�ګ
Δ�Ps"OpC� �!# \1b1�db��Q"O6	y��=cX��3��g�4d�V"O&��r+B�#��r� �\�V�<y�<{Ƣ}��MN�F���AP�<a�$�����@Nl(���AL�<A��8[`��䈈�l���b��y��E�K�蘨��3k�8�b�J��yR���vD(�EQ�L��4����y�
�	R�e)��W�>��ۂ.H	�yR�S&|�*���#8���9�"ʱ�y�&N�x)G��/6���[࣋)�y��]�Ynht.�7H$�����1�y�+����\Q�i�WVU*U�M�y�B8T�	�ՅѢse H0��X��y�_H��q�t�ɷU�\E�  �7�y��D09���π�!��P����y��ُxlN��茆/�n	y"�#�ybLH2m�3� �4 �t Z�J�4�yr-Z<Kψؚ�E����b��E��yb����!Ώ��4C��yR�M5"��a�Q	�5�%���y��� ڔ[$M�8*�(h��ڃ�y�kӀJo��1whO� D��y�bԯ�yBeB`����Mш�����+E�yR��b�����
��fÎ�2�A�8�yrg�6o��`nT>�vx��Ã��y��"΍3s��	����冥�yr�b���R�,��p!چ͓�y�f�o(~93�Z�u�$
�\��y�a�U��G�k��ԋ����yB+�
f0I�A���\w"#$���y�MB
�z�Q�j�/G�% ԋu��'ì�p��E�A�&��!^>4���'��.�t�x�r0h�&b��P(�'$��rp�G	V��tP�2Sp��'��3�L�'(�=��f_�7���'W�Q���� Y$ ��,��*��	�
�'�ƨ �V1
*�yƇ�#�z1h
�'W��[DA aT��0��r�	�	�'ְ��	OD����r����'h��`�̛-�(�h��%EED��'Dq�,��L�j���B��H��d�'Ϭ�p�F0�����M vO H�
�'Y@�Z�n��T.�����ٷ9'��
�'��1���v�p��N�3[�Xq�':q8s�ٕ���q���N�t!��'��˃�[�d��30㙹J� ��'�|ъ�%I�s�\��W�6�L��'��T�P#�)�@��$&A�Ps�'�0�	q�G�9�����E%<������ �a��R-���	*�'|/(���"O���u��|ʊ8��	�-���"OD0�U�D?4٢�ЈV�Ac�"Ox����9� KF�G�t���5"O<m�q���r�<9GO�S���"O4TڥeOv6p���'5;��!"O>u*�!`��t�2B+� p"O0�I�)�S.�|�"˓�W!�a�"O����J%�L��#D�"S�=�`"O��3�lT�F
Eb�_��""O b"�?VU�QҤR=d���"Oޜ1���\���skEa(ڔ)�"O�PG�+n�ݢ�	�Y�,5xE"OTt�Ul6��DAbI-br3�'R���i�J�>L�\z`�B�od���=D�l��C%��@T�� z )"S!D�̸��Å�	�ѡuLĬq4a=D�L�gY\غ����2Z�1a�7D���J��z�I�S�Z�t@ڵ�9D�D�##�c*��ҠjҚH�x v�5D�l�� 9 =X��M1N}F-�fK4<Oj˓��䖤q��(�A�*1�!	Ӈe�!�Ć��@����P |L���B�82�!�$�f�0tFA�*(������>!��@�-���@��3pz����ɋf!�dL#w%�iW��W���Q��]�!�(F�bp����&E�pQ�g쐅&!�D�4b�� ���N?"܆m���)��}��d����e!j}1�l�6!���9�i�<	��hOq��Q���U=J~D�C���0%����"O�����O�?�P7��--;h���"O<�y��U�w�C��W5b2��"O4YS����N���Ѝs���Z�"O�HC�o�7&�T��!�m��`1"O[�#��cv���
]��}ж"O�<��h�� 5�R2l��|{S������B�Q�[�	̺,r4�ѪR�RB�/V�.Q���V��n���C䉙^p���2�I;`�(���مC�C�ɸU��x�Q�ʹ)�� �7�U2�C�	�*O��F�?��9q���k �B䉻�䉪vg�fk���7�TO�B�ɴu0�u�$�7��� ��M���$4�\����^�(��c��Z�6�`�I2D�415NL�R�6)a��=F�
	`�f1D�H2�����
}*q��F�b�#+D��IR �2J��3˟
	�3�&�O�C� Y%��7}rNYh��
�$UF���V���SE�]��##��(�؇�H��ݩ�ᖍ��@#� K'F�h��ҟP����*f2�#�'��.r�Q#V<o�vC�Ɂ��у��)���T�|�B�ɘ6&��	#�R;`����B��d�BaAR��y�.���J�FB�	c)*(�tH��G��#�S��vB��1i��H�� t��db'�ѧ)�j�O����?���V� �Gb0�*��?`)��'a~R��1F$&��PO�[���2��y2��
�|�r#�F@nq�rc]�y��[31�&�	�DܬD^ڡ��I��y�.�
,O�|A3	��n$~���d��y�cV2ij
���k2]	�	���y2*M�R�@4RT�G�h�� ������!���'
L���E��r�S�	:$)����?����9�S�? 2��� ��P\��jJS<xp�(�"O&p�$�4��	R�/U! �""O��Sd �$U۰x��]>-��)1&"O�l�0
�?q�kX������
:��'��O��I��Eȹ2�쉸pF�A��p�'@��`K�g��5�"�ǿ� ���x2�S�i�ĘR�$=�A3��V���<���PF�J�-H�]�4Z��a$!�dR�5b���J��;�h/13!��17*�5�׮oӘ��ȅ�!�ݢjj��iÂ�}�:�{Af��Tџ0D��D�z��'��.Qzڜ+�O���y��ȀK��� 'R�6p&��th/�y��/1LɰB�.~����ϔ��O �� §�� �W�8d��H���ܑ~�ܨ�ȓe�"dhfj� �H�	�� �f]�ȓb-(SD��(�$<A��/32=%�XE{��tdZ�,i%�%�K�9<�b�fC�y��I�t�΄��f͜#�|P&-��5�&B�ɔX���צѷx6�y w@�+`&B�ɣ6����I�^t�����s����hO�#<���sԮ�����e������E�<�E�M�M��P��E�B� �a��e�<��KJ -��PP����(Q0�(Jb�<����7Ap�UÓ:3Z��+F�Ne���?Y�'P�;�ꌊX�D�dF=F>�����X-�%��A��kq'US`桅�mP\�d�9�^��g&��Yp%����	�m�Be����|3����ʯo+�B��1�,�c�E�!Y�� s%�ܾ=-bB䉶$���um�w�̄"�+ܟ%����D �;�{����`�"tEۚi���-��<E��GV#v3��829�°sB���!�$Y04Gz)�U$1ܤ��f���q�!���`��N��o��E"�%���	nyr�)�
N�R�x�Ҳ��8�.qr%��yB�ĸ5��`�61�`Yk�L��y҄�Q�D;�m2S0����y�`��j�r��B�T1[�05㡃����hOq��-��J�k�Z�I1�F��25"O>�A�D�QiT��b��s}BT��"O��{��J��(�@���~e{��'!�$��F���9ŁP=~�$;��݅2�!��_���:D��"5y�hY�j9�!�$�
_nݐ�T>+	����J<]�!�DԜU#�(���aXMم��w��Oң=��j���#ߓb��`�q�Pd�E�"O6]� ⃇M�$����4m�e�g"O���wb����rtG�!)B&	��"O��ve�7C1��FQq�d��3"Ob�)�"ŧc���8�$}8��"O����ΒBf��N� ���"O
$!&�j		�m}�-@�"O�$4���F����+{q2�¥ 8D���W"W�1OdA	���MK�����O`��<I+O?�BadΣ�&4���V�7� ����c�<)�՞m�6�G�0p�����a�<A�IJ.O|��2�O\:k*�$�X\�<qj3_I�q� ���|�<�s��FK�'Uax���<�{t����p�!�Û�y�jԧ;H�[�eK�&&L�P	¦��'ў�OZBPrC��=�n%i%�N2je ��hO?�!��kC��c �+Pe��kdb|�<��� p`�f���L���p�<� t������y��W�Xf���"O��R�U7�pQx��ӝ��
����O ��$ �[]6��p�X,D���1.Y!�͒;*Ҭ��ʙ*B�$)�3��NU�O�=�����>ki�U; Oʫ6l0P"O�ȉ�o�J1힎-�b�`��M�<���x`̤��+A. �Hb��K�<y�̠I��IVnÁ��Ӡ��C�<Y�(̰]�"���J?1i�ʘb���?�Ó=>��P_/��S�f�	(J~��ȓx~��#
� �:)QaJM@�Θ�?���~�eK�)��})�,�Wc�X�s��џ�$�l�����d�U��aBva�%�a���Ĥ	�ʓ�?�+�8)C��ȏ	�b@��4Q���!�h���� 2����FR�,]��ȓ8���Y�cX�%A�	� �(������ry2��nE���$	��pC)�5�!�$�*6t�K�㖸{�|-(WJ޺G�ўx��Wt ;v��p��U��Ƒ84P�D{�OB��y��D$C򦕊�����؆�ɰz��l�gE�>6:���ߊ=��C�(Gx��`����W�"��, ��B䉏C�H�s�]����3E*�H�~C��:�"]`��_'�p�8�혩>�
C�ɷ˨e�"A6�d��#��d�&�=açN̩�s���
p�Ӫ�D_����N�����'��'��|����
^S�K��l*��c1Q�T���8p��V(�5[�Dz�!!9�B�	�{2���k��������ý�B��*r�.	{A� vZ�AWoC�EpB�	c��PXc�D2$޴!��eY�C�I�|����!b��0�@#w��C�	 +5Ӣ/K�A��Xp�	�Q���|G{��'���HG](U�����n���)�q�!�$�%p&�Uj�/�o���/�(*i!�dZ'>��X����<�:PQ���0eg!��4R�,T�NZ�b���"�q,!�9g���e, �{�pơ�z��d#�g?Q��!y����g�8|�$X!(��I��?�}���E�F����P7E��#�I]dy�|2�s��A$3z��B̖ �p�X��vy"�'}a|H5c> yyO�6
�@-R,�y�)31|�T�DBI*;��In^.�y�f�pߒ���Ҵn=���sn���yR��(,dQiD�h�$����?������Op�g�'�"��W��u4x���b�5�&y@���'�a�T��I��} aLl��X�
!�hO<��$�(sx �o2m��T0{r�	`�'\�`��I@�,�;k$P��
�'���W�]�3v��R�M�f�`��'V"yk�D#)|!��ŧKV2���'�L�G�ӄ#N}��k #pK����ľ<N~�=�֣��_���Aǆ����;�@�u�<�R%��[��aeꐴ/��+#��g�'a��L��t	\ms���b^�9�A��<����"�z�x��U�s\m��I�	[i!�%kr�4Svc�L�H	�G�
�!򤉺1L�P�j��{ͮ����I$��	O��(��m(��vL�鄌ޠuO҅� "O��b<b>H�R�"I�؀�"O
�z� ݅*aPjsB��(^��Q�"O��i�*��C�R9�p��'E|İ�7"O���#�\�+�,�*��5VHfp)�"O�q��DG4�( 
���4=~��"O� �1ѡ@,E5:`���Ѣ>"x�"O0����yżhbCdK�Q��1�e"OuI�.>h ��!��(��t�"Oh��!ng�K���/(��A��*O����ސyj]Q7읺C���S
ϓ�O�(��B�W2�� �:|��d"O��+�N�n"l@p��O`�D�P"O��
c��>W&�a��l��y�PH�g"OJ,p�@�%�0�lH7?����"OA;G��vVT��*
;B�S�"O���`�"�z�T#߰E*����"O�(�)_&#�����N��Qw�'��|���͌4���ӡ(��d���B7D�x#w��9�r �DEA�q�(9��f3D�`a�+�Z+ �l�)�5�a�/��#�SܧN�̡#*\,g�
�
�Z�B\��+�v���*�>�z)ز���{�H��ȓ@� ��G�S�cH�Y�AJسX�l��0���s�� ��
e�3����ȓ6�(����oV�:�N�%bl��ȓK�6d�c�e=����� s�-��6쒼a0Cíf��;�D8\���ȓx�H-Ґn�]���E�V�z��ȓ>3 ��siG7uEr�"W�T�W�pU�ȓ%�r�auM��|�e��p�:@�ȓa��0'!�:/�т���R�A�IƟ�?E�T�S�C1����5�IAԗ,�!�D }4�k� Ë�0p��fצf�!�ğ�?�<l��MW����A:H�!���|��a�^/b�Xh5�B�!�Nhq*����A.kx
�I�!�պ1�fy*hT�88rc��8�!��P�_���W�[ ٖ���[5��'��O?}�u	�o)|u��@�t���#�/�w�<��# 3È�-Z:A<��uO�q�<��lY0ov�-B-̾MB�a��U�dE{��)�pGd A���!.�|e�P��=G0C�I��� ��mV!�e�הi+bC�	5~����ň0�@� 6n��|��C��"e����	[�:a�7ES�E��C�ɉxS���!��Y��!!1�B�I
V�)Ā��V�:�*�n>GU�B�	K�;�JG1O&
p�&��WXB�	�e��,��ĳa� ��Ȳ��C�	��lѩ��VJA��A�
�_\�C䉉Hpѣ�D!���G�J��C�ɞ'ݦT	EL�#p?�p�ˇ#eN�C��]�tD 5�+T��(ՌG3mjC�(#�,�`o�-�n�`S	5#	:C�IL�(��ƻ��@ �5wI*C�p�h(�"�Ͳ_��	�A��dC�I�\>(�������r��t��C�&b���a�<KբT��`@Ns�B��u�e��̩+cҌ
���9WJB�I�16 �Q�V���٠�j��r�B�I*@@H�4���k�hA���B�	��r����U�6m�H�f��oO��d4��T��~"��>|}�QB�䘼3�P�h�L�
�y�h�%��5�
+FC�
�-�y��[	��R�,V-�0�"�8�y�M_�M�b�C��;0������y�']=����Q�-bL���[��y"�S�{��l2q�>&�&ŉ��2�y��=�|���!~:� I�y
� ���t+��4ʐ�3�!�<#�]��"ODف��!)�hY�`
e.�adS��	ٟ,��KZ~P�p��.c��Ȼb��%6,C�I(J�L	�f���j��P�A�'�T��3�.�@L�g�	�_w�<��!F=���Uz|4;�$�!%,0��	�8"�L���C\��e��G�<��cКHeJ��ȓ�����P	"L�KTBQ0 |؆ȓQ���*B�X�C*����R�+~v�&�0��IC��س�˫Oh$)��q!�&D��  .N�F᪨����62��&�O�#ؐ(�!���T�kݟP�HP��Rk��scA˂2l@L"#�>Nʡ��<��*��κD^l�q5�MEt`���4�\lA�,� L�v�"�Ŗ'/:J%�ȓ%��iP'�E��y3��+y�����s|:S�Qs��5��D�#! ���;�RY3d \f��ٞ��D{�Z�HG��&H� &� �Y�B�9R�y��%X1Jܙ�1QHT�+$S��y�����g%�2B�d�dFV�U!:Єȓ�l �J�;�89��Ls�QK�m�<��M� q����G,���Uf�<A���l؜IE"̟]{��I3�Y�<)%H\2%A3��H�R�E٥�K]�<��/4]��9�d(Ɠ$�Z����TY�<��m� ���b,��;%a�T�<�3��G�A+��18ld��
�M�<��L�) ��"�30���s�R�<	g␪4O�	�`�G�yힵB���s�<Q�#ɫ7$�QP�A5*9�� J[�<���G.[̸�x����@F2��Y�<�7���R�"�³	�+��l�''
M�<Y��K7V �XC#��� �4�bW��^�<�gGS6| �12�����r�Et�<�Se��}HT�Y�JX���iBtțm�<i"EHL�M�g$��
��I"��Q~�<��g��P�P垇0Y��ᓥ�}�<�H��vD҅f\�n�q7�@�<ɇ�	�(4D5S��J�Kt0q)3�Ve�<�.	$�����L�7�����WL�<��Ŏ�H�����тj���)AI�<ѱC��x�@-q��QOZ��'�MG�<Y�,4e�\��G� 4lX��N{�<��E��IS"���L���w�<!fB�a9)k���+bx�H(�lPt�'Na�R�}�� �J�����+�yB���Y�x��_�vu���@
�y�GKf�z��E�{�p4L�y�"�[��bYNZ�a��O��yr���Lx,�c��(�"��y����t�.�\x��5q3�F��y"���0��HH��
.hD�� "K�yr��jZ����H
6�*�p�����y�@� U5n�K5e�d�`���͕:�y"%�I�X��b��V(�`�]��yr���9p��S��R��0�y���p�x�BXE<p·'��y�	�=J@�q�E�q��j��R��yҦV"j�,(2j�h� �U�
�yb�/E�|���\Ud����M�yr��B��=��E�?S�"���K-�yR��?|d�S%JH�s�a���M��yң�� ,#�-Q�B�亠KN��y
� �����q�ؤ"�&�9n٢�"O�]H�d��Y�<�3'ܡr HPq�"O�pe�%.vȐP^5��!@��'e╟8���JY0���
��P�%D�0B3��:rf�q�����Q��=D��
�Bґ"!$D:�L��}��H	8D���CI�TItH��>fς�Sa�4D���&g��*�����ݖ�	�dC.D��P�����p��',�Y��K-D�h�!��=@`��Q��+lp���/<O�#<�m�<f&���L�?�l��cKt�<q�͏l/����û�����j�p�<q����Gc�q��ɑW��T��-Qi�<�qC�Y�I�.Syb��S|�<������я�Z�xաQ-{y�'Ua|R�>0�tqP`Ǐ&^A�#ſ�y� +� J#�?����NB�yB�Z7*@#�����Yr 	5�y"�O�J~�QAa͐v{��[��y2b	 /v�`�AmKh�b�S�ހ�y¥7+o��H�δa^F�����y�%Y�z<q 盒H���Z��&���0>IQm�F���G:Tk8}
���0�y�b�%T���*T�>G�d��/��>�Ogç$L���·O���"O���<b캕.�,	�t�"O2����7P�CM8-ٮ�"O��H�	6-���3r�R�(�<�"O�ITM�7��ز3 J�PBԩc�"O@��jK*=ژ�jRA�/����"O�@�/KXR8�Q����-3 �'�1O���#�&�|!�a`�"u� T*"O�DzRi���Y� 4O�̰�"O5X�n�"0��Yd�C$7�Rؐ�"O�� Ǆ��oG�QS/�
�b�"O�\q2苩F�r@�u�.c�v�"p"Oн�Ч��6�C$�$��@su"O��	a~P�j,e����R"OpE�I�y�ꝲP���z�>8�"Od�#L޷k�^E�����Ub�"O2�D��:�ܴ�g	�|�G"O����G�F��U�V(Ss~]�"O��cWؽ(��ب���,l�à^�Ԇ���ar�<��oР$YD�V�m��C�?!0L�9BHB���!i|�B��1qW�-B�6�J����H�D�nC�	��Lܘ���6 �Bk�6?�C��7Rm���7h@;�a�$s�C�I.+���ȕ���٘�Ă:�C�I�/^�0����;1L�~g���0?!�LH�qL�Y�c��$b�`r��d�<e���,�S��98\�K
|�<)��AˠtbQKʜ7oЩX�DMx�<��DD���xѶ!��!{ܸ0��^|�<y� H8v��ȓ�M�!v����̞|�<�g�h^剒!�7`��$I��{�<�T+�$>�Mb�&���"(��Wm�<9&$5j4Jؒ���$B��i�/�b�<���\ ��{�i�x�v��D�\�<�foǞQ+Ɓ:�G��d�&=�Ō�V�<A"%]<�8��� 1}?xp�AN�{�<��eC�R1���"�6��:V�Eu�<Qt�5Dڢ���ō_,�|*AVE�<ᅮ� ������kM���ǈ\{�<� N+�b\�drRi�Ģ������"O�a�g��<���[,%��\�R"O�Qc�J�U��C��=~,�u"OҬ�s�PM��	����.Sb&���"O�I��ƽ)�� �ó_���"O�a���	P��Hӈ�)H,ֈ��"O Tz"�>H�TH4�#2���"O@ ��ץvM"�f@-z9�"O��8/�l�% �;6�tĉg"O�ИQA�$Y���cƍ$v�)��"O,a�	�G�"�yR�@*jGx���"OX,�w��?�,,��L5D��!a"O�P�*��*��$��B�q@��B�"OFxp$+ծ$�V0yF��fM�"O�=q�V�-�u� ����Y��"O�Mq�'ŽoH�	�7��j�"}��"O�r�dגq�HA�O	�;-jyy"O���b�6��
0(ܨ� �Z"Or�4*SG���uZ�I��"O�-���I�d/���	��p"O�I����3�X����S$<�0"O*�B�΋c�D\(�b˷"V�YS"O�\� N[#3�xH�n�0{R2囶"O,Ȱ���A���Q�G҈%6L�P"O�UHp��4h=���WdB4K�"O$���H3c���#�Ꙥ= �Dj�"O�`���4岦�nc΅P�A!D��d�]�f���{#l}w�ә�y"ަ7Z���"-n`���F��yR��w�2�s�j��'Pu�F'U��y�E� a� 0H&�E�	�bh��)���y�*��uy��W��D��%Gѣ�y[!!�ezC����\ys���y�	ݗA�p���C�$%"0{�-���y˜*cZ
�(߿L��"a�7�y��֮N����b����� ��*
=�yL�~\�x���C�T��b����yF�F��z`@V�J���"���y�!�!R�Q���i��3�aS&�yr.M:LT$��t��f�X�b����yr!
�AB��G�\�(�� X���>�yb��!$�d��BӸ� ��RJʭ�y��1Q���1�Q�CBl�,���y"O����!@�Z8J������y§H��$���.4u֗�����ȓ8< G)�6nE6|q�M��Rh���!���;q�ݗ��pQ#�Ǉ0H�ȓ3|�re�#J
��*_/:�P�ȓ:�4]	̓�A��x���X"i����ȓ~}��,��0��.�0�$@�ȓ|<��c!OH=o�8�u���\����ȓ�JUXd��P^&e�W)�܍X�'�$�A�d�/6T�`Ju`
��`S�'Q:��g��r�r�B�ai�'��h��cB�$�61�D�_�bH@�P�'.�a4hθY�tt7�Ԟ0h����'q��ү�!N�d��fʅ�6�H�k�'�<�@��	)�RfՐ0����'���h�#�!�fl1a���/n�<��'�L�a�%��H,���F�"�����'Qz3+ׇ$�E��E�:f��H9
�'�4)�R�.<lШFhݼJ��R	�' �3�l��M���C�(��p1�	�'Cޤ:�,��`�y��A<������ n����]R�Sꛂ\���T"Ot�j�*J�Z��Xx�h�X��Ke"O����aJ�Zu��#��
P�N�`""O܀�a��.7��������"O��&N FGb�0��VG��Q�"O(���G�-Ţ���0w:�|�t"OL���AA ����R�P;HH
�"O.��� �)����eV/�y�dg��p��يU)H(�� 8�y���Y�<�0LL�#2�����
�y�ߚU��$c�ϝ"���8ģ��ym�7Z<�Z$���c���A�*��yҤ�5l�lbT��'aL,D�I��y���?	�50b�տh|
��v!5�yA�-W����:e���5(��Pyb���b� � �Y'dYt�~�<��hֳ'� �0���6I� ˕.b�<�l��Vp���l@�wi��qr��E�<!���+Z�p ݛ"]��;�
C�<�J�}_p�׏W�"��Iso�@�<q`Z�C��rv얆it,��E�<a���p��GC)TnXⲢSB�<a6�[$(�F��.����	x�<��䘻�@���$@e��!F/L�<!WhҖ�k��O?&#zU�&TF�<�$��<,<c"́�0NFh�wF�W�<��� �!�0hw�,~�T�s`E�Q�<�2挹�h�R�ʤ�����D�<���-�����O�]ܴ���HZ�<�+Ӽ*?h�$�#VaDek�<Qb	G�M�-��B���|�+��h�<��E\<������9�J�<9Ĩ,�^IB1jŝm̾qҦ�C�<y�끐/�PZQ'ۜn)�VC�<Ya���Ktq�
�?$x�9A��}�<A�Kз��M�B�/7��#�a�<)��_*xΈ!�Ȉ�K'����cW^�<T�˳D�Fy��͋}��T��O�<Q���N�:Pu�Q#;bR���H�E�<�w��g��z%�"'�$b5��@�<a@�˯fd�h6���K��G�U�<�#�w��E)f�C�{����&MK�<����r����s���1�sJZ}�<���\9#� Y[��S�w�
q��"_u�<q� ? �ҹ��Fےqk�i� �p�<iS ���:2heJ�%ӣ��h�<������ G �H���Z`Ab�<���Ec�B�qwf�aq�ec��b�<�d� iBY��@<H�����g�`�<�b��Zv"ܚ`+��Ux�dF^�<a��Ԙg�Z���MΤ(^t	�«�c�<��- L"�d�F��.=@
0g[�<�5�٫zcΝ�b핤Dk0��%��~�<I�.к?^αH�!'z�f�i�H
z�<�A �@L4�Z�A�.`�>��pC�y�<1�k�a�E�&o2�=* 	�P�<Acㅕ_�"ų^�E�v��e��B䉃;�z�Cׯ<�Dc���Y*XB���n�0��
�*�#N�1�RB�	�}@2ਂ��8Y�1�@�76�\B䉴6\�]#�`�����m�9jT*������9�E�:jT%���6v��ȓtd����@�c����s�O2洅ȓ&��@��gZ@���y���S�? <�� ��93R��,��,&���v"O�H�`B�@�FmЧl�)j|Fl��"Of,{�+ [K�D�+��,hn�h"O�����V�6�k�KA dSY�S"Oc���+j��Tq���xԨ�Q�"O��bLQ ֠8�h�Z�XPQ�"O"P�W
X�0�f����ܞЋ�"O^0�t�ِ$���*��Tr"O�y3/ɑ��0�UDօZٴ)�&"O`�Zg�Y�A����e����"O�����DU���RA��&�渋P"O�(a%
8[�,h3 ),���ae"O�����'l,E�u���F�B/S=!��H�o��H��o["`r�04�!�D��{Ɉ��'ʎ����U&�?~h!��A�;��,�Ł���(Q��N`!�d]�]Ҁ�c ��MY4��N�!�dҨ;<̉K5��6άQ���9"p!�d>?��h�#�+̮��'ݼC~!��37��1'��]��u��'U!�/��� f�̈GxF����]�!���
M�`����f��5ZƉ�2�!�W�8� ��J*t�$� OV T�!�ċh/~��f��D�re�X�M
!����Tִ�R�A�0;���A�Եb�!���d��@��iZ�d����%Ձ\���B���(ӕc@(൸�n�y��S(�`�sf��L��aT��y"�J��x@̑�ND���y�C�:W��0 �vw�!ݭ�y�.�u�J�bT�V����"��y��[�&2�9��<V�l�AS��y"�E,1Ԅ��E��Ic�Y��y"[[m�s��GC_"H����yb�\�I<ʡ�F��K��XCeIP��yb�	>�D�O�@X�m`�dH��y�Nڡ9j��`�OW.h��#W�y��ڀ`j��p�랪A����ȸ�y�F� sI�ݳBͯ3�:msR�V��yrm�y�=��=(��X��N>�y2� �!�)��� ����'��My�J?!h�p�>�j���'�<DA�ɜ 8@�H�$��m.���'���l�?g��Y#���_��#�'M � �Lv�lT8�H�]@RP�	�'����҇�EVP�5i��j���8�'�ɐCO�X�nl�D恴�ܘ��'0�C�I U�x5b�`��� D��'X��õh0eP\���ۭ	H���
�';<�P�D?m��2c{8�T�	�'�y:2!�D7���I]�,�	�'�0U�C]&�i�
W"Eb��
�'plyBm҉(�V=Y��Cs,�
�'a"�A�F���〒�	�e�ʓa��	CV�R0S�����T�V�,���K��e�����̜Y��]ި��M0���e�� $�t����`����LL]96O��5+T��2���@z4$
%�N��J�2��L T��)�ȓa� �Z���M�}"V�;W4Nԇȓ1�0MU�J$#�
Q��%��=A|��W�~��2�.?i����/��5�ȓj{b����U��A�aT�L��5�ȓiZ4��Oſf��DQ�*�T؇�S�? ��0��ݒt�p9��B�g�\�S�"O@�%�H�?Qd}�v�L�Z�{�"Oډ�T��\���X�D��6���;�"O�Xピ5h�<X���v�,P��"O�}�a��F�>�
���-3�)ӥ"O,}$"�H@	(`(A5G�X�"O��IBo��slDehcf�KL���"O,@˴��%	$L�y5C�-�p�f"O����6rD[pAÖy!���"O�l���	�;)���&F�N-z8 "O�uau��<P�����&n�"OR���֫)(m5��	;�\Bq"O���i�/�Ҁk���,�0�є"O���0�6C�����Jǰ��t"O0�{&�('�`V�$�P-��"O�傐o��j�|x@��:W����"O"m+�T�~a�Q�)K��D� �"O�MV�
p[�esvo@�Tq^<��"OP�#F��A�$N�v�.q�r"O��#fl֦
�cWH�'��}ғ"O,�#���H����+c~�"O�H2��6���@�3Hx�}z4"O}K��B�,V,���1>n�E�P"O���@�*��MY��8�@G"O֌Y�U@���.Y!F�p�"O�Չ5�7���c$O I�8�A"O@�3��� G��R6��(;����"O&��֣ *x eb�)\>1���:�y�KD�nD�D�ʼSvd	�2�yBL�9v?�����Q;d%��K^��yb��y�r�*�Q*j�Ä��y  �J���]AbxղS%�"�y�EL�8��	��Lڼ@`�A�ᓺ�y2ɰ �PIZ%�M2����R��y�)�P�ly�ׂ$/j<Q%�^�y"�F4oWn�g`�.`�k$Å"�y"��L�41�wd�+\oҤKd"�2�y2!IS�`��Œ�h�H��$Y��y"%_�ibD�A��W' ��`[�y�cP�yR6�K��M-LAa�[��yr
�KO��@��ML
zx�T Q�y�'	�Q��#TA]�[QV�q�α�y���?А$�
Ü~����Ad��y2 ��*�q����}K,es��A��y"��=?�*��DV�z��$�E��#�yr@�����#A�P�;"�H��yb���7��(#�ް-@��f���yl�%u�~$�5�)v�(����*�ynDҒLAe�H$ ��y��+���yb�X
t����;tĀ���Q�y"��?
� ��@�yJ���M7�yϔf!,q���7VH��Z��y�a����6�SN�P�p����y�"͞#�`"֏8:��b���y���>[^T�9�d +0k�x�S�y"ˁ������H5`��ˢ*��yR�y�=����XW&q������yB+�/,�D+��[�$�8a���yb͎�l�{ ��7e���p甈�y�h��r�f���,YP	��
�yRA����u@ �0T	A�����y�,ΊL�0�"β)�Qg ��yb�GBނD
W��f����j��yα%d�<���cM�8��ሬ�y
� ���5!�K>rB G2�@U
!"Ol*���U����C���:]vQb"Oʸ[P�C*"��= ��q%�C�"O�� ��#ߠ�q��c��$:w"OHX��м͘���74ݸ���"O ��A�M���1�D��2#~̨�"O�-���i lH��"@*k&��"O,Ms���F�������OW�T�"O�@�f,ڣVsZ�3��'C8�h�"OP����5,�h��o�v6�	"O�)H����z���n�!'D%��"O��⃇�5#���p.Ez""Ot\�P�� ���Г�T��+ "O��S��f2����&DZ�9�"O.QU��+ީ0�-��C�ً"O�J��1ܸ��2����"O�4�&��63P���0�U��"O2L�iGYl���@�< �X|sg"O,�"c��.W�f�I�΂1�̴$"OP�+��d\TͩӮ��|uqE"O�"e�	�L���F�t��H"Ofi#���5ȝJ nL�>�X,��"O(��BC�F���I.ȑc���j"O�JSkE�.�@(���O��	*�"O։;��'fxBM�����xf*O��o�<8����#
�d�Bu�	�'���0���?T6HY��EE�/�(�
�'F�3 ��X�j �²)����'��Mɂ��{��!��_K�d���'V��N݆f����T?�|�(	�'�H	��]>�	��ڏ5��59�'�H�s��\9�t`aL��)�����'�^ ,;V��1xC�7�����'���1���Vر`P`�1+Z���'�XT*ͅ6=	 �@UȒ�'���'>jA�P����5�բͿur���'g-9',P3*�� +�������'٪��1�I(t{L�H��^p���'K4H ���R��t�ٺ0&D��'��xd�Sі�D�)-1�Щ
�'(R<��KQ!5� �Yd�['�ڼ!�'�v�C�^K�Y�#
��J޼u0�'8��@�����B �3YP�\�'�:Q�R Cc)l�s�eR�~��ah�'�> �v����TB��ݬHh>��'��L�W'̔v	�Y�!-H	B�J�
�'rDY�g�'F�F�"��M?Kz�K�':Jܹg�2P�ƴ�`OT76���'��a �+ؕb�H�{��^� �f�S�'�<����Nz���ÁF"88��'O�XF$�,1��3�ȍh|�	�'W& qqeO�[��a�o�;Y"P	�'ŴP��H�0Y�X,ٵ�O��U��'�T=�t��\~�au,��'c����'I�Dʥ�C�Q(����&����'Ӟ�)'D�j{-���,5hl���#�޸��6.5��i�,�=^26�� �i���M1LuvQ�ĥ:@��g[\�8v	�V���W�^�{W����zy�$bW��1˸0��'̦Bܪ�%��D{��D�@wI���V* �W# ���Y��y�e�S����C��V��Y����'jaz�i�i��(�%h�*R�� )CD��yB�� YJ$1a�0H�r������y
� |���.%F��cǒ�
����Gp������*jÏ�P���.Ӕ��2gO$�yr��/��<x�(ݐ'"T�b�N �~��'Z�T�4Jߙ^�f1���@1F#T<;�'�9(�Au�ؕ#f�[�8@y��'�JIx`���|!!��^#0�dI
�'4V�H2��>|����� �~�(�@�'KrXQ��b�����)V6q1��
�'�2�x��gq�!�6ab��B�'��E�lDJw��#�çZ���R�'7��KS�D�~PX�P袘b�'���w��$3����S&JC�y��'�D��^�]�T\�m�7�]��'ۂ0[4f�>o��zu��DāO���I�S�P2���$��i�L߸B8��􄨟�EZ���FB3t���[κ )|)��=D����*K����x�bO78�Ju�O)D��J�ǁIV��A̻R�>]�` <D�S%5m����oL�4r����,D�D���/�ƌБ��/K�4a�c�.�d5�Sܧr�D�FC�m�=�U�.ڒ��x$����U�i^X�BG	�X=jd�ȓ)n@� �2z�0X��W�4�ȓq��X�s��� � 1�,�
����nZ�)� �~�8�h`�/�h��#�^̚5`@�,$�9c�I���ȓ� �z .���aSJ`�~�Iy����P�Y�!�e�H�B�(�5q�H�X�6D����Ó;<\Աh���O�D�pd7D��#I̩Mͦmy�$	9r�4��Ad5�O"O|��� ]�+�> ��Z�[p:D�g"O��a ���'�!Vj��@�"O�T�t���~�.�pw�9w~^�y�Y�$F{��	��{=0�I��B�Qr����]��ў4�ቌ�Q�s�<[�#�]�#�.��hO�>�5���	f0}��I��~w@�a&�O�B���h���@L�L�}���^�@I��uX�4�<�U":W0���0�o���[��l��P�?��a�
.��ebQ��8_�,��� l�<	v��*��RSh6`=@!�m��hO1�����5,�f��Z)4N$�@"O�-�"V� ��!(�iV�����)4�S��y�AD�{�^�W?�:���j���yBL�n$4G�ˑ@�Ⱥ�-���y� �kI�a��_�=jԑ�4�٦�M��'��H�� K;@o|I�%P+7{J!:�'��ꐨX�.Y@�f��6�0y��dL8�h��<��F5VD�z�%��=d@Q1f"O�P����sĂ4Q�N��4/�y�oi�Fo�dr\��^�/�����Ye��3Rl"LHH���9*e}&���6�'\!�a���&�jb��E�r���X��$;�I���M�O�0⭓�+�iA�Tb���'.�I+���7V�2��? *��{�}�X��+�S�g�X�A�ŀ�2Q4i�qhG�{#=���T?)�L��Q�ₐ	=�BP��Ռ.��$%��)�g~�	�">k����K�g�����ē�p>	V��.7�0��kC,6o:�ôc�i؟\�\�� #�J�)8����&��i�ɇ�Idܓ�MF7�jUa��aJl��b^�'�r���)A9ST@겤�3a�>؋��Eo��	Ex�|�"�(!�аa�Up
`g�r��G{��W�,@C��=z����H�$����$D�(��j�9k��`�D?|�ã<�2
+�O� �y��AXj=���Y���u{"OJ2
�b�� ���;Mh�Pf���G{����'��U�R�/odh��� 턄I
�'K� �\?C~U��K�|@ ��y�'�`��ʅ�;b����0���@
�'>�����֫3N��!'�Ux1ts	�'�8+�"ۂ�5�UJA�jO��y�\��E{�O�-��f�6_V����L�q�z!`H>q�'��iRDh��L��'Xԍ��%�¦��t�)�'�a ��"&T}j�@�&�d$��	u�S�(ScM"w��c�e/SƊI��|��X#�JЗ
bJ��D��+T���Gx��)Zc�_��p�wdY2kΤXr��v�<!�E�-m�0I�U~8� UC��hO?牙nh.dB��� �F��D�D|�p����>�� T.U<a$lX�J;���Ä]�>n!��̋G����R����P,Q=azb�FY�sy�☻#h�0`�6Y�dQ�ȓEŬ0f ��*pNIR
�.-M�9��.x*0�JJ1?�!J��F,R�,�lQ�����v��'N�X���ǿ1G�@�j_+�y^3�:�c�i����E��y���P�bRⅹ;����ޒ�(Or��$ӎy}RI;b�	L�Lhdf[";�!��é:��q3#B�o�dm�gkA2w!��+2z. �C�;�E� k�	rƱO��h�}3Ǎw�D���݄��PZ�	�i�<yv�Ȝ�,�#�B�g_�@����h�<iV�F��1i �QS�Lҗ�^�<qEc7$��kT`�;H�d,{���]~b�o�O�����K�?�4Թ��a��!a
�'̈́�I�D�߮	3�F=]�΄H�'%ў"~��
_�L�.�1�J�-6��B&�L�<�7���xl�g ވ*W��A�RJ�<��EܶH�z�sBsǮH��j�<��eٺb�(�Q,T0 ��˳ɂh�<9�GȐ+㤤�g�5b0l�Ѩ�a}R�'cJ\��
χ-26�{�(�3%����'be�@�Q���+e�D<&���'(|Pv�V�{+L�*�d�9k���,�'z08�	#K���1�߯l<�����`�i�-J��Đ��D*n`�aG{��O���R@ ;r��l�![@Vh��'�v���`%I۠kN�W��\*�K�O
��G��o�6i����Po�l�����&��!�Ĕ4�܍������ڡ%���IS��(��(��i��-�����-�E%�"O�n�|�`aP2  C*�Ԩ`�x�G&�O	�0��+O��Ѓ%A�6��A�'��Γ{�!�U-��F)^P`鎧9�����5>����s��q���&"���Gz�i6f�~�Vo�Y�r�3 ��9��4��	�t�<ᱪS�#��؉FMR�h�G-�?yq��s���
�XA��a&�
:Ѯ@ǥ6D�葂ǂ-G�U�E�0 ���!��4D���W�H:@Z���m�1V��a��%D�ljC�Ub�����͡:PT��
%D��
��_U]"8(��ǜ3�,�X�n0D�T��]�͈e8�̅�U��]x�O0D�0��FB�� a�h�4���h�-D�t�E��_����������R$+D�D���!'պ�!��WPV!I#�'D�(y� �4@�x���M|HK��'D�R�+m�Н� ]6��i���3D�� �A�W��&O@r4r��D�R�5��"O��)B(�V���$�|���"O�L�s�(H � ����0�6"O4��W(Ȅ~�z���OB�R��)�"O�{�$H�W�% ��>�>�"�"O�l� ���keNΎyyX�Y%"O�(q
��C�:iۆ̔�Yh�e��"O�,�PΛ.y��*��/N%�3"Of��R`ސ:��Xg��_�H�"O��Cd <o;�K���b,2=�"O��;���W/�h*�%<P��"Ol:vG+H�p�[+�$ ����"O��n��2���7�IA��"O0��(D�~4�m:�@K�A
d��A"O<L�_����#-�@6"O$���X	dZ�3���7��@"O�Y����Ti�	XV'���e�"O<E@�ا&-�g��-^l-r"Op7��56<�%F�QL��Y�3D�d�B�l�"U���qEn��&%&D��q��Dp���@0u���D�%D�4!4�Ԁ�X�h f��,��!y��$D�Xtg_Ҭ����j��YK�� D��q�m�Z�8�g�\���i`�:D�PH$)�0	X)x��#V�ȹ2D��8��;^��;�"�be>ɡEM<D��`-�%��䲆gI		�;�:D����d0 +���(�+q����;D��c�,�.o�lЉ7$̥0�F�"��9D�D��GN0(̌� ��%��:D���f.Z7}��e��ܕ���1M8D�LZGd�p���e�ڄw�a@g�6D�i��+����%�Y�v���"D���P�������q@,��0$5D�t��19�p�q,��@!�y)�<D� s�IݴW�AH'a�c��)�� D�q3i��Mr9���ߌ^��	�e!D��*��/\Z����J������<D� ��j�����^��r$l:D�Ȓ�z%)P��[�N�Fh��拟�yr��&�v�qd�imr���*�y�#���4=���P�\Z�I����yb*�I�d�@�.W/�U�����y��"{�`	D��6Zq���W��y��x��c!ҩ<]9rl�Z�<ɀG�)֬t���6X�H���M�<qR��J@R8�c��2�"i"�e
E�<@�����ǖ�(�|!��	F�<�AT�}B���'À)�J��N�Y�<���_<��X��ƽ2�� �[W�<�cH�
a�1
���A�4�QPIw�<y���2C��Qpč73�^�A���l�<95��:1 \|�R߬R�H��@n�<i�������Q��/�����!�k�<�`KOܭ�"�M�l뺄�g�W`�<���
��Т`P$y��i�̕b�<�a͝w1�UB$��/��Z��@{�<�]36���³'���� BLs�<a��>Q��₍F&54 Y��EBn�<16� |� Q!�m'i,ܒ1��R�<�we@���L�w#O8r������NT�<&\��!c7%�gʖ��'�W�<a6kǘzzla�G�w��܊@�N�<�F*�;�6����Q�J4��!WH�<� ir���:�-�� �4Ql��1"OJ鵠H�����Zl>L�"O4����r�����R$P�qX"O �b��K�,��K��yD���"O�i@�g�O{��C,#I2�k�"ON`@�AM4��z�@�"z8j�7"Oh��#���p�$D�+���B�"OlpbpG��@���f�ξ�<Hz1"O��j��8 @�ZQb�?�L�;�"O
(�`�,u�����ġ=	�`0"O$YA��)H�k��I+N� }�6�'�舉���g.a|2�M< �����ϵg�`Pb�d ��=��W�Hɒ�! @�O �V@Y/W���I���0��Mz�"O��c^#� �5j�J��a7��%K¬�5�׍�"}*W7$��i�)ɩt�Ti���c8��J�)�S}"�E�A�=�b��I:.}���Q<�H�J��ݑ(�ʓF	��|�'Șk��'M���,G?	��#��ޣy�$�!��iN	a\���+P
9��4jV�K�m��8���"n�����c؞h�`$W�N"���J�5�<���N�Ld����~�����3�$��A���M�����+�r�`7h͌C��tS0�`�<I��D�G��8(#I�X�tT!���<Yt�K 7�,7��)n�m�R��
�S�.|y��"FH:xx���gK�	�P���G�:P�QX�'قY�Oڜp,:����.��jm�H���9��<I�j!�gy��J�X?�`�w'á��	���+�O�I�푔�ȟ��h$]���1�E7������4G�iqh�"RZ��$A3������	?-&��7kE�v]<�
I�S�i�(���rAM��D��#OZ�X5��@B�+َy���S�<9���
�T�Q�퇊	ٴ9��!�D��'W<l�@�I�Y��F�T#Y/C�|���q4�,����'<�!l�J�Ş.|���2O�#����P0�Dp�/� ��9?��ŏ�sX�#}�E�݆�0��$3[���jʣ]��i$���ʊb�g�E�GN�p��ɷo�z�rLڰ��ƢȨ��)�F�ԭPC�~r��:��!!
I0I$��qǄ�+}FEz0'����d�><OBQB@�H��lJ��}ڤ�R�ųb�Yp�O���FEV(�m H<ѷM��,D� `�<��K��rTM�Tq�$�[�'��Xa[�́@�+f��˲C$�8	�P P�� ΋g��'&� j�� ��AF����" �j`;Ed�"(��9�#Z2ʸ'���1�٤a0H2��F��蚜7�5S�
'⦜+�b��I���P�>)DE	����'n�=J���y�h�����0��t����"gq�}�1�Η�yiL����I#fWx�0�oP+7T�]��|������R�' %�C�,�J���W'M�pM8sO6:Ղ��Պ=di�D�x"�w6���)�ny򨍙y%���B�%J>:�S#�R���<�S��'O4.�c��ӟD�ֈ���M�"4����*F�bH �h���ēT�����jP�Rp������$��P�5�L-M���q�ɕ/J�q4LK�9Ⱦ�x�*�5��Ob��c�*Z���x�a�	p	Y�&N?t��/
"�B��x2K�;>�4�%���,81釣
��<T��#��\a���=�h��,O<�I4� ��&Q�)
>}�`C�BF�L"��Ű>�D-ȓd�r%C�E������A=ь)��ְ'V��x�)��m5�'N�I��S$��I%MV��eǂ�%ؽ9���'wf,�󄂷-̕id,V%qj4E0r�Պ)@eJ��U�s�R�\�̠J�E@�ɼ@���Q���I�/rnr�ђ�FF�bC]��'~B�#�����Z'�F(^�1�~�Cs�FDs�i^�6�(�P�a^p�<�ۙJ<�)/֡�xA�g޳n����4@қ$�v�����r�����v��h�BU.D��Ȓ7�^X!�D R�e�B��D�J�9��6�1U!ٶ)^T��W��剋'�Ly�5B�+W�@8��co0��Č�i2����	�Q�H�Q�$J�p��7_�b�j�y�a/$��Ƞ��>e������L�H�PUM+�jX@px���0@��?	��7Q�ıu%C+)�9���"D�<ʳ-λh���R`�܉0����h�OഛF�*ʓO?�ᑉ�+[��8�R55P<l*D�q�'�j�
����{��(Z��US���Z�'�L9����c���iÇ�������'^����(�>Yv�V��:��N�a�<N��q$K�g�\2p�׵yHf�cW�;4�� p��3ǁ|�5��lQ9��d��xB�Y w4��mZ4���IP�� `��Sz��̮4_��b��O�
	{Dt؟��Ff^j� *�KʂpYE��
b0�yz�i�rxi��*�@ؤO?���"W�~&0�h�"=p����`�'�du��a�x��4��Ǖ
FS$�Q���y�|�'(Q�Tƀ�>C�5��	���杼YE�P{���2~+��{�S��e�,?qO�c╻qbX�<��- Q#.]\=��~�l�ɠ�=$�`��EJ�Lߨ���G�D,ҡ��%����F/���E�zU�ԫTm(���?j!$R
^�!�O�n��"@#D��$�zU M����7�:��a �O� ��ES��`���<�O��x⤎�*��r$U� �-�q���>�QDZ�XM��za"ZG��*���	8>np�'�9j$��	�%x@��C�>x�ay��(QD��b2f�zJP��F@��(O`ʃ��)S@ȴz&V�y�@'?�+�,d�:��	ӗF�1�ƚG����O�rXI���N|F�����%4���-j�-k'��h��'���
J����yWF[;G/�}8�	��y�h@@`�χ�yR��G����V��qr,���J���n`�H"'�G�{ʢ$�P�	�`�Ը���~�ء���-�&����
P.�U�Bl�d��負�8oG���WO�5F����&��	������&9���\;�-����d���?�LۢJb40�̆3�z�{@g9�I�52Y�`jF"�# Y��KY�+����y5*a�4Ȓ�[�R�qb"(k��H���J�:��UD�$ ����)Nx7.i�����O"���շL��!ցޖ%\x����'����,J�4T�xR��(�����Ѻ&����pCU�%�Z�J�Y��#BH��[����2v%�n�Q��d��K�P��.�,��0C	���� F�e��ם(Hz8̨���lȼȡ�Y�q�I�U�L�YǊ�9��S�0�Y3���T��H���&<r���UL�*���n�6	=i�c'˸Y�P��r��<�`�P�%;~���%�Վ*���S.`��@!�ν*�,'�<+�P<˧O!����P%�^�1�)S#!
D�aѰd�qj���W�*B��)K��Q&�J��i""X�B!�0�~R�6y.�=1�E� �� �?�p<��$GpR,@9[������3�.��U�&9�HZ�&�!)�N9�q�	\�pI��U�g�<��M�2�Q�ī��>�$kS�ޠs�Z]	aA5}�ؼD���bb*z��̳g�fo��$n��/(8���銽_.�� �2�
�SR�D+/�jܻ��[�
`.��$��!�8
U#�?��ɘ�C`钱9BH�U9�#,��>biyVΘ%�B��A�=��7��,/��睬jd�d��k��ziN*4�'8��B�	53CJ<�QL�Q8Bh��B�p��a�&�ǔ!@%�E#p�p7�]VhF �!��P:Ht�A��u���'U(�q�"ĝ�T��P��/��=�
�;����!г_
�;$勧7�D!W�P�i�lxf :��C#�ԦRu����-�	��J@�'��0�t	��0%������f���N>��ʎ�g��˖늒O���#s�jݡ���Y�3��������$����mB#6R��Ȇ�
BҩR��Na���"�⟔�F=���ߓ+'��Y�Bd�LIqʔ\��9�*@�:�b���@1���?�S��h�PjZ�0�$3��HG+PB��.f�`���9�D(�"B=w7.�䋆Y�x-���iP@���I�2�>O�9;ր����hAحb
A��"OL`Zm؝I�`yn/������>)���^7����ĸԞ� �B�Uc��>gF!�$�|�E���	�X�03��<=!��΁b�lE�Ԅr�"�ґ+��7E!�׾-D�E�P$��>��Թ�X)�!�$��(��ㅤ��2,�P�JרO�!�D�Gf�Aa'R�f|4�܉>�!򤈺�x"�Բh�����i�G�!��>��$�G�}�0U6�!�L=g�ڹ�6�B:dT��	 �V��!��ӁI�4���ê~6Ni�Ě�e�!��6 �^(��j�g�� �6��d�!�����tk��:ٴ1+^��!�d�?^�@�J� �����]�!�d�XW0�1�N���!YP��3�!�݀1�\�"��F���U!�$�,��A�j�2 ��W,�F3!��K�(���x7�	'��H�B�~�!��<!@ �9�bZ5Q�%���֛a!�P�V��Ց$�Y�7��qd J�y	!�� ޕq�E����w/҆ 
��W"OP�A*ֆc�|;���G�|�"O�|���S�bC.Su�C"|4�<C�"O��8����]~��7'��R8B��0"O4I��hA1+*l�������"OP����*l�l ����)>D�����
�=X2Ep��i� �Ά��!�D�?��Q�1�T�d4�x���0�!�ʒ%��� �2!l�C��*�!��H�j vbŕ���1�AN2k�!�$��!dXI� �6��� �Ş]�!�_�/�d���^�P���c�@�<s�!��X/�P���̎P�4US7m�VT!�dƃ,�$p��2R�b�+"��
d3!��ġ����I��[h�0"CD	5!�$O�1�� �C�)W�tDHf��:�!����T
p��R��9����m�!�M�8�̈�քD�8�T�̚$_�!���&NV���.��=�.L��MV�l�!�
|w ��!��?��k�M��
f!�dہo X����E�@��P+�I)l!�d��X�����(tٖ�y��W!��/v��؉�)�\k��a�Ǖ-Z!�*�Z�9��N9�Jd�%�9�!���@���� 
3�d���"�(�!��F�"�K��U�rś�>�!�$�"v*|�8�☟x��=�7���!�$��/L���t���A�rYG�U#N�!�$�/_�0Y�=:��%����!��ۯL�y� $Z� D`b�"�!���!�,ˀ�
�dܹ+$.�+�!�D�n$&���� D����-C�!�ۼ0��9�ĈZ�d�lx���+j!��D"j\�ٱͮv��@Ԃ�.%:!��gɤ�QrDpU­�N֝�!�G�ƨ��E�!�&Q3��|�C��*/��� �O�V��LYH��C�ɠ��8g��h_�4�$��X�&B�	w0v<�ra0}����@k�9�,B�Ig�t��iA�vu�����R��C�	?�NQ����xS�B���%t�C�I/x>T���  �~ȃ��s�bC�I N���t�ѩ`^��"_	:B�O�)����V��w�B�Ia��EOR�S�
�(2b�4s0B�ɤ#��hfH B`�)�Gl�m��C�Ɋ{�B��,��V��A�mK�M	�C�	!�(Q�M^.!��M��ƒ���C��;W�"P�A��}�}�ԁ¹<�C��&'���@#�,?H|sQ'��o��B䉝�"���lE�
�Z��7铩B��B�	�\���fI��=��/�~�fB�Ɋlt�q@���[������,^B�=^>p��s�ܛ^|���4IY/}m<B�	����Ӥ�5޺I���5C��C�	�XzF���l}�숕�T�N9�C��4$(�i�ͿuH��m�$v�C�	�T|��H�!"��ᆪ&^��B�)gޠbeg�aS� W�ވ9)�C�IA� 2���U��$��f��\��B䉿IH�li�n,#`��Ş�`�B�	���ا�'`���ދO��B�X9�0��i�!v"\�E��B�I�V��� �)`��p7��3��B�)� �ZW��<� �3$��m��ti"O$\;�fZj?�AkpVcZ�+�"O�<�š�<�����Գzl��"O*݃�L=4�T��� W�PK"O��_EA�p��#�0��p�K�H�<	d)C���A��؏�t �1 �^�<���P�t�Th0%�ʄ��\�Q�U]�<�Ӭ�6�L�a�Ъs�f	���v�<��'�-m�}Bҧء0����C�q�<�W��.y��&!s����4/�l�<���Jp-h�f#ŀ�H�m�<q�#���xЙSJΕ��@Q�n�<����Ҽmx����H�:�Z��Aj�<���`
��q�6E����`�8C�I;8�$(�.d����+d���@���RV�*�O��JG�P<J����s$�5f�n����'~����,��6R���ɦfdƝ�u�@<l*Ļ��ǎ[޼B�I%07"�#u!ǲ-�4츢E��4�X��b��J�$��A�\i�O#�l`T��d۶��O߇s�HiA�'o�E��h+R�zmY1G��k�n)r&�)�"�U�<���(�gy�jFP�Pݓ�'��(@ �����ybGȻ��02SA�jiVuV��v��S�) 5\ؒ�&5lO�����`�����׸#%<���'1z9��I�HHp�"�i��1[Ȅo ݠ�� ��B	�' Jm� L6�I��IN���p�y�E��}X��T���r��i# Ǫك.� X�n�2��<
p!�D[ <���W菋6-~����*RR�-����x����'�@QE�,O����7_�ɢBN�!�Part"OR�� LARJP����
�0��3Q.E,	�(���I�Ą�	�f�옃1��4H�X+E�	
�����@i��$�Aܹ�?�J�%E�<����`������Wn�<1��.n&�Ca�T�&���n��؈�EhN������c%	�;S�x�
_�T �o3��'<P(�$/]s�ŞɊ@�C b��)a��6F�@�D{����#R��D�4`�bd�HC�
�7e� 5m�D�!N>)�S(����I�K���#GDf�)�E���6m]�Z{�"����$������	U�A��ɇ�3B�n���ɳ�F�:PH	�.؍(s��ViF�i��D�<�J�)��xRh	1)r½@3j�~yB��,h�D�B������G��p>!�ǀPlPqSdKZ�ǈ,&"Q�vm��z�A8_��O�0aU��v�Və��)Y3�(0�C��NNP=Bd��[TqO)�gM��)�ʨ��a���,��VbX�z]��H1c�2�h���J��n ��'$��j�/4�3�D�~�U"���6=�8ҋT}:\��_�Uj�A�3OJ-���>���ӂ<�(Z����S����*��i�2�3� F~���D\�)��q��'[O
���@S@�4��r�ݶ\�dY�5$��~	0O�݊뉁]�t�*O,R�*E.OLDe�D����'N\C���@��=���A#�ua���w�B}��F�)����xR�M'V$����%`�O��|�%R"rvpI9�"樌�H>)�nA 갤�@-62](52w��F� ��tp4爆x���2&��?(�~�:�H(}B��{Z�c?O��pa�Jђ�9�0G�ʰŇ�
�d�ɚ`��s�̊Tp�剄
1#$�	Nlt�v�D~���f�ѲA嶅���'��LJ�#�O���l[�!�(v��61��AY�TĢ��p"QH�D�8��Q{w�$?�&	X�y�D�e M.-x<��֤�tx�L� �,(r,ݺ$��h������X�q�*�MٜO]��ZK�n��'��d��UW�S�'�T�7'Q�Z�1�� &��!�KE|2`��z�U�	յ_��T��e�\rݠҡ�;s!�ĉ�/�V�Jt�5H���A=S���(ԭBF �^Ϧm�'� �g~�N�f�ЕZg'�*�R4�g��>�y�eBڊ�&�9B� ׺iܶH�s�@��ܓ�I��R݅�IKD�h��H'=��3�ڨqh��L�h��M�e'��{��1MO c�pCҠ��{B�cŊ>$�(���J��}ڲ��Bv���,0�f� ���nO�r�<�?�z�c�IJ����ƾ&
p���3D��Xa����%i�%�\�vl�Q��O��Q�ޒW^p�O?=� Z�ag-
�rL�(�c͟0@�ݰ�"O
(Y��m��)y%��	�R9aF�>Y�
�<$����j_(Cc�@>*���2oI�9a~�����@���b��E���w�B:\%�}�'��D�E� l����D�a!�8���$R�!b� XV��~����~��A�Ҋhp`p�!g�<��̕=WTM� ˇ*����(����S�AT��d��>E�d�1ZaHլJ�L�2-�6N"@!�A6��lĴ¼���'�:I�I2�8�v�>�ay�A&)cҹY�H�Yp�=8b���>)2�,�H�B$�����DͺH�0xB�A�B�ɂ(���8��:Y�8ɺ׫ŃXyt�=����.k.V�;�6�S�x�<��kS�|��$�`�%D��g���Uۤ��Q.̕G�PXt��O�h5����LiL�"~�2js��!�L�4�h�e�1�C�I�{YL���)a#��I���˓>�����ǕtXJ��䌑d�ܨ�c�O�^׍�u�a~R��;db�4���ٴ5���1�
���f �f�񤟉'ǜ��f�'<Ƒ�W�,�Q��hR��k>0�DԿHl������17��1�n6D�\#�"���/^Bz��, D�HY�̛�(f��c$�`�bH)�l4D� +G
�&h�ѣ� �|�| �47D�h{��ݭ1(l���<��`���0D��b�E�x�TCI=ʒ���N14����ͮG2�"��^�Ж���n���j��'ZDM��F�	���SZ�5!
˓hZ%U��'��I�c�LĨ�&ہ]M���egB<BJ�B�I}��JV�;(��>4�6��A�>���«o,u"��F�}��Zv�-§5T|���գI�Ƚ��$�H�x�ȓ)능3A�`|pJuI�
Q�|���.غC��)��G T���P%�Fi�g��*��XK�T�� cU�U�TC�t{�	�e�08�\᳁ح�V��"���W���U=���.�XX��A��I�w,��8W��5!��Zag0Oڥ@vc��܊d�����DbC��0=r�ב)\}1c�Ү(�B�IY����2���� De��-U��'���J$]�L�Q��<P�m8��	�>�ݪD��~�,0���8{!��ҙ@�
���?=��=Hm�oF>�)$��\�N̓�ك6�扨���!��W'Q��P�NB�y���"��3d1���(^�)�3�_@n�i��Ijld��_#;�����-��hX�&,O6Kf˸jt�(���W/o��'���yv�î_�(�fB�g���j�X�imP����ϵ^�֔�Ag���x2��;��{���.(�n5{C����(�j=kc�%A��3�8U}\b?S��.��$wB��2p��s� %D�<�Y)�b����@�uݸ!#,���yRj���Jǝ|��I�![򵪇�ܧ�2��!�d�FH�#FD�c����ތi�6�z�	�-$LOf���h߳��-��X<F�i{%"O�	h��B(^�~�ˠ�J5�y��X�er�[�f\%���`g�4�y�(×^������Q*H�0e٢�y�jǺ[��d˂���L,�-�uD��y��0/�)��-B�J�%��HB��yB��~7,@���C��T ���y�k��-�xr1`�F��P��yR�١'�\����+�>Lcᛠ�yrJ�&���W�C���0j�/��yb)���*�&�Ye3���ǆ3�y��%��lw�)Z{\�`ץ.�y�F�<;����GWx�AG��1�yb�֗?���M�05��F�9�y���^�ʸZB,� AJ��y��#�y�Q;�,�9���=���K���yrI
�E"��`�]�J4J����y
� 䤠t�ɜj��x3Ѩ"P�@YC"O��0�ݤ ����/)	��'"OZ�0�L?t��ġ��V�Q��Mڐ"O\���H�Z-���e���0"O\�F [%"N��21�a�c"Ob��ǫ[�gQ����U(bM�5"O��ص�G�P��6J�"���R"Oh"u�LtRdz�ɒ-��0�"O�����x��Fj�<�U"O�P��a��t��'D[e��!�"O ����\ �@�7BFнh�"O:IJ�"��F]@X��C�(M\���v"O���n.2E��k`l�Ix�Z�"O$	�/gA����MU?<ȉ�"O��k����Tb�i �h
�%B6"O(�.8.�B��w����Գ�"OFAh�Axړ��6:u��%"O�D���ɉ��� �O�Z���P�"O����% �Q��عF��@)t"O:��fB�!�b�{J�	�
�"�"O��cb��Ÿ]c�@��h����"O&�zV"[y?��z7�>h��1j�"O,�ڒ����NH�2	���ہ"Oz аJ�M�J�z����\�`�p�"Op�sG�	>$�b�X�Y��y�A"O0����:m�@ŭ3� "O�5ZB���6D��Do^6t�0 $"O�-��M�%��&�RC:4�"O�x����2d���@�O�Q��"O�ѩ�-��e��4A�)�-!T�#�"O 8���S���0(H& Rz7"OXh�2�T:/�D�2e)C7P� �"O�lA$�ќd�yj����.L\9�"O�8���F� *L���O�o��5"Ot�
B��5<��h��x�@�"O�,�k@ &[�l1Ġ��r�8�"OnT��<z���dz�A��"O$0[����kk\�2��>N�Z���"O�QPD�V��l��]B�,��"OP`���ַ!z-�PN�6x��"O>�k#�{*!��F��'�x�'��)�3�?a�bL�.�4;���W�X�3�;�\�/(�<�G<��Iƌed!CR)^4�.8
�b�_1�IJ�(d�x�)ҧW0aU�г3�%Q�"^�D��p】V493!�8}���^�|ң��7���Z�hE�t�Y�吼=��q��<��F�C���>%>��c��g�����z��������Q�*��}��/�u> nF�+h����GX^��B��>I��,?3*�2��x�����f@�QHR="�d���~���(1M�W$#����w���� kq�0=+Bݙ��<yεXPmL2��O�����ʎ����K ^5V%�Q苲hzfe�B�M�#�BS�@�##}*��c>ՠ�� ft�K���m�8,����Yy�r��(�b9��1s�Yk1���)ta�u�'��Gy���%T�2V�7�a��牸i6�T�a/c�"On��(�(��@�91����f��Mղ�:�����O�aCe&2�$Q��ݞ3��}�-\>2��}4j2�$8|e���6H��j��G���|B��͘	; 1�F/�&Y�r�7�ɩ`Ў��C!P3i��i���蟾]��@�$��H���C8O��R�̛���C�	τh�8扡���b>1�ƈ��P�4R�Y�R��`�:D��;�K�6�̑��0�B��Ň8D���W�q~����hB�rZɻ�G5D�h�-LM����,#6�#U�?D���Q鑼&������2�%��!D�$:5Ȟ�;�,iQ�p>��� �9D��B"I6d���!HC�P��c:D�� �
P�+7^��Q��]t<�ȓ]�Z����H�U� �	_Ʈ5�ȓm��RBOM�B9XQ#b	ňiyTl�ȓ}���c�Cz�Wټ\ T"OA�e˃�):صSf�F�uؐh��"O�`���(�j�1�ЉP�<K"Ol�Z�L��:|��0@�b��T9b"O��$� �B]d�/ֆQ�|��"OLЧ*K%o`��PpH�*��PH�"On�:t��/�:)8�'�s���"O��4��rX5��'�%y�Fq�@"O%��NG*��E$0F���"O�퐔�D\y�V��=MV�� "OD(X@K׭L�	���^3�P{`"O��"��$lhu���
��a�f"O��%雀5�6LMTB�hD"OڨP�ZwԴC���(\�YQ�"O�H2�#3��uq`O�X
��"O�}"o�M�֬�&n̾�t��"Oܙ��:t
)�p~���f���y��I�j-��#fP�+H$�#�nU�y��ۭ9��)8BP&%�^ɓU�� �yrfB2[V���.� ��kb`��y�d
�5l���˷j��4#qm@��y򬕽EvP�S"�^"^}R {Њ��y��V��f,#��k�8�i����y��҇6��m��O^,b�Ktퟲ�y����9�@�K���h8����ۗ�y�#[�[��<	"�a}6y��d.�y�g�z	��ʰ��RDV�hrjנ�y��ýw�ك�H�?Kϸ!�a���y2���^�q�$iB/��(#!�A>�yR��4�桀��=�"�
�.���y��`�B��q�}�X�P��0�y�ɯU\����r;<�KЩ�;�yRO(8/�Y���vŃ�Ȗ�y�O�KFb���EѴ��\C�f\��y�o�:ٔ(ȶ�@"���y�I�lq��P�A�2�Ľ�anE�yB��<-�����A6_����1��y"��*yH� K��#]�T8�@��y"GU0i����k\"K���p���y��cA������EpĹ�@ʛ�y2䂙=���(G&��y;7l�y�[�z�!�v��vY@ᚅ P��y��h��=��e@�`�(���L�y� Jm`�,�T.áb��k��ک�y�cBu���*�L_ o;�86!�&�y2�@�<4d�xIE�gdh�pƗ��yBHʻ�M
�iP$x��U��y� Na�(eр�X���I�p옕�yR�0!t���ACzdP�����y��_�L`���>�P ��yB.�6�8t��D�9^���(p�o�<��닮7T-��B�z���$E	a�<��^�}2�I���t����}�<���ٯT<��4��:F�2��Z�<�Ɓ	�`e����- L�
��R�<a3lV�n�z��"��*%�y�<!t�HLF�����34�h �hJw�<����>u���D��E�\`�b�x�<��C��A.P	3%�c<����y�<�Ư���ƥ���%>Q��{�<QJ�;OA��`6iw����Lw�<� �Z�(�D1�5���$"}����"OL�KtDI E,*ez���;.QbD��"O�aQ�`�#8�쭈��ϋY/&�#"O�L)e��R�|�bf��p
j)�'"Op��2/9z=�%�#T�#"O|�cRI�/B�YR.E�~O��"O�{Ã\�_V�L���^�����"O���cFS�g
F-9"*��x�T"OvP2򄃀O:��
�l����b�"O�cC�^*78�m0�M�c����"OkT�@09�����ۛ
�ʑ�"OLui�j��g
���6^�,�"O�9�ۮ`Ңq�Ba�7t��ɒ"O�]��s{du��B��B�b�p"O�T��숼i�(��6���v����"Oȸ�,M���I`@D�"�Z�0v"O ���NN�H!��Ӑ`L�h��Ţ�"O
�+�/�6^oz��`\;\�L�e"O�@I5�W�V���u	�%uM�@�w"O�e8�����A0�Y�GB�h�"O�Ds)3,����ԈW�t76Hh5"O�`d�B����Hګk/R�(�"OJD�O26qH���5;�P30"O��ASe͆]������3"O��Q���(Ҁ{�Hӂ!����"O4H$�>%Ԙ�9q�� @4[�"O,Sdn�8/�2t{�gӜ�ti"O�I@çA9�`@1ᜁVL ���"O��RĊP:z-<� ���0i+0�se"O��N	RЬ�`���@�"O�-aB/DU8��ȡ�C���R"O()YŮZ�'�X��A�B,a:�"O�<豇P�Z]��Z�7J릸�1"O��ե��K�U��:	{ �a"O*e�A�TR�&͛M�6.�Lِ"O�}��ne.D�	;����"OD�{Q�̂L֖;�K̗?��"O��
a\4�hi�C�Ğv����"OJ�0�NF�
�40�]9X��	�"O�`����.6-�)�3f�'s��Z�"Od ���=H��s*@�J��"O*a� �в7!L��6��'�0�a�"O���@N�#��]��)_��p���"O�L{bJ�H�tU(�8G�~a2"O�ACZ<dgB��T��W��{�"O���E.���߹�tZD"O�( �CW]���:bʏ��y�"O4hZ��_2F+Q�ܑ)���"O\d��(IY:�C�+\�vYHe"OD�k���oR�)�½M t(�F"O@�@tk[�N��Pq��m�Ɖ��"Oz@�@\4���A�0	����%"OZ�(e���+��!=}*|Y�"O{��J25ex�x��\A"O���Z}�,Y*GZt=!�"ON@ t!:?���s���!2�P�"O��Ā�gH�t��d߫kBPC"O�1�D��5*֒E"��#r��"O(�G��
��A�,�S9J(b`"O�t��
�t HWa[ ��	G"O4��c�̑,a:Y�Ԁ�A����"O�kr�׳Qz�Sr�d����"O� ��T��bfEG?[����D"O�+�Eےq��i�� N�v�ے"O� �58p�Z�	S�J��ԂZ��s�"O�}�#U/Q��!bDt�pU��"O"�!���
! �F�K��8T�`"O@�˃LTD(��C��H�Rzl5ʰ"OLR���7F�6	�O�h�p�"O-��{
蝉&G�n| P�"Oν����[u��P�K��!�"O�E��叝7s �R��R>,��"O0Y�A@�W�	He
�"P��Lh"O��@U(��iI�Z�ƚ=�l\`'"O����W�W�^H�CE׮Ǻ��g"ON��C���`o��8�G���m��"O���&A�#����c�:]�� ��"O�(��/t~���U�Ͱ_6D�*f"O�q�a��s����*c����"O�*'+�;1UԽ;qj'S~r3"O������S�GK�Rd0��"Ol ���o������ �h֕"Oj� ��!@�P�ǮL
V,C�"O�he듅��MHR��\���"O|0��R�lN����M%I����"O����"V�&X���X</�)P0"O
�%��WƖ��V�.�2 "OPA���9*Rą����*6�"O�8ڣ���gȄ�bdC�	���yE"O�}����gx�=05C�&]:�"ON����r��H�t�W
&�.�q�"O���f�V�`S����F?�R���"O��c����Q��	��6]�2���"O��kt_�V�D-{@�H�ID���"O�����;3�E4��%6RёB"O�i2$�GD�f�:��
>$���"OxAbT��3��݊5*	8"��"Ozh�@O�9%g� kT(�� & }�"O\��1N�&$)i��琶*��X��"OJ����`�h������[6"O4��&��)������-j�ʡ#R"O�E�d���yb BG/�Aʔ"OJ�za�[2.�B�!�7c˺��C"ORM2���!>���!X�,�f���"O��TL�3*6�sw�ǥW�n��"Op]���L�,�,���+AX��q��"O��Bq+�)�B0x�J� %����"O��C�ɨfmDћ�	�C��z�"O8���;��A�JP5���R�"O�t��X�J��� ĢTt�"3�"Odu �� ~�l���+��|[�"O�y���\�*gH[1�[m���Z"O&`���
�&�ʆa
�j=@"O �j��Q����5��b��	;�"O���ϔ�Jɒ����f"O�՚1DX+x%8=�seϊ����"O��H��L�W[��[�D��D���"On�K�@�n����/c� ��"OX!����i4�?�0���CS�<	��
�(���F���t�<�1��-e2��̂��Cʗ7�^C�I0�d�cą~���� �2� C�I57ި{Ud?R�q���[��B�I�(ļ���*Ձ$U �"��Z�F�B�2_�}b�hV>"�'�" /&C䉛ZB�    ��     �      �*  �5  A  �L  �W  �c  �n  9z  &�  ˏ  M�  |�  c�  ��  �  O�  ��  ��  W�  ��  -�  ��  =�  ��  ��  &�  h � � � � �% �. �8 �? �G �P �X u_ �e �k �l  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����I�<�q�~"�{b��J{���kG}�<�"�>N���2���˳�c�<��έ<ٔ��ƞjq�#\�<Y0�U7t��ՏW�E�z�8���N�<��!�&Q�ꍪ  ׹ &���g��I�<�t�A\;nM�a�
�b�Hg�H�<�٫0����݉c��J1��I�<��j��&\V���@	`T�m�`!�]�<!"(��:`Pd↩T�fd�8fA]�<)��-JB�X���T'
�t	 D�Y�<q�(I&2�b��k&<�4���i�Z�<�,��R�8���^$� <kŧT�<�ׁ#���5��-T� B��W�<q���e��E�W*�,+x,p0V�<�Ph�3J����BΕ�t�ʙʦOI�<	#�@>KE���2�!�j y@f}�<�6���X06���O<|n%��@o�<1慈gl���l̶F�0�ɗV�<��/!��n�)I��ģUo�}�<�#KQ'H�����P?vq��Pwy�'953�@l�x�ѭH�%���"O� F�aF�ٟZ�%�G���"n�C�"O.�p�G\%>/^ )vD�q[N�X���Q�OD!��9Lt�RaHŘP<�4�'�:��-��H�h�E�E��]�
�'@P���2-�M��I��<Ϛuj
�'2fII���9�,(�!T�-5�))
�'d�Dk&�]Bo�p!È�#3Jҍ��'j �	�F�" p�Abʹ.�l�'0M)�[�+.d��nχ �N���'�5J�b�'mi���L�0nJ(z�'.��A�G�#���3��+W�,��'ў�}�$%Һl��tB���X�(N�U�<�6k�9g�B�"E�Np��mZ�I�P}B2O4��D�<E�2�"�h�a��?A�~R���f枩���D��6�t�Ɖ$D��q6�O�d	"u@޵3�: t�!�	�<!7���O(un�H(��S0���A��!�Q?*䄚F�ĈR��;f.Oc���%b�Q�>�*��yڕ%J%j	��j=}�td�ȓ1�x�!qD�02�L�i���
�f�=O0�#sip�2��4,Ov}yK��F�ʱ�o�!����'��F�Q�@��V�{�	`%�	�z�h��ēT�Ԩ˥������R�c�DF����Z0n�>3��c�b��H�C�Ii��=^)��ڮP�Đ�E,��<��ōk�)��<��iZ�S�v��,�/!db�!�
�R�<QG�����"۬e����&ɝX~b1O6Q�뉨�Y�$M����$��ؐ�RC�	П�!��\�z�
��w�r�w�/D����R�C7�=��Ƽ����M8T��bo�
G�
3�"��(gܤ" "O�����Z�( scB�fFf�a"O*�!e�]�aV�
�ǫ 0PQz�"Or�+�.ΓN�F�nN�7�ua"O4���N��l�!���q
�<��"O� ��L?A�Ԡ[���'嚍��"O�}!#JL�6׼����XZ�&��"O��`v���!��v��'�P"ON�HfD�����f
R=Zv�%`7"O��kl�4Eǈ��S+��:h�0"OF0:�*��MW��؂�VD�]!E�4�S��y�m�j��*0(�:2]�0+��ۆ�y��4�rݳ*�
غ,���y��A	ɤ�j��ފ�X1���y"h-fǈM�tE����d2a*�y���&e∨��`ѣ>�b�a�ԏ�M����s�!��搆9�2A�& �h��p�"O�B`�K'RC�uX���4�vu�"OҍQ�Κ�м�P.դ]6�@��'��'�X�*�OL��X����})�'S=�Շ��V�Ȇ^ �hR���?�S���4p�,����I���$,6�y"ѽN�2���J�>�X�q��ٝ�?��'�P�c��N�0b��J�9h�`㓎�eA�,��.�(q�FT! ʎ�t�ȓ*6Z�Z�M<_
&��W�D�����	G�đ+S�
m��R&|���1�c��!�_�g�����d{�M�����!���O���uh��L[�4�v��!�䝰gyY*3,�1v�R��5L�B�!�$IX�jP�'�6^2�Ò�Є`!�$�"TB�i�%n(�Id
S.S!�d_jق��"���j}�@PJ�8X�!��j���Y2Ca~ ̘�Z�!�� ��j�A˷b���ӵ瘽1��)�"O6Pa��V�	ᔅ�H�#H2%�"O�)R�N%> I�P��w.0��D"O����Ǆ&�Z�3�IZ�6!����"OU�QdE��E"t�Or��t�4"OXx�'F�fʪ(`e��fp��"O���d�J��Q1g�9�����"OD�
Tk �*� �B���)s}*����4�S��y2��d3�Xu�Í"�����ˎ�yb	S;��gm��&�����W��I]X�`��0���=~,�����Ԝ��d+?�!(O2��\!Fʼ^/�P��En�<	�Ȁ�*�x�gד3�x+0K�N�'��D�ā�����ao��$�0��P/ܥ�yB���v(� g�SP┪������1�S�O�8a�n¥5��YyTh�3w �Pa	�'�6qy"�=Y�*��SH��lA�(�I�̆�	:��U1�a�?`������؟}�dB��o[�����:aQ� 
B��"" B�ɳ[<Ĩ��H;\�t�T��:}�?!��I�R�}��kw̹p��P,!��MZ���qʔ�uvR̲C,B���z2�$Oe�%�C���������.8q!�䞕)~R�Y�ٰuF��T�	k��hO�H��4��/���Qd�d��E�3#Vaz"�3��0Ԅ-y7g^�M��jT̎�s��c����ɽ<��4�0�N)I��)��kN�T�c��F{J|�]F��d��HDź�r�G#U�!�Qou�L �L/3N�A��V�!���#3��
Գp*M!�� ^�!�$�?V2͉�A^�t����!ȚX�!�Đ�_�!�<~Y6a��Y#�!�䈢+�F�(�C�>N=��T���8~!���H��u����7#�ԴA-$k!� �� �䝻Xw$D��k�!1^!�D�3O�,h�
Ȭ.J60���ţ4�!�$C�<m�L���:D�\�o�!�/6��A���@0�C׆} !�7�R�RE)��X�E;4,@�!򤜏0($=
��:e��MI�jެO!�$��T����^�
��X@�Y	!�àA���
��+(Ou`���,�!�$�q�F�0脚d<��Œ< �!򤟦j}��� ܈E<h)Ƅ߉X!�D̔U�p
�·",���7cĸN�!�$�(����`TZpFX	R�@v�!��G�?Ze�C	�qWbLA���~1!�U����*v�@i*A"F!��Q�<�p���$^D|`<�0OB�!�$��µ����Wu�e� .��!�D��Y�t)�[�Ep
�@��[�Q�!��� wx\����2B� �bT�@�=�!��1�rxB�DP�k�.P6�T�!�!��K����o�5��	#��/k!��9Za6��*V�gZց���G?N`!��"��k#�ѷ5NL�Ș6DF!�Z3L$y�@Dr:LAXa�_*P4!�d^V�T��}��!�ƫ�?0!�D';���Ba�M ����#m�!�Q(�B���ɝ��@��!\�!�ҝQ9Flh�(}�]k7�Н�!��;���BG[3pr4�ju(-Vw!�dC���H[#��=VTx�ćph!���w�2��#�P�����-Z!�� l�x��,���P�m�0����s"O��R��yVd0솽w�� {u"O:�QC��=�����J\:�8)�"OrQ�@ʌ����Qi_Xvte��"OrTH7nĢ���2�i�V�|���'���'�r�'��'�"�'b�'��ԣֵN� \�B�؊,�V��C�'"��'���'_��'#�'��',�k��
S����ɀRt``X��'S��'�b�'r�'/r�'wB�'B>@���s���3�	I��Qu�'Q�'R�'���'���'`��'_�m1C`��Ix����ެ0e@���'.r�'\��'���'"��'���'?�4aUfȆcŌP9�呄P�\|#��'���'�r�';"�'"�'�r�'�2�B��H-[�jR�K"�@)��'���'���']��'�r�'���'��Xu���Oi�51�)ıw��z��'��'��'>"�'b�'���'�xUҴ䈥1��(x#��{�n�a��''��'�B�',��'�B�'�2�'�8ǥI�G�QBw�5Tx�m�S�'T"�'���'k"�'��'���'0l��GJ^�[�$��X�\�ݓ��'�b�'���'�"�'-�'���'hJ��ŁGHB�A��S�V�3��'R�'�"�'_b�'^��'"�'Dq�*h���O] qK5��'�"�'���'�2�'�d}����O(<["e����;�G� �
� �� �'��_�b>�A��O˂.�PH2#�>�h=sJܞ�T���O.�n�i��|��?yb��b��f�NѢ$�t���?��T���8�4���{>���'��S6C�0(�j���Ҷ����b����Lyb�ӎF���j�H�����4ˆ����Y�4q=���<щ�$��1�w�f��pꓦ4~	K/$q���'�2O �ŞuӰ�ٴ�y���d��2��/��D�@�I��y�:O��	��ў��柼hR$�7Q�h �/�,��8 @c�x�'K�'��7M	�O 1O��%���6+hI��:hƌx82�!������O��Dh��'-�$K0��8#��	����4;�T�B�O��$]Rd�(�)��?!��O
��*0��9P��&M
.����<I.O,��s��x�oТ'(��[��C�u�2���mk�KشUt�'r�7�8�i>�R"ː�d䜽y�%N�6*L�C�v����˟ ��� \�n�g~B4�����,C��A)�'�>&�����)�ǚ|r^��ٟT�I蟈�����kEEM�M��ȩ���@��黧�~y�cz�p1��O��$�O撟�$[��	���!LR��.�"�
��'d��'�ɧ�O�>����=K �b�N�y�f 8��� ���{�O8��r,��?����O����|�����4��̛��O�b���O��D�O��4���;��V�ش~w$ϖG��}vE�q�xm����vARnӦ��
/Oz��oӒ�m�*D�ۚ�e�M��t�ӥ�����S ��	�'Oh3�K��?i�}b��x�:���i0�-�Z���U V�<
��cr�!s  �mjҨ� o�v��.O��d������$2�iV�'I�&�ْ ,�&BR&2M8�ɠ<�d�O�F�|:C���M�O�����N�̈)1��D��t�$A�.��;�'��'o�	h��}ʨ(sǗ�U��]�.�7Rz��Gx��gӎ���"�<A����	ɸX�!I�O�vW�Iv�]����f}r�}�J$m�0��S���*�|q8��f��Hz�,�9�P��"㌶U:�F�<�'f���c�	�{(>l�
J�Z.hu��kM"�RD��ß@�	��t�)��sy�,v��h�!Z���F�KuZ�2�J!P����O�m�^�*a����@r�ћ-�4ҖL�.�\�;��쟜�ڴJ���ܴ���LZ2ac����S kj�;�*�L�Nl�V�G2'�P�	zy��'���'��'"^>�!&�	�D�80��J�~���M�WH��?����?�K~��sɛ�w�: ����;�Pd�����H��u�c���nڢ��Ş�D��4�yrd\ PuE�f�W^5B+ ��yG� jIxe���䓧�<�d�[�M-�+���'G��h�W�\[۴>��xR,O:�Dҙql`�Z9)6��+8f.㟐��Ol	n��M�`�x�H�$�l$�rI����ir��1��D�.&��6Kz�f]'?A��O<��K�+�ҁ��h	�$�d�٤���v�����O����Of�d.��sw�j����&� .��-���ޭ�?I²ih���'7"�oӐ��]�ÔHS�������Z@��M#��'�F'�[:�6��� �T%X��L�J���h�Ih��tOF�g�]%���'Vr�'jR�'G��'��	b���2i;=b���?����\���4t��� ,O���&��>n�K�fғh��[N.d�,1�O���Ox�O1��H��T4o�UB��'���:@��j\�Dca���]��H�'&�@'�Ȕ',N��R��A�Z��DưM
�9B�'�B�'f2���X���۴E�q��G1m��l��D�ʌ"U V��6��aћ����r}BB`�^aoZ#�M­�>*���신7	�mr�!	Fؠ��4�y�����!*�ҹ���C���SE� �CWE���1�������*�<O����O��D�Oz���O��?3�L�(c���;�$��,��(O���	�����4x��M).O`�l�j�I��&������D��JN&s�<�I<�$�i�.6=��0�v�k���g?�M����2�(b!�0sxy6�P+p������D�ܦ�����'�2�'@ �uJ�	
�qٵf�"*.0���'�S���ڴl�\����?9����	ʱO|���0�çK�VI�W�B�U�������
ߦA0޴i����	0����G�3��QP�2X���3��52Ϡ�h#���^w����I��iޥc�˒ ƶ0O:n�$6B�����ڟ��I�b>]�'�6-۪r�T��BD��>\��]m�ޅK�f�(��d���?��[��J�4Xh�}���@�X�u[#�샗�iQz7힒VH�7�2?���J��I:�$K�hh�\{۷ }P�p��$D��6��<���?1��?I���?�*��$����M;�����10p �¡��5��K�~yB�'N��hoz�����W�73$22AB!.��ck�M��i��O1��81�li��)ǬPI&�+}�@R�d�(�D��d�0�ڇ�'BF��'V�7M�<ͧ�?���^)Dm�ub�����A`M �?����?������ۦ�#W�ϟ���蟈`���s�R��r,K�1p;���K��L��	���� ��t���K�k��'T^m���	vQ�'M���reI�=W�j�O�T�;#J��dW��?���߮S�̥a�	�}iFH��@���?���?a���?A��i�O,aZ�ě/y��u��&�"c���"L�O2�oںL�Ь�'�7M2�i�a2gI7Jr�8�7b�"c��HYGǲ�T�	��%*�4u0$��4��dQ1XE�����<Kt�ÍжHC�H`�"Q�Q+J}ʠm�<�2�i��i>��	۟��	�p��#rF5ۓm�fU���R��ٖ'~7-B�|ʓ�?ى�4��iݘrg�'N��u���R���?9��J����OΎ9z�`�#-��+K	G]��"��MDf ��O��G
���?Q���<��i��
�l�r`�_!5,����G"=�	���I�h�i>Y�'�6M��0�P��+f4��E#>�ؠ(���D����?��_�,�Iğ�	�4�3,.)vB�y���f�>�p�����M�O�mzZ�&���v�	�����@��y�6e��o������܌��?q��?A���?�����Od����^h�<��כ"M��8q�'�B�'��7���=&��OhDms�I�%Zf\r�e	0~����6�Ƹb�F%�t��П�ӅS��m�u~�d��^b@	�KKt���ua�%@����p՟�T�|U������	ПX8U%�1a3NE�!$��� ��˟X��ky�hӞ�xF�OR�$�O��'J�n��E��'Q�����\E���'��|D�F�u��e%��v�N�JӅÀi���BTP��B����F6:(�شX�i>I���O��O�	�gO��&
�;W)�'w񴵋r`�O��d�OP���O1�6ʓT�����=�r��AB� W˛'% ���'�r�oӘ�,1+O$6�%e?��1�$g
��)2�Gk�YnZ�M�����MS�O�Y7��$��DS�L�S��=?���0����i4n�̗'iR�'?2�'��'i�	*ht���d�&�ʵz�FFrѐ��شf�������?�����<	��y��פ-�"��'A�{C~P�C�K3c��'{ɧ�O��} �i���(o����w�	� gP
5�$ �q��UQ��p�O���|���Im��uMٻ0�8L�U�T������?Q��?�)OhEn��:���	͟���:8h�	i7⌵c;���@ޞ't��?9QU����ݟ�%�p��M�LPY#EÖ >����n7?�F��-r��%h�'x�����?���C-t�.][���,)Vf�`�	�?Y��?���Zm�d��y' ��eU����{��q�ą��!xӫB���?��=Z���'��i>� Ds~��B���qĞD������Ԧ�	�4]<�f-D�V�f:O���d�ވ��OJ���4[0�,�Vj���F�2�|rZ��I�P����H��ҟP�b-�~8�Ro��o(J��|y"�c���QA�<���'�?i!�M�W(	� �6*Ӣ�+P�_�8���'�M��'g���OK��Y�E�:X�HM����^���X�	�K�\�8{�@�b2�.�`�IPy�b�	r�<:�˒�Y�\>B�s��?Y���?���|�)On��~������%�N|{4��OJ  �eα���ɣ�Mˉ2�>9���?�T��'���Y�Ј�FD$��X� �'�M��O��#aMA��b����wY�A��h|��iQ.
(w�p�'�b�'��'p��'���s�d_�[ۮ=J��
.5E�E�%B�O��d�O6�o�	�F���,�ܴ��:pvՑqDZ��Qse�dI��x�j�oz>Y[桑٦5�'w����n���p���' ��u0�C.��	j*�'��)�s���uJIlb*xX�B].g~�)C�(�#���E�%�	쟄�OM�Ȳ$��@�:dJ��R���B�O8P�'��7��Ӧ�`N<�O��t�!��[c��+%��5�N�2,�6]녽i|2��|"�i��@�<�]1CF�[�͐� s�f�ğ����������b>E�'HJ6�N1m@�`�+W�nht���d�Wn�H���Op�����?�Z��ڴ1 `��Wc�]�dx��#+�	�i�h6���V^6-)?�G#?Q�l��Cy
� 
���+ˏ$����FT#o8άG5O�ʓ�?Y��?���?y����-8��"( ��T�0훳%>��o�cpm�IҟL�	n�s�����e�F�B�p�L�!Cjl̺��ь�?i���Ş+�\��4�y2�]86t�0j�
G�d�#+4�y�cC��D��Ʉ>��'��):
1�:5j��S
O��}Q`Ɉs���ܴz�ʡ�,O���D��Đ���#a�B��c�F� c�OD�lڭ�M��x2�ѩ:T
���@I�t�P��i�
������:x���d�2-$?	���O��D�W5��sF���@ �Be���OB���O
��%�'�?����$����(_,wOVՊs���?aC�ib2���'s�~����ݕxn�Q%)L�\�1��'iP4�	꟬l�.�M�� �M��O~��R��4���!�C+B�H1M��P�xVh�7oR�'���ԟ��	��0�����D#L��FO�7=���@é�)U� �'�x6-�?sTF���O���:�9O�2aӳ3f6�ʇG�8M����Emy�'n���=�������$��eI�*�yMQ� �f�Ӱi��˓j��I&ï�\&�<�'l�����,#}�4�B�cJ��S�'�r�'m���4]��0�4 }��A�����m�ɠ�e�-3@\�9��pśf���wy��'A�F�o�nh¡Z�|�!�&*F�A���	�fO>T�6�,?ig��x�j���-:��/ZS>�x2lСBq`�X#�j����˟H�I˟x�	蟔�
QeN�n�Fe+�A�E�d�0�B�?����?a��iN��aʟrmo�q�	<o�̋�&�a����-ɦI�&��N>���M�'�����4��d��*y����T�I�(��
o/~��u�^��?ᄩ"���<�'�?����?�0@��_�c� P��,qhŧ��?����$�Φ���ƍ����Iğ��O��pB`m$:f�E�d蘄_tj�Ot�'�r�'��O��O�иc�D�qC*Y�BnGi����	�<�JTǄ1?ͧ{��d���h��Ғ�ʰ<��a� �<7w(\����?I���?Y�S�'�����)
�_7��x�$<9h����)����I̟�B�4��'���2S����>\oȡ�ֈC�*�J��%uJ�6�L���Y#��	�'d�Ɂ�Ƀ�?���%2�dݜ:7^��aę�3]<�1T7O�˓�?!���?����?�����b�2�b��D��,3����;s�lZ����I֟��I�?e�OP�%z���^�PZ�H�� PoPmcɊ=en�mZ�Ms�x�O�4�O>�A E�i|�A�ai��O�d�8��H� y]�$�P��h�'+�'s�ʟ�	�d�´�W�Ŵ!�ȕr!��
�����	����	Ey�&v��Q�T�O ���Ox�g.U�,��cO�%�v	��7��O��'Y�6���MII<�S �=z�PK��<B5�i�UC��<)�=����M�S�|�����$�ObTJd�O�����q� ~O�U�H�O��$�O@���O�}��e�Ѧ( �����Ap>J(��I̛���Q�"�'�6�2�i�a�� E�$�~�8��E�v���
e�dB�4{���� �	u a�`������?=��*�4���ƏA�t�vy��i�Q��kyr�'���'�R�'Sb��^�K��mw(��/.�F�-O.�lZc|a�	����t�S��I�	�tK�y`s�I�D�zM�@�����O7Z`�)�IR�M��`eJ�3H �@
/t���E#t�~i�'�x�`�$l?�L>q*OrI)���|pfU+@�#f6�s#�O���OP���O�i�<!��i��)���'�fI��k��7+���%MV�[��0��'�b6�$�ɬ��d�O�6-��9��J9m�T��pDG����l�g~���a��M�'ſsu�Q xך�p�k[�m� k�#R�<����?A��?���?��DB
)4����CԵ_=�`ص �7�b�'1r�cӆ��6�n�$��%��p��6��eBSGP%>w��(��O�I͟`�i>m��Ś��m�'5��pA\(@
�Y$$��2����u�Y�)ƕ���EC�'�i>���˟X�IXGRIx6�Q��d��S�8���	ן4�'�n6��������O �ĵ|:��_�a&�ш����<���A𱗟4�-O<��sӀ�$�ʧ|H�� c"ÈВ�ᓡR66A�����^�p��4;4�i>�r��O��O�Q�7��(>�9E��6^֡j5o�O��$�O��D�O1��ʓKR�#Wqk�̈́�#��	2�(��o�>�Y1U��c�4��'��˓�M[&��f�:9�qN�W��iQ��e ���y�ja�t�xӺ�eΞ8sa��?��'RT{d9GsNd������к�'P����˟t��֟���h����(��l
�7H�0���%R��n��c� �����\��~�s�X���3c�P{0�hĆ�>�̰"��,G�No��%�b>Q��I���|�V�a��"Q���r�cW�&0�`Γ�^)����$��'�'�L:��/���T�r��<�@�'���'�BX� ��48ll����?���@SpġsdN�mf��&��	8�<���B�>����?�N>YUo��G|��+�cO����C˛K~Bl�#:�ڝ������O�؍����Ba!�D�N�?�PlrP.L�S��'��'����ş��a�J!)���C�M
"^^�2��,��4"&MY��?a'�i��O�ͬo��C�n����(#��&�d�O&���O ��g�`ӄ�{'�ȃU-韪m� *���>|IB8��92��ū#�2�d�<�'�?����?����?��I�6�2=�тڇG� �W����D�ڦMhf#�����	ǟ��ҡ���8j�'�9�(�B��3P��ğ��	T�)�S0*�H�C'S"eM�I3A��U$h {�=~ �T� �H��O� BL>y.O���&L��/_���'D�7t+��Ѥ�'27�=p���D=��A�&�K#����;I��¦��?�Q���ݴj��~�l@S�H�S���ˁB�ܶ4KD���:7m6?��lC�����B����x�+�R��`���M IW��5�d�d��	������)C��r�ܱ$��q�'�R�`�>}��?���4��1�������A�,7J�@�S�x��y��\oz>��gm����'gy)��:eEİiǍ_�$��<��mȀ��������2�	$%8d�б`��z�S�P�"<Qq�iȸ	�R����X�	^AF}G��7���z��?���i}��k�b�o���S��#ږ1ۗbӣ���@	p;��b���h�恨<�'F�,�IC�	'V����Τr�^,knX04���͟8�'���T]�@۴d��Ӆ
�D1��]�q��
 �ű�?��{՛�D�s}�'�a�㊈�1��#r# 5��C��'���Ђ$F�6���"bg�-A����~���?��+� �)yA�T�<�+Ob���,�R����]��X!Mܠ�V1mZ<[�`�'�"��W��]+ބI��ɀ�+|5�W��N�RU���M�%�|J~����M��'���#�OK~���/��tj�'���B1�q?yO>�(O���zމ#C��$��,��D�% �$Zą�Od���M������_ަ��V*͟l�I�p��`�,e��Ke⅝r�B��'i�F����Ɍ�M;��iu�OLؒ��<
�d-�`�O�Zs���R���Zp�D%v�RDl��'D�r��ɟ,�#oT\Z� �Qݭ	F�a+������IƟ��I�`G���'�d�C䖭�R��&�	�Dtsp�'	�7�W����On�lB�ӼS� ��5H��X�$�81�� �$���<Y���?Q���
%�ٴ��d�7-8͉�'9�NQ*��S�N&F<�!n�"�`A���4��<�'�?����?���?���nǤ�#% 5~f�=Z�'���Ŧqc'�ʟ��I�� �"E�#j"`4���L�'�j��*P#|��՟<��M�)��a��y�A�	[�	�@��\�ڌ""�
������QU��O���I>a-O2�81oԒ5�H�j1|Rb� �'7--= :�"c��j@L���	sB%q�Ě��?Q�Z���4,��� q�R��� i�������	!�M �� eq^67?�6I�('��SM����5�%Y�x�JW�O}��PV�|�\�I��<��ǟ��	쟔�R!*�]P!���	�M)Z���'G��?���?���i��ta͟ęl�u�ɜ}& �t R0}e*��&J���O<���?�'�ܴ���>> �d �Vf�`	�[ M�d�gͦ�?6+6�D�<ͧ�?���?q��	'1.�,�71\QZG��?�������͟��bb�<����ٖV:�Re��:\<jS$A�	"��$�O�6M�j�|2`��a�����) vO��
ՃP�,���Ɯz��e��$�C̟$�О|hO.k��1c���
ڤ�[ :�"�'C��'��DY�0�ٴ��P#o��+���@�Tj�L�2���Ϧa�?�@R���ɱ>�����h��ѫ��׫�:���ʟR�ͦ��')r�&Z�?E������J 2q��@�j��W:��2O��?1���?����?	��򉜒
8���þ��|r��E P1l\E�u�	П��Iy�s�������'����B��!0m��L��?q���Ş*/�=B�4�y��M#W ���Sd�AN� v�H�y"�J>SԜ��`��'Q�i>���=��I��M��l��(��^�Zh��Ο���̟L�'w6��%kl���O��$�@82���A@7T2p�k�"⟜��O��n���?�H<I��X�<��� t��9�D�%�y~��Q�0�@΋!�O��	�hRk�%f�`t����f���֊y�B�'���'���ퟠ�2��:�¯,yz�AX�$����P�4g�b����?�E�i(�O󮝵H>��h�
�8Qx�B�s�$�O����ŦYZ��צ��'�,�{�D��?Q�q'˯ഹ�so�R���`�E�:v�'��i>!����\��ܟ|�ɎYk>ip�%X�v��̠�o���\�'}V7��W�˓�?�I~�� ����an�C9��(&��� �����[��ٴB@2�x����K>z�֜����(@�����V/ ���g:BE�	�R�Xݨt�'�1$�ؔ'�昱U%��=�F�#�.�P��9e�'w��'�r����T��:۴HB�b��V��\��Ǳa�Z<�&�6B�{��4:����Hy�'C�v*p�\[���v����b����1��gW�76?�7��6]��I<���߉;2f����/q��02ũy�$���<���H����t��"��w���I9Q'���͊��?Y��?A�i�:���U�x��4�� � �c"eŕ�z�+�-ք�@e(J>)���?�'aJ ԁ۴��dH(h�� ��1�^	�0��Qo�v�;%���?A-3��<�'�?����?�4�̨D�|p@#À�Kg��1g���?����Oͦ�ɕBT�l���ȔO�J��1�ȢU!���Ȅ$}Qr�I�O���'1��'�ɧ�	Q*�&L[b�J�}��g��W�� �Kֺ6䬵�g����.ui��Lu��t�^4q$��F�<��[w\���Iß��	�T�)�ay��u��	Ԡ�9Sb�)���-����g&G�}r���O�!oZr�B��I.�Mk�
�	{q�ţV�H[H* h"�M���Vn�`q0�al�"�xpR�kF@�?�'�@<Y���F�J��
�~<JX�'V�	��I����p�I_�daGe�RP$
�rv���ul�rZ�6m�/7�L��?�H~���Mi��w]�M�����v�bJ�Y�����8�m�:��S�'{��[�4�y ��hYL������P�#�&N=�y��ĺm�J������$�OB�D�����A�7G�y��<�h�$�OV�d�O�˓R5��fP��B�'?2��G�
m�U�\�y�<��EIG�]`�O���'r7���p$�@�u�	�FU8oܸm�Ab�E4?�p$�8Es\�����.��JvB�dˮ�?���#��hK���.jJ	�#b+�?���?y��?��i�O.�(�"&�P��E�Ar�Ҕ{���Ol5o��j!�	ڟ,ߴ���ywC�@ҵ�u�>XV���D����y}�n�lZ��M�%H��M#�O������KQ5��uօKв�za�n��'�X�'�"�'�B�'-�';d�z�
��LpY� ���@P��`�4FVB�P��?���'�?�U�"T���h';�rܐņ]�s��I��M�Q�i��O1����$~)���4��0W����+��IL|�ٴp��_;40 �O>�O�i���蔿c�>0�#K�J��d��?����?y��|�,OV�lک#0Y�	�]Pxp�G�ig�L[���"N(e�I��M����>���iƊ6M�ʦ1�f��M�.��� �:,�3rR*<��n�c~��H1H������'��c�9����gG�B[�xW��<����?���?����?i���a�ԳCm��/
^pöD,,yb�'�$m�N�Z���<A��iF�'`�\��&ʼR���pg��eŦ�S2f/��צ����|��e��M��O��)Rɛ�M��x K�8E`�ZPq�����'�'��	ğL�	ڟ����I1���k4<�K��U�xS�x�����'	n7�צ�����O���|�ĥ1]s�0!\�r���!GXU~�%�>����?�M>�O�¨�1hvZ�3"�����rR/�7!!�}��E���4�P����q_ƒO>(�E芐/��uť: �%�@��O��$�O����O1��ʓ)���akv���%`�)p�G����'�B&g�D�O��DLyr�iC<��D�د N��� KM� �L��W�s�^o�A���l�<����2F�?�'#���7�<9P�Ҿʈ[�'�	ٟ@�	�������w���Ƨn8�ƙ�f(��Ebn�T��Ǻ<����'�?I&��y�&i�
(��'�:��p@N�W��'s0O1��m��m�l�`�XX��S�/u~yS����;��I�!!<a�"�'7�$�d�����'�f�jF/uW�=�֘u�Ny�'��'�"Z���ݴ<�VH[.Oz�dչS����ɞ�q���T.@6^Z�tY�O��n���Mst�xr�ז{�)ZA��a�<�3E,ה��d���*$���I..�1� ,���)���Z#���zď�z�*Y�ls֚�D�O���O��8�'�?ᗏ&U3�p�#_����oW3�?qW�'Vx8���?5�i��O�3L�T�"�ܤ[}`5�&Ǐ)Q��D�Ѧ��4\����ܣu������b$H�R��ti�����#D>���g��N[�y%�������'7��'���'�<[��2&qr�үO�`���U���ߴcց!���?i���R!�Q��?��;��*�bհ������\�Y����R�<�I��J<�'�?I��r�\��F�-�~ ���0Z�v�(��?o�~��'�v�Sq�������|]����D�đ��	�`tt��0 �ݟ���柸�	��Uy"�p� ʓ/�O$�� C(r�1�6+C�Q��!�o�O��nZt��M��I�M��iv6MQ�1)�"�vajw�H+�H��K{��!�X̛D �?�&?-��3	��@��X�l%�����]$G���Iԟ4��ڟ��	����J����å@�GE�e�aL:j����P�����Iş��ܴ(��Q/O�nZi�In�j���N����T���	���N<�5�iV&6�r�j��gӢ�	ݟ��&�Ɣg�r�ZF�iZ�Z!gR���iV�'�N%����D�' B�'CB̋`@3nz±Ia����a��'BbV�л�47�A0���?����/x<P5!HS( ¬��ϛ�iK�����������ݴỦ��)م(��Y�$D]�~�#w���_e�]Di\J0b7��]y�O��@���h�rc��� u�F+�6%*���?���?�S�'����g��4�BKT�Ցb���g:L����H�޴��'N�˓�M�fBYz�:``�* :�9c�O>n'��k�B<��z���X���p�?��'�b��bD��m�`I�##��n�S�'@��L��[�c� C(D��m��%-4�������M�A
����O��?�(���K'�Q�n��͒���9(�����׈tS»i�R�O�O�6�f�i:�� @�ōW�=�J5�ݭx��jA1OrUJ���~r�|�[���ٟk��
k�@�r�$�9!k:uBrg�����ퟀ��by�rӌ}`l�O�d�O���3O����%���ñ-� �rf�+�	��D�O4��q�	�kr��Z&Mڢ�����:5��	$ EC�+�<jBU�|���O\U���E�\�Ggԗa�Ƭ:�OO�F�L�����?���?����h�����&*X�co�y�r��@�������M�`�Ο@�I$�M��w`����+P�L����c
O�F8@}��'|2�'��6�M>)�7-,?i�gT#���)I��1�U{�b�s����*��L>�+O���O����Oj���ORT� �,��I�"�2#gPQ�5�<ap�i���0��'�'I�O�	S
Oc��Bf^�
B��ق�Q�&��B�&�iӶ0&�b>ʥe�&�����M�X��L��r�l����d
r.(�'"U�X�'8$TBp� _��4H�D�!1
�8!�'z��'v����V��`�4P4�����l��䦚2x-��k5�tJ���it�&�đ[}��'�2�J� ʓ-h`ftI�l�3L��:���+�6-/?��ӗ.��;���qc�Axjd���P @�(��o���	֟���ϟx��ٟ���kF!5�BE�6��)QJ4�?a��?1a�i�(��On��i�@�OX��A"��?��e�0�#Px2�A�I�I㟜mz>=���ʦ��'/J�!�ȍ7�*��耍 PsC/Tt�������'u�i>��I�t�Ii{� ��?�61x&�(!��ß��'p�6ϸ����O �ħ|� ɒ^���!��'$���c�
w~��>���?���xʟnX�œ�ws �a�i��B��uZ���%<Z��@����i>����',�&�@���5}����!�Y,G �A�,��P�Iퟜ�I̟b>��'ܨ6���x^ hW�Os����A�B9u�2�[���O����ܦI�?	�V��C�4]8�Y7a�:V�|�3'E
>U�PҒ�i�$6�ӌ)�`6-<?i'!ܺZ�t�]y����c@�iR�]����y�]�L��������ƟL�O���[��?3YT`����%��$emw�l<(t��O\���O$��H�d@Ӧ�]�%��l9�-B�Kvp""��3}Pڴ]��&G �4�6�)韾-�Ůc�&��Cr�\�!c���$\ѓJ��扄� aP�O~�O���?���v�r�ZIտ� �k% Y2G8`���?����?-O�\oڎ2�'�2Û�\7|T@�,p�������([5�Oh��'�R�'��O�)�G��g�n��B�L����QR���£���K��s�5�S�J��U���A��Zb4	�d��ev�sm̟��I���	ݟLE���'����g����x��$i*N�za�'��6m
�c��d�O��m�n�Ӽ{,�)7{L-0�V��ĩ����<q��?	P�i��x�6�i����RX�P��O�NQ��G�o�4��匝u)t��JU�	\y�O=�'D��'`��=c�\X�'�<!�JDq4D���(O�n�Y+�I����	M������fЌ(9�=�%O��q?�C�i�������4t鉧�O�ܡ{��x֑����	���d+þ9���Ϋ<Q�ͤV���E��kyB�P=��I*�*��+�+2��'��'��O��I�MSF�A�?9k��UӠ�(�`мA ԩҋK�<ᗼi��O@M�'��'���Z�{ߊ�:�OB�=�dP�#,F%��u�i����d`�f�O�N�&?���$��r(�� ��0�5j�P�Iߟ �I��(��Ɵ���r�'(�}0fo֗0:iac(��������?Q����/T#;��I��MI>١ ݀ug�����C�8țhٖ�'�7m�����%8D6*?�� � &�zЂ���^	���\�>���I�Oty�O>�*O��4cb���,2'-�A�&|�e�6i�VI/3d�Iߟh�O( h«HҾ�)�nR�P�$�j�O�'�2�i���O�rܔ��\a8(b�*�+S�=!ʍ\i`nZ��4���j�'��'ud��flϳ=��A�N%|��yk��'���'�����O��I�M��F4S��x��Z�t;u�L�R�$@#-O�5l�k��\�Iɟ ��D,!�<��-A�3M�%�r)��	���mu~rK*O��x��Q��]5����ǋ����b�$Α��<���?���?I��?1+��p�l�� ^���[Ȕ��Ն�mږn���'�b���'��6=�M^j�`|�bN��/$&��d��O��'��ə,b7�u��x��P�ta�4یu
��x$�s��I��Q4K�@�J��uy�O��Q�#�<<��3:_�`��
��'B��'Y�I3�M�d�V�?���?a��1,��ly �J� �4!�晈��'�����dz�t$��SԲ )A��I�I@�\�$4?y���^�"��4\	�O��U���m�!n���AFG�%�0�R��$V�xq�Iџ<�I�$��n�O���cI��Ь\�b��E.G�~R� �O�U�p�'�"��
�杝/�Id�P�d�J�`���I��t�	��M3R�0�M��O���2k�����,eu^��Ԫ��-�Ђ�	JSn�O
��|n�iY��'l��'��0��,k�z����T%D�.���[�\�۴S��%J��?�����?�����P��s�΅S"J}��$��4���;�M;4�iz�O1��}�P� �Ha�I��~� �����𭟔A���"jj�IG�'�J%%���'?���0b?DM)T�� ��$�&�'+��'(�����P���4:��Y����9�2�\�q��dz�Māg"�Γ��F�d�ly��'f�vCp�R)��f!��Շ��/�m 1jÝ~6�7?��A�(X���Q������a�� l�PI�A�*��m
ѭq�X��ӟ<�	��d�Iß���䗙��yB���  eD�1�
�?9���?q0�iF̼(�O%B�f��O�h�ծ&�p�8�g��OМa+�"�f�	��hoz>q 5a�禉�'G4�I֌mY@p��$��h�uj_--��ܑ�&��$�P�' ��'��'@&�I"���dC���LH��W�'.�[� ߴ\ Q���?�����ѨW@�8E,�iXr�M8��	�����1�4;ω��i4Y9z�`��A�]	�ׄ�"��@�ĵ�L7BLy�O<������.9�G��bJ(`v��#$��y���?����?��S�'��
�i� #�f��@E�	)��R�N	�'D 7)�	��D�O�-Ӂ�+6K>(��m�*O��m��O���91�7�7?�ƊǒKf��2�d��gy� DBU�i\ 䥙��y�W���	ڟ���ҟ���ן,�O��-�v�S�;^�c2߸*���b֮t��i�e��O
�D�OL���D����!�˓j]$]�h�� �87�a�	؟T&�b>�E�N�m���&-��G�����|C�)�`҂��t,Wj�HqT���<�Hzŋ�0x�� �e�M!@����/BNճ�D_*f�Ry�@/+���R�eW:^��5���+}\!S�*�1/*�ur"CP4ZǢ�XF5�I�c`\�q��@B��<������A����O�/��[�i��h�z= T��z��$pH�?���jV(�J��!�6�K��X��"=f�T0����m{�� �0S;�`��G9�@	8u`��7�ָRv%#*T�qs���Yθ�ꈦ"2��`��o�e9���x�&!�|<��̬Z�RXk��G�~�`�!⯛.שּׂ�e@e�.�$�O�u.�MJ�Lsd��b(�逷$��!��Q�	$��;aG���=�s��y�]30I�[��!��u�I����'+F�z�Y?��������1L��
f!ȃ.<=ؗ�2RX-IL<q���?1�g@���'H�IZ�4E���Q*��2�j�6��9˛����h� Ħ��	۟��I�?1��Ok�H/ �Ycd(�.J��(F�Dc���'�2�Ā%�r�|rY>��!ko�e����$�:m޸U�	�J�l�ӟ��I��@�S#���<��,�x3�ܸhJ09�65a`ېpқf+B�>��O��?E�����I�ɛ�FÌh��O��He:�4�?����?ɳ�[�(���\y��'r��ø_g:)K#d�<z��GM���O���$�$�O���O|�����Qj��2�ɞ�dd�	�/��%�	9^<���Oʓ�?�H>���&Б�+��#Ø�Pc_׌Q�'߀�ʏy2�'��'Z�	�b��@!�V�"��HBU/f:P�DIDA}�T���I@�I럠��;U�h���'�e�D��#B��$j��]������͟��'4^�	�<���{����9�PX�b�8?a<T�c�iJ��t%����� 2��>�)�)_zr��DN�ES�(!DH@q}��'P��'�I`���O�T�C
p�a`S(&2A��M�7�~7m�OJ�O��D�O$����?:k���f�8<p"��](s�iF"�'y��>�8��O}B�'��De�;Y�%� �A:y���n�y� O����OP����O��O��S�p(r��"E�P���蘹:c�6-%?Q���M����?���rt\��X�u�D<rc }�%�C�֦w�$6��Ol�D�aW�⟈�}���T�e�jU�s �15�P�փ\���*h��M���?)���W�x�O��كB.���:�0��/nl����
� ����O@���<9O~Γ�?)��dr�8*"�ɯf1�{`%�5��v�'D��'W���!H2�4�.�$����U0D;.|b���-Y��� �}Ӫ�D�<	q��'��s���	ڟ���VR(*�����ݪ����왨�4�?���/������'\�'�� 3�b�=a���J��>����k?��OX��?���?i-Od�ʳ��	J]$	xv��Y�x�I�x�$���	�$����u�ܳ2>�m;� �Qc�Aҧ�B5�M���D�O4�d�O��Db"Y��3�&�겉�>ax��F�G�u� �c�Q���	柠'�����$�'p6mB�	�Z��y	�K_$���cя ��O.˓�?�� �����O,0Y�@��E)��4,� ����.6�(�	���'��=�L<�֯�s��C�W�\ �$ �%��ny��'�
�G[>��I�s�):@�CWY�l�ꕞD��� �1��OL˓e�,EExZwa��#��lp�𨄎_ M� ��Oj��([����O����O��)�<�;'yhd��oϾVp&����mZ͟�'c.;���t"Ѯf�QU+ؔ5�	Bc���M��ɡ�?	��?i���2*O���f�����C&�~}�B,�.�t�i�O��)§<>���OU#7A^���� )Vx(<k�iCB�'�B��g,�)*J���g�;z]�%3ӊǖq� Iv�.�OPA�~z��~�Hԙ�t��ˍ�F� Ё;�M{�Dƽ9/O���Oi�O����k�*~�Rwǀ7y<�S��~�I����?���?�,O���p�0I�9B�k��I��d�3�T;,��'������4�'��s��=� ���4
�8��egƯj��dk �i��S�\�	џ���Oy�l�
l���S�xҦ̪QK�-a@�4X�땼W���?�����4�����t�|�;A �9�ɸ�����'(��'�W�Ā�ǂ�ħ�p�Xg�|�B�ু[�,�z��v�i���|R]����ȥ���)q�G�Q����� �3��Աi0��'��	�B��4�L|"����6�@P��X�+Q�@�[D�n�'��'4��'���yZw�%��n�U�8 A���p`	�4���_�F l���	�O��i�@~��Q32
����c ����4 �Mc��?���?����'3�s�0��k��Y��$
�L/ �֘��i�@`���v�X�$�O~�$����&��S<\��牉	��eD�=�����4�?Q��?�H>������/�L���Ck��ܣe���Qm����ߟp�3�`yʟ:�'��ǧ�;hlv��8��J$2�=����D���"�N� R Š"�E�r� �-ӈ�D_�7U�ʓc���n��!vP,�$�!t[:����<C�����xrH���'��]���ɟcKv���-��G��Q���)�ON"�ßp�In���?��'܀8�叾dʆB i�6d+۴oxF�'�b�'��_�@�E%A���L<����
��O����"�MS*O.���<Y���?��N�̓!xB�q�K�]�\4p�K�Nܾ�"��i,�'�r�'��I"$a������E/o���psO�$�\�(�1 mZ�m�şD�'I��'���y��'���ۈIG(��'�A����ԋ��};�&�'�2X���I���i�O8�D����i��5��=SSJ����j�	�S}r�'[��'�r�"�'���l�'LZ���2+ÁrG�T�񩘹xӜ`oZy��O�7��O���O2��y}Zw��YP�}z�j����|�\D�ݴ�?��и͓+��s���}*f�D�'H8IV�G=;g��C��榹� ���M#���?1��r%]�T�'z� !eM(�r�87��</�D��r�:튴0Ob�O��?��	�5f�X�e
*:����ܿS�]ݴ�?��?9���W��	jyb�'��$М���'j���z	)��M����'�2�'F�ȹ�����O����OH�#�����93Ğ4np�\���ͦ5��7W(�8��O�ʓ�?�(O���ƒ�:��bf��6,qa��>6O�&�'d���'���'��'�2Z��k�h������6g	�X��-4I��P״�2�O&˓�?�-O$�D�O\�D�,NF�X"��*R�S$��j�`��5Ov��?���?�-OzӔ��|RF)۳l�V,$�8`���`�ʦE�'�_�@��ʟd�I�M��ɵg|�@X��_�����Ŷg���(ܴ�?a���?1���<t}R��O4Zc�P� �&RL�,qjN-fsR�qڴ�?1)Oh�D�O���D����O���N[�h�p?���IANG�Imϟ��IVy2��4-�2맨?���z�iƉ���R����%[9r���OJ���(��ӟ����a����y�ٟh��/[�?����bQ���z�i|�Ij���:ߴ/��ߟt����D��C�<TI�m�8(ȘY��ۻ= �f�'�R�H����|�iL5�ʴx���:4�aI��r�VB�p6��On�$�O����N�	���@�ǋd4��I�q*ГԩN��M��D�<�O>�����'%�k�� �
u �T�Y�'�ui2�o�:���O���ڜ.L���>���~퐈ogn���mҊT�Z�s'�O���'^��	�|��'A��'#���|l�/T&H𚤁��~�����M���>	�����[�]��UP��+,�N�x}2Vۘ'��'��P����C��h�zE�cB8(R���>H�N<����?N>���?��M5��$�R/�h�4ej"�� �������O^�d�O�ʓڌPW?���k'
��)�l�@�*�m1vP��[�X�I�,'�\�	�p�᪓Ο����2{Q&e���T��qD'������O,�D�O6˓ĠX��������J�hA��g6PUK
¹Gp�7m�O*�O��D�OL�z���OB�'-���s%!@{%Tjߧ|�H�ߴ�?�������"�%>m���?��s�J;0���*�kʅ9��ř��B3���?��{�`������t��4̈́�*����.�����M�.Oƕ�$���ay��x�d��^��'j��B�c[�|�NPqdDZ�h�4�?!��t��� ����O���8��Ŧ?�����
Y:R��x�4w���·i���'0��O��Oj���);��U"B�Ƴ�>�a�&��i`��oZ�^$(�IG�	{���?IV�ГN�.��m�^?r-��Ѥ͛��'���'Jl��9��ڟ��Kո���?=_�1���}"��n�w�	��@�M|����?1��nz�P���L�h�F�82��TCL�9Ŵi~&۝�`O���O\�Okl%Be��^�w/�WC�4*����2�8��Iy��':R�'�����8���P.)ya�Z���;&o2��'���|�'�"k�n�j���� ��ʥ�;�P��'��Iϟ��I��X�'z*��sau>Es���s)T�S ��tUL��*3�$�O�ʓ�?A��?y�a ��?i� � m �*�içj���b�/p��	ܟ������'m�u���0�i 9:QpT�Ǔ�(���n�)�,nw�'���X�i�B�>� 2�E@Ԇgi���҄�e��@��i���'^�I=X�l9H|Z�����)��U�p-�2;l^�@E�
'6L��>q�2d�в���S��)Bu>t]1PA�H}v�p!�˟�M�*OV�ۣk^˦�����d�6��'�L)�p.I�`�p٨�e��%$j�x�O���8l���d�{>�`�׎ ,8չ��7}
<e�^�M�V��u���'2�'��4�3�4����Td�C椬!G�L�I�ā���অH�iRߟ�$�"|2�@sT�pQ�]�@�hC �V�W��$�d�i7BX�<�����	`y��'���T�f`��`�#��)""G�$#���<�Ճ�\`�O1R�'�2�Jdl�����%��3h�t�r7��O��*��]x},�~z��?L�$�!�.]��
�0FD<���>�$!���?I��?)��?���7T�0�姒460�ЁA�/��u�-O|��?QM>	���?�7�A#*H^�!��ү[)Ή�޽(�N[u�g~��'E��'�b�'�dM�7՟�d����,��劤���Z�nI�p�i���'�R�|��'��IY�O��\2ݴ�j4�DO�=ȝ	��>UA�$�'F�'=�V�h�v���	�Or4R���5|���`��ۗ .�{�V�����ԟt�?�����'�aqbfA�>#� $A�z���4�?I��?��q:�}����?)��?�'$N:�aR�]�ʭ���wl��kP�x2�'���F ��DЏy�������rh�h��f-���3�i�R�'�k��'Cr�'���O��i�M���
Iҍpb��inY�a�{Ӷ�D�O������1O���X��N�V���
T M}6� ԼiجػЪj���d�O����X%���w��k�Hdv�t�d���Y����4�򀡉�Ϙ'�"�Ź8��������I�X�I#"�0�L7�O��d�O�&�O��D�|���~�CT�]� t�-���j� 1���2ĺb���G��'�?����?����r-�ą�ELa2%��1��6�'�Z,�1�#�$�O��d,�������bTnz�� ǥJw$��U��j�&��쟈�	P�'��\�Ǒ�<phȸF�
��	�`�,a�O����O �O����O�8��D�}�hͰg�ܽ�2$�)p1O\��O ���<�5�fe�Χ4ĸ�6
L2�Uؓ��<�8��'b��'.�'c��'o^,ӮO��SO�  �U�ԅתoֈ p�V� �	�����[y��� *}���ԓr��N�� � ���qb�@Zڦ��I[�������<U&b�r�#�=Dpl�E�R�)���aq,m���D�O*˓o���&����'���"ܗO{ڈ��_�u8b�B��,.�Or���O����IK���yU�T"�J
������ͦu�'J�P�$�gӴ��Ox"�O�~�W�4aE5Cz!�����h�mlZ���V�v#<��tB���H�W3vl.݋6�J��Ms"�бU����'�b�'v�4%5��O.��@A�Jq��C!Í�!������3g-�S�O-B�75�2cGa �*g�u$С5ZJ7-�O*���O���F�i�ٟx��l?��Q�!vRR��( ���B�
o�
ۼl�<����?���G ���
��_v�XD�F^�Ry U�i�r`�7s.c���	X�i�m��D�2Ub���)��WTVm��b�>y⤌W̓�?)���?�*O.xK�B�(1���:W�J�?T��,-6.4�&���	֟($���I֟`�h��=��s��L�Y�٢s!��KM�b�0���t�I|y�N� F(��p��A�D��7�����ߙו�4���O�ʓ�?A���?�r)��<q���6�j�psh(|��y (�	����'�b�'0"Q��(��I�Ok�Γ[\-:c�VX��\2��Q�Z~�f�'t��������d�Kh���M[2/�f���`�A�Y3*]�P�Cڦ��	���'�X�h�~���?!��<h���'I?J���h��/&���T�T�	ß4�I�r�N�Id�	hBҋ��0�*u��A-H���G7�V\��r��e��4�?q���?��'J��i�}�+�W����a㗉V@�p�J�|��OB=jf9O\���yR�I�R%2��`OՏ+��5ӆf@�L���r��7�O���O���}}�]�t*�쐪n����c�P<T����rlZ#�M����<����$5���,��B�+|��iJen�> X�A�EF �M����?���'>�ȗT�h�'.��O��x��X$m�N="`��#="l�R�l�'P^��O��O��D�Oܩ�D� G��p"f�:"T���o�����	pƌH�O���?�)O���Ɯi�r��:C��Iq`��&-C��
�Y�h�u�e�t�'e��'1�U��D�E� �����ea����fG�u��K�O���?�/O��$�O�Ĉ�zK��t[�&��+�W�"�A0O����O����O���<�%��|z�iJ?���Yp��	w��e�9=�6S�<��ky"�'
��',N]�'4�=
���(6��a8Q�ܵ.r��� �>Y��?����D�+&:��O��[�z��Ȓg���^x�� hk�7��O�ʓ�?Q��?	aMQN��OJ(5.J�^�"u;/�6Z��"#�i���'��r��x���'m��O�����ߠ0|q)K/�ԩ�U��>���?I�C�^������ ��WJd�h�ΐ�✦�M�-O��fM��i�I�`���?A�O�N�$xޒ���-E�kʌt��g��'�#T8�yҬ�~��π ���$LnZ�P�E�,��HU�i�:��!k�T�d�OP�D��i�'X�ɺ%^��K�"}��	�����[���`ٴ2y`���?����?���'��	k�슚rA~�K'!Hu\��ne��D�O&���Ox0��'A�I��,��v�e��0bQB1���x^%l�ϟX�'�<�p���i�O����Ot�D�'M��8@�O�5���c�Ӧm��l1����O0ʓ�?�-O2����R�
�d�<���K��f�!�i����%�y��'�2�'��'剮\�:�����Ra|��u)X�Gm�=zQ��!��Ĭ<q������O����O-CF�E��A�OM�&B�qA����eY��O����O��$�O��N�b���2�j�S���2F��P�i �g��Q��iA��ڟ��'@��'j�����ybdU��l��
"^�n58��U$6��O"�$�O"�D�<�#(Z/=��S���X�E7�:7�	 K8����\�6��O`��?����?qri�<�M�P�rǋ2Z$�A�_e��2
Ӣ�d�O��=6M��U?��	ٟ���/��XғW�I����B܅f�.U)�OH���O,�D�%}%���O�����	�4�l|i�%�=^t�$�e���M�+O*�i�P����ܟx�I�?���O��
���0a���}��+jڃW�F�''�C��y�J�~���O�kR �K���p5�X
��tش4��$HG�i�'\��O.듔�[	�d|��!�Y��}jSc��Xm��7�"<���d�',>�{�ǚiIf��$��e�6�5Ci�v�D�O��dSL��%�'I���`��;���G�˼�	 �%̮U���l~�I�"��)j��?	��}�V�q���)��U�o�7^pp÷i/"H�,
��듴�d�O<��?�1v|��R��c�6��� K�p�\��'N�0	�']��'a��'Y�U��;3,�SG�R�F� o`��s	P��Pp!�O���?y*O��$�Oj�$��4+�M(c�	RfT��bŢR<�+R1O����O"���O^��<����;��	�QmlĈ6OB�Q\(Ѱg�|��Z��IBy��'�2�'�@�(�'��,�c��4����k
�\���X�m�|���O:�$�O@ʓB����U?��i�i����'>O(@��D�[y�|Yv�y�|���<���?���}��͓�?!��wT���  �蝛�B��y?Z�BR�i���'r�I08M��x����D�O"�iy�!�E�9� U� P�H)(��X����Ο@���\]��g~rߟ~��`iӳ���IV- z=PMJB�i�ɪ@��4�?���?���}=�i��3�k�m��P��(w��@�b�h�z���O�5�`9O`��<Y��$�̷m00
EjBJ-ĥ!�`���M��AJ�"��&�'a��'���+�>I+O�mcfKM�=Tb�;O_(��3'OΦU�B�`��$� ���U��kьB+t���x�Z�+_^�9�in�'�rH�:_&�����O��	��$�Z V|8�"�+�6��Oʓ��p�S�T�'��'�$��! �Kd��5k�@U 8�ns����=1����'���`�'�Zc�8���$I�x�"UZ��M�:���OH��<O����O(�D�O���<��L�`Ţ�Oky�谅ݰ6sR��a\�x�'�R�|���4̧C�@\�LX�T��� �VD��ao���IП��џx�IMy�h^3����0m"DyYs����Ed\+�~d��4����O|˓�?���?Ʉ��P�T��Oֺ��%�	<i��A�k���M3���?A��?y)O�i�Ct�t�''>!�F�S396P�s�ִ:��� C�m�j���<����?���O������T�b���oM�0���R�N�mw���'9V�H���[���	�O��D🪡�`(Q7#uک�4�'�2�SDP}��'N��'cT�Z�'���'��ܟ�D�p` �C�L��oǤ&E����i剷t$�3ڴ�?���?q�'E�i�}��EF�Pߘ(r���*	~L@�yӲ���O$9��0O|�d�<ً�D�N����W)�a�Ф����?�Má.޵o㛖�'a��'��t�>I+O���`;*�pa8d��p�z��&��@g�s��<�B��;���"`�T8�Ƭ�m(�9�E�i�'���ݦGA.���D�O��I5`Vڅ�f��5R) �B	�,`7��O.��O&i��0O��Ο,�	؟\i�aY�2a�I��J�C� ��c���M��a]��xTX�h�'��Y�l�i�y�3�&��s���">�2���>y����<)O���O��$�<TS>v�8�5�L�d�c��L�^S��@P�D�'�rP�@�I�t�ɛ\LB ң���X����C*+�5!B�j�h����@��Ɵ��vy�a�j���S�BS�Ʉ��X��)�K�s��7m�<a���D�OR���O*���X�$ F��'����!{��䣁�|�*���O���O����t�'^?E�i�E���ha��9c*�M���zKyӼ�D�<���?���M������$xK�MZ�KE/��-af�B��z�[��:˶<�rюS�������<!��v>!ȃ*2^���D�g�<ijnɠ��P��#?��Tz#	'�9�,�	)f�s��!>�x�ЂK��c՚�9P�S�.���B� 3�L��"k�!-b��䆐�j`:�c Ǝ�s��A�=�ؘ�.�5+�Q`�m�;
4T�ፆ?�� �r܋
��dK!�W�8h%�2f �H�y� �� �����d�����f�t�.��+��?���?��!��ƒ�P��$�J�Vn�R-s2�)h��E�Y�(�[�C�O�i����F71��'���i��V�nԚw̘�(�� ���rެ�8�	�O,�+�ˀ�ȸ��BRq��_jZ�sd��)=|u�����$��r�O�ў� ��S�\�(0Jm�s���@�"O(���$��:���JJ�d���'��dx��4���D�<��!�d��%��bU)�a�1h����&�C��?Q��?Q�eQ�N�O4�d>Z��X;��ŻR�J�@�$S���9^	�-Х;�h� 灇kx�H{���B�}���8\ƅk��$/�Y��V�.��0�&��ax� A�%B�3�`�DM�oT����)'l�d�O��=���.$�2��"@��.��Q[2&�7�yR�� ��iI&��'0H� q�å�'϶7��O˓{�h�U?��I75W��턏_v����B.?����I���`��������|�#kʑ���j2ߌ�jش2QL�жD]�y�D킲ᛕ5��u��ɆB�4Mc��G����a�ͦM�i1]z�ic��0'���D#Oz�1�'BY�@�6�IJ����� Z��xro<�	a���!�Ы;-j,�t�Ĵvj~D5�:��ݴ_#lp3�����@p���fx�����䓪N�o����M�d��c�2G�6h�6�� FBQO4tP�`Uy2�'r��p�B�a��9���n}*��' �����*)uni��g�x�ФOd`��mO�����[f�OǨE���W�c�]��
�W���H�4�I�O�b��?U�3�_,��!��i��fq��5� D�ȫ���v�:dC7+���P�SG=O�MDzR��.���9��0?�]*���0az6��Oz�d�O.<�"�D�\ ���OX���O��Y�X��E"��"t�ɡ��{�@���-�=6:���F	-bP�d�9�3�D�E�]��h[�]��;5�ѓE�Z�Q��k�j����(b��8g��|�͛i��\�t�6n�yjt�|�4�	@~��S#�?�'�?!�r*WS6=�� ԞT�ڕh���:�y�fۚY��CaɃ[��	!k�-���m���)�<�3.
�f�JQ�w�*I�H�׊WNa�hHWO
�?����?a��du�n�Of�dx>�`��!y�z�1��H-�|Q�%�"s7�B�I�N�F|�����DP�ש*��!�(�`ءkX��Δa��ȃ|7��"���90��-�O���+Ϛ �LL+`�\ӧ"O��U�e4�A �J�>7�ъ��
A�9y���R�i�r�'�9`���z�x����;��*��'l���5~��'N�	ƾL��|��єE�@���V�o��@��f���p<���WK����I��\|S4��3�$Շ��+p]���/�$ŕ5�j�s킺KU��sy�!��-J�\ ��
�,Y�G�rA!�NҦ͂���?��37�ȕW��I8�)#�	�U�Y0�4�?�����I��0|�dG��fL�ҩ�<8I 0K��l�d�Ohl3ŝ��l&�ԔO哘X�̥��OΚ�P��S�lք�'�^�
�
��S�B	��P"�h�"U���X����J��'i�){Ð>!�ӟ�I��M#���OQ�x�i�%L���D����$9��|��'����yB�\$7���y�oظt_��A��[��0<��iu�7�+�d
4����nZ�h�
P��C����'sr�'릘p4�D%���'e���y  �(je��d&�4Zf��~́ RE��F�.	Ae⃸_"���|�e�V��a����%BD���历t3:�X��-K���X!D��%30�I��L>YP�O  03�NO:^���醮�?1�Oz���|���$S��Z3@[�%�٩wH��!�ME�\�/�mþ��f��Qx����HO��Ry�M=�^ģ�L�[��-`��$���Bo������?1���?q���$�OL�S�<1.܋#W+~�49@��Z+�HI���o�-�Fl�$�����2�\a9�=�Fe�ĉ�/��5:�(��SBY+s��O�azb�Ʃ/�j�2G��CGr����D�N�����?����6�	7K�Y{qO�9�r��7/T�4�^C�I!�n�@�:8�T�?�b��j�O��m�X�Ŷi���'������3B*�РeR�m���:��'�  2Q��'��	(tn�|�-�'F,�y��� �"��*�?�p<Y/U��
�@H�q%̇��AyU��I�ꄇ�	�2�$4�d˅W�Z �e�Ðp�~8+ )ЈG�!�� �y�Z�B)G�`kFy�G�C��!�$�����JGZ@Ms�n�f������7�	�o�r���4�?������$�j�� 0)��;tC�6@ᦼ�Em�zP���O�Y
'��O�c��g~R) �tHDH�Cóa��x���.���W�N#<�ZG�$vj\��ͭ~A���GAJk�$ޛ[���'#��'<��+T?A:|؛�o�S:�=ڑ�$�O���� ���+O42t��b�K{5�qr�'�\"=Q�D\�Df��`�V�u�[QJJ:\M�&�'���'���ѧ�Y�D���'��'��_a9r��i�Z���z5�uM1Ouv�'Y�PI��M7�n�k�h)�{�e�.��<�@)�5U�r�*f�W.��)Q��E��'��)q�S�g�	4
=*y�+�Sެ��T��.H�zC�PL��dD�����a�&<�x�t�"|b�`��%/������	<&�B�I-+����𠃐3FPQ! �MȎB�l��R�.T� };u���jB�I�`�M:S!����s�I�.o�8B�	�-	�mJ"��dY��``�55JB�	�I���1vޘ/��E�wG��pC䉏z�8��3L��x����d�_5iHB��
a�\�
�ƙ�E_�hX�dC+t\�C�ɪVk.���/N�Z�l_ gz�B�� 5QX0�iݴU����`	�v�C�c�Q"`״V����녅d�zC�I1m��UÕ *g�<�@�;/P�C�ɣ!?��"��U�v����_KӎC䉆7<nh3�[�b�%��Nٻ:�~C�I3JH��A�$-�(B�#�?H�PC�I�T�z��MC.o٪p1D㚗:{C�	�	�l��䟩 ��̚�i�6K��B�	r�ĥȂ-Z3[AZ��嚨݄C�2U�42)�:% x�(��$dC�	�?���ä� h�
�7��DN,C�I�f�U5��At��S����7C䉖a�l��W�QE�����O,g�B�I:TV�P�Ն�4^�z"��4،C䉿"�j�@&kK#2t��z#��J(~C�	����c؅TV䁑�	 �8B�]D�XqÎ�3�(*�q#�':Z��5BA�uP�P@A®�
���'����Φk:��GMD���ͻ�'�&YR$"�L�>i�v�������'�\r�{�X�+u"Æ|��h�'\��ydʉ�,醁�U�2װ�X	�'�V@+��-v��%~�d�R�'P��#@O3rt@�SE!ݪ{�����'_ޘ�$F�y{�E��mè%8:�R�'v �c�J��wU2��E҄�*���'N�4)�rR���cBY��2�'�&DCS�5q�`y�q��4c+~a�'����kI|T(�۽U:��
�'���'�UY���)ìB>T�Bp��'<���O�Y~�x�"!Q^��	�'�����K���"�I�P���a�'�&U��59"RX�Ԯ�K�l�9��9�>Pѧ"�w�'�>� t�L�=�T���PR|JE3�H6\O�}9P��Q������#!D?GV�xz�G%2v�&�X:��Fg����W�F=Y�h`pS�ҏ�*H�E<��¯W
* J�ML�:�l�?�+ӯ�|�����O�o�H
��I�J�z��ȓa�R���� �z%V(�`�95�(��$�M�q�S�ǪBI��M�‪|�'��x�ucß� ��gV�<��B
O���UH��hܪǮ� |���re�	��e�֍>d�(��b�I̓:l�yB������DK�,@%@��p<�0�,�@�� ĲP� �DФ= �螉P{4mYaΓ4cjr�O$M��2LO(lu]�
�b�s��]��1q����
Nt��!g��#Π�Q�Fl��+�V���K�}*T}��f�A�"E)&�^m�<��U(3޴��g��JۚQ��e�
�X�6�][�f����	�;ض��S,;ΔΧ�ē"�$�c���jGR���� nx���,'$�a��)8�1�*�(0�L�ʤ ã[�a�։:G'�@����2�'�^��$��N�1��a�?��`�f֝�axb�YL��3�S0�]"MD� hd�� �"�b<yBՀfp捁e�Vf�$����z�e0.��d�E������AF����3_�&����sL�m �
�L2���.�L��hw��@RTSlM�yRo\�wG��p���
���x��Q?eu�tzs��*w8|L���'��Q����j�D^�����/�7'�b!hF!E�C�!�DN�_l�ؕgV!J����P�g�,��֨��c�ę�{B`�"�p<�`I��,p��eg�6c��s�hG�d����{K�'��;8y� J�%&��%�ĊG�w!�@qQ*�e��Y`�
O|̑�̒�-ц�yD&�B��ժt��{��\
nЩQጯy�X�-�Oq��=
vIɋ>��ܚ$/0�l؅"O~�^�����UKƇ*,�w�/H��� �5d}��JO�;�q�>O��h�6t~r��$#���w"O�qpQlV6j	�F�׌�6�x��
'WEfd�T���/�x�Z�b��u#�8>������ F舅�	<_��a�em M����[�h�@x��MT$� b���!� B�I>q03P�V�$�L<�V$%B��b�<�R,7��+�C�Q>��n@8Qמ���w�v`��6D�8����wOxTP�f�"Z�d�U���:پay�W%��$�>�=�r��G�S�5 �G��;������!��ܢ
%T	B�]=�P��H:b_�,��J�(�b��R! ��I�+^պ g����A��ۆ%Y����=&.q9��/��e[P%Ӫ霨b�Ш~üH�e�a:��9�D� a�AzÓ�j8z��$��$ۗO�)-����'��lK�'����	wjF-��� �S�Ӯ����*bJQ��kg�1W �)}�E��������v�.�a�hC#,�
����?�Yb����4`��RM����T�Q��>Q#�^�[I��`i
#l��3ũ�J<Q'��uѷI={3Z�kQꑫB�$ŀ�OB��б3���V-�hp@C,h|��g�\}R⁋$�y�<�Q�|��/ļ	��M��	�R����`=��L�c��P�p�x�(Oy�i@'�D���ף<{����G���"���/�8��� ;��R��>?Yq#n�v���NݝD��a�ǟ�ק��S&F^�p�ũE��ՒCÔB5P1��c���kP��/a8v��R�ߩ-�x�3�X�Fu���kWȟ�ԧħj����F�ݼ������D�Q 
u����O<�󤍡W�bE6���g,��ŕ�M:��'���b@@6v6芧�ŒQ����D�mp��ڄB��"����Ѧ$џ��Vb*}V�=G �v�ҲI<�� ��*�2�J��� ���  ���'3�O�i�m[�F��y����kEְ���'٦�i�왼7�*ٸRl;K|�hӔeJx��|z����V�F�ڔ�[���T��{����uMQ���$�R�488h���N7P����j�	J��3��~�4G�#\n�v=��0�ޅ0�����E�0*�ڑ��@'S3¥E��+M8�� q0jD"9`����Z�F���,*?���ϕF��bs�I4d�F�J �L�'e>AyTC��x��i�!E3�5W�B�KX��>�Xw��d)N0lIC��v���T�c���S���e������28Da���E��,SrGڟ;9a|��	%)@ J��cj%�G/r)���`c0�2�Fo��� ��*a�Pc��S�W����FmQ )�p� 2 ��D����D8X �,�%]�t0��;H'����E�'�z5AA�I's�N��pJ���1O����p�h���Ѓ۾B<�����?����i�k�ylt�4�F�O�zq�#�Ɨ4�H� Hą�8��#Jx\	��"K
D]zթ٠��=�$�ַtH�$���_9t�J��P/*H�T���H ��@�C6�I"{��I��d����L^X,�%�����1k&琦Si�y0��s�2�&zHxn������=+� �r�ii��(�n�4 �3��)? I���ʨ2n&M�d�>y�����O��jcf�H0��[w��}��S�z6-�+^tl���'5+/�/Vd�	�o��  ¤� t���Q�(���S6�'��I��?��l���
"=���f�!��ð=J&�D�	�W�$��ԇ�6jH��2�Dü��H�wBY"�?qe��)\�e� ��=���⌄W��S�o�#?.0Q2���_(4�9��2!pF�g
sY���JS�� Q�g���O!���Ϛ{�
�A�AG�V��E�& ?"�mZ!r` �JS��,�% �OĿuwb���0-��b!] D�T�JU�ݧ~c���TI�8E&Dy�`��E�]���>O���6�H��!�V�{��Y����chA!��,^��^��X���kxaa���.Z�z�o?/:pr�hhd��ؑՀyz���W*ި&�
���F���=)���)fp�Ԃ=D�h;���X�R�j
�`i�����W�l@�5 ���M�$ܜ��a�r��/H9�2U$6pA���!�4)/�@D�[9	Z��DŁ�^0�͓�ት}�J����v$�����!w�p�i>�!1��;z��t9"��~��}3���<Vș�c^�g�h �3�O��������>�U��D���ς�
I�L0T�Zi�����䠓�V�����'��X2U)Y�I*Y)�>o��0�H.�H�S��	*p!M<'�P��p=� 4UX��.r�h}ɐ �MK�5"eNC�u���b�8O �0\�|賃�|�4�Hn$t�	�-`&�l*p�T�b��]w!�G�5��gLj
�d���7��q̨��U������G�p��D���åZ�¥k�LH�`�������'lH��;_�	��E$}��h�z�b_#�`hsG�  ��HV����
�`m#n��}?y�jO2c`iwO7�t��*Aʽp^�1Gx��P.���'�x��T&�-Y(���̫@��$�y�����	�A�����6C�<�@�� �R��I�y0�B,�+ގ}Ȅ�M�5*�,�F3H���ȧH �iլM�RL���?��fs�����7#�l��B���V�}AAs4�2��^OI+��0�O�q���
�`��mA!a�L~aj��4�	���b�UV���ڀFʬ��C�D'8�xS�]�R��T���; ���Q�NM�rayb��7��󧮍�Je*��W�G��7*U�'���F������2�ϐ[��՛s�S
N�:(m�Z�
�tgD��NqIǅH7E�J��$i@����E�Se|("&#��h��O��R@DV>%Q ��(0T����m̓>]R�p&��q���b��mA�`��4����6⎥�L�@�!�#,����g�'C@�q�@�(�����A/��4z6� XŋVM=E��R�����h�h�!�"�)gNV6A{j��	�	XԬ��"J�fdd0�ǈU�a{R�ܧC����JA�U��q�E��I�\���ዉOǤ�2"E��^�t����p@��`�xB��93���6�G��i��I%3���9�e-x\��D�,]3��0�ʊ  ��(K(p�R�0됿I,�	@�:9��ɮG�6M��*%@*d����i/a�xIX��Bx�������'���
�1FJ��R����(U��{��@�J�, �G�)��*�M��MKQ���E`��0�[�:���KYa�'�Č9��lN��[dō= �x<(5Fܸc��8��l̟���d�ף�0<��F@�@�%�F��[��ũ*�`C�I*]`�Rq�B>��	ӆd$QS��&<O�тl����p�o�&'��h��K�r�>��D�$RF�����I���i�)?Q�n%���ȘCd��P����3V�v@S�FC>"��H$k�q�B�&�ĂN��jEq��eg�Dx��ܠU>L:6��pԈ�8��D�%��P*D�Ţe�����V��R���\-X��
���c	Ǔ-N�m�g���d���T�>z�����&:&��H�޿�����@z�̐��372�໰I�*m/��"Qo�,9K!��@<�`P&+�$�#R��{����D�bU��à� �q��,Xq�@Lp� *��%,O�)
�Α�L`�\CP$O+c�X:�)W��`͘U�´}�&;�jK��#1��ȑ����f�4e����	�4�X#� ^�+.v<Q����m)6O\�z�DA%c[Rm��N�#+D��q�Ăy�4���@Z�G�$�R"��,n,钫OB< p(ѶR�l���@:1�2\(��H�wD�������"���"ӥr��5xC�	M����茔b}��$:��ʤKt�m#d��.�� �
�'	�!ӊ��I HиBŶjdq�BH3��N�h@ �1	 ��u��-���'��M�U$�xv�u�b�zt����[p�m�T�8Qt�勇o��):>@Q�l4w��i��`�Ns0��4EL�@qC�<����0���p<A�G�~�(�0�ȣ��Cr�P~�ɃLa�Av�@d��@��F��O#�� 0���b7,`����x7�5��� ��dus�#���j��	alϧߛ�f��8�Kݟz����0��6��)���Rq����*?2 ��sE�N�-��"O�p��/�j0��l@�i5:�3v#�N7�(��'��M�������A-FՖ�J<��g  6��h��'�B2��k�<� 4��y�F�T����r�<q4� ��lG��<_�$4��	Kh�<��0�H,+�̃�W��1��}�<���
;Tw�Ʌ��	�nL�d*Au�<A�䃍jG��ʤ��<�pPCP�G�<�C\4&G0x
���n*~����O�<i\�TAd�;����-�f4d��ȓe�V����e~R1�X�P\ZX�ȓ���j�,ۼPDҔz�J�iH�9�ȓ(0���@�pM��%��@ �"O��c��s}8��'2w�����"OD4	��-��)A�[�k��+�"O�%�eֲrhR)�p ��3�r�QD"O�!J�at8�h��	.���6"O�Upa���z���t�����"Ol�pMS	vt��7* @��A"O�q`KQ�p}I�iY�F�HdG"O"�8vI�K��L2F��%4�5x"O� 0�;��ϻz��2B荴S�`'"O�Hr@��:M�h��5h��8��"O���`$ԩXܶ���eB.q���a�"O>x'���\!�j4lǠ�3"O��/]��$൦�9���Q`�!���O�Q���݃ZWTh�i��Od!��K�Z;¹���V*��R���!��0Ymh�'�	YI�o�f4!��
`���q���X�� �$�S�.�!�䒩W��ƌ�`yzC.�#u!�䋥\���7@��n	��JK�M�!�d��fk\U�s��60�Ӫ��F�!�dV1w�.9zw'���z��ժ �!��$�v����U�,dP�n{!�$�q��8�䨝�`L1����5nT!򄐴5Tl+d��b��F�^5�!�R���!*qj ����5�H�l�!�γj�̡FA  �QCQ��f!��ɮ��$+M��ll�`!�?I!�I�,Dص�C-C�"������Nh!�$�7h�XHBWN�`��v+�4v�!��A
��eǅԈ��!��)L��!���kd,��E�̰�.S31�!�Z&j����`o�E(��XՂ^%�!�d��H+���J�J��ǃ��}�!�D��1H���C�F���	'��?!���n�"t`�8
�L]�6!��=!���(uW*p�k��\��i�.u�!�ۙh��=�ǉOg���"Q�!��
�W{�]��Қp���L�E!�dϑr0�)�*	�*��󰠇).!�D�d����>-���q�ι%�!�8$�x�9a�̤S��yf��<N�!�$�
,���'Ҩ �eǻa�!�$ޅC��Ղ�28���B�cի{�!�D��6
�Дm�!��p̍�t�!�I�\l(�R�j��G��xh��DA!�dU�u�̒��:�v	�ꊤ%>!�� |[����`�o�����N��!��S	J���6L�*�ʹ�A�(!�!���-�8y�3��	3�P	Xplդe�!��[t|y�RNK)a���8�5L�!�D�>d*��sz��1 �_�!��"HD�pNN�BB��ѯ?r�	D{���'��	�ƙ�^%�]kăO�.a����' �P(�R0_-,�b�LK�$�,��'�Й��kC��P9I5�� ��'�HZBGϣrU�+V�@8����O�����#���2i�wN$ �)��+�!�� P9vD��H�.Ve���#Gܒ*�!�ӷ%⢠��.��~xd][���\!�d��RÁ\.~T��ƅ�J���	�'����4�ŧ��=��%�Bd�R	�'k,���/� C��5%î���'���d��7[Yb�s!�ʿ>:��'j���R�#?~I�OKzI��'���#��/�����n�~R�'lf�I��J�ճ*�z��R	�'��aC�h�65��)ڲn��ne\	 
�'��Y��f����A��x���B�'n�8�5횵#�|)�Ad�ub�!�'DT驣aX6U����`o@�j�����'f:�	U(��E���}N���'Qv�1^?v��ٹюX	�J�C��� \b��q���[c�/7XY�A"O�����0�N-ÀBX=�1c"O���j�'Ec��AA����*�"O��� ��\�P�
�oξ��Irb"OB�����6�̝����+j���"O�hh�؀KF�tO�U�>�[`"O|�B&���v�	��,�9 �8	 "O`Y������C+]�W��
�'R��	�/j6()a�N��, E1�'�
�ӄx%�FΑ���"P)3D��
�W#����W�ڕr)!vJ4�O��'��ihd��z�z�6��N�$�Z�'�LR��Y4#$LT	sd�:L��9��'AF��G�Ѯ|
q�)L�#�'��dr�-R�hԀ�� �0�jE��'�ў"~2�È	&1<8�����F��f\P�<	ĐN�HJ�#F��`B�N^K�<���#�X��K#hX1��!~�<��Ah�`�c�b�)y�N����|�<�a�73d��z�g方
��y�<qDb�8'%B���@ ��ew%�t�<92�	�AT��S��%B���V�k�<��ȓg�0���j��u� ���h�<I���3d�>�q��2r�m���\d�I]8�$��#�"U��)c���4 V����%D���)I�o��]
Z�0M�u)��/D�[ri�'�<�33@غ+�H)�A9D�<�pe�-U���
��>��0iB�8D�`�tU�H�c�"����j7D��
��O6u]H������4-�'D�t��Ml�s�@�V7����E'D��R�	�"z�A:@)��Q���W�#D�ĺ��κX�h�#b�ϡ<��+Վ?D����Ή�	p�@�ώ5sr$��&0�N����C�W-`�@�E͢LD�.D��J@�6&���F��"�)[��.D�� � ��[�^�ō��`��a�+D���1B+]%H�Q�K�(]�q���)D���L��e��+ѐ}j��`�)D�d80+V�X$ҙ�b'_��
�&D�h�'g��v_�19�
]5����`/D�D����@�,���b��M\b h�o,D���n�3�J;�#��40ʷ@-D���.�1J ����W�FH���`5D�$�F.M�D6����Y�	�*���&5D���f�((��QlJ:S�B��d/D��9Į-K�r[�F�r��ç-D���o��hr�\��H:.����f6D�h�&!�A�L��iK�f��preo9D�ț�hSF��0`��4�P "�N2D���D�I�1��U�����b8���;D�p�U�΢ ��u�7�M�&x+�c9D���R�^�z�V0�e"�`@�@�7D�P�7O��J,���X�g����6D�9P���Iθ�W-�/,�1�F�5D�Pi)��0J�2�wAlQ���/D��g�4���R�I6RxJuʅ�"D�4�LJ�T��Sm�X�M�B�5w HE�ᓲ-�Ve	��W 7#f�9�Μ�%/|C��<ʖ�`�6_�6�+!���W)P�=��D�d髱nA?��
G�K_ȓ#���d^3c���I
�;��a�'�a�@D75�2�C਋�>`>H���{�<!щ�.d�C	ɶK��u��-w�<� .�u�$Li܀ 擨B�ȹ3�"OP����'i�p�h�d��)��#"O|Qb�.� ̮}�Ed�H�;!"O��z��P�\�����ox��S"Oe²b�C]�����K���]�C"O�ܚb�ۄ;a�!S�; oȁ"O.�	u�[7o���3(��[H�}Xc"Ov�ᩎ9ZH}{����P�"O$zKזO��k��,6����"O�q#ϻ��1� l1�-��"O\�JF@ZW	 �p�O	&
8�"OԌ�v��6)�*$sW�G�]�~8A5"O�43�V������M[,�tG"O��kDd��!0c�%F�d�@"O�z3g��V���`�$�. �"O`,q��_=SejhH�e�.Z�� �%"O8i����fȕr�/[K�tM�w"O�hGC�Z8��N�!�&U{�"O�9���Tc�D�#݌U�P|3""O���R,Й[��dZ���F3�'P��``��)1�J��w�D0F��P{�'��AZF 	�gL���8���A��~Rim�);����f,j���
ɱ�y�G�0L���S%�"c.by��ƈ�yr��r��"�0	ސ�!G�� �y����W�B\ZK]z��E�q��y��ǣY���q��լy�|Гҥ��yB��f��@J#�~!�R͙'���p>�5��38iQ0E�e���xu'�e�<��F�'���ݸz��I�V�y�<i��K��-�)Y=�^ybA��w�<)XM0�1id�An�����A�A�!���(y3��k�� �v� u�:�!��F10SN�V�SӪ�0k��\G!�$�)��(K"1�����	
pN!�$���@�&�Z @�mX�IԆCL!����I��:���b7-!��W =� �C�fPY֮�!�L�2�yc�ń�j�~���ڼ
!��.l|����-}�˖�S�&�!��*|��RA�J��j��V&a8!�䖧Y���uG֕T�ְ�C�׌I�!��>T�B)�CC]/,�|���\�!��rY���OXZi��QB���!�dɊ+!�H����Ov�D"	�k�!�D�2�������o �� Ц<!�D]5,�)�K�6	�ts���H#!�ߐQ���C���Mr�m�.k�!�� �n�f����	R��d
�O��&�!��G@��HA�Y�0yp�o�F!�*'�n�����5y������	!�F�Rs��Q%�@�5��� @l�&�!�ğ;61�3�	�����a���g�!�F�2qc� ��B�Yi��<�5"O�����P}x��,�pdB�ZT"O���c[��I	Z�}]t�1"O>��ra�|����hD�jN<1  "Ovl�#f
+x�@�9�m	�480#G"O���&L��B�:��.�p"�h[�"O�8"��N˾\��R6�X�r"Od�넩$d���pn�K�+�"O*X8fJ�(9c� ��V�[]�8�b"O:�cS�&6MTٹ7� WN�\��"Oޙrg��	Zr��ڑ�'D��sd"O� &1����2�y��� ?h��"O�� u��3�Nx��-T�t�1"O�A���9{s���nݖ)���"O\a�j��>�H��W���r�,D��(��L�d�#Fk��[�����+D�|���rP�H[����TJ*D�l�1b�P��Ԣ��ٵp�Z5Y��<D�� &#�ot����'q5\���/D�� BH��j���_	��9D�h��)ҷ~�Z &nV�|X��2D�4�ad��&��Tp��TaBU�	/D��W�׍, �I�1�\+M3`q�5@,D�"�� G#��I%�,n�8�9��&D��r�ڕiB`9�b�8n��X�2D� ����AW��d�<Avyb�f5D��2���(i*�XR晶hTip�N5D��`ědh�q3��m�L]5�8D�h���1]��U��,=FHe�7D�T�`LV�4�穕)�*���h7D�<�F�	��֕��%�/;�I��c!D�SA�2�
P0lҷ2Kh��O D��Q�	�X���@�Ϫ\R�)�� D�3s��K~��	���4=s�4D�`Z�m�}a��xQ̋�N0qR6�1D�HJ��.i!P ��ɣF� ��TG#D�,u��2L֍H�d��2����vL D��1���0��!��ɇ �@)yE?D�P�%AE�L��Qp1�ƁQ{���=D����o¹Ԩ$C�~(f`�0L:D������u�	b��ǁ>b���6D���mH>8�6���(�p�,��F/5D�P�%n�8N� �ɦ���U��Y��/D�lSs��y^D
`I�!cD�%;U�0D��y1���w��i0eA�U��E�;D�@�a���]��O h
��I8D��3���U'^yy�)CJ���3��2D���WD�~��(Ӓ�����G�5D����Z�
��HB‮	�ȥ	b1D�i�LK
V��D��3F�a��	0D����KS����k�J��*���
:D�0�m��^�j�#��B"ȁjf�8D�Dc�晑$�������_U���e5D�\iw+�/d�.��a���<�jMQ �=D�@�D � L�Ĕ��
�j���2:D�0±�B���s��U �z�a8D�q�Ȉ/B(��D;�L�a��;D�|�a�`ѐ �sF"O���Q�8D�$q�N�� �4�ӗ͒C���S�g2D�,9'��2:�|�Ȣ�P/4�*-[a�.D�h��P�R�<LW!P8I�*��l'D��#VEA;RD�)�"�=<2,h��*D��x1��x����T�ʅ�ҩ�.D�(a@�D'X�Ă�H4}��p�a�+D�d36M݁-��d���� Q�`Q <D��aE�1xp�����:�����8D��s'�˼O��������5� C%k6D���*�6>�P=t�ݢW�H`c��2D��� .��HzAD�Z�b�bࢗE1D�<PeF�;h<q����MAB�3UO)D�0�0�����d8�	)m,��t�<D�Љ�'M�עQcelɢ&v.��,D�pg� �:���,S(}l�Sq�*D��(a����@9�`��-����/>D��3 �L�}̨�r�G�M*�isAl D�� �y[Ggݶ���ŸP�ܵ��"O��}@|�C��z�<�ф"OhHXѮ�Z����(@Da'"O���S�M�&AZ�mL/A8<��7"O�=01"ii4���Y�;�:)3"ONb���B?PК���N��	81"ON�R�0|6>���=O�@EJ"O�M�3n�+���:#�ĵO����"O��Y%��e� �p��9I���6"O|lZ�̌=xj�2g�S��+�"OvH#�*Ҝ7��S�� ��eS"O�u�'�[�X�XH f�^�:Ӡ"O���v� ,��q�g*Χ%p���"O�b1J�'Oڌ`"7)λ��LR%"OZ�Å��b�=H�(H�0x�,@�"Ox�C��b,"�"�å8g����"O8��E�ݧ9ڀ�vN�'X�\��"O2p���Ύu�D���%�t�"O��{��pą挓 N|�lІ"O>$��)�"4�f�0�%�?i]�(2b"OlKR��$2?�0u�S]����"On�������l�֯E�NSh�q�"O�Tɇg�I�	�鈐r��p��"OJ�x� �(MV����C&�v<QD"O�A�����o΄0��%I)xs��*�"O6��@��&���$D�XC���R"OntX4��?fX�i�Ā.:0�kR"O�dR�oT+�T�I�ŗdz.��"O���å0�� �rbYcg:��"O�ـ��4oF~̫p�D�\Y��"O��B��W���C�ڭM��3"OD��#�Ɯ	�~��$�ʏ_\Ȳ%"O�! ���x�t@�B;sZ��4"O:1�Q>�^���J�Da����"O�k�gز6���rj��_l4b"O�Lڄ��D����F5oZ��C"O�I2�Nɺ�qbf�$Z� �"O��	�oZ�a�|ɣ��H3e�fly�"O�� ��?���(0$@���8�e"OV��D�P|<ra{&�E$Z�R�1"O^��.�;�p�ibN�.{���"OVaRP�#JJH�K��¼?�l4��"O��S�w�Dh��J\Xc��&"O�d�V�'M�T���`'b䩰"O~�*��;c߆���ݑ���۰"O��D��+%�Y�X�K\O!��?#�v�ЦB� [�x���j	>.?!�7O��!,�i������^�R!�DՖ
�^���M�M~捠CW,`4!�DL1�t}��ME&0k�I⡎�n�!�Č*t<X9�4��((~Ģ�&�i�!��4dz���E�WТI�0E�?�!�D��/D$��D�4��4��O�p�!��#8������ϥ?Pl��	@�6�!�d��m�l�,Yg���@�l��'ܞ�h�#En����7��96O��Q�'�����r���6 \�3G����'ۘ�)e�ә"e���VmA.n�9�'����(�a�,W�z%Rp
�'X\@�4'��LbЭ;CbҰ{2��	�'��U��ʊb�QZB.�!|�^�Q	�'l���f�!LL�:�I>x1L�s�'��qph�~�T
��ܸr�41	�'�:`bEG�H�@衏K�w��0��� b�a��$�\�X!CQ�y�t(�e"O6��js��Re��:[Q�M;E�(D�Höi�/�� ����:L?8�Y)D�ĳs�</5�8��T"Ja�ǉ#D�䠑O�
&jN���H'C���G'D�8y��ɌUPĕ���K |l����7D��:���6U>��!��]��bp�w�4D��80��)S���j$�
e�2D�\ұ��"�n<�gΗ e��T�.D��c�d�3� ��p쁴x����t�&D��K��̢���:�/�4/� �2�2D�W���a1�Kީ���0�C4D�({7B;����W�xo��V�0D�4���>#�45�w�;�J�"�`0D�T�Dس0m�Q��ݭ�Lx�� /��F���Ӷ%h|���ON���#C^�B�ɀ�ذqQ"y��	T��&�C䉿A��Ѕ�J^D�k�B��*�}r7��(�X@��o�
VI4B�I~Be�ׯ�=/��
ӉJ,aB�Ud����V+|\i��ʖ3�B䉰qX��4������'k��=�	çE^^9�0��}QF�5DW�^	��:!�Eya���Q�P�b��݃I����WH������6.�ޑZ5*��X��-��hfT�hA7���"��E�ȓV�,� *��2%�J$�9>ײ���Ш�&��0)�~�h�I4<�B�ȓH�b���I@�b�yP�Bα�ȭ��t����V���$��B?�5s�@q�>D��9�ޥՠ� �ܰ ��$��;D�XS���4�*|HԮB��$I��9D���`�5KDu�BND��H\��6D��y7.��6���� ĶLpY!3D��@�уh_�0G�.5��2�g2D�H"�O��,����ɻ4#/�Iuy���O
�B腉i���R��^3@I�!�,D��AT9��6� [J���$�<����/��4��V=w��+�ѡ5����hOQ>ik6��N���8�>rw}��	*D��pp����� (� ˻L���D(D��	��L�#fp����å=��0R0i$D���`��3LZ�y���x���ů"����p�
����\@�_~y�@�,"D��)�A�Hw�\ʦDދE�45��Ojʓ��"��?���mŠp[�G9&N�q+s'@-`C�Ɋ3�l8{T��s�܈	�3n*LC�	�"t�՘3�@����+!i��$�$C�	���t�Ϊ&�h0�6� �_>C�	9x�$e�!�܉[�va#L���B�	!K���ȓK$N�I��ֳs���p��	.E�D�
g	$��9��NM7_t�?�+Ozc>m�B��N�Ĺ��aZ20\�-�#�%D�����x1\��`��sa�M�4�!D����ߍa`N��f
J�,D��c��ݟO��e:3��%�:x���*D�l	�؛X	�-��B�n;`���(D�P�냑1�~T�aiƑ?8���)"D��(����3�T�ñ�:��]z�"#D�C�&�k&b$"�_8Vql�%�<!(O
�OQ>u�ecZ*Z6AX 'B|t` �A =D�0��L�$uE����C@�*epE*��<D��R�DWi���yFf�6V�۔�%D������	zF9����:j�$u��D%D�� �e�����i!t�Z�@��m"Ork�*U�R�r=��_�h��$"O ���(k�^�z�^�U��p��Q�H�	���&��Z̓��hѭT%�P3`� ~��X��#&L�t�O�B��E��i��~4~��ȓnv��Ap�̶4{B��'eJS�Ԅȓp�`4�F۴bCJ��g���t�ȓc���cd �;��2�EJ3
ވ�ȓF�½�g�غCS��#�T,:��ȓRP�\��.�h�qh@#	�
hNL��Ie�i����
�Aª�r��ݣH����ȓ}?]����wϒ0���g�܇�f�ĩ�ԤC������ &.��-@)�s��\ZX@��B�pBĄ�H�.d�U/��._P����X!���ȓ�l�"Ue�L:��3�eGu�ֱ�ȓ'J���#)tָIǄ�q_h���K�'6t���!_�Nz�͋2�8,�|��'�yQ!jڔo��q�a�������'�����:kT��Ю׿�
�'*�Ř��\8l�2��`"��L}��'��0h��̆]B����
;q�x��	�'<,`���$LH��-[�R��Dj	�'�*pI�Ε�o�(x�#ጥ*����'�*���`�%L��]�@bE(�\��'�ZQ�ԥ�$k�f��-����'�l�Si���|B�&� 4�`���'����C��+�*E��c�$'��s����s*ؔzd���(�C��<�!�pt�#�T����1Ì�@�!��a؆$#P�_�*m�L�!�$ e�^H�WϞ��V�f�H�;�!�$���A�����@���8�!�$K�c�$��&�<�>�s�Z�!򤍨%���
^�bDi����!�$#$)���O�=�	�ǀ��^��Ie��dpJ�5MLؒ��ҺvO�ېB?��8�O�!�퉲yr,yX�dQ+60 S"OX�@C��4b�T��B~h�`��"O,m���K.�
e{o�?�:��"OV�aj�z��;�+ҞbvQ�5"O��p`�	2	 tҳ*E�t����"OѡրG/�ȻJ�X�9#"OBh:��
�R�&'�-,� Ӥ"O��Ձ̊A�,V7�l�$��J�<�BT6FZj�W�a�>)�i�I�<1�bֺDU4��pGH�R���2PI�O�<I��kx�����a *l���M�<�1 D��|����+��4Js�K�<�p'�>򤉐U:,����E�<Yǔd�"���2���qSJ5T���׫��S���K4�>o����9D�$34��%l�pC���I.���7D��P G
'���b�\;PQ��j��?D�p3flׯ��-XvM��^jXI*V�=D�� �K�Y=��` Ń r�s�-D�XQ�j�;U&hxe�w4$ �1�)D��
5bP�(�J��"��%UE&D�x�-�Ј�;T��/6��Bi8D��C硉t�tĹ I���Գ�1D�D�`�L�C��ȑ�[�"F~(���/D��ɧ�+��Ӄ,M�{�B�C.-D���3��%3n������?~P,Y��&D�`!���#�"٣B��E���Db(D�� ���3/ E�L�a��,ڒ��c�Iv�O�^I9��@�'�F�`�7V�@�	�'-�:0KM�ojlyA�	�""y8*Oh���BS�H�8V����f��P
��`5!�$
d>P��О�*�@iR�w!�D��.��]6��drTȇ�:!�D�J�EK�l>bς�`�@�^�}қ�B$ĄtO�Y��!�zg�$�P�"D�x�fO2rD�DJ)�c���G?D�<B���S
n��Q&T�HQ^�{��!D����nF�R�q��u�hȵ` D��;��i�6*1C�1ugFYӴ�>D����_���%r�a/k�Rf�>D�PQ�ρ+W�ސЕOT5~�
�G�7D�4(�	@�JL�j �F�� h�a+D�|pdЁfP2x���N��Π#D,?��?A��i��q�htפ�)X�.\q��B!�DI�}�3��0�F�ʵ �H�!�N"ƺ�u���?��]EAPP!�D
 .B��t(R�Z� ����O�89�y��'�r�����d�I'r	��N����K)D�`A�����`�0"ߜ6D����N2D����K����`�ޛGJ�K�/����09��Tx��Iƭ��i����E"O��BD�/A��a�צ�Hy�F"O2� ��ށFO�ใ �4�����"OFUa��W(%ҙ�T@�0^��"OV9��̟?6q��Z� �����0"O�p���K�_�*����.5�ԄC�"O�1H�Q�h�ܙ���~T�J��D/�S�	�o"��i�k���1ʴ^�!�dU�!�H�W�qd*��7Ȇ��!�D h��V�� <%\T�p%ܘl�!�	��|qW�
 BP���P$!�$�@�:(Z ��0i-��BD�!�9paIh`&Ͱ<��%2��V�!���%Wmn,��C�5.N0�3��]��O ����b̔���
2Qx@�D��
I�!�֮J[�i�#/�,3�	n	k�!�d#R���
��,�kF,�'e!�$Q�Bu�ѹ G֙�"h�R��B^!�̮`�xy�2�� �4� �ȃ�=��y��ɍ	U�M�g�>0�0�y��&tĲC��	3H-��EVTҴ�H1 	4*��C�	�A��uŨ�4=�9PƂ?|�0C䉕-*&�*al��)ۈ!3Eߵ?��B��>k,��K^n�-�'��q��B�	,m���A Mz��(�*�����hOQ>AI���1w�FX�O��q�#D��zF��7�
Y�4J�?��0#�>D����ؐFy���1�C= �8s >�O��$x��Ktg��eU�%�f\qݸ�G��OdC���H������܊MPd��i=�C�I
td���Ќ]����ǉ�uPC�IS�� B "���,բa��(HC�I)\b�x����}���cI�A��B�	�0}��p��t�
1�a��7bC�	��,�r���F�C�%V�*�ВO�˓�0|�NK�n�P@���"\����`�A�<��P�����ѣ:�vȱ���G�<����<w 	�т -���A�D�<�G��Y�T�)B�L$J�9���C�<�`�8Q�.AȦХ\�h��i�~�<Հ�`� 9�T%$ko 9֭�E�<� ^Ɣ�vt���j�q@��|B�'e�O�I1?���m)i&��#Bp`����R�<!g�_?-T�mٔɅ D�>-c�JQf�<Q5	��VR�r�(�)�m�<�)N��A0��L�>�j�+�D�<iwD�
+�� 05�V�k�ĺďw�<�@I�4����!ƛ�|I"�N�v�<�g�K������"��$j�L�!�$T�j�D1i�Q�ve���@)5I�OVC�ɥ1�QX0�������F�J^HC�	�r��Pr$��>Z�%���o��C��6��� 
��@9�Ǧ5n#�C�ɜ1�.�*�a
�5���)Y���O8��O���I��9R�ș�S�l���̻+{!�ǯ0=nLps�YYN~Q33.z!��Iؼqr4̟V�R���Au!�Ъ(���@������Dޱ"l!����I �M�qN�8Am�#'N!��� 8#�쌳P�4�Ѿj.!�2L�$�a'��%��9-�0��'��%a`�ڄĀ�/K�5H�|�'!B��0�(�� ��01ۆ���?q����CUF*)0�m,,��9
��y��C�M:���K!��1��Ʉ�KtC䉦g#�����$vj�AGO��_BpC䉎pT���jU�u��QC֫�'AE��9�h���bv�0T��J�ǟ+GRz���5Ph�eO�"~���M�����b8B��ƋWp�9F/;:^Ԭ�ȓ\>`T�b�ƇY��Y��> ���ȓ6�4)�V��#�0��C<RXĄ��D�<��]����(,Ĵ
ܤ�ȓzW��ȑ�K���e�g�H0w�(�ȓa%�iQ6���pZ����a8u�N��?�ӓ]�|�
Rm��a�R.�%B�dɄ��*u&�Ɩ1��1 ��X�*v�@D��B�%�G�^�L.<�S���2a<FC�	�;�l�	�+7y���UA�s�\C�I/n��ع�fAu�����ML4@TpB�	��P9i��Q�
ff(�s'L�E�C��D�b$�B�;�x�S`ͦbH�C�	>tvJe(Vj��4�V.�LC�I(	2���ڐ����D 5<�C�I9.Gd��ᨑ6x��0k�$��j2�C�	Uj4��1��$Bf�{�(��	F`C�IR&x)�/�0OA:X ��r#^C�	�3�YJ��K#D;C2.&3(C�m|��� 'ѫ	6 q��!^C�	8���$O�0P{��_�Gz:B�![�|A!wI��iO�̠���5zH��D1�tm�u����)H��F���"�x���\��p0��?4xHitDM�K殴��jK�I#��^.V�ti�DI��r�L��^�V	��cW2Ѡ�@�W%;� ���W�'Ph����*->0&o�7=}�!��'%���r�C6@�%N
&*�,���'R ����۠|�x!����#*�q��'�*d� EŇC-�\B��)�jt��'G��Jg�ԆI�2�AL�oX٘	�'Ypr����I�65��֑\h�3�'��ų���_^��BA(V��r�#�'������! �@�b=eб�'\��PƉ�.{��
��*\IRٺ�'�(g������ &����Q	��� �\���.*�. P��6e~8M��"ONy!Ц�).X�x��dd��&"Or��ɔ?p|�r��R$(q��"O���"M�
.F���T`2"O$a2w��ksHm8�Ϥ{x�X �d#�S�i*'�����*ǭ}� ��cZ W3!� �T��ɛRov1���_!�dӲYz�X{��ĒrtUs�f�F!�D_�0�� �s��/]5|�Pw��V�!�F "feK����1 v�%7�!��K+^@q�t@��G� �KB�P[�b�)��X1��,��p�h��$7i�L=J�'/�lH��pV�`��
��d���
�'�fI�d��i�`��Ҫ3F_�YI	�'��0�Aǀ>�ܕ��֔.<Q�'(�Y��ը�9��-z�4b�'��i�=�(}f��P���q�'ƞhx1A����R$ H:E��5H���?ɍ����#~�.�i|�Q�2I��ʓ�hOQ>��I�"���!W�^�́�� 'D�ı�M�C�4s��אL�t��%D���sF��v�����%�H8;Q�#D��CbA@�z]��ٱ�P�=�J\a��?D��i&��# M�7�Έ@�H�@>D�DG��:3B3�%�(� �t=D� Y�˙1����\G���9���O���+�)�'g�@�aA�;4ܒ�� &Ahq��'�6U��*�m�@T�@!��	�h�J
�'�vb!a_IL� Gޛ8��� 
�'� B-\�Y�����dN5&0V$k	�'����#��Y�6|9��_tV�K
�'� �
�Ę9R�`����m�x��)Oh��Ȭo���bI=3y�q��ܶ5��'���'4�)�72�I��j?Cd<������DP[
�'��a��֐&ވ}(�$P!E\x�	�'�:@�ԧ8�qb�#�rO����'F�S�&��ȑ��0^��AQ�'��s�4w���7�\7&�dt �'�ZTɖ/��e�NyB�o<s�qJ>��H= ��1��
�p8���mƌ9��Oy�|��	��Rb� �F����H����+
��B�I�*ޝ���Zʰ@�R8]�B�	��F���"ėd,�MRS
˕B)�B��!��U� �ć]��9k����B��$��);��b7JV9j��C�I�]жYhI�u��aa��IZ���<�+O�'�?i/O��	D���G���Ezd���� �xC�I	k����Y�dp�'A��0C䉭o��x'M��=p�
�h� ��=	ç[v�x%�� �N���X�;���9��u1��#[�Б�QH�C�4!�ȓS6ѐ�ҥ'ڢ�YbɎL�؄ȓ\��5q�"���cO#V�d��Iy�'
x�:�FL*��@�W�H������)�Dd��3]0������>�(�����)�y�+��}����e�% ��dZ\���<1��D!�t0C!@"c�%�C�H�!�ď�|�$\���<( -� �]�s�!�ɋN(j��P�ɡN%j���υ=�!�d��,3�+�E��as��L5$R��W�'3X�x�f�1)� �����+���t"O� 3e!M�ކ�pu�� a���0"OJ�A�/�A��ሒ�5�lH�u�Iw>��%��/`s �bA]!E{`���!D�� ���GѨ(c������)��UP�"O̓���)d�:V�����`T"O�cݡ*�\�֥��0 �"O��!��;:����BӈY��R"O�l�3,��2x�iI���]���r"O�37��r��
`nT�<�4��"O��cq��!fJ��6(�`�E"ON��Ea�����E�RIju"OX��d��=`�$�U����ꑩ�"O.�1dD�MV��q6�� s�H��A"O�x�fȆ�%��<!c ��
��$"OJ�{�Q�>���N�$� �a"O���C.X
��p-P�� �Ih�O
8B��*;j<!�5n��t��9�'L�M��O�kϊI��]n�����'��͡%@�E�ة�2�ѳt���'��m�D���A��=��Q�-O�=E���.m��8�,ҥeB0:2Cј�yrH[u&
�0�#�WC`��oW�y�M�Py���$\9�@``����'?�'��h�t�B�L9�\Qf�2K"`r�+D�#���@Hb)�6	tK�����6D��Ն�2rFzP�A�Zbj`)�3D�pQe] N'$��V"څc�$�V�0ړ�0<���Z
\@�lK��9L� b�E\�<�Q�ǟf�Ԁ��:i��4GHq�<�P�ӑW�ݑU	9W?�· Om�<��P��v�+c÷+���b�N�<)��=R��,s7��.i~x��o�<�t�H:�QX��K&7��C��i�<�e�F �8L���$9Ӻ�IV��h͓�4eh�n3"�H��!�qME{��'¨Ⱥ c��PtcT�ݞ0p���'��26�f@�'�� |�$��đp�<qE$B/�|��dO��9����Qx�<�"!�T� ��ўB�@�bJ�s�<��D�dY��d�Vfz��Bc�Wl�<ѐ��#ꄑh lJ(&/�ţVM�d���̓3�x���x���U5-HZ�$� �'��>�	2L:�Q���+�"�B#�#S̸C�ɶ%���*V�#%rRA[�ς�,8�C�ɆR��8���.�B��p��`�C�ɴe% H�6�U�oU�a���S3"XC�I*w좴��jIhO��o��:��C�	�!������P�R�R%H��I�C�If8���脰3��"Ƌ����B�Ʌ&����'��p��\����R��B䉽> J%�(e��rB�:vB�ɬeܦ�g�]~����<SPB䉗A���R��jLpJ�U�j��B�	3���	B���&�بwnC䉇o�6�0$�{�����J�p��B�m;^q�+����jF�I+'l�B�	"�P���oM
���ĊE.�B�
ob^�0�����c��L�B�	>Z�e��G��0��y��#H�jB䉇q�j��ueC�9���C��CK C��	$�X�C�D�0�x�*5O�<�&C��'r����OP=a#X����EmRC�	%�|c����3h6��!�<DDC�	�U�����j*%�,Mg��'�C�ɴ�БBb�Y�&岭z���+�C��b�:lY�@(I��BH9)DC�	�f;Uha��&�\�kVM�ThC�)� ��A���g�J����Fh+�"O�p[��
elT9�(�9X�p�"OZxq��'�9@!m?D�
̃S"Ob$�U�֪���qF��V)��"O��y� X��4����~�(E"Oрq���t?�����L,9�!X�"O$��DH$�h��Aչa���Ȁ"O�d�
�F{BB�>�$�B�"OL�kcŊ�U�h�h��m��� "O&Ł�Ȝ�F�&c�a"O2e�m��q��E �E�3?n�m��"O*P-��Z�P�I]5 g�L��"O>�*@�D�x�Z�bRĈ-O��1��"OL�hX>*ΡS��ƕ{��p"O�J��
�HA��B��JS"Od|q��E�4݃�@�/G����B"OpD��E�7�ݪ��F�25��"O������Oi��&�	�H�06"O�Pkte���9��̷m��"O�����ſx	��*��H>H>1�E"OH��uN�'ZO�%��b2 �8��"O���Š�TA�BlQ�,�N�SD"O`��&#A�]�`�P��H���N&D�(9��A�~K*����+���Y�C$D��ж�	\,�u�!	�_��P�R� D�� �Hfg8��6`L2����a$D�����;���&2��#Ո<D�D��C�]��� W�ɭ&\�xb��&D�|@PI�3�с6�>5��4�(7D��6��	����F7�p�q�/D�Բ��fd�� �@�l�@��2-D�H	�3c�9[��ѯc�X� i*D�$I����B��t��h���DC䉇4b9
��@��Å�KCjB�	7C2�(pc [�d9
��Gm�B�ɬ8��DsƱt����XX�C�ɠt}A��µp���@sE�<8n��d�/u�=h�ֲ.V|�F/�31�!�$\?2L(H��Y$>!֨xd�%w�!�Dȶ�v�:4bM�Q���CfW�9�!�ưB��H��H�1|�xѲ��69!���%!ҵ����\��i�T�C�>!�d�`%xta$r,�ys���e'!�$��{R|��$yb�9�Z�j!��I1��F	nj^lЋ���!�DJ�`Zu3T A�K�b�́ 3Q!�䉒1b���ף~�J%5,�V=!�J�F���� �@���+�!��5"�:лf�@rHܰk֞�!�65jX=�Ƭ� ��0�䏢�!���"1J9���վg����Fd�&]�!�1hM��y�eQNmTl	� F�e�!�$��u�0}�V쒒/`�2v�U�!��^¹2�"O^��pe �� !�D��N�5RR��t�"�rU���!��^G�͊�eR�([ּ�� �2A�!�[;$%�Y�򠖰*d^���i�c�!�۠YcY��M 9D�;5�W�D�!�d��S�89�R��(a2%��o�!�$ŊU]�����Ŋ�L6�@�!��`Ő��C�}�B��!�O'i�!�D��
z��Q�Dѿ-/�u��L߬To!�Ą�W(04�� �s��9��+G 	a!��.�4���
[�v��ق��P!�� X��0+7de
j��B��h�"O�@EJ�dp���i={�J	j�"O��D�ߋ6���ڰi�r��$R�"Ob�+��*)��lS�fƵ)�Fp��"O�U1�gG�N�n�:�#�S�H��"O
 @eڹ>�94螼LX8��"O���ad�+4��1�� 4��@��"O6��R�K�������Xt�H�"O��P��йW��mS�͒+'r*р�"O�@Q�@S���X� �j|"O��c�)@ =���D%C N�p䉤"O9�F�7�*D�c$��~�*��f"Ov�	@�C�<�k&bS?�ؘ)"OJi6�N1�R��vA��<�~a��"O��RRL6EJȼ)��U�^���Jr"O����i k @(��ўAp�@"O�䂑�'bp�B�M
�>��r"O�Ҡ&� 	���[g�("+�YJ�"O�� Tx�l���C����"O���Z%r�ڱ��u��C"O�lJ��@wy=RףK"[Ͷ�sq"O�(�`
A�[��8 R�ŷ`��� �"O�8ҡh��ƹ�p�N�]sB��v"O����(�3z ����O�`�`�"O�5b��C�g�����'LΈ��"O��3�o���`�"�ޖ0���3"ON��B��l� `uC��Pt��"OF���vT ��ߠ&��Ha"O�*t�TBE�(��K
yV�z�"O|����|4�-i���TX�r�"O�1���^8&<�\�1QV�"O�٫E��92��i#�mL�T"O��cgԟaݚ���
#�y�A"Ohd��N�EDj�#�kK�3V$ �U"O:�����I�IC�kЬ!M�D��"O��2�X�L�\1����]� j�"O�������q�2ء���G��)2"O��0G-TTU�-�1lޏRȢD;�"O����k 4�&�	��7䵸�"O�ܨÝ;��{S 1/�(��"Oh0�g��.Y�2�B��e�6��"O�����ƽ
<��㘢{ǎ�Y"O�D�p���}�&Y��-<x��p"O�=Q �X>�$Ԑ!�W�8��Ěv"O4��$�[�NV��U%C��@"O�l�ЭJ(����ҥ�.�a�"O��a����J��6��
Q�գ�"O�!�DmZ�䮼bF�L�^���c"OӒŗ�2
(8��9��A�a"O*�"P��3520p#�6<�*)A�"O~�FIJ�!��I�]&S�,i˂"O�����˝j�D��0oڏ�Fa�v"O,( %Ň6+BРr�֝#�\a�"O [�Cڄ��|�����:�4�kR"O8�S��N�������i�>�9�"OD��%=�� �́��{"Od�a�5Lm��R��H�b��8��"O�<')L�z'�=CP��l�����"Ot�ӠiB%e�J k1�H�a�"d+0"O���nޮH�d$�#H��gt���"O4H�SBHz�勦F�k:R���"ON����B�^��p��ӼT�鈒"O�<b�H�= �����X�ylr���"O���r�]��;ѩWP/D V"O� ��:�O���H�E�6����"O ��$� �<Śc�N���, g"O-J��@�T�6a㖃޸����'`>	���$~@4���L8z��0�'A�)3�$w�IS��� #�Yc�'f����A���$	�!@D|�
�'�e��;�"L!d,�2hG64��'�(L�c��0h���s�ɸa�S�'�|@U��cl�����
'%ҍ��'�x�K��t�����Ǆ
����'SF)�5�@0-Shx�qE���Y�'�$(�G޷d��x@�@�O`���'¸	��F�2=�Y�𠍂~z� c�'�<��s�J�`YPM��A�'��HWi�%d ��W���TZ����'���0C�ʵ���q�Yxݠ
�'���1%ׁ�T̓����=3�0�
�'��(r��<����'�9�Z���'lX�"r ��_��� �>eXL�S�'ɦl)0�I�%|��cDG�X���A�'�(�ɰ�#b�-�S�V�^�
��'V�Z�?VT���CI&	�fX��'
�T�7�ȗ3�H�:�'].f����'�����e���`�J
?��5��'�ܸ�.N$y}����[���Q@�'i��B���I�s5���<ېxC
�'f�(ic�Ҷ�F�*�G�+�\i�'9j��eE-6���XV�D!ψ@�'��؉D*U?�$	f*�)ǲ��'��t�q�&b�h ��!�`���'�\�:UǛbd��30�.�[�'X�x`!G�)j�x����"�\��'��Y0И)�)"��E:���'��L���
e�,�kA��,�LM��'�����΃?��%aB+F��vTc�'������b�@l�"�E~k�|B�'�L�U��0.��9�sc[�r!f-��'T%q��ʔ��4y�`ղf��`;�'�����Y��qZF��a����'tD��7�
�oY@ᵠ�p��tb�'-,)QqI!�p�۵A�aZ<E��'Dj]q�aC/5�H��5D�3�j���'+ =���|�P4�J�x�Q�'f�Q�-��T&]�SG�z�X	��'�$��a�ؠ^7,,3�Q�#h�a�'@z��.�9�R�[cM� ��j�'G(`���� E�䅓�j�<iR=��'�6�y�,p�d���"�o�Q{�'_����&�	P0�Ř殌ir����'��U��N�t���<YYP�Y�'������վi�r�p���T�y	�'\��F�XvP�B犛�~���r	�'YQATw�&$XCH��j�8��'!z�:�ꓐ�\��H̪s�����'��s"'S�K�� B@�Wy&M��'!B�i�h�N���KALB'\*��'�27�չ�.A�rB��^i3u"OV��`A\#��ɑ0H�M�Y�G"OTD@f����"��-t�)#"O�8��+ �O��RD�.	r�X�"O�`	7��"#����g�X�~�4`s"O�Їg�,X�P��	h:|��"O�D��XΔ�x��5Ǡ�*�"O
X��#�&�n��F$���"O� 6<A!j�NH2a��V�3��� "O�Y2�o	����fشo�ЁC�"O�I2M����\��Ō�L&�� "O)�U-N��y�b ͐���"O8��4��r�̠�X�h��d�"Ob!3��k$	�F�ґz���"O@� ���.@qw��-g *�"O��+�%�8�}I��R	c��:G"OF9S�ڄ,:�9��f�u-�9��"O�����U�0<���1~�4W"O �p�lD)]�|�CEL�>0zf"O�����$��X�ˈT�Tq�c"O�9K�Ǳ4D�X���*�\l�s"O�l��6�h	�CCّQ����T"O�����Iì�Jm�
~��#R"O�p$b �^
�3��Y�_����"O���L�&�dЕߝb��M�"O���^�G:��˗GV<E�]�"O(�`�9^�T�%-@�H��#�"Otx3�%X'ϔ�h�L>Q�d`z3"O�P��

�Whp�$��$T �C"O�(wO4%�%닍$\\B�"OVRe�=w����iE���0U"O:�.J<SxI"i�h��kF"O�����3@�(�vET����"O�X��O�8��ZCc��W�.1��"O���U�?���y�/>��䫳"O|�2S�Mh�����`�Ј�s"O�E���6,x�X+�G�d�6h�"OPt�R	_M�i`�?�"�;�"O> ��F3Xʴ�ɠ�wm��p�"O��
���1�{�%ҭP�&"ONH�b��3� ��c�Ĺ~`\B"O�C�n؁y'θ¡L̤Ll|��"O���dE�J�(��C�Ғ���"O�4	&��z��X���/�:B�"Ox��/�ll+�!�-����2"Of�C�@*\���R!$i�p�"O���&D5.f
T�mW�W��["O0y�$��2�A�2��9:R���"O,��¦�sҸ��ۺ}��iRD"O�ipV���J�J��z{б��"O2(*�$��V9�!O�_�n��"O� ���6��u��Y-d��jW"O��y��H	�9c��;f�
�)"O�{�'�<*�8�AD7���$"O0)i` ��V�X@�P,CO@�{�"Oj��@M �(��e�V�ҝC��U�1"O�X#���9L�T��̡V�j�"O�-"�K�=c�a:�g��/P萹�"O�QHb�=f��0���8�1�U"O���jV�B#�ɘt&�_J� �"O�1R�$Ɗj!���i2��%"O��t'·�HdْGX;�ΨcA"O����i�D�|��4'G�s�`�"O�����.�*��ΆC`��"O���(K�y�Xx��7|�@XS�"Oj-#V��>`��QՋ�9E�h��"O���UX<K��*w*�� �PeQ�"O ,y5nȤ0?��'�Q�ZX�2�"O�$1i �4���qn��'EJy�d"O��b/R:F�q�ŌMV3�Q(�"OX��j�&�2�BPaޙL��"O|�K��R}�Ց�֙-�Ö"O� �9�@��+,�������4�n�@�"O���b#ƾ`
�kх�"i�|�8s"O�pI0nӤ�d��JT�-�Dq��"O�q'��8V���@��OyL��"O�P4,��sU�i�O5WS�,:�"O�p)�B��z����(.h' �x"O8��g)��@�xu��
@"?T��"Oҹ'` �?��Si��#6�#�"OF�s�'����(u�u&�t�#"OP�jdl�P�Z��BAK�M�h;�"O$qD�;/���2����$��"O"��e��X�j�A�A��!�"O�4�q�C`i�4����"O��9��XO��(��Y�"�"�c�"O�p�Ce��d����J�Q��XzW"OpXJ�H����"F��6�f@�r"O��G��o������wX8=��"O��ȐN�CF` A�F��$q��"O�Pb��g��ɔ�Ulf�`#"Ot�p#�L!~sС��nU����"Ol�it�UjN�5�V��u����"Ob��IOd<[�˟����"O��S��Se�P��U�+(��"OnqA�BL<U���&��d2�4yD"OTa8�X#	�} �` �C4���"O�����I��@񡇊{�-�"O��C ߮;Oԡ�S���Hj䑔"O(���,��t��B�t�A�"OP�S2�PD	�Dғ��R�^�"Op�'�+#�6���'�*�t�V"O�U�❁G+���`>��1 k�m�<i3S�_8aR��07��U�Վj�<	e'@�t����lL%b�=����h�<I��,d-l����5|

ɘ�i�Y�<�BE r��(���-wV	;�NT�<�a%Z6,3A�	�)I.�rF'�D�<����)y� ��#~sH\Ҡ.A�<�q��=@��,��b��n�*���{�<�S�^,H	d ʖnЛQh�*�˃Q�<	R�ۂ �~8��@��(�V�IQ�<ECH�V�h妓�K ��z�C�J�<��N�[�����ۤ_H�Є�WB�<���TR0�w��##�8IR �~�<Yю�#M�:ABօO k��mJƌ@�<�D�/�Qȏofl���<��A$Fop�r��� x,4*�,FU�<�!�<K�|y�����x$)O�<��ZL���(E��j,�BHE�<y�@�󼱑�+ذ*x�lP'#Z�<1�fףxe�H� 䉪-�|\�`-�Z�<�ĊO�PZ���g@��x��#��`�<�!
Y�r�I�ŏ�'~i� �f�<9�!J�,�6�B�L�`AiRe�_�<�5J�X��G�7Py�����F�<�B���gV���O1)�t	��M�<�WG�A�8�j
8|��U�p��S�<	jM A�l�Ӈ�6+$J)S#��L�<�G�rm��%�/�ĐcG�I�<�BI݊Bl��1V�F-�H�Ѣ]�<ɓ���8�Dp�L�I�*$�uV[�<Y�j^i���K��
i �Y�<a�N/UA� ���0��L��C�a�<Ѣ��+�r�H@d��uY�a�-�^�<	6,
Ip�)A1o7�P�@��V�<� :�x�*۠<��%�Ҋ�$F*��i�"O�`:v*�*�����/��( "Ov�)��;G���(�	9M�a �"O�5���5
���'f"�*X��"O|��3g��uE.$ٖ.5,-f�K�"O~T�D��2���$���[(�1�2"Ol���ZR��c�"�HD"O�����֢��(�,Dp��"O�5��3^O�q�"ǌ�b��}X�"O̝��^�'x��3��=��u��"OJ5�a@�C<\��ȤC��=bE=�D)�O�}j�̷9�<Rc��X��T��>�����1Oh���'J*�&�b ݚ@z ���"O�y��+Qk���ŧ�>s܌�@��B�O���YRbI�_�,��#@�*T�h	�'O�a5o�#QH�O:n�����D)O��*^-?��k��V�X�>��t�'�OP���MMLZ�K�a��=��|�s�i�\��	}�r��B)5��͙�n�9��b�<�>i�B+�仟���2��TstV=M^��S�?D���d��s٨|+MN�iʞ��&�8D�8J���D����Q����q�:O�=A���.L$¨UkZrB}qs��h�'��xb'	��}��/�,��٘�Û����0�S�O��� �T �.���M�B
!;L����	{���$@�6��y�A��:�B�ɵ,`���
 �b"�}�B��i�x�C�~v���2�Ϫwu�B�ɯP�!i9 �]"de�wRtB�	.?��<B���XY)���(TI<B�	�%BC����j�c5�K����4kB�@�$6�P����ԑp���\��`#f�ء��h�R������8D�t��/[��Z�z�-O����1�<D���S�Մ�D9����pU�	`l8D���	#<��A��
���=��f$�IR?����_� �\�;�*FX��#�D�?�!򤂑m�X9�eIִnVRYY�a�!�$��:�3�h�AQ�PS�V*Qt!�$�?j�x���`H*mX����j�!�'eC��I��V��P����:	�!��B�� �,.����ُ5�^A��	O�'��(��N��%���8�'T�)�|D��'/V�#ă�MJ����.T�t�r�'��<A�D	)��Qu��1Lq�H�'I��� �_�\F���c菹B(�k�'����̒	��`@A��;�h���'�H�+Q (J�Y��0d�<D��'��<Yeɹk��q+��4x�'�Ƥ�*/�:HS!/��v0�h�'�f( �C��x#�C�nl��1�'�hٚ�\���H��G�)��
����?	��F$w��QpdV�wM�]@4�IP~�'�4)�eCҼ�r�K7��� ��3
�'�2�1�@�;u�z���\ ���
�'b�q���w>����IܪL#@hYݴ��'6V#nڊ97�m�eZ�a�d�w�.��$�>qM<�ŏ�0G3J��&)X`�0�XM�<�l��K8xeJ�%�'��[MEO�	i�'B�h�1G�A�� ���\F�X�B"O�@��#�i�B�1�Hއ	Kڄ@�0O@ih�clڡq��Da���@Z�y8݇ȓ}(�ʑ"��XȂ�U����=�����T�Q�-���.�q����Wǅ��0=yM���S�? |�#`L�(�i��"��b8���0"Ony����'��%hB(�JG0�ig"O���E�v���$��
@,��$"O���0B�?j`�̈�薿Z(��C�"O�m��o�6_�Չ�A K�1I"O��3��3d�F�3�fG,	�|e
t��S�O�,t��w��~Ajy��	��O�~�E�	�.ux�`ġ^��"@��<O!�D0+'މ�  �A�V��R�|*O>��}R�S�E�����P@`���e��CD�����>q0����|����J�H2�Y�Zw��{��� �E�� "�P�m*N$r���sv�|�xb��JȢ�˞�?��C��׮��d&?����.2"�U���:��a7%�Z%`&�IU8��j�*��c��x:�'��9LjIkV��]9�E��?a�O��D��ic��P cє{)$u��$��'��$�ß|�r-�J�k��B	}�j��3��T��\�p:OF�p�ʐ��p>i��0)
z	зb?)�,�����Ʀ��&�"?���2*;��>�ӼD�Ζ �`g*H�_l,d�G�H(<AbH1S^a�f�#T�L&�V_l|���?遥ҮjAZ�েN�2���c���R8�Xi1��:��ܚJ��0 �q��̢VHNvE�z�,D���a��HڈӐ�X'Z�ssK+��r�����f�Y�'�<-AlQ�2b	�o��B��/ ����a	#J���&���z�hB�	%p�s��Zg�h0ČC!-}�B�I�
z����/ݚ��8Q��M28�*C�I+V��pF�\�b`7I����->z���=1�����s�!�d����aCԆЖG��ȩ�+�1��y���=�&�s��*�y���Û(o�C�5������l`���9l`C�	a��k��wJ8�[�]*�R˓�����10Z�@�j� d�4Y��œ�'7ў��x~2��)C���$j�6YHfq�Q� ��Pyr��	�X��Dh�r%G~�OF�ID����͂:)���5�
�u�r�B�G�&�y�+�,oy^h����?��	��?�&�$�S�O�n�!��e�Z��gA�|�H�i"O�ey�!��Y����@�Ty���E\�XS4l6�O��p��;b��e��.ת\xZ2��i|ў"~nZ�wp�K#�"J#�!�V灻$�C�ɫL&l��jS�b���*�c�J?C�	��r�����E�6AyQ��;>k����,�	�g��l��I+X������:d�B�I�X�Q��07Oa!��ɼd9�B��'�Ts�$�@EQQ�IX�6C�0]�D�:'o,yq&��� 	*���4ʓjN<;�G�3`)J���a��SX(,�Ɠ&�0�iw�G7D�2��EK�x��8�'ô�K�"�.pw�Hb@ݠ|d��1��OH����;m�Ҭa����&�U�ŗxB�'�����`* bn�y��C�BT�!���~B��&XfT+�΋5H�a ,֝�yaԋ(Y |X#F+;~DA�=�yr�G�B� S'*�J�i�W�I��p?�O�ef�� Y��-Z�È5�艱�"O���o��j��ᓢ
�Z3�pR�|U̓�ħ��� :���(Q��?=�j��/�p:!�D�L0�P�@�U�|h�c���Py�f�8e�fDp��� 1�0q�҇^���x�*Ý��M '`A1o�b�qBJ^��0�R�'�r�Z�l�(5Lhg�L���9���'��yۖ �6ZGt�2�ᓞ|���ݴ�Px
� ��1��OBp0%�����qw�'C�O�4��V�X�h fO^ȸ��%"O����/��\�z`3s��o	8�P"O�A`��Z1V�Z�8��`���!"OP삗dY<4����.��2���"O��b0����jf-�$[w��j�"O&T�f���n8���
��9S"O�}2U�9C��QB,��Y� �`2"O`hA1kQ	��0�p���LC"O�	d�ȉ.��q�-ܳu���"O`qc<*&P�����;<����R"O�����3H2���đ\�N �"OV�92A_	T�>�d ȟN�2��g"O��`�eWZ��7�.�\�P�"ONP���֔SmR����8%�tI�"O��a�"Ј]AS�>e��9�"Of��7�e:H��Q�uJح�U"OΝ)G��Bf�8���2++�A��"O�5�HʊX�yi�e�8(r�s�"OF��G%R�Qr��� �r��U�W�<���:9�����k5$,�ǂ]�<$��)r~ ����-5�YZG��b�<I�^�B���Y��C����kr��\�<y5
��O
�<����<����'��\�<��&��<��e�4]yH��E�V�<ɡ��P�0d����	���+w�<�ĩ�q���x�"�	n���W�WW�<��KL�c4�zV,^�@!,��hZ�<ylCL*L��FW��B!s��N�<�Gf�>d"�KI
N̰ �a]E�<!��� .��a$Y�Kv�a��`�D�<!Q$��a�@�&.O�Ԣ :�&3T�T��(�8i�����% ����*"D��s�G�x���`�V�a!�����+D����dϲd�y���vo��*�+D�컑�9*� ���R�k��+A "D�,���\�GƩ:���/!��E#G�<D�D�aG��nAм`�N=��YX�4D�\y��5,>,��O%��M��J3D����'p@RT�Ԋ��UJvXp�%0D�,�VLK�$l�v�?z(S#=D�d@3hV3���@'Y�� X�gB7D��V�P�o�)����l�#L8D��f�Q2���K��J�\�Q�9D�`�#�!���r�o	
��	F�4D��x��֧DB�84o�U�8c<D���Fc�I`�=i�����a�;D���d	Y
7^#����1���%D��00�	�C�:Y�b�`m�HCE<D�s�n:(5p@��mi�X�A�8D��ۆ�A�݊�1T�L"R�H҂)6D��@2�] ;�iq�̀4$~0Rp#;D�[4��L@s �6'��*D�����J�1䔻p�	���Jv�6D���B�2��(��QT0��4D�1U���g
��"��M��!2�!D��x��ַ$�>��c�_5N�$�<D�X U'�2M��H@u� �ve D�Vi9D�xX��I�Z<��� ��q�#D�8��쉐5����Q(`I4 #D�0!�H
�$5P��ȑM�
0떌 D�����)!��o�:(q$2D�y�M����|��J�h�\�g%D���ׅ�Zm|x�fU�z~�YG5D�� �Mنoaol��v"ӛ�LY #"O�	`@���<�3n2�&	bv"O��ڀ�Y~�)F�M�9��"O4l9A8j���aXt�p�i�"O��b�S����KH/O�
�i�"O$`��nx�D�ׁ~�R݋�?OAP0�̸���Ѹ�dҸJ�l���}���4"O>1i6���.  �)ݍQ<	�AZ���@�T'v3B���	�bT�`H��֎T�8\P��G�������0�,5�3,����(%�э)��@�A�Q<j=�	�'W�	+7(E,z�dz�2e�*���P�(Ő�K����O���p�]�e��aѶ����'��A�s�N8= � ���0*��K�4It��ig���g\xӧ���F,�v����X���=��"��y®�S$I0��\.MP���C!��6�jU�b(���<�E%�>S0�Q�苩q�Z�����~X����+{��x�w
�3Lnx"kU�f�)���-����.[���GNѐ>��?cN�i����tY��_8��O��$�Q��F�,\����dW��A�'t�i!�MR$K1§�Ju���4,a�a�@��E�Pҧ���F�I���D�VDP�uZ`�a���y��"MB¨pD��8s}0���Hݢ���"�б�iׅ��<��-�r�*��B�:�G�xX�p�wNܧrZ�	��O
�>�0%�P�h��q׮P6o���D�h�����8g��l�N#Weў�Q�6?tB�E�TeÐ����s�A�!���Iă��yR�h���T�M�'�H�Z�.���y�gJ�J�ؠ�=E�����	��a�4�V$�&�yr�s�td���	Bi�0� ۽�y��IN���a4�DF�0��e�Q��yRΙ�;먱`'F50��r����y��_�%>��H�����1�@�y�ɖrb�0aE�ַU�$P�@��y�dE,y�X�`����I�yA����y�׸U��$B;N��L���]��y�'^�L)t�R%DM8I	�&Ԭ�ybFL�f�4D�&D�Ia��E���y*C�.j�}⫝̸{�^����D��9�4�į��=Q��^�IJ�r0R� bQ!B`n��i��	a����U#
M��,N~k"��f�5L��t�?�����@"v�˿8��3� ڵ=����̊J�<Af�\>d�6�y�Ѭm	�5R��G�g]��{&�$5�g?B(�t_(r�CG�vr�YB�+�o�<�u�L
m�T*�e"f��i�ESΟ����'aZa}rL�c<�q�ߺ��!3�]���=�@�Q�1f��F��0j2�S?E�YXąʛH�ȕ��g�#�oЬz��h�E&�Gx�Oåp?����s�b(���Ё`	v1���G�`��};�m�� �]��[������H��� ��dΨq����0<1@oF�DŠ-{�t�d�7���K6��&U!��1���[�d�`��P�ҕ��=��� j�}���ºUb�b7 ny⩊��X�q �] ��}sEhڇj�����.���2�K���c��Y|&�q�L7 ��1`bXo�<�5X?m�F)����W*��V�,_����&m�i��{墁�o	��>o����*�յ�#�y���+kz�rD$�,z��Q�v�٪��?��!)��K�h�>_��xfe�)v$���6M�9Q� ���EJ�aZ>�Z�͌l�
�sň�<=Y�b���	܅Ef��"�`�-Y��Y���UPL>Q�����I`���-&<�P� ܐ������\�<�yB�KFl0a�ghG�s��p��#�%!7��d�S7��=���ג*� 4�dKB2 �5����|�r9�r��`��!�Ń'ʼF��p���&[4�a`/�=xt��C\ww���D�ʜa�R��f���="6h�a�X��jZ<>$<`�'����`� P�Ya �/�X"R*����!��ʕ�H��'���� ��?�p\�E�ͻb�ޕ3w��MX�S��O���a'��s��Δ��IkFk�y�'m�j�K7��m�̡rcg�mf �9r�l5L�V���3~������ ����C�n�ԑÇ<�I�|�h�EȽ-���QPIy�e�NV
%[��,5�8�'^&�Pq��"ci |��c^ `_f��]hE{4KY��&�,%����uNP�D�`�p�l�a{�� t���3A�x��M�h%�8��Gz͂k���9�l��&�	�r���1E�`ڣ���M#Q�y>����C2�:<�i��C����n5<O>(��閸yO���.u�$�3ʉX�d��b�6@:��x��P#=��(��	��/6y34c�`�5�#�?en��p:��wʠX�ƶ�@ARB׾`�ޝ��.�׿c�ʵ� ��0+R��?�AV
7jR9+��A;$j�� a��^U���U��̡SR�(����4���Џ���.7�֜�Wm^�re�U��ش9�$�J3���~��	8b����'5��A�G-��ēr�"��6�JzZd�x��z�N�aR�nƤ���h5�\R��,(�*�K5��8:h�v���G��٢"��Uq:�'����ք~��h
WW��V �B��]�s"���9*�'*\O�X f�+o���NM$5a�a����D޲K��A`$.�Ċ�f�# H��0���i�;A>�� h�/=R��G"O���	#���	��>4X��aV�y�j0�O�tIbXr�g≉|#q�T��*o���
3`��\6�C�ICv���E��L����c4��'28P�E��!��`xd�ӓ��D�D��~�ޠ�@��=f�剟~�j�!���y�&#��	H��׎�%6������}�͓�$$�ؘ!!\�ac�����"N���r�5񄇂5O� I�^�0,�ku��>!�~8�|"qB/a�FI�#*
�Q=�v�b�<I!��	T��u!�,��1D2C�o���eG�R۰zF�ݙ#����@.��c��<�N��s]�s޺IK��Z�#�B≳Q�ѣ�&@���e`�+[)�a���?��y@Rd�]���0	џx{��
6�,D��%�a1&,On�qPh$.L�M;�bk�R�����6G��D���n�2��䌏;< ec��'�q�F�a ����C@īO>�#F�A	HЛjP�k΄YPv�܌c<n�΀�Ӝ(��ܢ@��J��B"O�Mʲ"ֽL�l�����}$ �v옥/,r��4���S�q� 0j�>MV�O&�:B�;M!��DN3SN���"Ou !�tHx�v�f^d��O�qtDq��mKH�0FE@$9��$�WD�R3K�6
@���ĥ�?*D ȅ�ɐV�����	�?�*�h��^�t���(�; n�v�5J���a�*ZH����aj�.-�5GjX`),��DJ�Lބj�I��7<���j���+K��
�R��ЋV�ʈ�"O4�k�\>/TrQc�͆�3��mx��9%F�ɓ��V60�xH�	�7��>��U��y��O��n�4�i�oš#O�x�ȓ*&<i7�[6+ݶ�k��U�q0D�R�S6sְE�r
� J�Q��������I
?�!�V�V�č(�#��;��Ot�cW'���$ƴp&F�Hw�.#"�����qn�Ç�[?n2,2�!ϡ4�4 �&1�O<���	H��\�]>�hDE<n�x��O H�J�t���I�H�ܭۘO����/a&t�g&͚b���`.��B቗1~���� �I�Y���/ �r�+u���?��ΓPٴ�"ri��R�z�ن�J�I�]>�	"g�v�DܟL[�\��i�x�P��ؗ"��p�"��K���+�:O��Y�B�6�)�S
��bnX}���Oּ� c:���&զS���?)Q�,NҺ\���$Sߜ@����gyb��#9�BaCr�g!"�a��өnM��xg8�n��2���77T�*7睇/@LK�c,p�܅��2n������C�ѩ5��6'�0�VO�Z�:�$�Y{�@+��S�o���������	e���4j��%,I15�rܛ�.̬����Y5o��E;ã4� ���\� s1�Z�6:j�9S^C�ޙ�OvܢC��<����v �Wٞ��$	�,K�ܩH�!!�e~<�2b��148E#'�I����+_�Fϐ� ���)Y�H�cM����%S�����'�f��f��G,j	z���6P���/O���h�=hQ�X����"w�#~z2JY�8Dp�D&}M��Ҕk�z�<Q0,�i)�=p�Iߠ@������7ƨI��"y�*4j�
=�`d'?㞨zd#ي�(\*�(x�,�:���m���B��3,_�=س�"'�����M�(?�]�����<��)br�'uDY��GE�l0P�	�+§Q:���<(�p�ъπ�� ��y!H�?��Dz��L=�@��ȓ^���Pэ۴]붹�t[�i9�ɥO�ecU��6��O��p�E�!=��$��B.j����'{T�4�@���r��5Y����
�'*���'EŹ+̀qM0H\��
�'����Ʃ�T�|�kU�K���8%�\�n�nԄ��b+U��뜔>�����N�2a��ቷ_��Dƀm�h͘,j�j����#�K�V�B�,>�{C#D�\������v���Dh�bJ5��ӧ(�� ���2`��
)+g
��}Y�!r#"O�iÇ��!:]6XYC �ZM�Y(�jv�� �&��h��J5���S���I!h@�:c�л9���
�V��H�UML_���Ԥ�}8@ �uǍ[�Ό��I d�-Kp��7H����AE,���?a��A�9�8!r��2��_�M��p';�J��A xT!�D�/��lI1��-R�|p�aI�o^�I�,�\E0�'��S�OaN<C��>~te��
�1P�R��
�'N�0XQܭU�D�Sl��¢�,}�'X�8�9r���{�!M��Tqph[�@j�5k4/K��?YӁ͌��XaDXM�b��J���@���D���d^�1[6����Nle !�.�ax�i�>^U�d:p�|r�=M@<����ӷwʄ�P��y2#�i6Pâ���	���j����	'Dj5r1��ɒH00py�LƻFʑå��7!�@��lDS��H;Q�U)���$�!���0&���\�_�Xy����q!��2NZI����YT(���+п*/!�$"F�&��P��yBP���hZm!�ă+=�n�h��ɤg��)���K�!�D��UV�J?��s0��s!�Z����Ε�	m��RTkV�!� r�8��3��+,B.�j���7A�!��+d��5�nY�9F���FK�_!�D�r�Ly"��:m1��!�lO ?l!�D�<j���Qe�.�P:�l:!��F�V��l8��S�ߺpP&ʙL!򤑸���dAw�V�*���/ !�D۲Y~��
�|���q�υg'!�d�+B��Y1A��a�x�(�,!�ĝ� ����#c�*�2tL�3>�!�d�R$���L�lpj I��X��!�DA-�и�o�BwZ$�� �%1�!�,oHUK�ɚ:H0VX��L�Hr!�$Y*1��pq�䗃h'ʭ��g!��`Ԗl�&��$I�����C�*A!�ˑ@��wO�6�X H��=!��+y<]EI�=�Q��D�F!�	�H�4y�r�"B�1�@KT"!�	���e��*�9�@#�-D!��
F���(u��zߦ��C�L�:D!��S�l:�p���k��#5��<!��HL���R>0�ّ�.>!�$P>+2V4�a�C�?����L>$+!�d;Q��`���ݢ/�B ���6i�!�M�SR\=3@�&̀��5&��]�!�֓��I@��$����E��F�!��SW`p*1�ɱB���
:�!��[
C�E�����(��1�ɂ_h!�d�Ő�	�i�`pV8s1d�#]!���Op6��tE��KJDy�'B�-bi!�䗷^��x�+�>6�qQA@9i#!�dE�M�@���)�+��q���d#!�WD��Т��e�����ơ5!�dM*2��l��m�Qu����a"O��+P�,�
��Uf\�J�r��"Op�(�=��#������T"O����4�0<s���t4�Ч"O����Β]츃g��l�F"C"O2B#
j�A�p�5/�����"O2�FZ�(:L;EL��!�r��"O�@��e&,D� ��L/#�б&"O�40�c�U7j9��kR�H��U�"O$i:��
è�	�&S\<J!�� ��xc	Nn��3M�#`��"O,��D$� y�cfćY@"���"O��{%�ӲP��9A3�͇"O�"OZQ%T��4���U�W��]��"Oι
�*	 �ؼ�	��J�Z�8�"OF�١I)�p![�h��
R�u["O���V��.��@���N
3{Ё�"O0!`E�;��c�*ypΝ "O(�
5�Q�f]H��slЏ � ��"O��H$��R��	�K�-K!|�Ss4O �;�L������(�g��H���AJ�!*8��F"Ox���n^3젤
²X�i �_�LX�#ҫ
�f��I�K���3Ñ�i=�c-�~������<�d��	\?!ApqHƃԋ>�bl
��ڻ3�B�
�'�\�ī�7�2�`Ġ�|r:���аl:A��)
��O�8PRDOۡgH� S�����KBh�<�Ӯ�*`bEZD���	�@��GM�䦝�"EM�N�\H�>E��4�� :R����8�AOէ$���~��{0��:In�42B������'e�U"�E�?RT`���
	#��J�8�� k��#����՘;L�!���!{0d:w�Ć!�ܑ�Wa�d-Ԕ��'^����&{6@˲��(5��D#��dZ�,������Ӽ��OY��B%"P�cK\|�1+T#�T��'�X�!F+$?�I ���P�H��۴�.�EdƳ
>ӧ���F��{��X(�A0E28i�\=�yb��O0����ޘgf�p�W����D�S��c�EK���<0(T/Ki�ȫ ��,,U؛��V~X��gi,
��i�Z�]CďF�T�˧*�`��񤏥�4S'"�D���VQ)P�ў@�#I�5�ЍD�D�ĭPƮ)a�"G���t�Ī@�y�⃿, ��%�y9�@��%Ȩ�y�ˁ]�E�=E��S�t*��E�wq@�0�� �yrc�.��� �� dL�E
"��y��	�k6dxQJ��eV�y2a�D��y�'ˤL&�U u��4\�ތ
LK�y�ҏ:wN��&͔P)r ����1�y�PAFQ#@)7J����t��y�bG�m���-D(�'nƹ�y�-X�9 �&�?�
,�G�.�y�N�Z�Pub��AKz�cX��y��Ѻ<�:�
a@�*>��,qCi���y2	�!� ����42벀�gn@&�y��>��ܛ�F��&#�ia�d�%�y2l�J6�-`@�߻�����ߧ�y��C
j������=A��4�5�U-�yr�ͻ_��)'*<�\0��	� �yeΣ�6���%�(�`��C�=�y"@��Z�qrU�=)�LHHSL���y�B�h��<{����`8b���y�I���B�r�f-l�b�5���y�H
L6�0�p��"�1�R�Px2I�&��402H�d���#�O��� ��"q�pI�ъ?кM��Qo�3�	K��� ,�0g\����F&ː��DO bt�-�R��Ox8y֬ϤM�~�Y�F<+%>�ڰ�,F0�����O6ȓBèپ���@v<�6!Z�!�v$E�a�剄idX@�Ț���]"@B�BG�Y����v��q��$ �nS!<9$�@���r ��+�!��U�7I(�i�W'y��3(8T�TAQ���b�d]҇`��:���C5�ԗ3O ��'���I4E��yG��5;Q��a��S��̑�C!�2"�$nz�m�V��	����P���6�f�1�glN��(��+� �;3�V2~�]�&$�����>Q���AyȀ�@*A�2k���zh��|�AG�?i3���h@aB�"`�)��7(�&�1�eʻg68IQ��.#�����RWV����R��a{2!��}ɨ��A!�-���	���V���,
8�M�2��SF6]�+y����Q!7.�ذidS�R�ݸU$�@���I�9	�<!�'��V���;� ��U��T�	�q3h��bĤ �J%�"(Q�I(xz��\$RdZ�/T�)�U��ყt;d��O�EQ4�[&
�� �����Ӎ&N�a���u���|�kS�FƏ�ZH��̹���7@�(���9ZL@'�
� ��yycD��
T���䁀w��pi�1J� � ����'����G�NXځ �hΥS���c/OGu�4�,OJ5��� �i#,ҕp*���U!+������	m��+��K�.N؁� � ����F���Gr�dۢ�]x؞8"��ә&��`űU�tL*a�R�p�.����,	N$;��� �;שR 
�� ��V�z6mP%��DNOU��!%�մ/���[1����<1u
U�)���;�F��y�kM���G�؉-�p)�@��f��`�����<�"��
j^<r�+G��!ܨP�<�1�rA�#������,Ph$qA�|�\(Z|!�$�2.�K�bU�rq$�	>���!NJU���׭Gd0����>���� f�j�(2��i�,Dz�#��b#���ҏ�6���.�%u=�ʓ�~$��O���`s�	b��'��0�
�2R����+�b<K��Z�A��83��'T��_6���J�&�%�ք��	(��B^+��lz�B�ɼ#SVM�Dú��ɼRϐ �N�p��<+������&9���>1��ưkp�b� �GY�u��e�E��:9��x���J�	D�?I�G,�fǜ�h�,�}5xi��?D��FGɐ[{2�9�A
�Lg8=R�!��ks��O�dB�B}�g�	���#��5?��$´�J.+�C��(���P�B�6~�o�!^�{Eh�  �B��'U�8ɴ��BHB��*�KZI˓���r�Հ4��ʓz
h%f�
�r�p�"��Nu��ȓ� ��Qh�e@h8p�A�k�\x$��X�D�)6�&��p���y
�!/�?&���I�c̀CA$B�Ɇt"�]H�B�4��9e�MIi \W�_E���+��p�~&��V��"�����Ͳi��JG�>$��K�G�)a���b��*(���Q���|~ԵB���(T�}��FL�\h:f	Y,+�6E�p�D�<�Tl�3[QTu� ��<�����g��a��
H��dr�v�<�c �'R� �����}1L������I�|5F��㭎>����<v%�����!��Q�P�;D���N^ ���G^-T��#��[�qOr �1�3?���պB���h�KU!J�2�q�l�o�<��(S�S��q�$��!�P�y�`�c�<r��
(c ɰ�l�M4�1�
Rc�<��$��=;д�UhG�qa�Ei�G�c�<�!�ިG����	H�dE���p�<�7���j�´*�k++�P��jGo�<����"�9�B;!��dB�Mh�<�ae6G�v�bG@�P����	�i�<�B(Ry*��6%q�	V�k�<!�����A��6y`|�2`�O�/S��a %�'2']ÁׯE�<���K�9����vH�ik����I�l,0�\+j�RPAׄݷD�OPXE��O^�+��T�|v5�1��f�.�YC
O��&�~L�b����#Aj p��L�	b���W!D�E� q1
� Jl�ඉ�7�p\ӏ�	~ �I�L<�A�#B�{^X�30�d��F�Ȝw;�	2���v�FE%D�8��@F�;⪔��[��BW�<�r.��7b����\�5Dj$���i�|�
xt$X 14ȃ7k@!��+nj����>>��]p��/K���f��=�B�Z3d�P���{�U�?j��P���e���"@J��?��hջ9���{��n�~�*��=/��PpĬ�8t�f0��Ǯ�0>y�᝼3]逑́�33�\��f�T�'��hd�G5�����ÛGP���"��9�����F�R;!�ā.|+dM�M�629��ycΎp>�ɴ���Ȧ���:<��@�K�J�OW.�r�:$�-s ��e�i�'�d�Q�)��i���C.zs.A�H'����y�2�����gܓe���w�>���NE���%��	�d��h0��/�D�i4���.�	[���4T}���Ga}��T�`�����GY���&��0<a�NH�g;J��H>��K�N�1d�(���#V�g�<�$FŧP��|9��P�<|�ƅ[K���{ �z�{��Ti�1|�"� �8}��8h�-M��y"���,P��	4��t� Pҥn���yB.�1����Gm��k(�� E
��Px��	X�? ��C�A���aw�����%	.8�!�D�#��@��̈́J�����S/ax�#6i,DB�|��[����ǡ�)D�Tܺs��7�y�*P�-�NL��_�2�U�������}/�d`6)J
��)�'Q��SR�"k.���V�N�>e�<��W ��	�f��> �	ׅ�U<S%�>Rn�8�X
N~�=�K-D"��f�C��V#�*���B=[�p5�I��r���@ ��,/���pA *�
|;��Z��*ea,Ɇy�tQ��F�'w�����!�a$>�I��m}V�zd/���Mbt��~�<��Z"[�J�r��:9zx�H�i�]yk��{��رՂIg�哠	�Ś6�@�jo�}�F�޳>2C�	D�a�蟔C�nY�/��J0|�'����7.�|��ϸ'th��'�1)��U��-r^����Ovb��t	]2{�
�qu��
�VAB�i�G��=�g� �O� �	�,&ɑ`�C<c�F�rr�'�b��`��'D��j��)#�\*$!B�X�Y��'����0��$2v�s�bŐkZJ��I��
��E� �qO�&0x���u�dlS Ay���"O�$���%)��Q��\�8mr�!�"O��1��ƸP��Dё�b!�A�!�d�U^H�& K>B��T����/*!�D�,���3̔�7�"�t��{
!���-oR�!��9`�L�x�J(k�!��V sC������ Qݜ�ۂ��48�!���=k�^���!�����f�I�!��WG�rTb4��!�
X�祜�!��s�t��7MI;;��R��H�*w!��N(m��ԠT�5}OPuQRk�0o!�Q+�H����~��ì��H!�d:�~h"��G5P��U)���"1!��Dm��;`��/a���!OY�!�ԯ@Äiq쟼3,M�ĩ D�!�D͖8��͛�"ɚv�@	����L�!�D�l3�q��+z�(�W�!{d!�$�WI�H ��6ib�8Z���#|�!��E�k����dC\ b�*��s�!��]nξ=��D��.��gɏJ!��	�Xm���hȘ4�J��g�ب
�!��+��O(f� K�@ �!�d> ��,�c�88��Uڣ�	�eq!��}ހ�`�*B7%D�Uw�ɥ!��1�h����Q�mȭ
�!�܇:Q
��c�^)_iR���BB�]�!�F�%�6i[f���cNT��!�=[p!���^@ā`Az�Pp���@ ��6�(�\X���'�<q⃄�8�̑Po�69��ڴNB~��ֹ+��ȟj��ဇ{Q��ad՚�H��V=q|��;?���)�F����.tF�!��X��kD~�,Ք'`�[�QP>�� 	מ
�����K@�<���"�	���� hz ғ�L>�ǦܮLåa�0��Q��>a�@Z����A�8�~�'�Z��V�L1j�X�E�p�T���=n�� �F΅P�)�'J��c �I��YCv�T1vlq���[��`[�x�ՙ���:��'	�Zmk'*WqU4��጖��y�@��6v�p�͓�j���o1�������Q���g@�{ʨ9�cJ�|�����|�����?a�D���8���:9#J�5��"H��S�`���#�D�^�x-z�'�BA�7޺&fE�j�^��spT4{��3pB4k��	�E��X�RQ��,�<U��j�z5H�1�U����*��s���G�T�B1�����P�����0��F�]�q0���cI��� A)-o���}<��IzO~���.��xd�O�bUŸ#��M�ӵi!F0��А�8:�1��P���	��%��(iR�^�eL@�UJصY=pʚҧ�6ہ+Uo}��M�i�b��;OP1�Ƈ�*AO���N�"~b��ft+td·Vj�c��@�v�x�qfW1BF�ҧ�g�i>��I5l��*�WW�Р��Y_�0YK<Iu�C����h�g�? �`aΔ�(&���ͮd��Ia�J~b+C]
��;�"���SČ-U�D�sO_'�l��]�l��{�h<yu#7?�|��'�|�0�-�6++�d�&��	V�@�*۴��a�vE�,�F�1��WZd��D�d�]+Y��Y�i�0w`d����ڜ)'ر��jޥ���I�M�ɑ
ç!#����ږk� j"�`*T�ȓH@�eڑˉ:F�!E�F}�̆�E.Q*Tk�(�҈Q�n/�����.2�ޝ؀��Z)� B�>�!��ǣ]Hn�a�G�8L�~�
P�R!�HI�M;V( �}o��`!φ�Y�!��N$��Ey�����^-S�Ά#�!�3V-�,�uG߁o�h���f�!���X041d��&|H� K�%T!)�!�ć�^�䂅 )<$�p�i��o/!��0r��$Ж+G�h<x)�*D�} !�#� e获8D��k�6P7!�DJ�U	���-<%��xd+�BQ!��GApUC�(�2MU�7�K*@!���A�$�#��2�q�	ƍw>!�J�)a&�ӥĊw�t���N��!�$�?l���ro8C� D�J4�!�d*Uwr(&�Ӛ/4�0�h�@J!��W�!+Z='�H!�B>!�<AQf�B�LL<X�a�3m!�$�^dF<;��A�s4���UNJ�P�!��3����֯G�%���u뒹E�!�$��n�.QR�ӆ}�b�+S)!��9T��B�߰@�̸��7�!�d	�b��P�]�}�S��ͤ�!�d��Z�(��e� xleT�Y�7�!�Ą�w�H��"jrx�T��T!���	���3%�1$W\�ٴ�&I!�X (��]Ʉe�).�8��8L!�,^�%*�B	 m�(r��#�!�ڮ"Ĳu sBܪC��P ����2!�I�w�ɲ�!����#<d!�$�'���
�s2L}�f?G!��DL�t"p91�:!�Ao�n>!�� #u�]ّFY�S�����֯dF!���j"�� *.$�"��6C�3!�D�4b@}xGb�&o��h�'#ߙ5(!�dT�@|`@��Ӽxg�i��|!�D�V��R0�1�t샲�J8!�d�4��!o�"�8x �ꒈ�!�$����(������"�Is��=�!��!
¸�o�#~��w���Nb!�2���H�E�$i1ׄX9{�!�\zr�Z��H( ��ܩ�CLl�!��@x�qY� �;��@H�ԪaK!��G�:��`i6�����ђ(�:O�!�$�,S��C��ءB�`19fh�:�!��%Z0�m��j��JN�٩���?^�!�d�m�8[Ɔ;��j�&�+.'!��T��k�==����)�8�	�'�am�>0hd`9�^x�'#�8�C��B��C�U	9�L`1�'�X��u���K��h���"� �c�'C�ĸ!L��8���3��]�-��'I����M� ���r��an�H��' ���GL�@s��3M���	�'M,�x����2)��Ҙ3�|:
�'�@]I�Ώ�6C�1c���!
�'	�=�EfֱV�T��T�(���	�'�^t��(?�p[�Iӱ������ x�@���[a��t��'�%څ"O�MbVDP�Y�ӰKGڎ���"O���Rŏ z&�P`s�Q�|�8���"O��`A

����A�D�	��"O&K��H�"N4B��(t�[�"O4�Pđ4#j�� ��$Z�ؓ"O$J���+Ni���ED`v�bU"O�Yd�ɢV��Q9o�6wRu8G"O��7iS���(p2��)PG�5#�"O��3!�89��n;�$8G"Od��qE��Y��`1D�,TM"$"O�lS@jU�Q��qq
y�^��D"O:�;���KX��)a�R�&U�(��"O�� ��և
�.!���1'[  2�"O�aS��H,����םk��M��"O��h䭁7���Pgǁ5%4<Q�q"OB�k�r��S�Hͷ"+�qs�"O`$�u)��k�*a�B���P�*O\帔hԐ]��Ͳ�M�l�0e�'2:Y`#�M��]آm֜R�$m1�'U��#­�V�"U0e�K;J�] �'"�;f�؟ar��G�.67T���'�J�Q�3a?X�Q��V�|���'�>u�%A�����|>H0
�'�I�B�"mۤ�.=pf��Y�'S�is����F̂�ц��	34)�'4��w��oݞLif��\��*�'<�����N�G�Q;sG��Y�Ց
�'ʞ{���<]�b�#����g?T8`
�'B��	�^F��A!���LPA	�'T2�
�6#�ؑkʴy�	�'�B�Y;#��!h㙆P2u�'s�%��'N�
W�K1`ڐgZ�[
�'��EB�%o�2�p1HӴ
$jTS	�'��	�E��(�� F/ғ}�>�b�'a9Xg�K\}�(�t��q��'v��b@֟l���[��A�e���
�'�,@�m Vz���T�nd
�'7�����H�c�f������o����'���4#)X��� ӬГy��r�'���BG�O2,��2��j\H9
�'��Уbˆw�,�I��˃fU���	�'��[��Ҷ.\���
��
�'b���	�1�|m{d�����!
�'����,ƨ�1�$�0z�X�	�'��8%��Z��$zaN�x/��@�'�+cm���t AP摌C��q�'^d�D�4tY�I��ܜ=�� �'j�����?�$ta��-5��]2
�'�f�3���0T�Z��Y�1�*܂	�'8Z(c�Y3T��scפ^�p��'��l�Ê�YZ#b�X4ܬ��'��hPW�Z�~ @��R�J*O���"�'X��$թ&(0���C�"�k�'Q�)a��\�&�����Lq��''�!!'K��m���x�V,��'�.��'�j�
��t`E�o���"�'��tQ��7w�P �*���VY��'�
=R&ㅿ���;��%v� ��'zNy�/��`0t�R�C�~2e9�'ۢx��O(-&}z��
�Ƽ`S"O
|�EoȩF���YH�9!�T
/�!�d�|�D�"�\� e	�f��>!�D5}�\x�Be��r\�� �fN�-2!�� 4`��Ȋ�?�J4�D�Ì>g���"OB�f���{�Ə�hT�h;""O�4a�ҭ T�AKa�Q�nf1#F"O&H���ğ=٠3��K5rI���"O ���Phy�h2��9*f��"O�,��k�%a�&�l'���"O4��4��#mH ��-�P}	�"Ol�+Q�1��$`��@^�LȠ�"OF䈓ℭ[0x��Q44���"O%ǝ�t�AQd���[�*�i'"O޸(Ӆ��%��	6KФU� �#"O�ti��;}�J�qd�R�H$�"O��K��Č!cJѐ2��!4	�4"O�r�L��:�n\��	-�\	�"O�҃GC:rmz� ���\��a"O��ڒ�J�Ќ��JC�"��"O
�
r��[����ANcn��"O�$�vn���2d����Qav�*#"O�U(�,]?|](d��OA#�\H�"O���T��lBD����-���"O.�ڤ�
Sz��E��"v,l�;�"OJ��f	�3A�K���j���j'"O��p�g��$"⅒qeV>�"��c"O@ � �E5iLԡr�d�]Q��� "O� �V��M���<O�a9�"O�px� 	�|�9�PL�U�R"O8[!��[¬x6M�m�Z��q"O����O�T8�X:�ŉ3�8=�A"Ox���Ll���:p�($x���"O�b�Q�V#Ux1�H#8eb�;b"O�CV�_<޼�+�ǟ!]dĈ�"O��*�苄)��hRF�0hj�*4"O�� Y�7�<)���dF�4�"O���o�~�$��`l�/P�"u"O�M��IF.q� @��l*���T"O�ma�e24^$���\�x�"�I"O­�Sf�f�ʅ���;��:U"O� �!��W�qˣ��62���ȡ"O+O�&D��m��I65� 1�N�<q���" I�4g�����Q�<�&�)|3���c�u�`�RAJI�<���Ր;z�X�A�;.^ �� OC�<�v���2Δ�a >?��#�Kd�<�W��<b���AѨ�8c�� "墍\�<y#B�.)r8 +��A�%h.I9u%�[�<	��Fr�mB��ð2�(`�F̋Y�<u�**�걃�+�+v�x�2w'�I�<��b�LXP�Q
S�0�>ڧ�VO�<��Lzܶ8jTLDB��2�L�q�<1A���gS���'��V�<e�bh�y�<���(
����wN�xZ6Kv�<���ߣ:����'
��<�!`�t�<��A ~0�$#CfJN��6&	w�<J�9�&��%O�uw"��GdH�<�&�U+N�(���>	��d�K�<��h͍tR��F�>Ke��8G��~�<��S��`�Q�,��
�*)�G��w�<Q�+�(&�؀��ش�ڜ��q�<��j�^�l�J��O(�%C�D�<���-٬#&T�1��5��D�<������A��C��}��mB}�<1e��ma���5Δ �P�y�<A�3/ń�I��u�K4�LD��C�	Ql�42�$_�h�D��vC�)� �*�/�,?L�⃄�=���"O�$��Ɣ�K���V♚:�:*c"O����C���!^J��i��"O��2vM7i:į�N�P-ð"O�*0��O�j@�n�0S�h�x�"O�\�' �X�i���6_���a"O�S������K��M8b��,҄"O���b�@�z!Yď� ��@��"O��G   ��   �  B  �  �  *  q5  �@  L  �W  �b  n  �x    �  x�  ��  
�  N�  ��  Ӱ  "�  ~�  ��  ]�  ��  "�  ��  �  N�  ��  ��  ��  w �
 � � �# �, -6 �= D HJ �P �P  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e�'��O��P�]�۴$G��d�q%"O����bN�#K��X	0�O�#�yԮ���v+T�4z��s�����yR"?�EP���2.�R	��%z�=E��\Ȭ i��3Qlh׮�	.���<
�<����$�`�(��@�ȓ|�<��TL
!��qC!o2䭄ȓ~��s�X�\]��9�E���F�<I��^�C�}�R��-�h�J�L}�<�A0ho��+��ݐ%�]bUC�^�<���ɸ{�Z\y���6a.�Qe�Oq�<1t
���A�G��J5�-�3�o�<q��w����EQ�*@�p�S�<Qa�,��ms��Q$i�QzREY�<9�����A�Ђ8�3��R�<nM7w�jǁ\ۦ5#�E�N�<yt�g�zQ�EcKU�Z����q�<sK
 1rT�h�$��B�O�l�<!$�x�Z���U�����M�<�V�h1�\� .jV�S �G�<i��8�V�+s"[,hn��UaE�<��_�P�S��$t`�(;���J�<a�C*!�$�r4�KZt��҃�Q�<eب)����.��{3�����P�<A��]D"A�Di;c��%�ЩCM�<�B�<.�j�D�g���RbaDL�<��!İ<0��i�H�k�x�$�Q�<	�mO�
a2�*kC���[3n�H�<q�M&eP�(Q��^� ��%&͛]�<Aԇgގ�Ƞ��$~�$���s�<!�H�E��q�4�
,g�<	�c�q�<#Դ
���(d*�E�VD�9�!��6x<y�&F�(9&P��G�!�D�;(G�̨#`H�4�=�� �!�� 
%���J�]���"����"��,�u��k�O�m2�gӝY��Y�s��A�h�
�'�0	p�ˊ�F��0a¥�;[`�'Y`!��N<�lh!��5dbh0�'�,P	ĩ�$1:�p�0�Y�'����yB�'S:�H�Ļ9f`	:̘�s�0��'j�)⃬?m�F�h��
�|?V9��'��qz�aT<1��:p�A�CO��	�'�+�Ë�~'�$���;�zL"
�'��Ə�|��L9�H�7n�)	�'|RD1WA˞_@jy2�$�+�Ib�'�n�*̇�<����P�R9!%� q�'q��siW�R��´��Fd����'�i��xg\��4�<@�rl�
�'HQ�Rf}�>L�3BǨJ<��	�'{ȕ`7�W]< �;Cl�����B�'A�	��S1[p�i!F+0B���
�'� Თ�ə	�:��5Kڲqp�]b
�' ��A�(�.l�<m2��:o�0̘�'��`��GP	����B����)�'°HA��E����B�P�|p�y
�'�b�(t�b&]q���C����C(D�ph���jz T�V��pe���2D��q��T�Z��)Β��uaw�1D������v�ز��ˊXkĉ��.D��"�%D�wE���0kɊE�¥�!�'D��sfl�6�Z$��n�c����Ո!D�x��(U�!�2q��͵6�b9Z�#D�t��,ǨSY0�C'�L�P��5D�ș������][�᜴|�!
��3D����_\愚g�*}�*��*O���$�wX����F�.m�rA��"O�'ڱWy8��䯓<tf$�"OP�[��A0r����M^((CA"O|�:�%�4/:y�g��*A����"OZy꣪�2���J7@w@u�"O�x�© ��ic�ݴ>5\0�P"On` 쑺l�Ȅ��eގ,{�)��"O�YbW��g�2K"E�9P�"OX�ɠ���?�p#��Z�iA��"O\L�E���7������ݙa�, ��"O�Y�bEچ)a�)
5/� � �ZT"OD�Qt�Y.m��x�c��?HK��Ѷ"Ox��W��KKp,�Ȅ#8;6M�"O�a���2�64J�E��xB�"OH� �c��5�Ҹ5PĤ<9�"O��	''N�E����	����6"O��p�3��!c�枠E����G"O�uf �F�{���w���"O�,8�37�ڵcg�"rx%3�"O�����Ь��o�4-gP1�"Od4x��L�t��hC)�E��!w"O1rnZ?}y.��0���+�"OЀ��F�zCέ������A�g"O.�Q3��%L���ʒ%�NEҵ"O.��K����M.��pa7"O�h0'×8x�kgiE?���8b"O�����Ɏ/H�� �Ֆ$��S"Of�5cI�p�(T�v�؜^��"Omx����scH�q mA6W��H"O^��@'D-lX,�!�ɡ:\NU�6"O��"��;�}5*ӃA+����"OV�
Ԣѹ���1'!
N�"O��`��#��eۇO@� h�`"O� d����Q:W�ޭx�M[�:P`��"O����1�n�P֬�>r1zB�"O��s���یq؇	3{"~���"Ot�{�J�%��A��zB��"OZ9�&k/u��hZ��J�;� ���'���'���'���'�b�'�B�'�:�+�$&�Q���[1@�����'/��'���'ib�'��'B�'!�`���FH�,@��GJ#w��7C2�'�R�'�B�'�b�'H2�'I�.ٶBc� �"0Z�5$퓇���'7�'���'y��'��'�"G[�g��}y�O�}4�ZJO�I���'���'�b�'���'B��'�bϋ:0+� ZA��+�d�穎����'Y��'���'"�'�B�'���B�*��h��^'
J��j�!6�'B��'��'���'!��'@2O��c-f�RK�5��H+v�(�R�'�2�'�B�'PB�'���'���Y��@IY����F�,:�R�'�"�'1��'0r�'_��'��C�@! ٓU팦n\�0�싗8_��'�r�'���';2�'J��'U�٥K��
�c�'_Q��ka�7\?��'��'���'���'g��'5L�Mx|���
z4`�	T�r�r�'s��'�R�'b��'�'��&��ȴi'Ζ�M�ZG��
�B�'��'���'���'��6��O^���FM4\jb���';"�� +�=�T�'?W�b>�7����-���Hf�
t��P�G�x� Y��O��mZY��|��?q��޴.Ԯ� �2?�(��g�8�?A�����4���h>M2�����M)��c-�9[eH �$�5{y�c���uy��ӠD�������x�������*�4ZE���<����f��.�.�j��CE>Ό�i猈[�����O~�Y}��t�3sy��6O�CdF�}t�Đq�ޜn�X��?O��	��?�&�%��|�Lp�Y���ކ@�Y�4��3i��p����3����E���"�6���ċZ)0���.���pl�?�RS���I���͓��\5h&�[�N��ĉ��+R���p�e#�!4Vc>q�u�'W����xo��b���s��Xf(�/r|�|�'r���"~Γ��H+3��" ܊�A�I�	/�*��/�����dH��}�?�'RpЬ��#=Jq.��秊� ��Γ�?���?�s�^��M��O��,�J��&$^"�s�`�% W Q�� ��PܒO(��|z��?Q���?���7�DZ��W���փ�RiN��+O(9o-�2Y��mޟ��	�?�6
�ԟ��I�~�!�� .���Β� llB�Ox��(�i>�����Õ�@̾�ۡ��x6����Q�_����iy�n>Dz%�	�G��'�	�n��Y�T%��x)�lC�b�
i�t�IƟ�����4�i>Ŕ'��6��ttx�D����ѥI�Bk׿0�C�c�Of�m�R��+q��ޟ`�Iԟ����;V�¹iY�����ކ"�`�[b�����'� �e�?u
g��d�w��P1���"uR�@�P�Z.n�쁙'���'=B�'�R�'J����hVy=���o
9&�Ɛ�B��Od���O� oھL�J�'s����|2 �p6��S�c a ����&U�w�'�����D'�3i�&�� � \�7�|@�cI";E =����Hl�r��'1� &�������'�r�'�ֽ�Ȓ��z<-Sz�h��$)�?����dئ9��c���l�I�d�O�0��n�/�0"r,R<m(���O<y�'-��'�ɧ�I�':�Pmp��/�$t��	=A>fx2�C �6q�����@>�%�D�w�:���.T.`�Z �B?n.���Iߟ������)�sy�`x��Ńs%]5n,�,C�X	��!J���ų�^��Sݴ��'�X��?Մ�6RA@q�u�E��B��$	����3wD�Ѧ�u����+���
iy�h
\�,l8�(K>s]�$��i��y2Z�p�	�,�	�0��ڟ`�OG��9c��5a�q��'WI�hԇl�B��V�q@��D�O�ʧ�?����?ͻ'�&QS1k���ǧ��n:�{��?�I>ͧ�?���=ZP�ܴ�yR͂	nW�p9Ao99�x��d.�yb���T������4�<�z�4���	�hNs'��<$�$�O�4�?�.O�pn��E#Ҹ����4��9��ِ�ؙ8 e���>q��?1�W�����$�l{�F		�4����\44�}
��7?)�CK���9�Ā[�'������?a2��e(�
"�d�����?����?a��?�����O���nG�v��K�E:Y�ĄJ%�O tn4|��'	�7- �i�5Y���'�r ku�F�@<���w@z���	ҟ���7��)l\~r#�g��	�5P��(�%}��s��	���h��|�\��S�x�I����ʟ\J���,n`!���oP^���vy"�y�x)��O����O���󄔷07>���
T�)^N�9��Fd��a�'@r��I*Q��b�n�hR��9A��ɯbGެh)O�a��Ĉ��?Q��,�D�<Y��H���m���[��Y�+S��?I��?���?�'����8��ß�HwMƔpX<�-��Z0�U4�T�������?�^�(�	[y�l�L�@髒��/YNRQ��FH�a!4�i���!��e�O��D%?-�=� n�#�T+�m�E�<*�T�I�;OB���O.���O����O �?��h�`H��Q�B�f�T�qu��Iܟ���4rL��*O��o�K�	%S>u���F��IT�Ӿ-�@c���	ȟ��IGh�lZ�<���6J�|
�>D�|9i��GuN "��,W�P�d������Op���O8��X� q�����5��!�a�I�Q�����>ʓ:%����8���'�RT>��� �Zk0l��k��WN�$� Mc����^y��'R�|�OT�`@�R�T�B��;��� ��tE�(E�./�8�O���L��?�q�!�$_;���i'�]8O2Rm��c_�B���d�O����O���	�<V�i����e)R?ht�(�4"�., G�۪X��I%�Mی�>���>�z� V/R3R(�c�e��n�d���?%�?�M��O�nY3X*��)����$��$�V4��jF,g��4�� Jn�$�<���?���?9��?)*���KC�|��{��Ϝ|Ш(�n�>�<x�	ޟ`�	\�Sޟ������5��
C��<PV�C����:�?1���S�'7[j]��4�y"BQ?�h1���U�ΥUW��ϓ�v-ON�D<�Į<��?a�+�n|(gɔ9�p��MH��?I��?a���d�Φ���˟���⟴�wC�aVplP�"�;G�d���j����I�����z��	l�P�mހ~�q0�@�(� ���0���X�|: +�OLS��ݠɛf���4K��
�c	D�Jh����?a���?i����yŸm���?1�iۜ%�d��d������"ݯ�?�3�ig�u��Q��I\�I՟�]?mn�Z&#҃ZG��
���p��	�������x�a@���̓�?���:=����=�ZX�l�N��l�O��"/��'�x�����'b�'�"�'~����#H�B�i�5�/yd�+�S��P޴	)4����?�����)�Ob�$�36�8�� @ȶk��Œ���9N��?����|����?)%(�'[�dԨC[��R��]8f���0�Gy~�F_�p������rt�'��ɪv�.	�$L�r����Z�w�>��	ş0��� �i>q�'��7�ǛGP�M�7Y��ӷD4
i�-;������������?�R^��	ǟ��I�N$�*`LD�o~�8Z���f�0 ш_����'_��z���I�O#G�S.&��&��;�d�$��.�y��'|��'b�'�2�i�?4�,�J�(	�ʹ(�M�<q�\��O@������qUkp>I�	�M�N>�r[iM(6��5%����!����?���|se ��M3�O�\��A/uX�١�/,rqѳk�Cs����'��'��I���	���I�t�M:S�9)E|�Q�T�U��������'�j6�^3)θ�d�O��D�|�7j�v�PG�*+b
4�Ip~"g�>	��?H>�O�VL�#v44:u��S��M�Gb���Q�醊S���|:���O�5�H>Q#��{�|���"{*$[�._&�?����?���?�|2.O2d�Ӆf< �xW!�4p���+Z�!h�1`҃�<��i��O���'�2�WV���@$-�}td]�qگ`�B�'�F<	�i��iݹAdl�?u��\�����`�P�Y�~�Nؠ�$s���'�B�'���'G��'��Y�������P*̰�� �s>9��4�������?�����O^�7=�`�q�ÞC�| �支v*X��R
�O��b>i"�Eަ��F��c�5{�^9i c�b>p Γ��Q�7N�ÖhL>�/O�d�O
L8ckΏ �$$j��M�v�1���O��d�O �$�<�2�iO"`�@�'���'��ݱk޵P�r[��n���b��{}�'d�O�H���&�������V^�1[�����%f�N�@pb��L�S�O���ޟ�)�Dߒ'1�p�g�^�]M@��_֟��	ޟ��Iȟ\E���'��Q)��t����f����>A�w�'��7m�t֊���O�mo�b�Ӽ{��(+\��CUŁ&s.���D��<���?q��=! u��4���g2(q��b�^�#�I�P���af�\�B�5�Ĥ<�'�?���?����?yV���9" ����2/�P��	U'�����Yá��H�	ޟl'?M�	u�\�ЇS�E!��F�/ ���O(�$�O"�O1��@ #�� pY��P̄'�(��T{o.7-1?� gGU\��Iu��ky�F(L����%��alЁ� �8 Q���?���?i��|B,O�oZ�]��	
ZS��R�ݲ@�DU�V(��f^d�1�M{�"J�>���?a��)2,"���ln.!�]sK�T  �ܱ�M�O�-aQ��"��T�w�Dl�F�:x�ki�0u�����6��O�$�Or��O*�?���8 �𰦊S4G�`U�ܟL�I̟��42�ș�'�?��i��'J���!�>;2��dD�&&Q	��|�'F�Ol�e
�ia�iݕ�1+{���m�� Z`l�Ap�V��ɓ/��'��I� ��џ��Io:��2(Љ	8tHS'95~�������'ތ6Mˠ6r��d�O���|��'s�~i "I� nPhR֍�K~�Ƥ>Q���?!O>�OS�ё��Y�J� x����0J��*&�9�k�i'��|*G��(%�(��I�|�\�KG�Բ)Q'%�ԟl��㟠��ݟb>M�'pd6�M6
�P����WOU40��bn�O��d�����?y�_���+:��%��]G� �	�O�,�Ҹ������̦��'ʸ�y���w�*O� n4:s�3q�$5�` �qq09�5O���?Q���?a��?������m@L���ǃ�J���F܆f�ld���'�Ҕ�t�'�:6=�R�	&/�.).-��,D�cr,���$�O���2��IH06�7�s���U�-Ҥ��W��-��
h��q'�@�b��`�I_y2�'���+�Vl1�|�6D��r�'<��'l�I��M���������O�]a�	��z �ᡲi�H�8����'�D��?a����qu�1��a^-���T
��_��A�'%���C��.g�����~"�'��p�)X��z���-�^
��'�b�'���'��>�	'&��M�CA.s>���A.�@�	��MC%�����Ҧ��?�;Y�bd��"٧v���Sv�\�&�z�Γ�?i��?�Cd��MK�O���U/�?�ڑm��GG" qD�SI���6)ܾ(7$�O���|Z���?)���?I�_�03q�L�S� �3�m��p)������I&�Qyy��'��O�R�C�N��k�ʁatH��B�ߟQ2��?����Ş@t���%�H�l��-۵��+��,�>hR���,Oh�ⰄE��?9;�D�<�)؜L�H��pȔ�3���Q�E3�?����?��?ͧ��$Cͦ�s����s�D��T��P��nMa�H�����ٴ��'�r��?��Ӽk�MMZ~"51@Ύ~�bh���&9:�޴��ē�W�2uk��M�Ғ����Y�����O�s�a� [$���O��$�O��$�O��$%���":(&�X�H�+�v��8g�'��'�r7��W���Ob\na�>� D�6�Kk�l��D,qX�Q$���	ğ�Ӑc��<m�Y~Zw� �����7<�l�ue�('2n5�q�Q�^]b#�d�	Dy2�'���'3���:�:Q���H�nΰa5G�C�'=�I�M�u���?���?�+�&�IvKAmaY#�8u�5b���)�O��d�O�O�Ӷ ��P�ag��^䰹1��ˈ{�eRK�~P��!?ͧ������a� ���,̷�4���Z�$,��?���?)��|�7���?+O�!�S^��Ĉ�mF��@�}ƪ8���O�d�O"���<ͧ���O>����
(����!Rvb���O,��� D �6Mp�|��;�" ��' R��hnn@�"֯	�� �OP�T�I��?����?A#�F;�?a���?���?��->0��Fmǆ�n8K��8*�����$5�h��Y<�?��Q�������Q5F��D�&pΙQ�Z�r�뤂9e����OD�_1Հ�4�����O�	��Lh�l�I0thGH#7�����+K̺�Ɂv�� z�'1��&�����'�(��v�܍omT��Akް'G0U��'>��'�rV�@޴jWj�����?���W�b���q�\����F\
�;���>���?�K>A�K��D�$]�C�U����M~B�;B��PQk!�O��@��#r��%Q�$��� �:98�uXs!B@~��'$��'2��S֟h	�
��.!��LJ;�H���՟,@�4 �Lq���?�q�i	�O�n�7��P��F/P�h�d�dq��O.���O(��"�x�t�/L�׃��Ȩ�af_?"��d��nETa�N������4���D�O���O��d��Z���#�������"vhUh�C�<qf�i����'�B�'���y�#r���8VnR�s��t(��ꓢ?i������Ap��Ш��&��`kf/�3i�����e��ɽh��1r��'��1&�<�'S�蘕N�D�F B� �T@c��'���'����Z���ߴ#Ԏ4��>W��̇'c��lKr���M��ϛ��Jr}��'�b�'���P��P4�L���� `�x iF&8���d����<,*��i��9�onĉA�(��P�\HI�>O�$�O���O��$�O��?�Kp&��6����q珑{TV�'$���,�����޴���/O��l_�I:*����*0��g�0$���'��	���� vQ�oi~Zw�����د\{��rA�e�`��d���~]�M��Nyr�'1��'(�#P���xw�̖T�6hQUY�p��'L��7�MK���?i��?	/��Ӧ�2�t{��ܝ2��x9�O\���Op�O�t�j��n��+��X��@7nAl���mK~�O������W��y�)��WѾ��`@T2?����?���?��S�'��R�9�'N]�kqH�-D��*�@k9��*O�8lP�����T ��R��B6	�}��my��Iݟ�I�?0�l�J~��$6��Y�Sc�)\�W���	p�Ol~�X6 WH�D�<���?!���?����?�/����@�
w�\!`1��h���ÏƦ)��������ҟ<'?����Mϻ4�DI�G�:X��0SI�:�,qK���?�M>�|�����Mc�'A(���C������U%{)� B�'�>�:��
J?K>�-O���O�y5G��(�D�@&O4�YbF�O��O����<�E�i`&���'���'�� s6�G頥��`ǩI��ͺ���s}2�'I�OF�k�nԞOM�����@�ˀ��g��`9Ѩ�p��@���z�q��ϔ�$�VEG/q�:PI�Ce�$8�+�����ߟ���ȟ�G���'u$�ck�e$h4`�f�=3a�����'��7+<-���O"lc�Ӽ��]��Ժ�cb_j��<A����D�bL,6-;?9&f����)]B�? d�H��W�Q ���r���c�0 e/���<����?����?)���?�"�_���M�bā�h�$�� ܫ��$�ڦ%�q�����I͟P%?����p�F �`B�"� g�^�W�T99�O����O~�O1��<�4[?Eâ�u@Z'>t�xZW��
�P7mBFy��Ӫr�f@�����$
J�a�HP�FrP�)��	Y��D�O����O��4�&�U����,U�,�	A����"9���8W%9S�"��L⟘ʯO���<�w�	t4����~
Ҝ���I�8@nu�ܴ���B�=)�C�'m9 ����� O�L R	�X�Ti�%�Z.-����O����O$�$�O���3�S�FlˑL��I��HYg�T��'��xӆ��1�?���4��D�T�[�ֈv�,A�e�P�Z��ThL>����?ͧrh���4��d�7}����	z�f���*V݆P˓JC/�?��I6�ģ<�'�?Y���?15I���(0��C�)�䣂�?�����$�Ħ�Xp�I̟0�IH�O,���2��	 ��/f|�+�O6�'����?�S�,E�c�9EN��W�F�h��L?U�R@��mX?P�8���������p�|�+B����l�r���$��1���'���'���tZ���4�~��w,�]�"YS�O����D΍�?�������H��`���؟��P���YP*��AB�V���n�ȟ��I�R]m�h~rn��J�t��}���[(o�5{��-oЅ9����<�.O��D�O��Oj���O��'�0�*�S�u+��౉�(P�ޔ���i] (���':��'
�O8B�z���(U�
���	�.X���*�2?G����O��O1���(��a�.�%;x1ֆ@8L2$aU<I'���cY�9��'V�'�������'*
h
5�H�H`��P>�<*��'�2�'��Q�B۴A�Y����?��$����"mH�2<X�ԏL�wotT��(�>����?�L>���� ))f��ε�D�N�t~2N�k4�b�i1�zT3�'�r��LPM`�F�%1�X��G߁~Cr�'M�'[�sޡ٠f��=8�I�.4��x���Bٟ[ٴ~;8����?aбi��O���لi�0kG�l�����g���D�O����O�H�-}��Ӻ#����M<<��d��̻U��h�ǁ�J�O��?����?���?a��=�J<@����-8@��*G)�1b6nʓ0����J�'d�$�'UV�Ra�+X"$��i@=?ʡ*��>��?�K>�|zVJ	��D���aT��	���ܚ`.D�۴t�I5��,3!ܟ�$�4�i>�ȖJ;*fP�bk=~�fI�WLğ��Iӟ�P��ٟ�3a��uyz��bk��q{���+<�`Ra�^>�9�c��2�C5�(�4�̩oZџl��蟸�	�J���
QcB�����ı� ,dͦ-��?I�  R��i����d��f����\�^�"�2Y�I)�7S����O���O����Oj�d)���wv9kEaW;{�<����7*�0d����	�M���N�|j��D�V�|���O�dm��L���\���R�'������A�~����l���ӑ>�� [�.`����bROQH1��'2P�&� �����',2�'D�e�(�� m� ��M�*�dA:�'��U�4�ܴ<zX����?������H�,�k� w֠IjQ��&��	����O���'A��#�N.c0̽�e�?v�����W1�p�cܯ��4�F���s�,�Op��rț0�`��C�"/�����O����O����O1���A����G�C�ZI�S� A�c�
kL�0��'�B�`�b�@�O���Q�
��)�rc&z�$B0�ĬV"Z���O:�R�fd���Ӻp㝕�0��<��`�W�����	�bw�#+��<Q-O��D�O��$�O����Odʧ]+0�	E�Ⱥ>��܀��	�lZh`�%�	ޟ���o�s��������ˣ^��i�d蓹F��H���'�?����S�'=�t5��4�yR��&�n�B�2e|=r@�%�y�F%Q89�I!��'>�i>��	#��y��DY�yp3�߮mn
a������Ο��'��6�l�|�D�O*�d\�q ����-�xak�ds{��ܲ�O����O|�O>D �@O���Ί����FMi~¦D�!����:W�OU�=���:"��!$�p�N�/!؉�w��:���'���'�����\{CQ����%��RE����hٴW�<%�)Of�m�f�Ӽk��
�&T�5X�BUt�P��'��<i���?a�s��-��4��ĝ�)�����'.��	�H� u���1�OK�!j2����;�$�<ͧ�?��?����?�b�w���x#e�J)(MiV�#��ߦ@��U	u��t�������kkX���ǟ,�B,ލ��H&��1@%��0�MFyb�'�"�|�O�r�'��fһ(� D�e*��<j������8�&��O���A�?y�2�ĸ<iOG,�BX���d
Q���?9���?���?ͧ���\Φ�(�I�2Ѭ��o��i%��r��,�B�z����4��'Ͼ듡?Y��?��%�\qb#���U��݁1��-d���4��D�k����'R�H��&���t�z	z'�\�<����D��r���O��$�O����O��6���
���0E����]�*���Q���˟\�	 �M+�Lް�?a�!5���|b�_%?�(ȸG�/�Zp���L���'��'��@���8O|��ȿQ~� 0E�W��Sʘ u����p'Ҕ�?�1�%�D�<i��?9���?�w *<S�͉4�Z h7B�{���?�Ԧ��'Uh6��_�l��O����|��U;"�$[pE�v��-A"�I~�&�>A��?aJ>�O���%�yZ�i���3#x|�uJ=^(���%����4�B\��?]��O`��k�?C����7'Q�c�QÅ �O��D�OT���O1�*�E��6�=A�0��0C��9*B��R&E�H�l��'12�t��⟜�O6��Z51?V��cAʇgq� ���|k��$�O�m�2~���Ӻ[a�H����<1d �IW*�`�0_�+�����ey��'E��'�"�'�T>AWɖx�̸���u��CM�MSGCԃ�?	���?yJ~Γq}��w��5� A��3�%�ő�'̸, c�'p�|��t��/I�;O�qj�I�|�≪��V�FHf��7O�DH�n�(�?9�D&���<�'�?�+)7�>lZ��6���ͅ��?i��?�������q�G�M�D���A���uD�x�	�[��(SQ�1c����@��`�I U��Z���c�� !��٣f��3Ǌq%+Ƕ�\JN~���O\�x]TD��� �(��ކK2 �����?����?���h����I�-.��9��G�x�F}�'ʡ-t���Ӧ�C���L�	��Mӎ�wm�HمMB�4�F��"D�j�ٚ'�b�'"���꛶���1ke���J�P0 �/4�"��S�̓O��|���?����?���f�1�Q9��Ż&(�q\�hS*O��n��&���ҟ���^��	�����Z�r�n:f��,b�4��_����0'�b>�Q�7�X��E��-/�����$�o_~B�_�Nrj|��䓻�D��*�1�/Z� ]\33�Jd�.���O�$�O �4��ʓ9��ʕ;CX�M�����τt���ӫ��yB(jӬ㟀��O���O���P�9�ep2J�7�ƥ�  -(���x�m���� ���䟈�>���<�hx�"��]<]R�:2�{�|�	�������I����U�ǸFz�X��ۏF���'M=�?q��?�u�i@���O���g�n�Od�#�&���@�u���0&��O�4��� ��{����x�R V6#xlX���+��d�J��h��p�Gy2�'��'7r�E�)avXx�kC&�2�i���/���'���0�M#����$�O�˧��1��[M��MpsmQ�,z�)�'��드?i���S��Ɩf12���-}U�u���wnly`��A�tQ�9P�O���?!��*�D�S��  $EJ�dJ���;��d�O���O���I�<A��i�y��S5'�V�[B�[�/DJ�iC�4G;��'��7�)�	���$�O�����/���uC��%�b��O>��$�7�-?�ċĠ8v��>��Mŋ�
�IdFaD�Y�`�3�y�[��Iӟ\������	���O��
aЕK8�a
�.ր��@c�}��cI�O����O����ئ睶}��<j�K�xJEy��a������'�b>��5����y͓,e��8KH�c�dBŇ�&Le�}ϓb�$����O<i�L>�.O��O(iҶMUj@BqB�1��,�q��On���O,��<it�i��2!�')�'��9����(Qf�*A䙉n��l�q�|��'����?�����j+h����ߟ�@�� *ƤK�bx�'�	��l1��p����Bӟ�pP�'<~��h�2MB4!z��8h`Mu�'���'���'+�>��ɼ�l|�����o�6��K2��ɘ�M��a������Ŧ��?�;[��r�M^O�k#OL�5��P��?A���?!4�@��M�O�ȓ�6�
4kq�dYP�"�$e�g �<�O.��|���?a��?A��/�����u�A'S<g;�q�+Oxdmڐ��1�Iݟ��	C�s��c�ܟz���$q��@���A���$�Od��2���4� 9#�F��d�¹� ���zz\aA��3���y������'|�$��'O��������� eIB�� �'r��'���4S����4x;�@X��h;>�@vKۃA��Ś� 
5m�V����P������m}2�'Z�w�&� � ��⌶o�Z�*�#�S����k�@G����U���9cWH��a'L���#�/E���!.}�|����@��̟h����B���:��Aj��_�B?`Yڲ!K��?���?�5�i�4Q �Os���~�O ��4
��<�Ƚ��GU�-yV���1�D�O��4��Y�@�n�^�@`n����Le��Q�K��D��y��س^���j�	oy�O�"�'�(�(U��+t�͌]v��`�X���'�	��M���*�?���?(��8#���4q��ԏ3*A*`���ӨO��D�Ox�O��:�(��6hW|��	�bA"d�ܽ���R$>��ioK~�O��D����D�VP!C��7*��Hd	<8�����Y�V�R�3ִ�
�J��`$0w��_���03�'��fӆ�`��OZ��*��\Y��[i#��v��c���$�O.�+Á}���$W�[�Ǻ?��'��q��PY �a���b�r��'N��V���3�jOJ�	
��ɤ=��R���2�M��L2����O��?c���k���@|�����O���%ȁ�?����Şa��Mxߴ�y
� F}AJ^�XD�b ��~R�A"�?O��[Gd��?�'E6���<�-O�� *�,�J�o��v:a��'7��,4��˓�yr���/`0���պk:�DH�
Y���'�V��?��������[�-�{��а+CZbU�'����K��+"0�*P���
^���*��'��퀡[/aT1�n��)�a��'��9�Cm$~W�3Vm\�Y:]���'�6��KǠ��O�o�{�Ӽ�g���-%f��+_-�
��׬�<����?!�-L� �4���@�"!�1��O2*0�ŗ'���������"*��|�P�dE�������]%=_qI�G��d𦝚�Qy��'�I;FjZ�-� &@��N��aCu}2�'�R�|��
]>t�TAb�a޻U����M���sC�&nV剞*6����'��}$���'��T�S#4:�X@Vҥm�5�񉼤M�##�?I�FY�z�f�y��Kr%*e���?��ik�O���'�R�'�RK��8�� (U�J�)2�$�i����Ȅ�Rҟ������S5��Iq��P�$@����%,0�.�O�%*�k�-)@49��#<���X B�O���OV�n�3\F�'?@���|����X`�tC�w�&=
���~��'�����T�X�k��擟,�����D|�P��)��	�䴐�J�<}��B��O~�O^��?Q��?A��)9mhȎ%��	ȺPp���?a)Oj�l�P�4���ʟ(��B��,֌H�P\���Q2�3�瓱��dIL}��'/�'����XR��y���.��y�U�d^�%�X�%�.q���'�������K��|��B�;F��p�ZA%0 �(؆	�'���'���TV���ٴ]��$�� ���aۯ3���;�f �?�<���CD}r�'��T�`�ތ��u�#�Z�^�"P�U��z��Ǧ��''�8 �?��՜?Ѹ`�8d�,;��E�~��\0O�˓�?���?����?����i��7�b}���Ay�d2�Ķ>���lZ�/��4��֟���u�S֟�����1��==���Æ\1@..�S��<�?�����Ş	@`��4�y�ݠ�8W�2,��Y:f�O��y"!�sk"!������4�����E��AiE� �6}9�EQY����O���Od˓^*�f��w��'���'J,��C�&sCR�N�90E�O�'l��'K�'8�<���?����v�N٤O|8�-��x��6�(�Ӄ}��$�O�esv��:-�Ԃ���V�&�����Oh���O����O��}��t���҂���U�* $a^�1��͆*J 2�'�t7,�i�m�7�8�,i��N�r�NT1Gr�\���4���E�nv~¨��Z���,�t����lyJ�$�/>=�J>�*O�i�O��O��d�O��r��è>.l�7�N�dT(I�<iq�i-"xR��'�"�'�O�R�_�
�209��$@d��d�>����?����Şh}�|x!B�8�饬��)���j󋉧�Mr[�HQ��_H��?�$�<��Rb� 4�Y��N|��n�!�?���?A���?ͧ��D��ݱE�ǟ�1j�9h��xqa%�ms(Aٟ��޴���?Q]�P��֟���,;�*�k#$TYE"�+cX0��nɦ��'��a�"�O�J~���:���Ғ꟣P���@Y��ϓ�?i���?����?�����O�H08�`�M�pXƅ��69�$h��'r�'e�7-XD��O��l�Y�I6ҕ25�$Z����LPY�l'���I��S"T\�oZF~ZwX��i�m��#/�@���B�l#�2cꖙ'�R�OF�	Xy��'"�'BR�\�m�L�����Ye`�I��T�b�'>��*�M���6�?���?�,�.)�7G�&u_H���M�Y ��8O��$o}��'���|ʟ����
�� ܓ5�G9� ء��΁"~�H�2n�=\����|j�Od��I>��X�@�RAЫ�i�����l��?���?���?�|�/O�oZ	O��l��"�k��tI��S0N����ן��	��MN>	��(��Iǟ�M����ة�b�(�T�x�Ëɟ��ɞ%�Vl�^~R��06b(��'��$؆k<�\Z�fK�؀���oF+7��<	��?���?I��?	+��qi�	9>���`�ɑ�;���ܦ�µ��џ<�	��,'?�I��M�;we u!��z��*q��,Jp�q��?�O>�|�Bł��M��'�ZX����j�p#�%L�	�'�����N	��W-߭��� R�B�9��A1P��<~�ڍ
�h�4Ȫ|�������@�̊)��C-ɀ͔AKj§6� � �>=��q'O(S���:�(�*f>Z��ǤF��ڲ��<KX8��&�&H��T0&
�<�Z�Q�,��ÁY*n���y!�pM� V�W E�� ���<H6[��/+&tra�K�cir�PB�kDx�P��O<!
V��աXĸ�S֔���F�W�Q�ĉ�G��Z�/��t�ѕЬ�����(G�{�j��!�
j��	�2)Q���@k�)�"2.���c~Ӧ���O8%��D� �N}���f)���^6m�O�O8�D�O��������Ex��c
�Q����ʙ�x���'I"Z�<�Ab�����O<���VM�Ff�*\��,���'v�*��NW�I̟��	)g��IL�I]���lZPac�� ���#��Ц%�'?��%I�.���OX���ק5�@Ò^�Q���ȷMr~ �M���MS���?9��U�'�q�� �CB��I�����hԓ&�8���ix�l��z�>�$�O���,Y�'L�I.E
�C➹�l5�#`����Bش\v�����O��0J��`���!�~���b`��e��ߟ`�� ~u��ʬO�ʓ�?��'�����A�j8�\*��LmvT��}b,]�'�R�'Y�G�D=ԝI&ǐ31�( p�#.�7��Od�5��E}�R����W�i�J�`����a���i L����>�P�����?q���?A+O�)�3��\��BFm�������ݵZ��'���۟8&�d��۟�adAZ�]��D���_�N6�3�	Z&�&��	ڟ��	Dyr��&�n��"x�JН�B؀�nW(>�6͠<�����?��[X��h�'�N�u��k�z�c0`G$Z$�i;�O��d�O��d�<yt�������U(Q�pg�Y�V/��1�� ��M����?	�N��{R�UH25".ׂ)��� O��M����?Q(O�`W�Uj���'���OdT)�u ]��;��,�GY`�'�2�'��$S��?�P@Ɵ	S���T#<H�\�$i��ʓbp-�5�ih�'�R�O~�����"`�z�+���ə��
�M��?A3&�1��'�q��1�v!���ʅ�Rf�2�d+�i,��8w�u�����O����^��'+�I��t �J�;�D�CU��~��ش4˨�`���i�OH6)�l���$)�Q�#o�M���?��J8顴Q��'r�O�I8�+�K�5e�A��	*��'����|b�'�r�'fx5�f'߼K��	y)B��X��� g���ć�N�H$��ߟ�%��]�/3V���)&�Ȁ���X�ZOz���<����?�����d��a#���͆D��`�a\Pq#G���ē�?���������<q��T:�\������z�i2X����ʟ���`y҈�Y���S�q�$�)�C�!O����AC�Xo���?q���䓝�4�����QR�� C��v�E��E�-X�'���'	�Z�x)���ħf20�8�ѽ���!C%�2$��	z��ig|�T��ҟ���L��эE�+��AdO�~�z\��ig��'���1S�m�N|�����1�Y���ěU.������c���%��'���'��yZw��2��+|Y�9�%�Tr���4�����qV�i��'�?a�'�	�Q�}�&l��.1��& �6�<	���?)ї����4@��J9f:Ja�3mDЩmړi�:|�I̟��	����Gyʟ��!cF?[t|����R#J{�Be��V}��
�O>�gF��L��MR�b̊V���b!���Ms���?a� n�k(O�SZ�$�!�� ���4o� 
�N=	T�<Gx�n5�Sݟt�"��+��[�x��$M+�l���X�0N]oy��~��2�X
��U���*I�u8��h9�Ol���O��?��L�=-�	� �;!ܦ(�B�J;-�.��+O���O6�d��F?��"�bE����	_��X����yc�C7�ǟ��'�BNf)�)A�1��!K���7����,� %����'�����O\ʓZ[�m��$ !��:���C׶hN:��?I��?y*O�X���g��(����s�_���ç�Q̌���4�?YH>!/O�)�O��O��(��Fs���jS�նNg̕8�4�?�+O���ݲI}˧�?�������(����r���� 倾/��}'�l��Ay����O�.�W�:����#�B�ҷ-�(��Z���G�U�M�_?��	�?e��O����uJ�0G@�}��Ǵi �I��T�	7�ħ���eX!ᄻ|6�u�D��,����VNfӴ-؅��O��D�O��D���S�4��6�d���' 9&--����)��C�6�Fx��I�, B�0XGA�^1��1v�ǅ�eo͟ ��ӟ�ڡ��byʟ��'~À��Y���S';M�x�/h𱟸�䳟����A�Pg��CA;rή��Vcq�p��9~jʓ���k��_�TzE-�Hܺ�@D�Ro�{w�x��^7����O����OH˓;#|���CL;�<�cd�nT"�!`ٍ8#�'�B�'r�'��i�%�EZ
�)@�M�% �<�Z�N�����<1���?�����O�d
�ϧWVA���J6c R)r�N��}�LL�'T��'I�'U�i>)�	 �69AS��10R�ZS�H;t��O���O��D�<q�a�;7h��؟<A�M�V��˦i'/4�@TF���M�������O6�$�Ox�	=Ot��-�����DoD�y��ti�>���O��#3�	J3V?����8�S$0��y1H(u
����)E��	`�O@���OJ���1���OXʓ��d��p\@h(bDĕ
�x3��9�MK*O���dE�)�IПl���?M3�O��@�H�n+��,�h�ڴ���՛�'D��]��y��'��V�'ff�=h$ӊW��]E��;AfR�o��lt��A�4�?i��?���J+��Ayr�9oT��b(ߖl�|��A�X�7�M�_B�d;��-��Ο�Q�K��r�n|��U�Z�R�SG�'�Mk���?a�X��T"S\�|�'�r�O�)*��FL��$��V=f<�D�i�BR���#�i��?������ �P��, Z�>3�$Vr�\��i��(��b� ����O˓�?��b�48� �N��<�0��UG��%�'��'���ȟ��l�:��a���<5X����*�F��`���ġ<������OV�$�O<�KF�F�
Y��ˀ�F�Uf	! ��<����?�����۠MW@�'�p�(�E��:��Q!HiZMo�Ly��'	�̟L��柠�%�f��X�.S3d�e� �<>�������6��$�O����O��tbf���W?I�	3ˊ���Ȋ�m��(3m�.N� ݴ�?	-O2�$�O��D����Of�
�0�̜0�l�#�F�ydߎf�n!nZџ���Hybj�e�H�'�?����s�6팝�B�I=\�q"b�!%��Iԟ���ӟL�	k�L�IMy�ԟ��m��; �²OőQ�X�#��i剎�e��%��(���?]��O��Ǩ?.+�O�\w�4����6B�Hm�ߟ��I� ��I��9O��>��*M"7d���Z�^�ˢ��f뛶��7��7��O����O��)Jt}�U�HJ�-@�.�f�sEN Do8]�u��1�M�����<������8������"kD0.�e�9S2����#�Mk���?9��A�y��[�d�'DR�O��ZE)C;��M��*̒V��(���i��I���a�j���?����?QE)��:��q7�8,Z5Y�ċ;SěF�'���H��>q-O��d�<y���s+����QBk��(�TS�V}".*�y"T�`�	�����Py�`�������LQ�4�(��!���a����D�>�.O��D�<����?���z���l�f�h�cs�	�KU��N�<!��?���?I����d��B�&��'n>�A���7�M��d܈\leo�Ey��'��ş��	����bn�@`E� Iu�J��D;;&YB�Ç���D�O��$�O�ʓA�(PW?M�� Ie� ���S �މ)㧍=�"��ߴ�?�,O����O����y��d�|n��Z3v�dh��M$h_(3w�7��Ob��<1�i�m�������?��e����m��?/��	�Mƥ��D�O����Oj�#�	eB#^���SFGAe���g+�O�˓�}@ �i���'�2�O�f�Ӻ{чUEg�xj�j�1a
rp
���Ϧ���ٟ$�fa�,'� �}��	�
�d@
+�|YC)�%�C��M;���?����X��' H�H
(�j9(q��ެx�W/pӂH��7O����<����'�D([�AO�2|����_-z̘RS�{�b���Or�e��Kw}�W�$��S?��/ ���D<>5�8CpO��I��@yC�yʟ2���O���9>��;T�r�	aW�(Qr�Ql����@�U���D�<����d�Okl�.<c� O�m3hS�B�.1�6�'��!˙'c�''��'�"V�ذ�/�(X��N���J�ht�3$��YʩO�ʓ�?),O����OX�d�"�r%�e�b7
b#FL(Tx��#9O2ʓ�?I���?�(O�hkQ��|�Bˆ�x�8���5��I��M�)O�D�<����?a��V��`��[cI>DMD���X��tl�������Iџ��Iş��'T�H�B�~���T�t�'��v#L�y2�x��с��i��_���Iğx�IU^
b� �!^[�A G�"�tIT�j�Z�d�O��z-�p�'T?���ȟ��� 9�%�q�4!�VE+��Ҥt��`�O���O$���2���ty�ҟ�5�L�w�,|���gql`h��i��	.3tt��۴W:����@������
�*7b}��*,Ue�<�GQ1�F�'�f^0�r�|���ۋUW��F�
�q�+	*Z�f��!8`�6m�O���O��	Y�I퟼�"�
=?< �k�ᐶF�TC��<�M�@*D�?�N>�/��˓�?�G�n�̅K�C��ns��Z��¸ �F�'���'�fU�>��OD���p�ƃ��lV�C�3v/�!Fo�z�O���$��O��D�OkLO+  2��S��*R| 1 ��t�F�'Pz���**�$�Ob��7�������U+U�]i'dB�WЀ�� U��X�G����'&��'��Z�����l<� EK�V4�┪19���}��'��'���'�.4��G.n�3�a�[
I�R%�>�bP�x��ݟ���Ay2��$,���ӋL&L��4삘N���:5N�+�O4�D>�D�O6�L�$�	b��1NJ6Ww��)3��e�B0�'W��'oR�h��N!�ħz��%��:y�ĉ��(�~�h4���i�2�|B�'��b��y���>9�J&*u�0	��9$�U�%A֦��	ޟ��'?8���K3�I�O���H&s�*�!�FΕ8����F�$<N�i%�(��ʟ�§y��%��'G�ޕ{Ԍe��E�F!�z�o�{y2�B�4}�6�]}���'��T�,?Y�g�;l}�ik��Ɇwj� �P���	�I��H����ڟ'�4�}��,�1<a�m��� /���4e�����M���?9���ⷙx"�'^�!xghܚ��ҍ�D�%�R�|�0��^���|r�i�Ob7�^�{-�p+f�#`��S%h�	�Ms���?Q��]����V�x��'���O��U�]�d\��2 �:(��f���;[�1O��$�O2�DW)	���!=S��v�&P0�o�ן`��@
<��'��|Zc��h���O*7����M8jT�®Oz����O�˓�?q���'9�ΘHphۿ<�1J���"Д  ��x��O��<���O��$4&+��{��+��p�F�/K�(��'�O�ʓ�?���?	*O�8W���|� .H����Px�Ċ�� �6��@�x��'P�'"��'�,@b�O��BS�( �بR�2p�	"dX���	����Iay�bϔ�,���"4,<�]ん�	��r��Ŧ�E{�W�$��z�$р{��0q�'I�b`�p��
*�V�'��S���H��ħ�?�����L0vf�����	�*�X�*J���D�O4���=�v�QGd��@0���f��b7-�O��$��F�h���O����OR�ɤ<��r^�x:�f�.b�R]`f�H1���n�ݟ��'��ub���t(�n��0늲7D� m��M�K(�6�'���'����>�.�u�`�"i����I:s���E�ɦm��Y�'p�'�"`Qk�H���M]0��y��0[.26-�O��D�O~�8w��O��d�|���~�k��na��5�Mnm@� ���
xFx#<������'e��'w�Ձ�,R"ަȢ�Jٟ�
�Y�C`Ӛ��_�Jp�$�Ov�O���|�,�,MM2p����,�B}��]24�'��B�O��d�Ot�$�<)��K
�*��;s��W+W����Q���I����	ߟ��?��aș(�	5"�JlM#FK�:����|��'62�'�R�'�,�(uן(�r��V8J�Q�ȝ�i��Y��i���'2�|��'
�	�k�6-��d���$�͖v<%+QT�|����8�	]y��'d�%��^>��I0Jr -�%S�dC��:��>c֌p�4�?iN>����	pȉ'&,D;�n*GYrH���*��)p޴�?�������.9r�&>����?;%k[V�D9+�	�.} �{�� ����?��a|0�#A�+4̌����0��mZfy2��F�7-�_�d�';��;?y�j�)ZӺ}��.�	�A;S�ڦ��	����#�>���OÞ=gmJ�xbШۏ_��Tz�45�:)Zu�i���'�"�OS(O(�dƸO�� �2��$MtM:󄉫6�F5n�7$��#<����'7 ��fJ�=S�5Y ��	<F| ��m�����O����w�������O���g��p���C�2�10oZ"E���$�[����	�@;-��|i�tAѸ�4�X��M�i��,ZaR��:�����O��'h��%K��R9�@�GD,H0Z|PJ<�N>����?�Ħ���ǟ�Ҁ�� ��ݑw ̪���'I/�I�'<��'"�|��'	��΍X�"�hP�  Z�u#�#G�w~��䋻��"�(�?���<9#&ʟ:�*��V�_��y�"O�,����?Tx�[7� 7]���`��ԮBHJ �gP� <��0�� ����%�c.%����Q�<��(��_D���wg�.|a�q�eI�p���Z�I.8cT��e�칡D.��c<80�`�4H	��f��1<,�yf��~�,��g"l��Lc�#^�i}nhKgj�$UH�P��)u�H�cɩK��0�EE7U����G�������5Ș�2s�K*��'L�jD6#i0ٶ$�G�8n�|2(��� w��V���/
LPT!t�>����Z��AJ- ���P�S4��`8t��;.\�!PN��s��'[�\	��?9��i�OX�����`�4*�c̵z|���"O���k�3׎����-b��'��#=A�f�
b��]	�*ѳ!(X��FY��V�'�2�'(���(Z����'#��yg�G�M������V&��6E��?Ȳ���I5��d�6U:
0�r�|��F�{���g�$���3��71���Iܤz����'Ih`p��L>���
Z���h]6B�F���E�?1�O��8���t�,tg(@"�G�0 ~�����M1NC�	1
n�Q���c80���10 �vő��Sßx�'�-�`B45#�M	�C� 0>~�R���=��P3�'��'��`r݉��ß�ͧF���s�O]�!��D�Vm-L�DJH�0��9+�k�\��x�	ϓ�|��'�U �hZ�E�qs���bH0f�ta���"Z�"ϓe��"��=�ڐ�	�Q��p�a�D���	T�'V�O �����5=4`H.�/�d�@"O�qX��!����B�U�N����������yy��S.T)��'�?)d8��YpFGH)2��y���A��?�o�t�����?��O�2����Z���MW����!db	�J0����3K)�ݻ�9O��S
�	^��%8e)Kp?�0O�8<p$��@�떏Qj8��ؑ��O��<I���a�\���nPt1�j	�H�1O\���P�@9|�b񫎁z�-ȵ�"�!�$����!�]�O�Z$���T�cb:as������'�Yɧ�e����OB�'$�N���G�:!�&�Q4����A.�G������?�����/�Ir�Oԕs��i���ɱ|e���X��Mr-����}�$� ��[,�B��e���S�^���"R�A�xڊ����@8��'����Q����7ҧ�*r(�c��ً'��r&B��h��x�#Әl�|$���-c���l��0<)��,m8*	 �^nP­`b'6�,ͪ�O���d_>$�4�#�U4���ďPb�!�� ��Q$�>-����!hC�1)�"Ou��K������OI�Y�Ez�"O<�c�̷%��ɲ �Ψ\K$Z�"Ohx@��zC��Qd���B�"O M�r�0�zp����0[�Ʃ�#"Ona	/F�7,�{�`�Ff A ""O��� �Nv��W@���C"O��س�H���:o��B�d9ʢ"O�LP��ϵD��cD�����s"O���M���`g�4;:�u[�"Oz�����>Y>Ua���q���"O�l����:WFp�r�2�&�a�"O&c(PK"���T�#�,�2�"O4(;��JvɃE�܏l���a�"O����&u�,���&�*��幅"O�`j�I8.04�A �)��iS"O���r�	a���Q�H	�sv���"O�*B�ܺtA�5�P�À_!P"Ox� �-�Z�BFCȝ`�b�k0"O�݋���_#�P�UKߦS�����"O���@�����ũ������"O�<�P��K�@�TfY�s��A"O�L2��A�U��yಃH�C���"O,%�U�J��8�q�֠A�*$�'"On� 5&˿}�)�P$U�h���V"OD�e΃{�����ȫoW ��e"OdAY���1)S�V�&D�zd"O*����+u(d�Me1V���"O���VdV<c��̫�	�F��9�"O�!��;8ZRՉN�-�f@R�"O�e�� ^��B�.β��I�"O*�'O�B! Dr,Z�S�6x�b"O�pX���l����&k��H��k�"O��j��P=�zUؔF�Q����"O��q�W��5i���4�4{B"Of%����+��鰉�0k�ܵ��"O(**5E	x��UI�i���+"O�\�N^�U~�y�6(�'SBR���"O@���gԌ]��s��#&�"��C"Oܕ�A��n�(X�I"i�B���'f�e3�Kaʽ�C��>{>��\�o��� Kn@8s��&ZA��Ac!�wѾ�F}2��7�>�!���2S��Y� (2�ԧ3D��˃*�9;����MʞF��p&n������Vu�S�O�����Ѝwr ���M1����'3�-1B�V,+�z��F���@�O��P�k؞�#�m�U�,D���/;�6�+9�O�
��iӊ���O�=O��Ÿ��˯2	�(�"O�MC\e|~D�a�1�ܛ���K�'� M�C铫b2��G�N<Ll���\9n�rC�I�.�l� �Ȓw�T���C��:�>�LN��Gx��逭\aL4K�-�'(�M*�Fy�!�$Q�.��AI
�B���!�.Sp!�$҃;�\ͨ�ʐ!? �*3喰KB!��,d�� q��U��u2S�kX!�A�*� q�o�7r�T(u��n�!��@�c+�tA)J�bW�(8pO��!�$W�^0�4�@O<`qՎ$�!�D8QJ�[���(2��b��+p!�DO+.�� \�&���1`��g
!�߈uS����0Ts��W	�!���Qt~��i��lkWs�j���'�V�j¦J�$�⩑��A�c�v���'�"��	�$*o��R�D�H:����� H��~�4kE����"O��륨�\�P���Cݜ��*��'���KM�����آ�����"Ĵn����(D�j�T@qL4�PD	�m�t/:�	�	�dI�y�����)ͷ(	
l�j�j���V��4K�!�$�>{ϠH��t�bf�6jr��s�v�r�r�G��N|��ѵl�j��}u\.A�ұ�t  D��r�ϴTc0!1CY;lH��b�,�.-��MI�n��)��m	����b`z��%EG������
��@�Mm?q0�L3\���O�q�4#RC.�]2f+77�p��'�*82a�'��y���+8�L	1n[(ǜ�ʘ'T�y��Oza{b�G��O�j`yf\?I��Z}ۀy1 J^�3�*�`��?D�X��g%�M7!�*	������(q:R��5��+%���LB8yK����HJ(�x�HI�&ިj3>�C�%��:��}��'�� ��X�+����FP�u��n�	hΤ�1 �p�F�@�BA�mg&̒��-�I�io6"=� -��@���ۥ�Y�Ժ�"MU̓]T��&��a�@Y;r��� ���'�l��V;xU���G�-t�~5�ȓ<�H�Y�$��θhT�Hc���ܭU��{7㔻&�5ϓ��O��5�w�p�Q��A�6��p�дq���c�'Mb�Jb"�?4,|[��T�Ė�B۴|	�������븐�֍��:��ʓ�<ړv�b���	�+�̅��ԬY��I��!�+3g��Z��#"�/��웠�R;��
��C)b�!��ߞI�.����B�j�@V$N�g��9q6��=�qO�9��ܮ$�NQ��B�:=H�ę�Yo��"�>�8��=��!��C�,��B�I�"SpmqRꖻpf]!��B0U��(4	�&Ge��k�%R,Qٴ�(����;Q�p遆f@/j��0⣆�����}���ZԊ@��4�l�?r
���'��g@�+  �1�%�,x'��XІ8ғ_L<[$�� )ʦ� 7�-	�DI��4��)�6�47t��#�#oC��9eV�wt�����_����m��s�f�x3H׬�p>i����$�B,��
XY���ly��c�4Q*dm.+3�jv Q�И���Ô$z�q���/�1H��E��y�H	�h�	��"o��I[�lM�\��@�0���<�O^.ؑ��ɺN9�n�1���A��(aZHu s��J&aR�Ըu�LFB���hz��9Zr��BP�<1��I,fh�ۂQ�S������D�'e��16�ؽq�����f�(%� �����0#w��HFjF����z�LZ�<���g��9ER�)�)�,�`�� F0���W,U�B�|���� ��6F�8Cr�s����d�1,�� .�t��dj	�X���	� c�(�B�#��K�r �f�:Gn!��H�z!7D��~Ԧ�@D.�8-��0��02��Y�C�>%?M���L�1�`�]�d��WŜ=z�>=b��Z�B�I�$st�����
�Q�C�Ơ~��Z�X5��ɫ4` y�hX�o��e��T���\�'�ԭ�a$
?r�.a@^. Ҡ�
�c���1�!zpr �M�#j��b3�ح&ܒ�� �<���Pq$�v��h�%Y���>y�I���<z���r�蓰OU~�d{m>��#i�jo �IE��?�W�R;=���LLe��#�]��܋v�܈��C�* �[�+v�|H���M�>���>r1bS��OȄj`��p��ȅhd��QS�!��lcd@��E?B�����'2�PQ�) *R�	zCH�g�P=���NqF�be���wdxr� �<��o��D{"�'$C�\�n� X�K��0<�$(	�e�|rw�
`ނ�ǘ�U�� ��IJ�f!Pe.��-���Z!� Y�Ն�����`���ۖp��	���S'@|d�'aBP$	� ��P2HM<,��t��iC-@F�	&MI�.fp'�U=n�!�D���P}���V��i�Κ�|AdI���,Pj�'V�	�𙟰� ��
V>(5��9s3rx�E�6D��s"�1H��u�c1g�X��T�Tg�Z���J�&q"�' �ˀdE$uf�hT���v�	ӓz3P5��ӥ%�����M�,���`B�N�v��J�����Н��<�&��&KB�0�������	�<���Q���bR*2$�|"�$�9��]�ա�2z��hH��f�<Y����*�e)�^(���V�B��QJD�4L���O��,���	 y,��y"͞25��s1%	,Mh�B�	+ �>upCr՘�!� Ieވ "3�C'g�8�#S��>"��uS�8,O�\��N!+�:�j���h�hz&�'�i脢*dj��P�������LtA�%d]B.L�@�!��$�nhz�
O� �@x�k�=A4�M��&�9�F����>���]{�:�(#�1Ho|L�#�VѦ�>٫ӎ�"�F����F�8��f) D�D@���&2@Z �?���D$$L^m��(�E� �m��?�>�������f���;b�xèE�w��)�	m�(��q�q����a�d����] t�`����~"�ǽm�I�� �?aa	Ր�(O�5đ)2����c$�+-��6�'&��I����`.���cʸC�DbhK
��-�uDL� 5������/a�7M��E1���������a�)]���S�I�6nO�y)�س�l����	��l��'�>���8����E��q[Dm:B9��j�̼Yc+U�Y\^�ŉ���r�"�ݹq>B������|*�۟���u"W j�ܜAb֬����˃P��(c��w��ز��$$� ��Ӷa�>b R1
DF� 戩*O��
A 91$�'��'r�l����b�p��g\+Mڒ�XS��R���c�!=�I+Osꑒ��>IBj]	6JX�ׇ��4�����ϭ^!���+�-lmnJdm_�k����J�^:B݀V旣�0=���Z�l�҄ˎ�`�R�y��H=���)O�H��$f�佰ROU?4��S��S6���T�N%"�D)���P9>C�	�*Ġ �b�$@�>y3��n�:P)$J(t�6i ��C�wc��֧���?qAЉZj���B�J�*��9�J��R,$���'���R �����@�1s�,b�B�@�뎜%����wp0��:��-�\w�0�8g�Ddb�xz@W-I���2C�$���Ï2�IMKġ��2�S�d��Ǉ��w�t�ؔW5G��X��8!rn����IpTq ����S��'LO��9Q���_�i��<^�a�ܝ�Xb��A�ͿSUH��ɸ6p@��g�u���W$jB�c���0��u��ჵq!��P��]3���:G�0�PsO�R���@�G�B>�q`S+uwԱ*A�-����	�?^�>��uML~M��
�e�9��`��I�e��Y�d�<�� �CI �3peIS��"5J;m�r�2��G� �0�#T��Os]��D	b��Q�EW0NΠY�4�T�/Y�O8�p�JQd��L$��M;I����k�RV�H��Κj%^%`���1�Z���׆d����i�b�C'��:.��ؔD�?� ��G�i:\G�E ����|�q���K�!��_�~��#�"�zK ɲ4��$P�^h��cHb�)ڧ!�:}sN�(>���C��[\����O� b��U�K~�CA�v��&���!��mB ��I0v�nk��)p�ver�H�Z/6��dC6Ynu�ȟ�z:�{��T�.�u�EMS�P���uÆ,)��4aj�q*$�۳5�x��0S�O6h�&ɋ�{��lyuD�6�@��"Oց�Ł��:���+��ΔA��u��"O��Hq�֛���B(�\��ؤ"O�]@@�@H����<Tw�L�T"O,`Q�"ȅD�pE���!6�rh�U"OV�[V����MV��Y�v"O�EEC8M!f�@)K��Ȳs"O�q2���:��55 Zm�H�"O�LJ�m�=}TT��3��xB"O�XIC��#W�ޝ�PnW
x�F� t"O� ���"abt�lS�'���ڷ"O�IPǃ��z�4��-V�1��ʗ"O�0�m
$'����t�V���(�"O݀�eێD���0k�����"Od�`.�?8��4�=dm�;"ON�ЮՁB(x�#L�)qE�c�"O&HxAI�d����(Ӎq�*�1�"O蔈�Wl"&`�H� U�.��G"O��j"�G���Y7��h���[7"O��R5oĩ*���MӉ*�ơp�"O�p��	�op^�P���
��ձ�"OR z��	�k�2�4�̸M���P3"O�"�[�1�f	l<N��4#�"O���/-r�)���B%pP� �"O�TfN :��.��tX�T�"Ot �G_�h�0P@5��X^ܨ�7"OFL*Umm0ii�I]�}(����"O���.ab��vb_�`"�[g"O� @ՠ��C<�6\r�gP�%B\)�"O�H��"l޽sa��jͣ "O"�Q��:��J�%��f� R-7D�8� L�,�Z�ʀ�Բ>�)@��2D�l�%c h@d�z�萁0g2D����-J��hوf��6B��PJ2D�|3��)����☛rn�t��0D�Hn�� ����̘�
�J,J#�$D���OR����ee��[]9W�$D��9�d�N@N���#[ ln�-c��$D��E�G1u�i;-��dL D���A!DP�*č[�Hq��aU D��@���+NX��U�Yum�h�s�8D�l��Ls+�qJ���&v�^`2U� D�p��8}a��QKR�z����?D�x��"�#�՘oΘ{�A�Ԯ<D�L['H�"WF��V&�9;N�y�1�0D�����Z�Z���PŊ�%6��A�C1D��х�������ʊN�R��N3D��5��C���z�쉾Z�B��'3D�����Û���C��@̐�.1D��#ŨW�s��t{E�GF��&�)D�H蓢B�\�h)���4΄q�-&D���VC�;'������h�vX�'�����K%�"ؙ��@�U���'�a����#�d����8N1�
�'֜!�ٓL�(�P�
9N��'^�J����T<`���9���'�@���p�.e�w��@g��@�'Eּr�@�g�R� 뜛29&qK�'!��R ş%\���xK	%P0Q�'��S�-=��*b�ק,�R�y
�'�ZpɆ��|�4:�HG�{5B��	�'b���V'��Ȝ�:��M}�s�'��Eq��|����i�{@�'�^�*�QS f�X��Q4q�Ƞ�
�'�����9
���zc��c<8|@	�'\Y'�H�e�&Q��&QE	�'�<�'	٘)��q�Aא4C�)��'�x5�@c��xF����L�$%.@�H
�'�<8#�ˈ-nc��r�l+=8�
�'�����Ί!Q��;cKOK>��	�'}5Jw�O(k��<Qr.Ԧ{�
�	��x"��� �ҡZ��8�̭�"B��yr�˙�`��!�^�<N8�Q7G�&�yҥcM:�jЅ� hmq��Q��y��	�T��A�/O��𩒢ڪ�yr#�,C��QVI��B�D���>�ybC�p�3�e)x�FB�,�y�N�5V �cb��I&�(&��y�R�/�t�`+�i�ݸ`(��y� ��*er�ɔ�_,��+=�y"��35���ò�G=[\S$ǚ7�y�C�|�b���N�$��h�*Ԟ�y� �s!�l9$F�g&yst�]&�y"CX�	��)�Ӈz��, kY��y"&i��t ��X�jw�(��(֜�y2i>ą�{�Tce`ԑ]6���'�hCn�#�����cޕT*J��	�'r:9Zr/
p����Z9�^��
�'��p*�ɚ��yi��V��y�'&���OL�jT��2�o�@$��'qX����M�T3b�ԝ�f��'����&O2F�a�遠j�
���� ��`a��Z$H�0N� 1���Q"O�}��!�f]v�q�MD8*��@"O4�1�V�oj����1a�p�c"O�����=0�� ic)�#�"O��x�O�3��@gj=
��c"Ov�CtgK&&l(����<O_X�"O\�a��?P�T��׌�ll4�bQ"O@L�0�ݥF2��d���SS�t""O�$���ހ�N30{F4	��̼�yR�"��݃G�1$�� �,H��HO��=�OR�p����.�¤i���l�����'_�\&K�uդ��3d���h�'��<�qE�y���"�K�`<H�'�����٨]�d�=03l�8	�'~ؙ'��/�|�C���-���!�'�&ȃ�,ޮaq(� ��.1�8��'�,x��$�0$��0���٩(d��'�B�:��J5/�����G��ys�'��|"6&�$ODB	3@A��h�r�'"pQ�c��O�D��b ��Bm:
�'9�u��HI���k��,:@q�'����O]�L��{�nT0J��Y	�'/���FD�-�A�)3>����![�����'{����E%2`��ȓ99`�q��]�4��,���!EG�}��+F�B�(�, ���q&�Hs� �ȓ1�jm"vd@=T�,* 
,Q�`���K�"�.ǬC�V�$�����"O0y9t�V�pI�yr'��!Z��R"O��w.I2U
�*���^���"O�@*���q��)E���H ��"O��@'&U���q�P�j�f���"O"�B�aM!d��D�i�l�F"O��q�g��Y��C��w� y��"O��YDMH�py���M�����"O�ۤD4��h�周u����"O��!'��9���!m�` 
�"O��Hkɽ �y�f�5uQKr"O����Bm�T� E�3w\	��"O� ��
X;�MȓD�b$���"Ox��#mO3y��p�E�BgG�8�"O�P�"	�4!�tl2��[3I�497"Obl��H_06��q��=͢���"OV�1OP	p��x�VD�4W�4`$"O4�1���4�� 	�;MU�1�d"Or��-͊�t��"2I����@"O"�S�gк�J�y w��XQF"O���GX�y��%��Z!n�I���`�O�^�06
 2H_��k�O1S��<�'��q	0��,vw~H�a�ހ�4��'c��M��-��0����	)x�1���'�!#�GP�z�]�Z�4���B�<� �A�U�Z-↥�3n��w Ju�<�Ε/=���p�$K�|�hUno�<��n��m�����!":҈����v�'Uў�'N> Yեݞ5d��ѴI�V�Є��c��=PJE�!�q��ɸy��5��G�L���Ɣ�I?�1�R%ò�(���[Cn�*�����U��
L/�rĄ�Ub��+q�O=S{؉���]��(�ȓ ~ W�:9)`��a�N�1=@��ȓ"?t�y�I�I908L�86@\�ȓ��yX���I�i� e۔"���j���8anF�,��ۣ̎����S�? THԧ��o4ȡP�$��B�"OB� ףY"cR��[����
��Z�"O�ѻ��
1�>D@&"ϞH�J��b"Oj%�A <Kb���_	vh�=�"O�Ir6�	�IX6���e�\]�"OlQ����<r��@�Зf����"O
�3B�X
E�f�S�2�v�"OZ��@��}g��r�T�+�60�%"O2�x1
Q�^(��р@����V"Oz�Ɗ�x��,J�'�QqU"O��Y�U�U �q�D��./lT�b"Ox��N��p�5c��$��B�"OH�*�@̦p=�ܛ C����(�"O^���͇\�����ǎ4#���!�"Oƙr�#�8�<���T�d����"O�`z���|��12U��7w�u�v"O��x!
��\��D:#SQ"O*liׯI
gFL���țk�&Xi�"O୲CF;1����"��.�
���"Oh��é��Y
t`)��1gtAPs"O�� �7��rV��j�W"Ob�8`��1���B ��kK����"OrT�]"+�� �T�i�~tiF"OrqPe�H�#�^X���w�а+�"O�g��0����+���� P"O6i2q@��5�9H@U�$���)'"O�!��*��,�g�H����b�"O��I�O��^�|����T-{��=B�"O�D�Ƨ�'z��-��6V�\k�"O4��A.
��-��%7b���"OQ1an �8�`
�+1J��"OH��AgĖk6���w�aN��q�"OD�#̄N�4;0j0L��Q&"O��D�%h4��r1h��1��"O��*�a��[q��3��	!+X;�"O�D�fO�jUh��U�, y�$"O줪 ň8����cZ�:�`)�R"O����C'`�h�#�%
����`"O,�1�N�5x�0�!��۾K����"Op�s'(^U�3�
ͬ4�
�;�"O�-�7(�"7u(�& N����"O�᱕��!H>Y
A��3W�U�"O��y�.<�n�LS�h�� yG"O����M8 ��Z2˒�8X��"O4 ��H4E5 Y�@��-C����"O��q&�-|=Za{v/",�x�"O�̱��.K�ŁQ�1 a��"OZ��EM��(� ,�B���W"O�H��fΝM*�"� -b��X2"O����"�%(����p��E"Ov����ۂ�3���\�#2"O �dD@.l���AFm�@`�f"O�`q��	[7~���@��6��Ы"O``J��I�va�Q�M;*�j�ä"O����ٯ^+��j�gB7/Č��"O�9#���
�^�)q�$DЀMs"O(� �!ϒI���r���z� -�"O�1�@�7 +�m�di���y3"O�}T�Mа��RHF�h8C�"O�x�5��)�����b���"OH��oE�w1�a�ǈ�z�Ԝ��"OL����T�i�N�b2��31|��QE"O��q�i�!�����݉#�0�@W"O�4 ���;@QH�G��j��p�"O� �m+uZ��M����oef��"Ol��!��<5Qb�␄�"j[Ÿ�"O Y@㈀I����DM�!P��"O�9Hr���c�'I�N8��a"O��f �H�ܵ+R` #(ȭ�F"O�4Y��s�2��#AI	"���f"O�Թ���=c���Y����"4,�"ON�[1�Z_zT�,�"2�q"�"O�-z0��A�}���:rP"O��6�٢���>�;�"O�� N[LLI�q�T	Ut��Q"O^5e�Nj�����M\�/*Le"c"O��A4m�+�~{�\ɀ"O�l�e�ڤF�8�yw�S&g�P�"O�H����	'��+��͈Q*���"O�m+ �L��r�Y�|�
t�s"O��$��4�"�	�/��=AVY��"O�!	���m-���
�H	L��"O"m�Wފ<:pq"Wi��EтW"O�rV�H��)�JTk��M8 "O^1��Y�v���L	�v��A"O��P��r�z��B:�b�Ru"OF\x�C��HZ*ܠ�)ѬF8D��"O6CI�y���*W(�,:i�p"OJ��	6<�p�a_;��A�"OZqku$�<#Pe��!� z7<Y�"O��Q�H�|��|1��Z�,��"O8A#��Dh�h��/�7\��$"Oj�2*��	ɺ�PƎߢS f��"ON�����T������Q�o���!"O*T3��a�1u/��$�Y�"O�Z�įUV��*D���0]�"O�M"u�5(�� 4��Uո�"O���3��#w��#�n��)�Xl�"O��'�QD�x@mI�8�,��s"O�ybF(�(�
`+ژOȨy��$%D��[�o\�d��ZF�W�[��E�Ќ8D�0@��' "ֈ��'�	Ŋ0� D����_�}�S�p*�
�?D�x;��PCE�M)�G# 3���;D��)4h�F��L;�$�%%���s,:D��!�K�A��i���Gh��p�4D��jB�W=Yds�ȩi��My�2D���E��P������qN�eC�/2D��� � "$ J](P�y�~�i�,/D��R#ř"}l����B$~it�"�.D��XvhN*,.��Á��f�F�r�!0D��"���;���s�Ɋ � I���3D�`r�� =���cv)H6V����d0D���q�O�H`��DoS� ���/D��ZU.�1@�|� �Ȣ]y�\sq.(D�h[�F��Yҵj�h�S%�'D��y�e�C��\�g�T=�=�v�!D�D���ߜW9b�j�#�8 �Yڔ	?D�ԣS͔T�J	��ϑ�r����c=D�p(���'TVl�����20�t-pө?D�\vF�FxMa��E!R�45K*?D�lcc���lqR�PB'���[�D;D��a��M�_��H��_*I��|#&�:D��z`O�}f�"̟6���ˢo7D��ʅ��YF|�����	`��5D�1��Ȕx(�ڟ�΄q�i4D��(Q�\�j���e�{�0ʅ/'D���#��`��`��Gx�q�1�#D�� �uѷgA:R�8%��lБ8��(@�"O��z���|N�!�e��24XR�"O��C�dǗd��F�Z�_b�a�"Ohp��L�PȰ� L�G�
�S$"OZ1�hE.?X����"���P�"O4��e-�8�0k�&(�N�KU"O�QIs��g��5��K�~�@��P"Oh�aЎ�{�|�˓�%,f�� "O\HJa�T���I��*A[��(B"O�9y�� /�l�|P��o���y2o��!u�;��ܨO 0�O��y�U�Fݖ���@��Ze�fS3�y2�G�{Z�eˌ.i�1�D��y�!��fp�h�3��2r�Z7���y�k!Oπ�
�E0V�\顶C��y�����i�/
#8����u�ǎ�y��;m��5K���z�����y�iR#|j���`��%z�� S�$�y���/q�0�+��,�ubҭT��y2�^��pk��"���5K^8�yb��;8px�4�O��43c׀�yB���"��G�8}�"�:"٠�y"M�"	1�1 �n��ph�G�2�yr H�H�xi���5��)����&�y�e�v
zD�� ���D���y�-2P�(јg�����A�6�y2�1N�Q+�(�v�T���'�y"��K��1��l��|�%���yr�G7��Y��H�]��C��,V��PJ3mHai��x5�N�d&�C�I&-��is�ѯ1��$����#��C��1p��ZDo\�S�X����֩3}�C�ɡ"��8aK^P�|��٢�zC�I"s�ԓ��U�ED�u����V_bC�I�8�|��`�Ǆ%z��,<`C�	�(���P�!K�T�jS�ˡ�PC�Ia���"â<j�x4g�7"x�C�Ɋ�`RD�^(`	�
թhٲC䉘*הȰ�-J3���h�'S�ke|C�ID��!��A�	c��p�,F7�@C�	�,�(l�,F���s�D�"C�6&��$L>/)fA�񇆬2�B�	�cƬ���.��3�Fd�"B䉝z���9�*�)*W���CD�%��C��+/ڼ@ҋP�q��;�FC�FnB��<#r�쉐�ز���Ia��}�TB�	'R�8pf�'~�A���g vC��/�����%.�#U�x�r�:D���bƜ"���[3��kS���7D�0AF�E8<��d"��<QڱzF-4D���'�R�M��;�`�Y�Ɓs�e.D�T���+s�R��P�65�i�f�&D�DٶA��5x��BckɷZ�d����"D��S%�yj,ݫ�
�4ْL"D� �)�}��-0�'���{� ?D���D��7�,XZeН:���3��2D�d;D���s���ƍ�8)��r��1D�<��),��{��N�Ovx"�0D�Tb�Nǰ|4�	����ewxx��/D�� �1-�QE�ަ^�(�3��;D�#熋S���;�-ЮyC� �i$D����Rvȹ�PmX�l��UF"T�D*3B�9n�2)#���;��1�&"O�)k����zG�j )�F�vkG"O� 6��Յ�,c���$գ3�=
�"O� rS�>?� ��7�2�\$��"OF����ܕ70��#�C!�%["O�����(
��9b��$VD|�a"O|�#s`@$F4TVB��r]�}�"O�<�� ��b6��cZ�D>F�P�"O��sHK	uz)q����[��0�"O�$�&mY-�>��Kͅb5�tH"O�ٓҦ�(ڂ��J�L�|%�s"O�,[AOߘXr�3	�
^���"Oj��d��;�X��Jey��"OF�z���7��8*����԰d�0"O�]9���g^�0�%_�#� �1"O��Q0"X�2%<Ј�M�=��D"O�z��NM	�܀'-JX�i�"Ol1���,�=��"4Oe��9�b���XF�PeB[�.�,�ȓ%��`6� .%c���?+��h��?9�T�K�c��`�f������ȓ �p�e؝3����`�7�%��L��Urg���Z9��*�6���k��cE��:p�������e*D��ɐ4]���tO<P=����-&D��thͬn�d�+]&+��sTG"ړ���*§ �����ԓ�=ے���_Ghh�ȓ�*��RB�;�n����;5L��Z-��Y�Ā����с��8��+I0ȹ`%}��$��86<�ȓv�\���?+����q�˄p����P�
��ƅA���!��S?!����M]0�%���Vg
8���K�y���ȓ5��9{�.ԏa��|Jc&�h���ȓȑX-@�%�d���C4{��ՇȓFPu�U+^�o��@h�-\R�!�ȓ�r`1�K��d�v�ѯڥQl��ȓ5=��@�F^�L��Pd�7h���K�� ��E�X͈��)�4o r܅�(�z�Y�4o���aB<;3xa�?��N"L�f���[\�tA�g�by�ȓF��a1!��V���[ E�T����u�f���NUij�At��$a�怇ȓO�TE���?W$�t�&C:�>�ȓ'��i׈J�R�b��x��T��۠��cʘm��$/X�,Y|��)O���d����m��
_�+�Ԁa`�ڼk)!�P�e+Bu�r-^�� �H0�>�!��M&b�bAڂ@�>X}��z�I�!/�!�D
�A1��s�eۇ�L���^-'�!��@�`�����j�;S���(����6R!�_�v͑ӅG����#xȆʓ)ciSf�^
�Ű��&lB�	D���h����vp��i��`0���0?ٗ�u��M��m�3�*�����o�<Y�Ȕ:U�&43CksJd���`�<قѤc����A>^�`I�r�<�%�H(���K�$ж���5#@m�< m5rZ6�PU�6��Dذ�q�<Y7�5o��[���K���aJo�<a��؈`ZPp�`0\��r���i�<qd�g�c�k�^}�h�o�[�<��W�sT�SB�\����	D!�Z�<��<��8���j$,=%d�Z�<��!P)DV+0�P|P�C���!��@%"p���%��	|.9eݶ!�� ���Ԋ.�<|��8gly*�"OPi��$T�[���O��~��_�����=p� �zC�N���s�f_8�"B�	AF\���Y<�(�%�-D��C�	�OO<	���՛F�F�rq�,�C�	!8e1!˓�D�I�˕�+n�B�I�.!�$bB�N�T�9w/�,e�|B�I��p5¦JY�Ax%���J:C:B��\X��#bL?t��	��=3Q�C��%H�zɒ�_$l�<xe#P	-վB�ɁUi�H@S���#V渠d,#[XB��<|�n�(��|G�hIs% 0FPB�>�΀��� ?�n��ïC`�C䉜C�����"���w�3nC�IG�	�F��R��T҅���K��B�I�E�R�V�}_DY2h4:�C��9?h�4�2�
(���H�nC��:e��i�J��&N�����R1�~B䉟,���QKF)I>�
��2�C�I	#u�kteV�K�Tu ��k�B��!G�5�r�Ĥ6�f��-��PA��� B��sd��%I.����C=_�!�N�s�&�.Y`��e�!T��O���dB1�ְr1Æ64ڴ ��V��!�d$Qbf�2��
s� �R"	˪%G!���7�j�/%(��0�&�o��q�'{�$ë�>E������Y�z�v`	�'��9X�c�*(@Iʤ��"ۮ���'�HH���J)(���S���|YxO>1�r�I>L�<	�Ǆ��zeX@%�iςB��V�D�pE���y�n���n�XB�	r-P��ب�V�U��C30B�I54�çX��2���W"�C��P9�ؒ	Ɂ7p��g�A&�C�	3v0�K����Z�8"c�Ӆ%��B��
|'fD���+~��7 ��+�B�38 ���ݺ�>��c&"��B�ɨ=��\�0��6 �2\���Ԟ
�B�I3iV�Q���8tt�
�ֺHB�I�GI6�3����"��;�DB�	�'�v��S�Ηq(�Ape�b86B�I�y�0�!�H�j��rL�wJ����h�x
䣞�M��=0�� w��败<�	X�'m�Ɉ)�����Y�Y��EI��C�	�^�&X0���^��X��aA��tC�	 ��QBg�t����b%�V��C�	<tvi�E�\�{��ؒ@e]
��C�I7�8��R�$fa���E���[�FC�&d��@u	�/uL)���8C��8����(��4�pB
�Q'C�IK��kvA��Gd�pR�����B�]u�M�� �7:-)���!�C�I>l����-�X�$\6q�C�I5E�R<9��%	�m:����c_�B�I1�8���/ƞ)-�!!�̋��B�|�|t���O��)H�	�Zl�B�ɖ<�n)�a��t�D���]��ʓ�hO>a�)��Bi�Hڄ����R�v���I�θ P�!W!��Ee�<K^���#�f4xV� +(j8�V�B�qֱ��/ ���_4]3H,cZH���t��ɑ���z�d�+d��>	�J=��h�J�[�˟�i;�*$K�fЅ�e����dվd�4�	g勗qc�E+��� "��7AP2|�.e��
�yB�z�U��G{��C�-[��I���:^�ΨU䁘q�!�Ē/��}Q��S�;��B�!O��!��ĉ!Fu�ҦO:_����dOX��!�䁀}��Ӡ/i��m�L��l�!�Z#ưH��U1T=2�3�j>?�!�dI8�`Iʡ��q'j���)DA�!���*.�Fƈ�9K&t ����u��'��O?�"f�!^��B��CK�*���E^U�<�v��PP�A�Rlހ�n��G�H�<�m�2R0��c��X�H.J��QF�A�<Y���F��Xr����}w�r����<QV�_7@`����%���i��}�<���߀G�Rа���af���z�<�R"X1kc���$�
s��9Q�+\�<G'#�^�;� Z�$ �����p�<��ObA�&S4}֬�j�<q����? �tCNƌy�@3�d����<	�W�&��d���Bz�h��[k�<���׵/D�=q�eJ�HƖ	x��D^�<e(�|��1�$�n�\��Y�<�v�X�H��Mi���	k����%�J�<��'��P����ՠ,wc\D[�a�<9��Td�����\���_�<��&
Q��a���M:�����[��8�I��،�c���xy��%��@����t��CQ^L	�u��0����ȓ_�9#L��:�@q�5ǂ��Z���<X�+@�F��PJ���ȓ#z�Y` ��s��ճCL8 �ȓN��-�ҩ�7�8 ź�G�z�<)q�X�6�*| `������)Ym�E���O����́*[Z9q��?�r�'�T��)J�=����>�0�'���HG2/���ρ5ogL����O0uy�jۖ$���hui��f�>�� �'���|\>c�擪lM�@�G^�|bOG%�6��k�P�Y��Ě@A�!"��j=�ȓb����,=Z֘����	->���ȓIz�1Z� D�Z4B�z�E�C.�u����=��苽UbH�V(�(h���ȓR� ���;+�8Hـ��gO�I�ȓ_�(�hU*�7�‐�E,!?�Gb�'w>	�f��!�EH4e��zhI�� !D� �7$�ř�EL�t�bI�* D�,y0�dD�U U��v�PQBe=4��!4oܩr�@A�g�g[Hx
��x��?!����ɢf�$9��[�n�'"Of(��UjX+��ւ$
�m{B"OԜif��E��tP�	!Q"O��7�	Vp�BbG�{�b`�"O�P+GFB(�vՃ�Il�~ ��"O��3B�T!S$}�#��l�֌�r"O>�ʧc�!��U1�
�F����"Oʉy'�:@�1� GՓr�l���"O�E0��V��r�eШ
�@qb�'w��xbOG�t:sB׳>P�����(D�x:C�2���C� ��%�,�E	%D���w����}�eӯi6J�P�=D�4S�E]s�pA 5j�>gB���E&D�����]�0�
��c�z�ڱRǥ<I��哾,P��#��	$�.��D\P~B�	�
�|�sB�^]40c#NJ�FodB�	I�,K���.9wLa �K� �C�)� ִ�QŔ�m�ĵ9A�ǡ!/�y("O�*�@�n6xKb'Q�}v|�u"O���J6O%`��.G��""O<�P@��
u� h�K���p��P�|��)Z�'GD�K�Γ��v��㬚7N��Ax�'�ґ��G4!���nY�K�J}��'nΑ��O�'ؔ����=�a�'��Y�B��ɖ�]>�3	�'�b�IĂ�l�,���2Z�E��'V��s�䍽_��Y�+Y�3�` ��'�z�*
��1j��~����'ebX�6��z߬�Bb	�~`�"Oʀ��7u����F��sϤ��P"OB��cE��jR�7�@q� "O�)�%k���F �Q��o΀�#�"O�����=
Vv��ǡT�Y��i"O��S�&L�r�B!BL���"O	�� ބ{�]�PAI�-%�!�"O6��4��F^��¡��(-��"O�iK��H>y�BJ�ϑ"$t�"O�X�잠jǆ�A�^�}{�"O4l�~a���8>ձ�oǎF!򄎍g�|:�˓I mRb 
3	;!�dD,12�Y�.E%&� X���U(5!�d%�m�K�6��5�7�̓	!�I�W�|�ݴA�R�Z��_�7R!�Q'Q�̡a��ZXP��u��/S:!��E�I,��R(�c~к��^�>�!��>\&I&�N�敱���j�!�D΄ea6y�I׾R��C��5�!�$O!L�9:0j�kM��`#[�y��y���%U~0Z���N�bp���2�B�I�A��`����SJ=QR >
3PB�I)xt�g�_X*� !�P�'�JB�ɜM��H��WUu��2�-H-/!�S�0���#����bQ-�t�!�d	�9�X����D��!�w�� fA!�d�>�Y��GH�d��IԌ	L,!�D�	x� �Ǒ)P�a����E��h�D�.r�<�w�];"�*l�pc2D��ZF�A�,:���"<�����2D���SB"���l�Ct���#�:D��(׀8g�B�p��V7F�V�
:D� q`⊩Q�zU����@%��6D�d�g�ņ1H�8�0
.249�cA"<O"<�C�֌C3~��֩�z��`#�GV�	o���O=lqaСՄ'a�@�@�]�"��	�'Ͱq*f�ʐ'b�si��]�� (�'jr ��萧~�"�C��]ݖu��'O������â�S�'�8�r�'O��z��)>��s�
�h�I�'dwm�����"�b�c�'�$)�GI_�}�� $`��bd��'�%��,���PS��8�8�'��q��+f�ЃglO=kL���O�Z �'¢�ZGG�0��4�@��uפ�r�'��bG������Lܑ`p�uc
�'����.��R�U���Z�\���'���;c�1=�8�k���YkRE
	�''ĭ�'��:p�p���1"���"O¹�� �����(�h��"O>a� (� usr11�08���1���8LO�܉�B�'q��׭O��j�"O��@D��w��Q����"�z�"O� "�S�I�mQ��	���RR�"O�����z���h��Ǚ&z��R"O�`k��ٿX��}�V-ϡʨ�0"O6l��#t�Q��m�8����"O�"��B�r���R18�����"O�-��	R6eZ�ʓ�ˆD.d�C"O��C,ܷ6,��c�ԴN>��#�"O�$k�M9Vtۦ*�\��"O��0Έ�r�;�� k��A�"O�9�tJ�g`�q�#�L����	}>��1��lt������>�Ќ��$9D�@[��ԆO!EŐ��A8?ɶF�j���ҝ!�:��չVL䁓�4D�\��Y$s����P�S'��q��%D�|ۢ���A���y��Ԍ(�r}{t�7D�� G(��2z�SӠ5'� �ӆ1D��`�b�,�FPq`D�m+DqS��0D��(�I�f���sl� %nF�3��"D���Ѧ�> 4ٺ��X3��%� �+��=�Ol(h��0��h��Q�	
��s7"O����^&�L��M�.�ة�w"O��ÃB�<I�IhUGȣB�*%��"O����!ȼ��,��.����"Of���"-yt����"Fj�_� ��ɂ`\}����}�Hy���D@��C�I�p���ؖ �B���f,�:H��C�	Z2���G+Kh�� R��A�Im�C�	#��b��=e����-�FC��&CR�"����6�@���	�d�NB�	Zh�0t��K�9�N�| RB�	�WKh4��̀��<|�%�ЁW:�B�I�b���aM �E����o����C�ɹU$~p��g�-;�}䚟"��C�ɋ5�a�b:"�5��Z�KO�C�	�H\���%U'P,HKZ�G)6B䉪AM�$�"n֥
��p��Y[�nB�	�J~�H�狚<�\z�B��fN&��'�I�@q�����M�@������z�C�	8<K4��&��(���^�W� C䉋<���%�{�B�1�NڍzOC�ɕGpL�
@�*C�\�JP�ׂ^�C�	�Js�u	t�D*
L�!3G��LݤC�	T�@�[������JʜS$�C�	J�H]sqk	�oz��v(G�Vr,C�G#.=����0 �R)��+�(c�&C�ɭr
̩�靂!e$��gC$�C�I.�`��0�82LO�Ae�B�ɛ(I:pDC?y;�M��LG.kw�B䉈w4v�Yա]�3MN�84��<��C�I�@���� �'J�6([ց�3
�xB�	3�Cԍ\'%����B�P�i�(��$+�ɜb�̸�g��F���P�͇sf���%�ɷ$2���ר_,���yKʉ�XB�Ih�0cw͑�y��u��ʮP;rC�I)5��� ̗�<H4Y����Y�HC�	�?��(�CKI�Vp�X��-aXtB�2��lV��n!� �g� �BB�I�MQ��x� Ěd�-ȡ���B�I;�t��r��*T�e@#��YBB�#Z#��� ��MMR0�VJWz7��ȓzB���A\6���IZ>��(�ȓF$��۱���h)e*������i��e d!�
mT�)��t$�y��{���y����K
��͛�Rժ��S�? lHˢD�,�� W&�}T"O�(�g��?**�ԁA��	�Z���"O�M�O��P.<a�$��@�P@��"O"��S�1t�hg.RU�q�"O&=1vHD3il���#�j��i��"O$(���E3�
0���/j�hH��"O��B#@�P�0�����b24j�"ObYqE "Z(t��T+&��("O�1p1�����TA�W(a�CW�HG{�򉄟e�~u+TmY�04���N7I!�E�D���E�P��2a.�}�!��>+��ٓ��E&p�T�A��^�N�!��(�6�0�@	ӘM:��֫(!�D�Ҙy�S��*ULT!��(N�!�E�r >�)n��d�D6�M(�!�D�<&����nɶL���b�"x��O����;��ʭB�� KaM��>�|D��}��K1�Ý<����gD�|�ȓ<2�`Cv�:��)F"�1r� t�ȓ��ihs��B#8��!%��e�p���d,B��3e�� "���)F����ȓ
}���$�A�HQ�U��LRS�>���zR���

�B�����Ćȓ|\� 0V˃�ĉ���'
z���	Y�? nY�+ҁ�:�y��E�I�ҕ�ȓlR(�Q"�2H�z$�"�ܝH��܄�qۺ�S B�2��5��N�:0��ȓYź�ce@��9� �G�D�wq ��ȓ.MkP��<"%��t�� F#���ȓ+��3�!�)<���B��K�����H~��K�5Ia�At�h)a�3�y��	���gG�e2"dȖO�����d2����
�lS4�b�H,Ò�C�"O����S8g��*�ቪsH�D��"O�T f�	}�^��5�G@�`"O$�i�C��t��d��9GA����"OJ�:U�D�>��z�,�H4�S	�'XD�`�E4;�҈Y�C�zQ�QQ	�'�$:&bБ~���s�H'm.��	�'��@�@V�P]9Uܨk�X��	�'Ȍ���Kâp��0�ԯ��Y:���'���S�D�_�: �� (�����'
��c�vr���Îٝ$(M��'c4h!F��]`bec���ND���'�,݂G�Y[~�M��F߾;�>H��'w^h�aC�qĜ��퇾<����'\�t��t�Rh"0'�"e�����'���ɲmҬ]7R����Ö��y��'LpD9���G`^� ��!����'���!�!+����O�}2���'������@�Vx�	Ѡ��sh@���'�	)ad�	��]C!�ޤr%Ƥ�'�����1[����CM��byT�0
�'���@O�l4b��ܞ%H���'q�i(Q ��ݞ��b��.� ��'�:e�%G):����ХF"�F���'��(�RL�"JB����Q���'(62�"��0�JiC���4`,
�B�)��,Y(`XfmQ�g�]� �B���<���ߟr^�[��Ѽ ��ˢ���!�Ĕ,,� �i
&]��j�� M�!�D%��P�MB��5���K�=!�,\���)Ą@/����f[~b!��/8o\��w�x3�)��GE	#U�O���-�D!�3� 6�yG�A'cR�{��Z�cvYS�'��' ў�OW�I�$��=5��e��B�1����O~���
$���Y�`O�n!��F�IL>�S�͉�6YRP��5���3Q�+D���V�J'FpP�)P�s=�8��3D��0rC�W���S0���|@JgE2D�,�P��I�m�@���\��#�2D�pw��B���"�s�p²C�O�C�I0����dD�aZ���D��:;ɂC�ɚ*��bj�.��̲�X�s��?���ɆK#�P����:��u��A�	�!�C,UA�(�+��5Y�,R�@�"~m!��H�eծ���z+�;��!�DIT��陁#nyԐ ��8�ў4��S�'���
B@3���޻V��C�I8Ơ�$��>�fD T'�.f�xC䉚����1�ɭ{MX�����1}�<�=a�'p�`��ρ@�Z�x��	g���w�Z�C���J[��A��J�
�Ї�<��}���W�D�l�@�N@(<������6&pK� ����PB
��'��U�?����~Z�h�#&�V#1�*i�R�*�[�'aax�Ăx�j��B�NY������y�΀:����eͦ\�20Z���y�HUlp� ��]+S<nt�fnH��y��N�3x`�k]!}�����B��y2�ȫtM��"M�!0��S�2�y��*�"��4��Ƣl(�M��yb��.3�`�q��
^>d�mC+�y�
�HoVq�a�� ��IAU�՝�y��G.YiBQ�r'A'w�������y�j�&���8Ďִk��![W��2�y`�M9X�!�ߕd`�;we��yR�/dŋpm�Ms��Cq'	�yr�K^����c�(2��}Cv����?��'&�{u�0Z���ZBHݰ&�.Y)���'U�8E�E5*����ъJ0���@�'s����>�HH�T�
o ���'8���2�K�5�L�� RA^�k�'�bD`�� �ẶK��B<
���'�Z�x�G?�T�����2��!9�'=�hXg�³c~��6A�4U�\]J�'ޙZEo�6ir�� wg�z�2m��'v��[��2Q���qF#P1~�.}��'���1ׂ_�/	���l�y��b��;����� �S�803jϩ(z9��"O�樑,v��,ie(�9Ng��� "O��a@%��f����ć[d0i�"O>
nŨ	w�%�CH�-��U�V"O|��sEz*P�'�(��"OjI�6*J�o�${f�H�y��"O�=�b�@=�-+���-8�py�"OҰ*HȮ$t�C(F@���J�]� ����Ic�h'�[6~��d�a*�j��C䉝Q��I���G�&L�]���H�M��C䉬2 y�|i�i��Ѳ �C�I*2�ĥI��J.�Vb+�)e���?i���S�OHTj�.B�	*��`��A]�UR�'?f�g�,eD Q�E(1!(�'iĜ�҂F+���1W��.)�-�	�'76������sY�H7�
*�J�'d�9h�3�� &��1AIb�'^9�*�<��;��N$��9��'K�	V���1<,c�IXSZ�a+O�=E�� 46��E�E�L;=���kfV��G{��	�:$���aU�/�����)M�'�ў$�<i㫕/]b�`��I��Ȣ�C�<�W���\�*T��?Jǜ-q%(Ue�<Q&M��� +"��FϚQ�Q	�_�<�`��.	��U��5�b\���R�<-M��S&�¾oq�5;�ԜR��ʓ�?����S�O���AJ�)H��{�*�c��y�
�'����'�x��-zd
a��E��'�\R�],O-^P�#ϜiJ�#
�'Hdp!�hˉaJ6%#��G�.���'\r (F�ƨ.���P�D�����!�'!8pS�HA�Ex4�w��x����'6��A�NM�Xþ)�GҿoL���'_����-g��֦�� ���'Bx��u���2�"
��"�I[�O�H�[׭B1u�L`�%���[�"O�y�$���L�RT)S"���b�e"OR�rΘ;<��̐�o
(��p��"O�\*��K�>b ZNʈ>�\!�2"O�#�ꊕ��mA&�Ѧmˌ��"O^�z�21���4Y,m�D$Y&"OR=H#J��^��䡆�ʎ`I�̀v"O>l��Ǝ6N=��Ҷ�
�g��"O��	3���<�N�P�D;�����"Or4���׬`���b��7K�h�x�"O����ͬ$�J 1�d��UX��"O�p3���;=�(}���9_�=�"O�T���ʆ)l��{q�B+�g�!��u�*@�e��k,�xAm�>c!�Z�b�c�
4I\���e�Ǭ_v!�Ā�_��h�D�8�V9sD��<t!��^ oDlYT�j�.�z	�?7�!���-�h�ѥީ/��|!DH�S�!���O��mIb��6E��H�֍�E֡�$�	f���ԫT52��XAV"���d6�O:9huEiGT��WD�&R�|�OrdS0�[:cD����g��G6�`�H�<�ST���T�'.��a�й=�"!��hP^�`�gI�U���6��17H�ل�G8�m�U�@W�����e���j ��:XL�IE��D�1qbˋ+qތp�ȓq�,�q���l�Z��-�^��ȓ�"�{�Ù�a �8tJ(_�dȄȓ6Ϻ4h�kP��Srj��\Q�̄�f����(3;���F�
>�-��C.�"7�Z� F@%)Q&��a:b���4��b�:a�fͨ7F�z5R���<H�@�!2�T�i&-;����=�9�LC*^V(	֥F�5�����LP�5���zN��< �QA��=D��G'	��@@� ��E}9qƌ=D�����T�`�fL�:�9Y��=D�,�+�n�����4r���a'D��
��P�0Od��*y��a��%D��	��'�~5���H��	���6D�TkW�֖KѪeI�I��n��A�0$(�d8�S�'Gn���V*y� ���(@.P��i�ȓN�B@K2��'>�����Im����<�<%�E�q����"�[!�ȓ9���6d�p0BE Z�h֡�ȓnv�+��g�6��B�0�D�ȓhg�$�쒲~���D36�$x�ȓ$���"Ʋ9nZl���/-�����S�? �Eh�ˍ	�L�9%�nQ�$"OL9���V�+a�%cC�E�h�Ly�"O�x�B�9|��� �o��R刬�A"O��pA�����JD�9R��̣U"O�@)�ヂ*�v<pb�v��Dk%"O|���J��0G����M�2�leH�"O>�+FdS�U_(Ȉq��O�t9�e"OB�ɥ�݌)3r���\<3�d1�B"Odu����1is�d����P�����"O��֭��	;ڹ�ŁR,ib��'"Oh�˗͙�K���'�QdT�@�w"O*PT�dw�\��5TL5h�"O�ؘ�� �zNp|a��õG=,L�!"O����.��Cnm� �9pTv�y�X�LD{�򩃼J��!;NŨ%�����cHD�!�ְ%�\��  ))�"5�#��]�!�S ��ͻ���1v�$��ᆮ}�!�'� 	���J=`e&@HѠZ�!�+o. ��0d[�,�u)"J�!�	j�4�c�.A] ϒ'�!��5f��H8���d��+�HBv�'2ў�>`P"�1m �M ���r���d�,D�d�'�"3ΐ���-�2H`�8D���F
,e�	9�Ϻ��õa7D���r-żM*=h�*�-`��=��B4D��Y�#�y#���2�!��Q��4D��RG�G�P���b
�a$)��2D��������kb��ZА4S�0D��a@�V��6�c!��$=Lȼ*6'9D���
�>f���k3*J���&<D�HYtY�1>0��CC�8h{pn=D�t�0L��90�M���P�>�7�<D�81"�%�%hק�15�xPcFM;D����I�k��8�2AѴe2쪁F8D��Y�ט;�]�,9��&BmM!�d:S?���U�N�]��S Eǀ@!�D��/t����|>���.c4!� vp�(�K�P682CN<I�!�DZ�2.�)�O�o28��׍�!]|!���'�0���I�/��Yy!�gئ�R&B~i:u�I�
r!��ڬ�`t���/�R����O$`!�O�X�Ve��c�`���fh�gw!�D�P�t���+T��Qe�66d!�ď:p��) �޹2�D�wbÞM>!�$[+ ^���'�0���Ѧ"\8i#!�$?�n�WE�i���8bY�0!��LlG͉4aޓ?�]����/~�!��M�Y7�֏U�=�*���'w�!�D��E;�Y� MؼF��u�
c!��Z�Qώ	⥈V��D�B��#�!�r��K���]�m��n 0�!�D${�41���v��͇N�!�Y��1�DM�R�����:!�D\G�
�����g4��i��ă
!�Dշ!n��cr��w9�<��N�Y !�$�& @�B#I"' QY"U�!�$T��(��%M�Q����Q-:e�!򤟸p
���䒊<G�P�J�!�B�"�ڱA �d9ʵK�Ol!�d��2Q��A�Ň,9���`'�3AW!�D�4u(#-^4$D�E�ԀOYJ��� g�,dy�& IJ�� k�yR�ϐ':����J�r��J5�	�y
� ̝H�+�?j:ĝ�FAQ"B���ɰ"OH|�chU0V��W-���%�"O�t�v.Z�-�*Q��K4���`!"OZ�y��L�0֌��$�
�����"O�d�Һ'>�C� V�c���!"Ot
��P� �Be9�F�L��!"O�=�u\)
��B����(�"O�
ՈW;v(i��/=��H�"O�eR�7�H�GN 0��,�&"O�MA�Jx)6p2�˳_�A�"O�t�'fq�Z����P�4Д"O���%P�jU���%$ۋ&���"Ojh��Rh���i�bE�YFlH�"O��{��I/�uh� �2::�ԛ�"O���6L��qגLQ��4����1"O��k%��>~qd�РOQX́#"O�M0�	��r�mr� �/݄�¶"O�Qk&��	vըw �;B�Z���"O��'U
����WO��k��(W"O��z��	a����$ǿ�jY{�"Oġ;�����p&��v��8�"O8�
6Er�r�2BS�*:�Q�"O@)!E�8`� �	��ܑ3(����"Or`z�	�*��%P7�`(V��"O�Q�tW�9s2�(2�θT�phd"OD�q��K
:Ȱ�H�<q�.U�7"OT}@� �pn� {�&��)�֐��"OL�sRm1m��K#�̰c">誠"OD���N��|2ŏ�1�Ru�"O�<R����I0v�@��2-�'"Oj���$z����"Q=�6)�"O&�����/K5��V�3muh'"O$�EҊ	��4hF�O��rT"Oȭ�E�M'@�X��\�MH��"O�Y��ъ#d���!� i�����"O�5Fi�(:z�Af��iW*���"O�\9�F�:��t�O�4>thc"O�uK��Z�('�S9D�""O��!Hv�2P9�L٤:j���"O��⧨�);xpK�i���t"Oڅ�E���E�6� �»d���ð"O6��$�� ����QJ����"O�u2�@U*Ĝ�)@+��R#"O
�2a�ƀ|2�5?,x��"O�x8@a8Z�:�`a�]�?v��x�"Or����W�]!�L1d2Ax!"O`�RӃ¶#��suE�8o�����"O���EF0Y}*-2��Ֆu��1��"Oй!S��}Y�#�A�o}�	Z�"O�����\2xYs�+�>lh�-�$"Obi0�L�p�RP�����(ZlST"O:�2���"#�|EI� żY��a{3"O-�¬�h�`a1D�E�ԁ D"OD��MͰ9�4�S�ܺ%��b�"O���+բ&i�@d�7S�p"Of�;뎚&T��`'��]��v"Oh���X�gF����ʕg�*0��"O����Ѐќ����Q�7�<Z�"O��d��qg� Y�� �Wp�3"O�s�N��Y�l���Y�&ؐ�kv"O���c$գ0����@eGR�ެ�a"Ot<2��Ϧ	�4e�D��"O��(��=BuX��ȌS��ĚQ"O�@�r
�/<Fd5h�V��f�hS"O� `��aĚ��`�ڷ�'d�H��"O�A��qS�8Уe϶/QRa"Oh���.�<���`d�[���p��"O|P@	�*-�&���K��(��"O�՛�%�2��e���rtP"O,�C��؅V�P��Œ22�b�"O�Q��j��T.�i�!$Ac����"O�tR�G.w\��
#��i(0l2G"O�a���E<0z t��$O&G&�E��"O谪a�ΝL�D�10dԡd���"O@�rpG�L�CԿ"�qe"O�ՠtd�Sx$"�������g"O<�ڱ$�4J�r�3�%�8#��x��"O~݀�\6*� ��*���M*�"O\�p�
ZW ��(!���@/�Ã"O�Ea�c�S[h!�
�(�`�"O�!�R�3��I�W�K�-�4"O�|r���+����h[�	�=X "O�))�K�� Y!#.U.�`�"O@�'I�+U�x!���ʨU�T��"O�]�&d"_�Г엇1�2̈@"O-�2䋦GN��)ë��I"OX�R��F�z�d�	2� �0�x�"O�s�A^90Xl��J��g0�eA"O2	�fI�?^�zY�r��&z�c4"O^5�3Myc2@��ş@(�0��"O�@��6����<�t]�D"ONda���Μ$�$AEo&�b1"OD��o�7p��t��o�<b���"O8T���"o�ɢ�m��,��g"O 5���%'6�)CoK�?��P�"O`RaN���Z��^�T� x�"OBPku+�W������2oݾ,��"O��y(I���[��T'̺ݫ�"O�����(WR��p���v��X)�"O���ԥ\q�t`��H�r�v�r�"OJ=��%L=Z�@#�!�W�T���"O2���GIq����E�O�^�ṥ"O6��lѱQ�1�͟Yݲ�j�"Ov$��-��<��eB��f!V"O
hRƚw�`�q�[�yG
("O���ʁ�N_|��1�T4��U��"O�p3Ej՝fB���7�*��r"O�����)�� ����"O�T#qeۉr�2D󲢇.��#�"OB�J��� :�.Y � �=I��	�"O��� � �dW�|�S����t�yG"OR�QaNJ{.����N4��b�"O<x�#�
;�Hi��l$�
�"O �z��z .0���P�?��з"O$8h!�CE*�@ڷ ]�]!�G"Ojly��՚r�0�C�U�k�}Y�"OJ)Ip�U���ӡ��?u����'"O"��#�3Ad:CӦ�IO�,�a"Oh�+��]��2ȣү��-9���q"O���5��!�*8b��P�w2
��`�O~���K�S �X������&���!��P�\a���K�V�����A�!�+d(���AO�f�����~�!�d:,�6t�W(�3M��P�BO���!��з9Yt�� *m�L��/�**�!�$�1x�f�5��h�!w�3y�!�a;�)2�J���تV�C�t�!�Ę�Y�t�P�0{�2�bSBS 3g�|�x
� ̙s�O�B���Hw{�[c"O�4 ���F�R����9^�MC���N�O��mJ�=��S��Z,on��
�'r ����R+� ��c�(,M�9��'�qO��}��-x�c;|� ="��@+XK�|�ȓ~���AMS&�$�q����O$����f-b1�UW�e����2c�cWa~�]�|��F�+,�RŠ�o?02<dSbn;D��藃�*���{V�+4�X�[�O9D��@��/B}��+�>���+6D�H�D�K�DD����V-_7�c�j5D�@�C��'��D8��J>ʹt+��3D��ɕ/�?f�5:5(
�:;��ؑ�2D�����א>����V ��Mr<Z�
0D���B���� Ө|zH0(�/D��#` J(	���E��x9Ь� J+D�x`�mޞg&%���ªl� 0I+D���+�=SN�W��,�v��$D��3ҭ�M�-ď?f���xC�!�O�ʓ:x�=b���(6H�J�MS�R�hD��
�R!q`D@8\{(��TM��BN(��ȓ$���L�#l�BZrH_�<��ȓ"����� hd�m�1��YX(�ȓ}�&a[�K^�)���D.�qZ�ȅȓ:%`��.�#'�0�c���r�;�']4��w�^"���*G�*7V��p�O.��<Q�4|��e�PW�Y�Ir� �1����\��O2N6�H�F
"�ĸyQ%�)4]!��p,L8H���<P/R��N�78�!�B�U^�� ��>�-
����ў�ቯ8��0AU� �;�x�	��"kx��"�ɓ�H��I�v��Xu�4!��h�&�&$�(mS�'%џ {�؊A�G�	�+��2"5|O�b��`v�T�Wf�s�F$%�h�"/�O��ɩfbU�b��5&�6 �w�\)��B�I�O{$�0��D�mHI%��3=�̣=�U�8�ddH��b������٨	�`��IW}R��ӌ�IB�<F�~ �P�m+�w�H�Ity�ȯ>%>-Kɟ�ref�/������;8�@̓s"O@1B� oei��@��p���*���'�bn�M�'��9O�4��LLfh�Ja��?��AK�O�0S��Qo�f��ʶ�&���$_UD�Dy��I�����@��+��)TU�\����*�k�n��w��{��M`�ݩ7�z��e̖�H`�֩�R��M�'��`���iR�����O>�����~B�Ϊ(`N�b�>8k��#���8���/�O�	#�,�>��qLŲ.m|���]��G{��)��1��,	bE�e��5�#OX�n�!�D��mv)[�]�K� t�"$ʁ_��	����'4�x��0A	�tÂh��O�]�c��y�ڼiDb�k��ڈK���x�����M3�W�a~rl���
ds��D�B�N�sw����>�5�����ׁk#���
��"�Y8E"D��S��X��𬂯C��!
p�!������
ç^��z�N�$?���`A�0RӔ��� m ����CHڱ��*X e�	�HO?i�L��M{�|`Ƌ�9L|���#D^�<��!���l�i��EbKZ}"�'Ӭ����9}�Ȍk�eY
����	v��1X⩜�e��+���.H!��hʚ��f�_z$��ʅ�F�(�S�O� Tc���m�b�X���c����'����T���D��TmŶR���r�'�4t��o�rӦ��T,6I|������ (H���V�F�T��CW�i�jЦ��4��I [��(�6%G Q�X� B7f�B�	\��֯�I-Vp#$`:I��B�I�dpj8T��!XF���9ijB�I�-�
}�
��� H9��{�8B���-�
��7� ��0�����Ms2�!D�� "�2��=!��)!7>H�� O��=��-��n�@(ӗ�@�b�zQ�g��<y2+|Q��Ɍ�e�Qp 
=T��F���_���#9F"�/:D�D��K�A!�ʔp��c�M8D������/RуM��&�2�x�E"D�4���>O���3r���"]�-�ҡ~� 6�#�O��b�֙~�D��f*?���2�'Չ'���B�j=zO���W+��{�J�
�'�Ԭ+��[
n�YWmY&'~���d�M���cf�6% ���Y=N�!��S��� �rN�\�e��ўd��I';�$�Dj��Q)�hN1'�HC䉰�|��Ɠ[��sW!�)KFC�	%5<���j+��!��0�B��t�8 ��6@X	#�eɿ%�vB�	S� ��F˶ �hZ9R�ԅ! "O.�q��P�;=� �ѧT1���a"O�\�	����
����Ќ:��'剜	|�@y�!Ӱl��|��̳d�C�$?Ґ��0�T�XLh�"�	IT|7�=�S��M�ԃ��Q�bJPIɽb��*�T�<q�,\�O`���7:R`Q˒&�ş��'��|��G�@��ш�E܂.H�t!C���=!�y�
L {	b�a���'Z X�����y�Җ~t�8�� &="�BFB��'^qO��|:񏂚5D5c�+�k���8ሞz�<�t���#�9j����x�'ўb?��ьϲu�:�x�@F�����:4����*U�"q:���=f�tU�s�qy�)�'&cn��`��c��s3��S�T�?���O�~�������,Q�w��5���Te�D��:5BY�Q[�m֏)���!!2OZb��Γ~�� r��dި8I'N�Ն���O9����#�~!g�r������<ى��S�;��L�a눉{4� ٢�ז�dB�1qN�Y�������I�E�E�VB�I0����#���+:X%q�߻O�6��d8��9K�rQ��Â�$�BIF��Y\O����kx\Pѥ!���0`��1O�=�|�U)��CD�!3��<�|���c�<�ᎸJG��@�/�H^r�+��K^~�L/�S�'D� ���Bˤm��B�̍2*�N �ȓt�d$�pĚ�jnPp�ڢj�1���d#lO��G#�L����G`&���D"O(
 L�%p|zǬ�01��"O�ih/�'r�Ƒ0sfԄ��P˖�$�Şqa��Q1@͜h��Iy�@_����ȓ��dhP���hό<�MGx�'�J$cĜ1dL�	��Y��'?�d��2��a�1`f~d�'�"d�@""���(A��n��t`�'��X��V�Ed\qb� �'f7>(�'�%�c)�<O��8ه��U�����'Z&U	����t\.���&��Lp8��
�'����a[;$^�GB��8��B�	^a~����KP�k��ހsضC�
>$t�ŉ[Mp���� ��C�)� L�Rf+�5���0�,��"O�P�D#�nxh-��$#���+0"OjP0$�%j���w$��	�H1!"O��A#��{�)���W�9K�D"Opu���ľ��P▃\=�L"OP9�!����@�V шL\�x�"OfY��IE1{�%���L.P]Z7"O�Y�D�1 ���)e��H��"On@S���9Y���s�ıS��T�#"O�$Ѐ#�Հs�a�Y[�ъ6"O�d��J�:�I1�E�$fИ w"O�)�9R�� pХ�\�հ�"OHu{�̓Dm�1h�d
<q�z�{�"OLx��Eƾ( ��uW���qȒ"O�8�"��V�9�2k� 3�ڑ�D"O��xs�Պ ��0Ѣ��/�u!w"O�D������� E�5F6x�'"O�1��/V�F8��Q3E	 "���S"O�li6�z0n� �_�N�P}�"O�QP��s��k����	�4�y#"O���c��0=v"�'�+���X�"O��ۦi6��yXtf��l�h�(�"O0�AE�(X2�9�c�D�.����"O
�X��Z�h�xQ�)*�����"O�}rd`S�tC19F�5uk���	�'<6�c���#�XI�@]	E�| [�'��Ĩ�� >1��bc�+,lII��}�65���1)���
���x�D�1�x���K�Q��(��|iL���E�'%��a����$p!�}��{�Z�@�J�8GR`����#����ȓ^ځ@��<����R	�Z��ȓ2�J�x�d�[m 0�M��M���v�����L@�+�b�{�Hs�⑄�N]�99��K|���g�ѱc�*���AfLZ���4�*Y���Js�@�ȓV�b|9���>3��c��+�D�ȓ8{�I�D���:
��` ����nC�O]�H��jR*�>G�B8��[ݬ��JB�8!���Jӌ��L����ٕ~�lHI�g��gl�%�ȓ	�^���)"�>P��I�TI�T��*�4{���1���iE-SL�&��ȓnf��jWdǠ<��v���ڝ��y���v@�H�̩��f�yҲ���^�5��.�!����з=����Dr��bR�Y������0��ȓL~zP�g� ����Q�܅3�>e�ȓ&"���oH�w�L�R�SC6Y�ȓS-$�K�ʈ�x�P<�3 \ �"���f�`T(�� tX����"�h=����k��EAd)E�m#"퍟D8���!̪d��<Ԯ�btGA�Mآ�ȓ!���Pe&���f/¬	�"h�ȓz��iҡI[���Y�͒#e�Դ���R��ī=;VX��oWH�@l�ȓ.�|i�2o��R���a�&97�хȓq��з	7_�u9;Et���'���wnƕ����V1B@�ȓc�8Eǘ�<N�� �$ձ\�~8��L)�I��)�f4�ɐ��*|l��ȓf<�mԤH
da�p�j�t�&)��� S�LEB��'�8�L �-�
4���� %J��X�'�\��¦�v�:ɬ�'q�Hs�.�4���[e"��H�(���� ,�� y*zX �"O� \m2�-�5��\�Aˍp��Ȼ �U��,�a3*H���)��<��*�?`�����W �6��l�E�<!�͊6 �t�� ��.��)�����<yC�M�Dy�­=\O�����9�
�`vm�y��	��'�����O;3�ra�E YjN��'�K�f�^0��y�"@�lQXt���T���`�!�4�O8��f℃\Ӭ����)�3d��c
�w��Hq! ҠZ!��77L��r�8k3�I� �*X <@�C՚*�`��N�"~Γ^
T�
�W/7:��yqJ�i�Q��9������Ϙ ThY�p t��I�y|��i�'B��$��F����
�J��ez���a|��
#Ḑ�e�ӣD�d��k�d�5	�F2p�a��'׮���AQ�W��-��������䟁?��u������(�8PI�Z7 �h g�]�>m(q9"O2h*B�\�^��m0F��7o�@Г& �Ĺ�uH^���)��<�Q O/OK���8*����\p�<�B�Sx}� ��]l��t����l?�3`E�-��h�e���G�EU��� Wb����	��"1��'��r��>FP"��'��P�<��'�l���%�	N��Cw�I*���'��mV�B8'����JJ?���S	�'�d�"J�"h���8V癈Bh��'�~(�����<�P�됞w+bɲ���^;�>9(��W����S��0d�]�oK�!�$��P_x�T]�d��!�n2p�]��A'O���hQF�S�R('��O����6Kv��(.�~��7"OD�8�P��%��x H���@@��9�s��Y[JT�'�T/{��I�^�Ԉ��;M�� "pD�8l�
��d��E��9�m (���Q�F��"O��`c��)c�Ԥ�sB�`���'�ea��JSB���AMGG�ȓ�}��2 ���K�e��( D���79�O��b3�_��$�k��D�2Vz͙	�'�L�
�͂0Jz�p��@�(^��ao�+�<(�$癀�A�����7
�,�I.�\�șw��К���P+Rh�Ј5q�X	�']�L��;�7��i�����!ʗK3N�p§<D'�u��-L�T�d��'~2�k$�ݗ��	=l���Sႆ$"�KfD��4�4��d��9s2���}��!�L�$S� �i��%����T�\�1Кt ��H��B�J�K�I��q
�'�M��`\��� .� |���B�y2N��~�����7h�4��h�-��wȏ)7�e��[�I�a�$O��CBڇ#�Y��'/���P!�z�b���J*�0R��Έ�T�'O~�ҙ�AB�#-�����|�l���j�(� z�w����5F�h}� �G�ۡ�i	�'����Ռɍc��X"w�Y~��e����Q�0��H&t��e��j�_x��H�,�a��pz�
�y��M��O$��%HBaJ��׌Ϝp�D�	�v�<1��]�\;rAS�B���%C�+'H1I£�.C���b�ه^4�͂"�$>��bĬ�+S֔u��	�;�6|b�˔1n"ɚ�����RjȘل+וO
�eKpi��L�r���J�nu������� �ѱH�y[c���N��AcJ�sH��'�� c�؏wZ"�&#���s��06Z�� w�D�@mօA"�9��(+EtP:�Ɲ% �䑛wo�U�A�'X-(���V0$�~�K��5j�}���C; ��q�РxP`1R�M�^�$�c�A�@�1��E�"6����O�r�(Ѿ,��'��)��Y*6�����[�:��э��d��2s�O�iC�hj�DV+pB |{
V�t��4��2;�:æ��6v�b˓>���`,;,O��[��LUߊ=9!�E,����V�t���W��+�nK�#��1��ն`LL�>i��'�M^�0���i��(D���Ñ\��	1��t�M;�-�H7�������s'N5 �l����c7�>���I�F*B+�? ��K�*P<�3$]�|���H!� "ZM ��UJ�<T����w�^	W 4�����X���۰<�D(�2zz���g��n#s!�J8����j��x�2h�L�A)8���@-?���`5B��7�е� �"O�5�6
Ͻr��m �B��$� �Ap��S�I��h n��Py�#}�k `t ��������
B�<	D �8i��xK�i��;��ġíѡE���v+w��b�����H���G3�Y$F;Yy!��H���j ��n'���f�F�W��	���,���Vb)|Oi�DꄖVy�\��3a[�j�'n�2�ٕ �V)��i����NS�R�~dpG�(�6��	��� "�zv!���Ԉ"�O�rU41����)�Tҷ�Ա�h"}���0@|��70x�y�@Q�<A�jTXP@�`��3$g�`ƬZ7�RE��EU�dC�I�k4Q>˓��8;��8�����[�&����ȓS0R|����l�F�rQ�R� K^�l��u�rm[�T+n����O�]C�:�d��qmH�y�{r�֝۞T��g��������TO �ք�`l��+D���
W>Z�^-qg7p&��@�+�I$V�Y��蔯~��>E�	��}��KH8RP@d"�L)D�����P�����K�_&n Q4-�;}_�"����	N��~Bi�)H�M�1�[�nɚ�dņ�y�k��(JDO�Y�X�"P%ƍ�ybI�#F�=���'eĂ��-
�� Ϗq��x�?L�9��q�$��P7Qф0�W-�7=� 9��-D��p3̝���,��/[� ̼s'�&D�$����r��8�X?�)��"D��:�,�
1�����?zٔ@
C�>D��Hǝ3^μa�`�fN�ɛd�>D��h4(W�s�� �Q�Jt����+D����$f|��f!M:L�6'D�l� �$kVӃ��.��ܙ���� I��eta|Riؕx30q	AK D<�u.�0>)�`�.A�xa��L\�{��4S)����ۢR�\Ʉȓ=�B��� zg^9�4���`�|������	�g�O6�#i�|�ӌ�i�:���k���y ���G$!B]B�nSL��3+-i��5��Q�FĮ8Ѷ���=�Ъ�ZL��~�� �u�+@�؊��U�U��K$U�.�H�㉒V�R�3s,�Uܶ�sPJ�<�h̀6m3~`p�A�V�W��X�!�'��`#��`���I�$�N1�
�+���@�+���W$��W ��V.��+0^�' \i��8|�B=K�N۔Q~�H��^= �7��!��]G0-��&R�}��ɂP�ڠ(ƴt�DҁXa6��G��-@����X@:%��O�"�+���M7g�q�r�U(:� �  �J�5�az�j�A�X̓^j��h�DηE/���d�Q�0�~iI�״SC�|;��N
�`�ח�?)uϵF+����!����'���t�է,��"�h�Z���L>)��CX������@RU�2'ت�2ԐթK���	�'��<��Q���l� j��G6�?��l��$4q�FI�G��y2�9��xV��j�Yv�J�T&%Ё�ì�1U�L�1�H��b�'2b���<���iÌ  �tR�R�z�rP��	\�2K��j6$C�ɽT�.� �GD�wdA:\XK��ζi~<����dB������r��d�V!��? Pp��z?1Ǉ��=�9X$�O�(�x2�݆Y�=�`"$,O^�0��S��<kܴ
i��T\- 	� �0��K����^}��ѳx	,e��Oqy��W
A����Lr�I�0a*W������5�8Od=ڥK��`e8�4E���˷��G�b��� M 'X�]�I�(��H��1��dQ��K�:�Gr���
�FY����آ;� |�b�A�\Y��E�Ơ���K�O����N�R3d$���S�|�Hَ\N@ �vb����?�Px���o�2�90��4��"�+1hn��iқ���.�,��f�n�>�) �n�D��|�n�7\�
��Q�R0[�4XE%FjX� �c�$c�
�y�Z���
Z*:���.�-��)��Dl�^Q{�4q�ص�M�"~nڮ/,� {Ce	,���@�
x�O��!���z���	Wed #�UNJ��#KY'��I�l��lj��\X��y���K��ģ���en�(X�ě6k-���=a�u�'UN�u���?K�`c�Θ	9�<���9D\�%��'�MԋόO�����,L��C����h�~����]�tY�� E�%n��!�CA"�!��ŗd�`T!wj�( �sR�A$D�!����`�pP�
�����NS!�#�ڝ��I�O�
�����%!� w�y�$�.Oٔ"t�)P!�dӃZZBa*QkRC����c X�m	!���+z1�(I&r��d�q�@�K!�$�φ�H$h�03�� ��34�!���~�0��6.ǁj��\��n�>}�!��
Y�XXcCY�f���@�^�!��O5��e��H��S�Ʌ�e�!��Q�Pd�O� t�,�!�� �P�c�P4"i�Տ�mX	�"O�%8�mR�#���0D�٣[�T�4"O����BOS$�q@!4��"Ot���B�*�3R��K�Q��"O<�����H?��� ��Z"O���K�#b��S`�C�p�L*"O,}ᔯ�N"&���Y0X�hٵ"O6���(��:�c7cP�P�XP�"O` r�F�M��2�m��~��4"O�i�ӌY4̖�a6>�%lO��y��ا[�����Je��f�A��y҉&0���0�(�NW�����'�yBL�=�f��̩~e���b$*�yr'S�I�v�C ��8`�ĝ��y҇G-"B�D�E� v��yF����y��{��er��}b���(:�y�Cԛ3ʘ����t�i;�H�y�䞁,<���˜�\�*�:!�R"�yB	�t���Q�"��U�>i�`���y�%�u	<k�њ������D��y2�/'N�,rC Ս�&��Rh ��y��I6O��2���3}�e:3���y���7ܮ%���
5��(٢ �:�yҀ�j^��CP� ����=�y��`��aϾ�����&5D�p���70��d�68��-3@l5D�hj�藇:�%�Y�^��c7E<D�p�bF��\v���f�U3��L=D�L{b,ښ,h�
�'F}�)ju�=D�8f�66t�k� �[�4�91F;D���2��y�ұ� �U>4��#6D�Ъv]�K��Spd_�jt�27D�D�2�Ջ@(�1�?�ѐV�3D�x�1)�h�EJ�C�	��a�#:D�����6W��+"ݍi����%<D��3�IǢK1�\8�iO/� ��(9D���ᄝ�nM�A� �>�ꠘB�4D�ԋ�^W�����	Z����S�2D�3�N
h�N��`�K?v����2E3D�8��4�>���"ǖ{r-
�#1D��(��&Tg��9��ѿ7��(��.D����dE�xAK��6�zܠa*D��!!��DX�X3���8�T�r��5D�8sB�'A�$T�C�^�^sD3D�����ɣP��l�q��.���Z��1D�أ�hK�WX.3��D=D�� 	T�"D���a�v���y��^?Q��QBn5D��	�Kфej����Oe����$D���M�\�x`�R�(�j)�c#D�h����nn���e�!^��1Po2D�Tf�alHU{��+*.=��3D��I��3s(�ّ�E;7P	��.D���𤘋+	Rܱ�dB�y4F����.D�$1��Þ*��ذ��/�:��d�1D��{w@�C���� 1T�e!�5D��qnO�e��&� �Xc�'D���N�9Ʊ�P�S�<^�`���0D��١�.�R���]�~zu�WC*D�8����&OC�i�O۪|i@�o+D��x6��	"Q<�i���6�HA��c&D��&$%=T��Y����0��Q�3D���A�G�7k���*
2����!2D�`�І�F��XЂi_+���ڤ�'D��h��߅>����%�ڷ-{�)׏(D�� �I�F�"�S�]�xK�0��'��)@ �$*CI�&g�H�@��������rd"D�h[5鍽{�ޔ1f��<Fl�\���"�K� |sei=�H�(���n1(��q���$�ʅ��"O��� 6��Irp��H����oذ}g|Y����)��<�qN�xd-��/� w;��T�Mx�<��%A0��k5\6����U�<q���)���a�%3\O����#ˬE����F<�)�C�'�,���X/�L����fA�A�*W ~e 		�	� �y����:ij�l�6l4� ��OM�@����&�(��Ă$	B
d�^�13��0A��S�"OY��� ��!�f��()��Z�Qf��`�H_#��)��<� ��1��E�$�~5"(��G�<iW�^�x�<��w���e�����`��<�g,CzXr�`&J=\Op�z���i�C�?	X��q��' �U�r���!�� �C��"�����m0Bԓq-��y"BʒY�H
�k��b}�q����Oꤢ�� /����$Xk�@iU�4#2p�R �Y�!�X	�����L$T���ψ1(����Ѐ��*ږ��L�"~�|�����U P�j,$�@�ye�]�ȓ_Q��X3�ʀH��L˲(H2f�h�ITP7��Ű=�`���&����!ȝd���
ҥFX���5��	B�E&,���L1hQ��,�$�y��؟z3�]����3�����ą�y��,ݔ���'Q9#,��C��y"fɨQb�:ƂAA���p�dѥ�y�Nʊ��6�M6.P�@�K� �yԀ)��MΫ_�`�Wƌ�y�EM��J�ΑLHμ���A���'Iʴ���R�S�'9
�*�̜<?6�H�HD~�Є�"�R�ʔjR.��cA����FQ�o�m�ɱ�LE��Oq)�%ά0���Ɖp�IjdO�t�&B�ry�s�,�6d�!�#�Jg,���_���>�0@'6Z����i�NR��rA��wX����RM����R�h�Ԣ�=E 49�a�0u�i%�-D���ǤK
��[�	ξW!�PL*�S~!� "�Aؕ�M��B4�c?����t|�9Q�B�#x0X(��+D��dM>Q����F���~�᥎I���+۾Bjn諁H�[�vb?%�Odhk�a�0c��x�5
'd�HO^tЖ�&]�򙛣LA0m�SÁ�n�tQ���߸8�P q��<0l��I�� �ʀ�ߒW�(|`j�"F!��D�>&�lm�� ��D�J$1c��$/�=��"�Pn���Ԑ� |��\s<�󌅠>�f�34��k�(T	�%8�\ ��-����Y�L��:U�ܴ��D���%8t�	���%	��n_�T�t��-�S�r��B��!�D߄V��;�lK�(ؽȥ��/��!y�� �θ��`�	YTX���o��% � e^@U9�NE/,�^p��O�������y�<H�E�-�H��I[wZ�)��]�r�hR�̣i&t��Ռ�iq2��$�'3r��C��^����v��	aO�eb�'�;1)���2/����:�i��Ǻ:R��.8L��M���h��ǉ``�(��ďi߈i��.�|�h�o^��ZQ��N�-e�bL�a`֩
�ꥨ�'St: ����UA���d����V������^eo��za�W{Sv@�O=��]Y�F��|���w�N�x@Ư~a&މ|"�=���h�@�@$F�d�b}	�'�Y�]�և��QKz�+��gv��eˑE�I�fr���%�1��S�~����e
/���[q��*=�џ(��"�/��aҖ/�2|�������@cœj�>�����$�h5���|��]$�l1��I3+������<r:0�E囚g�\˓C��`L�j`��#u��j�|#}�K�P��u`�"^-vl41y�<q�H^4{H�r�)R=Fp�	��E���yy�G�)6�"�sTg_�)Xȭ'?�ԛb��)zc$���lڨ�`c�)7�Ћ")�kh�IW�#3��U��ʝ��=��!Vv� $S�e��P97#Q�F���	Y@��ݰ�O.OA���fw�3cF��y2�g>�3ǓQ�F���A	��y/�q�^u$_*1Ķ�X7-Y8��'�n��6l|�G��됇@��8�Ԧ�4,�Y)6��5�y���-b���y�m�.[�`�V+H�+B�B6l�����:PQ>�S�? 4i���2u�Y���S(~��M��"OHI넀�) <)��,P8.�>4�4L|�R	� ��ă�|��qArخ��r�z�"ܷ.q�C��c�X]�� ւA4���	��y�ꝌG�P���/?k@�ywa���'"����N�P�t$��Ӿɪ񙗨�f`�8P �I�C�I-+�.���O+Q�paF�5N��͊m�X����*O:�K��Y�TA5b¨]�s�Eܹ[� ��!/D�Ќ׀TZ]A���1�lӘ�2��@(,$��J!�'���5S!`Z@ڥ�9$���
ߓ\_T�S��^-(�
6�M�cOZl+f�4t	���� X�Be!�d�t[�����P�S��[ i�O�m; aL(�R����0�`�F�uY�2��2o!�ċ�ٰ��jVH��C뙉'�̋��J�b��OL�}��9�xd��M�હ���,�� ��$B�䓼r��K�F�MB��ϓ|B6����>��=�B�CJ��yI���N%fmb���C8����Ʌ�F�d]��Z���n�=Є�G��,2�!��=w�A��@��!Su�ǅj�!����ad�@�G�T��b���!�Ę�}`^��ŝ�D�{G�~�!��L�cU8a��O㪬�T@D��!�""�I2bo�7٪L�m��\�!�F!L|ꅩJT�i�aPSU#|�!�DN�!].@V������Y�K�>X����VP�0��\��@Ӗ]3�0�$stم�0o�*����̟��gJl��%냯K�l���Ǐ,D�P��/����$q�M���4��O q)`�ϒ�~�eϡR����G��A�O�B�QG�j�)�)��n<Q��"OHi�dI�0�$0�%gG�e0��7�O�@i@sJ�Yw~�Q�'Q��Pb��h��Sq�{�+
�TXђ�,ON�����`�*z��05	�`�E�5,�M
pj�aB�$	 �&�?I�Y��N�)v�/lO~ęU�(d�#��	/s��a[��r@��\�����ȍ=���0�����)�Ŏ^3j���[wb����s�,"�
4v(h�'۸��@k��`pC��P6z\6AX��
�.���F�U]}��eaנ��+C�|J��y[8Yp�w?ęz�^!6F)ф�v�p�(ӓ��`R�*f���A�U1~�~m�b�Q;��QwkI(�q��ו)n��î�p�����'{�nu�Bf�
>���<a�c��98������i���Aov�h���/Q��P���N;O�!�֌@
�Q3���*Bl]���J27زP�s�^+-`M���x��8K���$?��]�
�8�hy5�?ZA�b%��pf�8�S��M��ȂX�<Q N�Gx��r�����
R��h�g/>k��,<�y��E��CL^�1�
O�%��HD�RV� J��J:�L� o�m�T�J��ȠO��{A��#���ʖ�ĬQT���z?�o��A(~K��M��8:�F8��l��F.,O��IԨ��v6��48�]�ʲ�����[��0�$k�K�S!�K�I��= Q�Mcy2�E�+�8�� �a�~����V03�@���oFwVO���e	�<����4k��=�e,��R�:�q��t��}q��n��
���S5Z�j�@��S�\��e���I$�'^:h*��A� \t��#�Kuh�� �B'`i��@�z=�ԉ4�W��h�0�ӼYa�ѻjP�6��m��_��ć1�A�fAV5���u�B-v�ب�E�$b4Pc|��b@g�z[I+���V4��'���S�*�t�@SN��*]3u.�9@Z���:-I�Jܶ��V=9l �$�Kc���!!M1Λf�G�	��� Hg�ӧ������o#�#d�����R�@������z����0|J��ǺC�l����}�̭+���^}r���7����4.Qx����S�}��9"�)��;�M0��P�{�qO$�p��@	���S���\J�@�{� %��i�`�B�	't�`	T���qKʘbC����">)��N-�ȣ|T�<(��S&/��?hpP�,RP�<����7 ���)��w������E�<�e1)�2�+�$S�R�١�%�}�<�a��F��KvC�K2�a2��}�<��JC����j��MG�%��a�b�<���Y�FE6��dɚP�P�
Z�<��k�$��$C�ޛ0��@e�P�<��8y��@�<��UX�+Q�<� �10W�'%jl����ш,Z�`�"O�"�S2�|�2�S�6� �i�"Oޠ���n0��a�T/��Aiu"O�����ОMU�-�BgM �X	�C"O���nV�>�y�#HA�,��"OpP��İ*:�X��S�1�65!!"O�#AF�1vq��"�����"O��J�DL�ð��ʆ��I��"O�\Ba���B`Bn �?�luӴ*Od�Kg�[��=���27�8�	�'��]�df�/;Y �*F�%�"��	�'�EG�D�i����/,l��@�'Ǟ)Q�(���L��ō"e�f�#
�'mx /�fz.��@�>^�0�p�'�
�p/4
��p�G\!y>�8	�'��i��W�� ��g���49ڽ��'0f�	.$r)L��e>Y����'�(���fϨ��i�Dȣ;���'��ar@Z�,� ���5ː`��'�t�����]�T(�A�.[w�Mp	�'��,	��R-Zwba1�W_����'�j%0�ƈ�3R@� O�W����'à����/�8�d�E)�)��'u�x��"ε��*P
M�:"��'m$�Z�Yuj�R��F�2�6���'����cH�,���fX2%$ٺ�'�6T37Jͦi4"Թ��(:f�'�~-���$(�F��$C U�&���':a[�$��n���\ �����'�~i�e�֓M���1허)����'��k��>E|�a�`���_�4��'@ �*�͂c��tBӥ֟C]��a�'����`��7���z��;�8I�'�L�鷈:w�ā��$֪S���
�'4���V�^<�%� �I3��˲#)i:��Ë�1-����|Oȝҁ@�Up,M����<u?�]��e'
�y�헰+�����������L���fɊ�ohy��,�D5��ȓ<�p0C7HY�{@�T�Hr@�ȓP��%��^� ���F�e����M�����G3V%�-�"NQ��b|�ȓ*T�ƭP���ӧ�	����<�ÇGI���O���J�)V�@Er�Dd��
&��'�`7��؍�'���B^w� �3?�')�d�$�4J�f<���V\���kFA��E�,OrE���O=L��W%]�,(�hT�g�B1B��T�|T�	U���(1��	�fǓ0��	�M�d�8 ���@}rh�6i@!�֡@���	Ll�OE�Ub�H��%v�u��h^B�HSd�V���Rr�7��%���O�?�yPƋ4%�А�œN�	�1Ad�L[�@I�A\8�'���	ׂl}@��"l�,xԜY�)�ZQr)��'�,Ô���Mx^Ԃ
ç)�R��G��jѨw,S�R�x��Ż�~B�=c�P����+����O� J��p��cyp%%�����8=|E�X^M%�����۞r��d9�����d��K�UD��!7(�<a�kFy��IZ�a�J����w
L����تΦ����,��	�'�8<'?-8I~�6#�20eb� �q�$�6"
�h2И�0#�V�m�;a"��}n:�+	�{Q��B���=�4��/O�V������������|xX���S�{��@�b�*wU�  BF� @�h���OV��'@�2S�W�?����j�|_�<еJ�xg(%�@K}"��.U[��3S	I%���Z �\ �+ZGjX 5l�	C�D�$�����x�f�E�~�>q(7���>sPF]JY�@��`��S�p�^3�ݠ��Tb�ѩ��\:�!�$-]��J�O 7.5ry@p��
%�!��/1�X��AӑL��(c�'�;e�!� 
g"�9��L�S�Z���O�i�!�d�>.(*yJR(�8φ(K#��2!�� ��S0��?iT���J��p��E��"O�)pE�ڸ��q
���7����"O��!���o�T�ZB���8k"O>�`%o��%���($���mrX��"O�I��ŨN�@"q��M���ɐ"O�h��K��P���	��=A���"O�;��Έ@r�� ���0/2F"O�%�`����	�b�:"W�c�!�ٳBl⸒7/��>i�	�v�ͧN�!�_�S��`��-4hf��nE	2�!��4d!�Հ�m���P�L�!�FY�<=�;U6����"�!���I#���'��I�pxQ�B�[�!�P�R��A{U@V�H�P�����&&�!�dUz�>�o"Z�&H� ��!�DX%=��b��&Z܈c�.Sk�!��-_$*w[�byI��"!�=~�,���@e>NEZ$��'p!�^�@�Z�0��L����-z!��2�`�"�F�SH�!#g�<r!��3WO��j���a>��B#&�:gp!��w`�t%R=r{7JB-S!�*W�|{���-�T���F!�%)�����_�m{�@�fA�$)!���{���;rT$d ����>Yj!򤌆@�T�3b����E���]K!��[�R��!S o�w���(r��y�!��-?���J>|���T%�?F�!�d�.���g#R�tx�U	��aK!�D��_a(��ԁ̏P�ĹQ)B�#F!�כ[� �k��(��	1����m�!�D����4#P ��0Z� T�A"[�!�W�y��q����O�@�	㉈�!�L:o�.Q�q��6�D9� ND �!��0-PZ���ʅ
����Т�!�ĕ�GjLfB�Ut��qɅ�!�$=xޑ�a�: �r��6)���!�d�&@E��
Ԣ�F*h��P탄b�!�D�>|�t��$�Ux��<�!�d�F������'���ǂ���!�$)3��c��-Y4Re)G�N�/�!�]%o����ʰ*w6h`�R�y�!�$�?����ӛjZl}��`	J�!��͒Lŋ�̃{���@" ��8.!��LJV�P�b*��e��rr�̇%!�DÁZBJݲ�	�r���3��|�!�o���`$Z�t�0#� �!��4E@0�#���4#�aD�!�
'��4��([c`��+VN�a!򄛙R�&�3&�8nC�11�lS6rP!��VG;Pp��M�P*Z}��J1%�!��Ǟx	�B�3��*�jѵF�!�D[>Y��ģ���0FըQ��O�!�dNcs�HA`��� ���*�!�d %-���1&a  �0�RW��*U�!�Z�4�& ��LSX���g�<q�!�d:9<�5q��4v��y��Z?\�!�č��b{�M��	�R��фW%�!���}P� �`߇�4M(���G!򄀃=F$`%FP�d�8����ZIV!�A��� Ʈw�y �\%SS!�$������-�-a��7L����R�5�r�!mڹ�lI��y��֬P��D�!��}ɦ�9&ڗ�y
� �D�g�ʁgF` ���!j.�#�"O����Z�<M��$�UW��Y�"O�a����"'K� �C�<o6pI��"Of8{�C�>�j&�<`%pE�7"Oj��b�Ēx{�HE�]�5�Ekc"O�)���\&0�@8����2�`"Oz���ߋ�2��v��	� �r"O:����
)��|Z�#	Q�ؘU"O��q��#ҭ��E%Җh�2"O,���/�`����#�+)$ʬ�C"O���D� �TK���d`p�"O�)sW)��Z��#\K�l�"Oʴ�P�&�>�I��k�`���"OΉ+��ԇX���X�^]�~@BW"O��D�ϯU�����KW3v�� ¡"O����n7����٢#��	b&"Or`z _�
�xE�s��r��a"O���&-L���A��_1R%09"Ob<�'gq�0&j�1��I��"O5�$�B�E]�e*ѹK�}��"O&�xD
N�0i5d�xS��i�"Op�P"i_�1��0��P�'<L�5"OJ��t�V�H�� �%[��§"O�|ђi�"rHhׇ��pҐX�"Oа��C�$���ǔ$��u�0"O<���gÈP����2&�-�x�W"O����
�HO�Ar��W
)��iB"O*���ܧ|X��{��Ü)�X��"O��R%́�#��cg-��#�V�iD"O��qv��B�Ѻ�픛"�d�S"O
d�d&�6��X�M�d.�qW"O5rc�7>l5!���Ѵ(�"OH Z� ˕)��`+2%��[�t�"O��`��8��ph�a�z�Q
d"O������(���OR����"O*��uAH8^�~9��d	�\�R�"ON�"(�;��	t)�._�,5�"Oެ���3�j��'y�.�C3"O|��n�r~���`��;m`Z�@�"OB�+pD�>ڌh9�k^�r�z�""OD�[�N�7'��y��a�t�"O��*���k���U�/b	I6"OȰ!�f�,J�COQ_���V"ONI�S�ޟSs ����g��%"O8���K�{�������|�� �"O0TZ��H�sm����K����"O�%���()���F� 9�(d	P"Or(���f��]��Z�7�P�q"ON`��c�d�YC�k���*V"O]���H$"#j$��l�E�z"O8���ӎ{���I!0�d�a1"O�l�kȗcGb����kYr�qC"O֥�U"���Ait�X?�ũ�"O��{��ѯ2�@,	��̵P�0�"O�;���a�U�� ԛ=A� A@"O$XV�v�� 7�1|���	�"O�`�ǟvg�t�U �V��e1�"O������4C�,��(Ȱ	5�u��"O���#�X�{�����@�&y�D��"Oy#畑 ���'�D� \{ "O.Q�C�Q3
�� �wE�]1֕��"O�9 D_�"����]5x����"On\�g���p�L��N
��"O�FI
�phQ���
Ҥ��4"O� l!pa��	�d ����/��9�"O>�"�[:J�0�"��s��A�"Ox 4
�:|��1uDFb"O8�1�˞I���&��d�)�"O�n�*��Dh3I�����OժD�!��Ƞ@:ݙ�l�j���0��!��Je4���J55�Bu��D�!�ć�?Qr,�g��*�	`d�!�D��V�@кA��"*�j��D�!�dD���1,�!�F��UÁ�_�!�{G��6AN�/^Xj�!�H�!����@�Bd"\�f)`���4�!��V�j��M��-��`p�E/�!�$�L�Pq��C���=;�D�F�!�d��Y� ���
-'��I���P'Oޡ�d�$5�
�p��:}J�`Z�A��y��� i��S��O�]k��i Lӊ�y�Cݽ|#�K�,C�H�ɛ��V0�y(C�nhct䔤R�tH!d��)�y��]1�̀a�ڟ���
����y�%����9�ԥu����D �yb��r�ŋ�'o(D�5��-�y"'S���p�sJ|H���d7�yB�NFP��e�)<m��(�	�yRlZ�r�B6E���!�ϵ��4��'���@eD�1=�A+&Ɛ+lX���'�4��̗�xO޸be'�	r���'�^�J�V�9�rk�/�+�:Uq�'���QmѢG] �td�3
z��'�*B�@"�@�3JC%����'w���fȀP2<�B�+U��(�r�'t�����W�������Y��)q
�'^u;fE�9}�0�K"A�����'��	�n�?w����B��<C,�J�'����a�Т�F�5����'3���@�1��`"6��,&e4p��'��ԁ�Ɍh U��X3�Xx1�'ǾMA&���S�X!*����h
�'֌����+U8Ȑ�tO(u \0
�'�����.Km�D0�	^<t�X�	�'Bh%7��w�pT��9 �D��'p"����X&���#]&Q�;	�':�`E��q�<P6��C�
�
�'Ѹu`Qfխ	e�l��4�\�	�'a�})΄1l��A���W���\�	�'ox9��j�T|ma�\�_���'�x,���	
 W���b�� Pm��'J���e杹��,bả�f��i�'$�����6^����C&'���R�'{�E�biB�{�0��#���P�
�'�B\��c�%#� ujG�H4���@
�'�Ι*�@Z+L%�D!��-#�JiB	�'�xe����b�~l��-ƍ!�P��'"����L�e�h��2l�
eI�':Z��aش"*���e��j	�'l�idA�O���A�0$�i��'��4�P�	��+�F�#@*�@�'�D���Kj�^�"��Dh5��a�'JhH����L�Re[W⑴p����'Lb�"�	qF�]����#��Gy�<aw�'\��UrU'\-p���AFPt�<� ]�L��@��E���m�<�4��0�6i��[0ޘ��#�	f�<�2�����dE��)Nq��hM�<�+w�   