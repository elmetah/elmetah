MPQ    @�    h�  h                                                                                 �&J=Vq�8����ʝr�Y��7���_� ��5�q�OC��&�EuѲ�@w�^YD�0Y7	����gV�9;a�_��Y�����F�T������T��w���{�n����]��}�3)�x��_�t��C"�Ecx��� �+~!Q��;�rY/���G�ؚlC�X	$�̲�hj܊mH)	 ��
Sז�_K.^����-�c��fR�k0��v�$�qK�S\3ٯ�s��鄍*��'^�l|]ܹ����u2��Tx���g�h��$��p�)Ejc8���;�v�n��}�P��z�;�ފ����f6�}��O��՜�~O�ر&V��>\
yZ��#r�rݴ7p����祏Ҟki�� h	Glj��n�Z�����#8�F6�ޣH	����,o��>>	�|�:�Ծ�VSQ������s<E4���2/��J�􎌽7�V8�[Cf�u7h��@�c�Bx�>�gf呃V���/���H�҉�x�o��9u�G�?�:T Co����._>Ka,�}՛�L�
g�g"횘dK�%W�6�3�-��T�@~�늹�d���ii�Fx]���L�	;�P�GYÆOW|c8���),> a	sB�9��lU?�������Δ�'�h<�M/�!�:Z;r@�?��Sp�|���YAWmsP!��i�fH��()ě�S�k��ƱH��
�\���ގ�aR�u-��"���c���`�j���Ie��1Y2*kd�	|{��V%�?�I} �ZM8�(�J��5M�>�M� 1��s8a�c�{������}4��w�������+�ʔR��>tW��U��$�ߩ�p���
!gy���/��+i��VU�<��J�� p
�~	��ސ�Zf&K�:ȧc��v�恴'fHÄ��������ݬ��lBzj�/L�|�Ҩ�̟��q��������xkz�x-n�_�PEI�0�VV婿�4@ﰌ�P#
MDk�N�GL���^��1vf��FDN�6�D���B��ZZc�霈6����kD��&ϝx�_�P+�GROݶ!�g�^�P���L.��kƓ	!����~�W{<�&���d�S��,�>Nxoq��3�����^o�2ƴ�tF�>g�*�C��O�5k*P�}(P�k*V����yt澈ʽ��""��Ҡ`�4����/��Q��%p<Y���%
�~�I�YJeb���uI��#�
1�9L��?}�BF&jL�(s�� }�0�ϼ���+Q�j�`��/ި%�vi418Rmѫ� ��SO����قlVm��ß!�Hm=|�R��E[l�2$�}�B���3Bkk� m��رk�ڦ���iK�)��=8�[޶�w3N����-����oޮ�s��L�ID���1�-�Q�����7���ŭ������o��nzˑd�����n�:��Ȳ~�Ve<�	��9mY���&_����3[���
�j�(����q�͞�k��(��_��|$�|zM����v+ԍ��/�g�EY��ka�x��3�d�^�y=���r�]��f�h�����_��3?���B��^[�`��o�v���������T��R�Gj,�a�s����{_���GɈ��{`��4bF�A�*V�Y��VaM>�7��t�$�Ʉ/�&�g�&�6���t����i�RN]/#��#^���,i7*u7�B���a#wy�S��\�6,�`�^�8ՌP:6����B+���W��U��Fp;���)�?�~j�`�L�'��s�&ї�Yݚdu��W��+Z�\W��O*-1+��Mz}��8�k�2>.���׾�a�p`c�{ǆ�5�H����Ev�b��#��$:0|#?n�Lϯ1��~MwN�'�ڼ�c���4U��'�W9ew[R�l��&�I7�-(���6�9C42Hq�]�3�^Q_� 7�#��w�qhc�v����T����m	�0%Qn\�<AϲlAʧ��[������@�|*#���!�g�G��5�}u�B��� ��)�g:�6 �����k�MQ��)r��l�ԝ��,�_d�\j����2���Ym`�$���Z�*�h���l��$�����[I��x�}�EI�M�z������C:v�d�R��RU�C�w�9>On4�[�'v�Q��?��F��G�d~3b�Nz���~��=L!��A���e��ʫp�w_r]"�%�v��tx��ӏ�N�5��uL���;im�w�=�F��R�!<����^�����X�S<�+�:�L'R�;K��b,���c�<�Wn�p��Hz�J}����1���b�Z�&3Fw�<f����`�EQO!�jͧ\�+���60�\i�˅d6���|Uo*�^�l�ޙ_���; ����*H90
 ��"�]V�0�qh�р=:���-ܖ8�X8��*�'�]����4�v�js�WZAE\z]
��C�S/v�ID���7��D��bM�� �D���0=���\�[��I��X~�Z��=n�Y(0�A���*�(�r�|����d�7���6t��5���a02�3��PHy&���p�i�:ԓ������8R��Ee����!|80ǜ�F�ZF�c����{�]׸I�����h�<Jӕ�K�����&sR������˲3?z�c�;����#�cp(�^(��ݍ��L�j]ɧ���jO����;����eN�S	$��Pȣ~-��v����ޖ3��	l�?j�t�VrǷ��̩�Ŀ�/8�?L5���è�'ɀ�{(����5��ѯX��pw�^&0���l�/.x+�R����V�ǔl�1�ԥn�ڡ0��a L`WJ�9b)����p���dsc��q؀JPpX?��Z���W�2�UZ�ѭO6��΍������_�κ.k��lj���\jF�any�����$�M:"�:L�|MyAo�EK�K�?� X�9�0��d2<x�(P�aL�:��&}���{Bhۘ�/�S7H��X�Dp��.h���Q�W�m�u��16��
�6FT��G�.W#�14r�r�0V|�`A
�$���Y��h������~���@�Sc�LԢ ���ȩi~�(t�t�n`�)5wE���Ԧ�A�i ��G,U� ^��&J���
�����u�g�1w�S@$���E��V��'����q�D�V̶�7<���LL��!�ZB����9��#=ͪ2���,�
���F�f�B�4"d4���l��bV
�s��mҥ}	=�)��>���.����̺c�h鿇��F��̱m$�}��N۔�
N��2����Q�R��G����D��w�ū��z�*y��#J��?�o���EE"��
�j�-X�n�	VؓQȒ��;���W��fg'�����p�~J��5{���\5,�Zz^Nrj�T�r _��7��P��uŐ���h$T�jk���޹���ȾZ�F1^%��}����%go/�B>�8�|��Y{�VN�9� �@�.�T4ʶ�2�;/J�
Q����0B[>r���Rh�4@2B���B'a��2}�W�婤�-@tx��u�T.	G&���T;*-�J�.Z�a���}��g��
��b"ȱ�d���W:pp3��u���@9�Vd�a���Vi��)x��N�����drVP�j�á�@� Q�HZ,y-�CqnE�9�mU��$���!����<av/��b Z��������Ж�`�EA���P���d�Yf���(��ӛ��&���ƌ���3'\DHމY����-l,,���i���E�K� ?� ��`o2�y@��U��h>ʺ�}����w�(Rq��0G>� ��sS��u����D�4M����5�KS����m�#��>*��o��_��D�
��-Z
|��Ȗq�����bl�U���X� r�~_�9���ldK��Ƨ��vzV$�b�8^W���������gTVl*�j�L��"�﷭	���b��z���p�Rx)��zoa-IZdɋ���ˠ�V�e��{I�G��#%��RkN}����s��vEDf�F�����!�D�hEBq2|Z>�<���Q��`k�i��`�xR7PF URʴn�V��Y\����.������A��/���(OW�^+&�F|d&Î����>I`KqXr������2��2���t���g��C�`%��}�P<�(k�E*��rݶ��y���e�E����U[`��6���/�p���o<�W������_I�-e(���4g�Hr�
 LGb|?��=Z�j���(.�� �jjRi1�y�3Q�N�`>1Mޣ}v��W8�ϫ��.8ֵF�
��l�C���mk!�1�=��k�m�������~<.$xo��3���B�� ($�����!��DL)���8g����N;C_X�(m��U5B���m쇯�D*���,���Y0i�2�Rn�@�����
����1��ˌ:���)ޤ�	�z��ITe��!��`��Q�&��n踂�[��)��]]����:k^ɞ��nу��%�|?��zȤ��|����2��ʔ��@Q��Ͱ3q�N�/��Ƨ=�u�V,"���Lf�jn�@v��3Z�鏽H^6i���;a���v�ʝ�b1,�Ԁ�T4��RX�j����k�{����R���Eu"`�w�b����뱔b��Љ>ÚM��L;������g��z6qw�t1j���NX]2�IS��]�,1*��IB������ow�8S��K��D�`_�[8�':��D����K-��ϻ�y��f�p���㫯�?EȻ��Lϻޤ]��&�&|Y8	�u`S�6�=�z�5&�\���Oųp+�O~z�I-8�0`M����-Ų��a(g=p�T���C���Hp檻`����k��'�$uӐ|����G�1/�?M2�,�BI��7d��"4���'~�`2@R'�+�&�f#��	��9~��H���.��^�� �垓�P��s]�Q���"�T'N�˾�	.�b%ꭴW4P��j�ʂ!(����>�:�;�*~�������%°t�u�aܬz %Q��b!�6[�G�{>�k�S�L����4�ة[,�>�W���4qY��~�t!;���(�5ɂ䣛U�޳]��	���3��m����M�LB�A��E��v��q�����C��4���n�d������RǹC����Ud���b_g�z� ������փ����C��X�p��r؅�%�I������n�@N�����q��Z���w$�;Fzy��\T�ܑ9^��Z���_.<�a�:'FUR�d8�צ����hc�q���vp���H��EJ�:��;�%#����p&.P���ЀIN`�` ?O�O�KI\*u��t�6+��iyw��cP��A�/*~�Hl�C�_��;��!�)�6H��� "s" ����8q�N�ر����5�f#X����Ebq'Δ�g�4 ���L]׍�A�Qg]ŨH�7�B�μ%Q�D+f�7{4I��fb��( Np���Ӕ�O���6ɜI)-X����O�n=��0����2����.�����E�dD[��oe�i�5����|�j®�I�+t�a��lZ&�
��:/5����W�S��҇,S�iƍ!��=0b�ٮA�F0�_�Q{'�b�3|��u)��%�<�7��F�s����UZ�����W�lu�����d��Ɩ��T��p�����ǽ�]�z�L����ن�k�;\� G]S$4ۯ��8~^9�����z�
x��D�����t��r�%z��/���ژ�e@��:p��T����6���av�B�5���LB��p^! ��]s���X+)�F�k�V������>�n��ӡ��"�'pL{ZJ~.&b�W&�2k�n0�s^a���.� �XZZ%Z_QJ2�i��o��lj�6�c���0b���!6:6_��.F/nl�ý����F�|<y���F��$��"~�:�{+|��o>~K�1=��k�X��_05�2��k���>�ȐՇ�!.[��K�h�t��J�7�<���D�G����p��Q1Sumx��Lt����O�3T�\�G��#�x�rI�k0nh܉�
q;�ߜ~Y�[IhF�Y��~�FY@x���g�J{�ޣ0g���t�a��i=U)���E������ҕK���,L�\�����J �b�BC����~��B�1�U�@�M�@XyV���b�/��Z��:��^�z��V\LR�!�U����1�5[�>����P��T�lf��	�=�!"�\@�<�ո}ĺ�ܽm��N	x@�����.=6�S�wc��=���!"y��'$+�C�Iz2�e�V�=|'�����P�"�+�/���������"߸�M�ZT+�f�E ��EH���Yn�>3hR�M;�l��-6f������V�~EÞ��4L͏��\Pn�Z��$rE������K`��Y�T�a��Vh?�Dj�TN���q��Y�F,���Y�m�O�+=�o�3>��x|@���(�VI�p�[ed��3�4��2%��Jp@��3���I�[9��+n2h:�	@, �Bn������.%����<��xY���o�G���2OTv1����.U�Pa��9}K�o��O
]#�"��Hd���W�ɩ3�'ڂ
$@�P!ɖ���ͨ��i�!x�^)���ގ���Pk�üc�r��|պ,�0��ޠ�ih-9q~�U�o��&oI�� ��L[<W�>/&(�	P�Z�Y��C����C%�;��A���P<�_?�f��=(��g��6�aO�gDZ�|,\�u�ބ�>��-'�ټ���μ� ��T+�j�|��2���O��"���5i}֘n��8(�8�+a�>E�? ���sn2=�Y�ڞZ�G� 4��p�����l��������4)��k��욂w���<����
ץ��QO�/�j�ݡBUy�k���� ���~��H�s��Б�K�ԍ�Y�?vU���\}�Ic��4F�M���"lE�yj��9��Ѩ�H�<�Hg��|s�����+�xD��z���-$@���g�fi
V�A����C�`8#@ia�=NXIٌ���yJfG��0Q��snD
�!B���Z`���܏�-Bk��Ex�pPat�RE���=���\�/��.�0��I�b�<�0���Wq� &c�da�޼2��>Dh�q�y�>ӫ�CTj�2|�t�� g2��C�3��믂P�Xb(���*�[ݑw�y�l� 3��>Ӟ�mu`~Ϝ�1�/��{�u+�<�EN�[YQ�0�IrJ�eػ���?����
�RVL�[�?�Ժ8�j^�(��x �`��"ҵT��QSS`ټ�ޞ�v�>8Ƞ���»�<+֐�wE��l�:���7�!9;�=zŭ̈}K�;�D�Y{$P��<�*�ۯ~B!�9 �����pڜ���
).b8�ԇ��N�d��o�C9��R��}z���SD�1
�'����$��m�������%�]�̓�ˇ0UHJ���>s�$u�t�=e�|�\>2�_���&�g�sn�[�Eܷ $\�ެ��H��ݞ�c���3�՛�|Z_zC�̒W؝����ex��;��v����r��i*C�T#"=͖;ّ���=f��h��{��՚�3u�E�8��^ ��֭	�N�yv�+���wŏ�fTO�R��~j�<���S�+�{���ʭ�P� �`�q�b<T��䱱ϝ���`~>���*/��?�Q�^gx06Ltl��̟�RNS�����Q�,L��*k��Bu�C��?:w�CWS��6��|�`�p8��:,���̉�c�����]E��r+p�v��UW?�19�rDL
p\���$&��7Y��u��QY/!j�\�W(O`Z+��
z3I8<�h�$�ō|sac1�p�f���;�`��H+VȻ{$�ף���$��|Y��B�1�� M��/�]�ڲ��ba4�d'�[�R���f�i�̣��#�E����9��IH�Jl�)K^
� ��}�8��g�C�,���]�T���/�	�1�%ǅ��rGٲb��]gB�������6@�*�O����9#��+6iu�e�� ��x�](6��>�6��k�����"4�������,3=
�R��Ꮒ���Y���}�SƢ��޽�ע�S���8F��Ѹq��,�;n�M�>��|4�����v�sm��ډC�<��/��n�'ݬ���D���B��KhՒ�hd�=jbڟ;z����9��s���Ӆڞ<%�|Vp+X`rS	�%�<[�����	��Nݧ�+���bNc�#�w���FUz���F�,�V^�����$r��ޭ<�N:�_�R��Ք�Lv{c�b���p]��H�=�Js���Ö�`���:�&)z�����C�{L�O�5���\e����5:6&��iԥ"�~�n�#r*-*Y�l8� _-�;�A劄�rH�eM =u4"��<���qޤ��sI��|#K����X�0��`O�'�^�B:�4;.��FO��A�f�]�i8�R�*�I�,�UDf�7�E��b� 	�b�і������Id�(X�Y&��;{n�0`�8�M�'�q�ŝ��dߞ�&�* �5�(�ėB��)A�����l1	4�M�:���js�n:��4��D�(!�70���<[MFw3W{BC�׮��P����.<��(�A���`	��X���t6����鸠�ف1���6������#e��C�B�<]w����lN�↨�^�&��_uS?d��F�~� ��Ȋ)@��_ɟ3嵑�t9�$r�H��}��� � q�5�7�C�Fe��g삊�5)�%aQ঎b^>�LL:����+D������V~0�������nѨ)���3��k�L��J��~bǦ��m+Y�	�SsY��Nڄ��ϩXu!Z��[���ˤ��G�6��C�C���wT�Q�%_���.!�l��Ē�F���y5�r��$�g�"��:�˨|��;o�K�7d��0�XB�_02��22K�_���y�p�����B<4hQp5�e��7>�̃�D�!�S���.Q�n�m3c�g��� ˔ńhT!��G3� #��6r���0�}��g
��۽��,Y/Ӷh�Av�)�~I�@3mx��[�ϵ�~�T�ryt+��d:�)돝Em�F����N���i�,�OTI�����J[~F^���������q��1��Z@Z���;��VX�����Ov�g7�9g	�	��L���PޥR�6���Y�h�(4���k�|���8�
"�N��󬸘̅�i�m���	�Ֆ۔V��۲.o�H�j�cԴ��}r�����'��$���D9��jh���l�ޭ�HN��K�j�'ϭ9��������긙Ґu�N�ᚤE���"��c{n{�F�\S��8;	� �M�4fǚ��M�����~@��7T=�J��\kУZp��r Ӵ�஧�`��Xү�=�C�hZ�\jaEpv�M�Vl���vF'��޴H0�
�Fu�o%A>�n�|{��ԏ��VDt�������4 ��2�(�JK���n�'��[4�Ϫ�9�h��@G. B颟��i�4K�����۷��bxU� �G54uޟT�X%���
.P��a=c}"��kF
؊�"~?�d��*WpC[3�Ժ�ep�@�(�<�QyK�̓ÜiW,x.C���T��A�P&�������W�K,�xE�y�.d��9� 1Up]L�A��H����L<��Z/��^ ZL'q���8���ן��oA(_P�1)�Z�fY}6(@��,eO��-3�B�}5��\z����c��-�)+��nu�_����]�0����wP2;�8�:i��=�Hʰ��}����U�(��&��>�YF b9�s�n���b��5�܂8`4������O�|\��蒯3t�F5��O�z���
2u����J�X�aUT�u��x* A�^~�t��m�؋׬K����2�v0�Y���\�Ϛ����^���5l`��j���,�ăk���䠓w���0<.��mx_��z�-�E�)��R�V�=�ERް�F"#['@�5<N3���6�0�̈f�W�r�g��D%�FBg��Z�qS�9\;�T�{k��7��x���P|�R��"�DP��O���4.��WƤ����q��jW��&>��d�}B�͊�>?��q�����i���2Wk(t���g��tC�&�F�P���(�&R*���l�y%�A���X������`9�f�L/5s�P޾<
T$��.����I��te�o
��j=�>ot
°<L�tL?N�3�j]1�(�� �vVH���/�SQCw�`th0ޙ"�vz��8�j���$a��k����l'Q3��!!�d�=5�̣i<ʶIS�4��$��K�f���d�B|� ������]ٍ��)iK8U�@����N��o��^�|�K ��2���/'D`�G�"a��b���}<��B��6?c���`!/�gV�˂F��؟���?���`e͇T���>@V���&p���.zr[�Ȗ�{
g��b-ăec�o
�~��9��2|u�z��'�29_�>�� |��6]��氩�1�����ϟ�=�������.}�f�ξ������G�3�B
���I^�e�@��雨v��5�j��J�'Tj�RN�lj��B�$"��o�{��nĈ���`ы�b��<��
F��'+>��օ1)���5ֿg�6'��t�W1�:��NN��K]���,g٠*�EBPH6��xwJ�mS��G��`�)
8&��:�.;�uv�P�.�(���a��pleF���?;��j+LED���&�&¤/Y�E�u�&l
#���\7�O� �+�c�z��D8�j�����W�h�"a�kp1����I�����H��黖���Ah�{U$띎|����=��1��!M�W�x�-hi���4ec'��V>R��!C��� T��M�c�9��SHB���$9^b�� h'��S�����P����KT]����<	��%�Aݴ�zj��wC�8��  �t*��1��*4+��R=��TA�¦!ufR�2 [�t�XO�6�����!k	/�BO�b@��N�',�[a�M��곫�cT���(���Ϣ�v� ��=A��Y��u������b��0MqP�鷁��{��v��Ȉ^ЃM�C�����n�䅬)�G�����y�����M��d���bU��z�\�/��Lы������BpF��rά�%�O`�%caФ�rNؐV�c�b=���w��F0���&*��Z�^}_N�X�?}�<�-�:�5Ri#�M�����c�፲h)/p�H˞�J�#&������!���]&$�J�M�݀���SO�ν��\\��{�P'6!��i/Z΅9Ð13��D�*4<�lsn�_�E�;�!E��h�Hj0% X�".2���LqU�3�w����Xi���{\�'r���4v�A��q��YaAV�a];J��m���ē�fD��
7�/:�Hwb^pE �'}��y\�Ece����I���XOR���GDn�0�t�h����,Π^�T�Fdz]��v��+5E��Ĳ��¤���+��Sz�י� ��:��.�%��Љ�=�}[s�Գ!-{%0�鹮7ȀF�(����{]��)A��+o��9 �<aV�<0��@�W{֜��zr��%������ ��2t7mЏѝ�.]����W]Z�"�k�^Ć����5Q����SZ����b'~����'��%2� �������pU�tT�r|B#�����Z����s�0��
'+���ۍ���U5����`��AJ�^>���Z��`[f+_��a��VY���+��t��n̢ۡA%��мL��;JtCb�ߤ�u;��3sT�\©>ۀ{��X��ZU������C6�chΞ/��2�l��_	�l.���ldd�-A+F�y�o����	$%"ts�:�;v|�Z�o��wK�]g�P8X���0Me�2���:Á�c�����L�h�ۀ�7�	��I�D!*J����|q|Q��m�	���P2�{��T\U�G�	�#�fr�ED0��V<g
jȽ���Yjj�h|���{�~�I�@�)ٳ�p�q�8�Y�2/t�M�_Wi)FLiE(�����ҋp���@,����j��~�J�eJ� ��$t�tlr���1(�,@�s��6��V���@��d��0 �/��D�wL����K\[��j��t���7�½�90���6�3>�"u��g���O��Y�mc��	v����b.�C���h�c�_��H�ד.�b��$a`�?"�):��ov��n)�����؋:ܥ��H��<��;�ָT(;���ڒ\ʥE�4�����wnv��pT��9\;${����f�d������A�)~;#ձ��N�)\�RZ�N�r��ڴ#񤧁���
UZ���.hu;=j�U^Q�����ȏ��F"���R��K(a�o���>u9�|�A�*�V?ԉ�+�_��4 �2�CJ&���<s�گ[/V���$�h�l�@b\�Bd�m��)��o���(~��� �>#yx�6��G�q-P��T�_���.K��a�Xl}����o�
S�"Y��d7-jW݄3������@j �W�����^�WiU�Kx�G�����uؑP�F����h��2O,*��`V_�9'��U+kF�\��⒰����<�Z�/\���zZ��,U]�STB����AC�@Prw:�Uf���(���G p�W,g��1po�\���zE����-�� �	� ��A����+k] ��r�2�dU�����X[:�+r�}���9�(#�5�!�s>��, �Ds�ʹ�OB��ܽ�4�J����\@�oC��Z��*^�!}���:�xi�
�dh�ǡ��e4��l-U/��69� �h�~�/�J���F=�K	�s�O��vf��/���� �C<ݘƻl{�j��ׂt�ľA4�~���r��⋬�����xzw�z�|-�k��<
8؜ZV�Ys���xM�#v�W�fN�&�q؉�G@�f��`���T�"w�D@d�B◩Z���tSn���k�K����lx��P���R;��kӡJ 8�e.�
I������Ƶ��CWg��&\�d׊��h?F>:؇qi�W��L8�J��22�t2��gh�C�9��t�Pm��(���*����G��y`�j�6(�����f��`�@��gh/�V�+�<E�n��$y~bI(��eNC��ᵴ��
�.�L���?�u�.Vcj�$�(_g� �����
�kQ~��`4�ޔaFv��L8>Td������7�Fb�V�l���+�!ﭱ=���̾u��1���Y�$�&�r���9�B�|� Y�?��rڒ7=��2�)���8�͑��7UNL�6����y�h��Ev�i$�8�.D� =��V��X��������꺊�z���T�9��}|[���Z`<�Z��j�e��M�*�ٍE���&����饏[lY��~��8%ľ�U<(O�yۭєS>�K��|��z99�����y�aǛ�k�1���,���d�l���A�J<�=��7��(��&f�0q�Q���K3��6�.�^Ǎ;�L�6�Ov��s6�(�T�1wR��j� �_���<��{�~�ceX�v��`�� b2/�fαE���ߏ>����S ��{�P��gn��6��t�*���NI���Z�r���,��>*aťB+˘�M�+w�n|S�n��M`��'8A�W:"���P:������á'Ѕ��w��p't���?�d�E�L�8t�.�5&��cYI�u���ہ�F�Q`\C6�O�@+}8z�� 8�>��n���C��a�%�p�����Π��H����R�̸�U�$&�+|�q��8O�1@?CMcJ�ܓ��ڨ=n�hLp4A��'O69Q#WR8� ���~���!�>649/!�H�O����^�4� #xh�n�L�]VԾ�*D��2ST���ּq�	?�%=�����X.�S'Ga�����,V*�&���L�o�!uAF}�1 �k��S�?6l�l���}k32	ǽ�&�=�ԉOL,i��H���E%�Ѽ���;�bE���+�Tb%�ص���t���G����
i�1ML�[������v�DJ#0��>��C �]�%4n��^�G���#��Km�T����\d���b�p�z��l�j ���6���.:�Te����pa�rIp�%_���`�|�?& Nә���-��ؕ��Y�w��EF�����b^x3�k���;�<ĥ:���RD� ��3����Ic��v�ç+p�K*H��Ji���y�9���l�p��&.���K��zl��zO��~��\�C)���6�i�.z��"�L��h*��l�3�_c��;�!A�:hJH%! s�~"���՜.qT%����e�r���w!8X$��˖�J'�ߒ����4��،|�+��A��n]�JD숲��?����"Dܸ�7L�&��b�� ��}����խ�
dIچ�X�jR��s)nNG�0��T������l�{?���yd���{�Y��m5 L������ڼ�F[�=�W���G:@�"��Ф�7������
/!h�03Cޮ2U0F-Uu���{x��פ�
�QJ�t<�%�7���@�J����X�����O���5���ϹY�J��I⨪8�>]5����о��}�������Q��Su$�<ր~����b%_+>��B}�U���+9Gtogr� 
��y�̕V��62�+���e*㨼"Ҁ��P����5x�Yћ���%�^�<���U�+zӇ�S*V4�Y�X��/*nǼ顜^��MU�L��J�sb}�#����?�"sO�v��1�6��X��Zа#��n�Ao@�=`36�)��ޅ��i����_��.�}�lV�����F��y�I֕w��$1Q"���:x˓|9�oP�8K{�F�� X�<�0h-o2(���Tt������@�l��|&h��oۛ�=74 ��/�D\����wM�QB�m�������m�{�KT�6Gi=�#�*rZ�P0B�-Ů
��p��Y�!h_���,~��@�����'�4� jךtR0�Z��)�(5E�_��e�����m	,�ɰ����xJmnԺ���n������@�1c~2@�Sg�1q�V���{�ݙ���Ҷ����L#
2�F��La%�������[��k�������.��"Е��m����!�_��m>�!	)�T�Ζ�#/.%�M����c
�,�sų��|̝��$��\�:t�v��nD�P��>�������������z��ޢ�]���XΒ�E�]K��6��Znq�'D�U�~��;?2ؗC��f}Nn������[5~6�Z�����su\��Zf4�r��^!ϧV���<��e߶��wh���jW�,Z������*%�Fv�j�ՠ��|Eo�>P$�|�Y���V:���l�ϥ��46�2��J�����]S�[*␪<0�hk�a@}��Bߥg��j1���U��a��Em��YPx�8���RQG��r+��T'n��Ei.F�a�U}|ӓl
ι�"4M�dr��W��&3����i�@%8^r�_o��9'#i�1xdlJ���!�Џ�P�5��w�Vm�<�,ei.���5Z�m9���U昄�w���9�n�<�/��b�ٰZ"��_�n${�^Y��'ZA~D�P�C�P*IfΨ(�;<�b����J����u��\����u)]a�-X���$���U�ұo��)PO �m\!2��1����s�sʦ&k}g�t�<(�K��oK>V�� ���s�F��A�������4��k��Z�$p��k���̒������K�:߰�c���
�s�Ȃ����ڢN�U
U�q\ wP�~�
�����K$,�����v�UϴN�C������+�^�y�Sץl��Ej�Ȉ�OB���7޷@z�mf���<ˠ\��x���z���-���w&�7��V̕�����3t�#�Ҙ�N�U�����ӭf�������(�D[MhB]��Z�����ju����k�����x>OwP���R�R�h�F��"� |}.����Z�ňm���e�W�(I&�MSd�F�X>5@�q�O1�okR(��Ҫ2�?tmҩg)�C�lՒ�hP(��(�0*v���"�y��������Ϟ�E`��'ӂ��/�&���<��,�,:y+�I���e	7H�� 4�4�A
x̹L3m?���)�8j8;(�+ �>����3Q��`��ޏ�v0,t8�]s�&�
0�!V��jl]����U3!Js=�#��١Vʬ�����$������.B2= �h�8���2-��|�)�5�8��z���cN�BKC?�����A���D���s0jD����W��CwU�V����,@>�e�@��7��;j�xҨY*��!7�u�U����e���эt�,��V&&!S��0[)/$�q7��o.������ ��tǥ��3���|���z��b��Z�Դc��6�x�,m����8l���-���Y=^n�B�(�d�f����_��63�*ˏ��'^����Ļ��nv�>���"[����T��oRD`�js�Ӭ��ş�XR{薔ʾ|�1�%` b�̕Ak$�����]Ϭ>�f��;��p	�k@�g�p6ݖ,tI�p;�NDU��蝂 �,��*���Bnk���Rw�4�S������`KQ�8\�-:�b�+�x�ư��^�{����\�p⢘��?1.� ��L�L��=&���Y�uLz���(|����\~U O1�+x��zD��8m��J��M2�	QaPipg[x��s�qK�H\e9��;�v��jO)$a��|*N��3��1���M�ܮQ+�#3�C�?4|ŷ'�}�L^,R�0�������*��9jldHx���@^�� ��s������~��%@���T��ַB�	���%���@���������ª����'��*�A��*`��ݟ:u��ȝ� �_�N�)6� ��gŝkN{+�8������D,��CŐ�v~��mD��1���'���D��R�s���I�b��C��)���wM'�.�-| ��
�v� ~�[���TC�����2n{�g��9�}�J�������;=d��bK	�z\�&���q�DA���^گ4�DvEp|�.r�S{%:պ����ڛ�N����<vU���}�$w�F�m�Hy�����^s'��ʭ�<2z�:l�RHΔ����c�?��F�p��zH�J���T2�����&���k�5aG�̐O��Y�0\˴�:i67
i�"&����g����*�o�l��_�>�;�Aي���H�%A �;�"Y!�w�!q�I�D�P�m����k�Xߑ&˱��'����^4�Ìvå�Ag�]�k`��R��9���D�^7��*xb�b :_>�"�D�;PR��`qI��X���ɿ*n��0�٣��������V@���`d�)��vy;�o5�W���6aڗc�M����m���:������_п���s
D��a�!���0μz�-\F��K~d{�P�����R �Z�<Q
z�2 5�q�� �5C,��U>�z_C��(��T�
�*\���ۨd�����]�8$f����o���jS�����i�~t�x����PB��ɰ����<jt��rr���e'��п���¾�&@���M;�w�.�:?��'�5S0z��]��w!�^��]���n�+�R�W��V�Ɣ�	,쪕�n��S��ק���L�C�JjlbXSX�jܗڶ>sJ��_g����X�69ZK���-�|��؜�6���T�|��$����_�9�.��!l����cp�F�(�yFDh�2�g$L�J"j�4:S{|t��o���Kv	�A(Xs�0�62�qr�𮕁*�B�A�}2��S��h�#S۶��7�V]5�D��W�$y�rIlQ���md����-�q�lV7ET��eG��#��}r�r0�tUHn>
ㅽKLY���h����~Z�S@dG��x�g�������t�G��U�m)�$E���-�ҁ�`�,8��%�k���Jl���͎�٢�j�w���A1�vl@+S�,dtViC;N\����&�R�������L�t��A�ZcɆ�W��=�����s����1�M�C�)0�"+>z�(�K������V�m;3	d�������w.��@�?��c%�!��K�������$��զ56���)�Մ/Qw��"뚎Ӊ��=�~ѫu����O�ʱ���D*�R��E��R�1q��4��nlR���V�9ٯ;Z	���WxfXXh����wH�~1|�Hr��{��\���Z�98r��y��q-�����ɇ����S�tmNh�uVj�֞�N����F����h��;-?���o��,>+/�|,�7�`jV5�'�Ǧ�բ_4Q92|�J�W�������[%����[�h&z�@��BZ׍�����_Π^e̼�����xEZW�۫GvJ�rTb�P�Q��.A�aN;}7���כ
I��"�d�1�WAp@3��E�v�@�o*�Ų�"����i���x�����|Ŏ+g�PW��(�^����H,�q�J��U4�9��6U�������j�Il<C��/�ґ�G�Z]O�������Q����wA�`P�bE�Kc{fj&"(q���}���M���ӻI��
\Kx��p-Jt�d-���?a��4�Ҍ(�����w�h+d2L���kv,Ȏ���!�"}BhW��;(Y��	>��� ��ds����Ea��ƒ��3��4T���m�)�n���H�� ~���z솗N�K����ݿ
C���=�>���O�ɷ�U年�C X�~�� �ؼh�K?�z�E��v�e����eT,���0��-��l�Zjx&�*�"�4N���[�h���A�Y�A!x���zyu-��ɲ,���˒V��u�V�n�#�!�Mz@N��4��X�}��f�"��h�X���`DvVeB�ЙZ�E��P�%�9k�n�Hx��AP̈́�R1�[C���d䰛V.�d�ƵS�(vK� D�W]�n&�_1dM缞>0ȼq�*�*�|C��@�<2�At�*�g��oC��W�W�4P�U(��A*�O���V�y�Y��l������#�`j2ӝ��/u�����<�>_��o�t)Iޫ e�J-����ں
S�PLn��?� $�*jnkc(ՄZ y��H��h�Q��0`E+*ފ?�v��[8��F�"����t��i�1U�l�Tg�!��=f؟����'X�Ŷ,$<;=�����C�B�œ �"��S֔ڈL����)ۛ8&G����N"$"���8߼�J�����D1PP���sM)J��	s���]�@_V���8^��sH��_ ��������`�e^h�H�����V'&��L�_]V[D���}ІJD��4y�r� �oӹ�JJ�����|Ɨz/<B�����?���F��'D~���+�ڹ/��Na�@�=9�t�}p����of�T��Ao���3��Ǐ$θ^}���¶4���vӫ<�)/��{7�T�/�R��jN���չ��r�j{���������`"��b(�Dت������ށ>�iG֖�n�+�����gdy�6���tX1���sN?#d����=9g,�i3*WL*B�0�����w�S����X�1`�8w:���щ���"��-v�-@vp���2.�?����L��\�d�&&��Y�OuT(���@�|�\���O�4�+s��z�(y8(�'�F_����w�aO��p���8��̯�HUg�� '�@��Ei�$�=�|�J$�.O'1�=�M����#.ڞH|��?4�%�'��G��R��YR� �8�y��.����9��jHժ�#�^s߭ �y㓤�'�S���@��I��T.B�ֲ3:	��U%�4���N�N���ɾL�C^�E���"pk*E}�����[L�|Qu�V* ,s��I�P6"g��"��ki�ǳ�I��3a��],�ww�>������*�������t�|kM�ʆt�iڳ��w�����i�'8vMF�h)R�L_|v�����
дe�C6%��nV۠���E�>�ґ��
�o�~�ad �yb��=z7T0������k��
_�
r%��^]p��Cr?W0%H��m�u1N���ގ�N]�Ew�4�F�Ή��RMܘ�1^n;�!�'�p<MP�:��R�,���'��d�c���yepI?�H��J_q[�/���L�j����&b[�^���u���<�O��4��\Qa�!|�6�i@7҅jB���^T:*�9�l$ _���;���ƢH�P� ��i"��R�Sq�%ʀ����h���-ֆX�G���C'��8���94'������{%Ag��]l���B��5F��f�DR�67������boQ1 �*��=�����ڭ}�IP��X ����+Hn��0Lj����
wr�1a�3�dK��qB���15v�[���s%�r/��Ms���S:�;��Vf��ڊc��N����!��0iV��(�F��v3{�?wךXV��t��^<�p�-���̦3����Py��r&�U,/��b��k�/�u������L.�.�q]�w�s�a��y��5ʝ���S�dt�2�~O������>�������`t�}"r����@���Ij�ls��!���3�2`/�,�U�vq�5.�J���=Z^�+��E׸��9+��C��\�V���Ψ�E�n�P�Rq9�þ^L�J�Kb3"}�Y��u��sE�º+߀�NNX�}RZ��y�m����s�56��~ί���c����u_z�+.���l�D���7�F��Hy�^:��U}$g"�T::.K�|�\"o��BKq���a��X.�J0��2}��)'�e���[Y���=h=���я�7*�L8[�D�m<���meQ��m���ӊ���b1�T�IG�V#��r9�0�{c7
~�V�&�Y�hM�X�1~���@ T��,���I��l໌t��^�Pn�)WA�EY�l�H�������;��,sĢ�[�����J��J |�/c6��t|���1َ�@�r�'w�Vĵ2	�d;�	���Fe��ƗLY���<���f�a��ŝ��?�N�Y��蘾�$و"����3�9޺Um���	��bGW����.۽���$�c@�>�i��h���'g$2c��0u��,$0���+�Jr��4gb�i���V@��Tu�p��LQ۸�&ϐ�P��2Eg;J�lˈ��A�ng'��mX����;u ��92�f3�r�9tL�U~,�9��C�6i�\טZ\_kr����ῧR%�����T0�/��h�B�jMG��9�B���`�eF¨� ^��������oo�>Z�|gF���lDV0�K�"Ǘ��·4l�f2���J�-��Z�/���[ Zª��h�0�@��1B�(��dL�� �����?�S��O&?x ����$&G�����T�5��B(.<L�a���}��	<3
�h$"���d���W�i�3������@�����eU���
�i�"x�Y��t��^�P�3�CF��1��uo,����nP�D98�U\T���\����$D3<~t/-��ձZ���]ߎ�$���då�A���PC?�F��fŞ(,#	������KƮ�!��\���kQSχ�-ΤڼZG�K�&�g=�V�&�c�2�o+�&#ȩn�ʜ�&}���(��Ŧ�>! N�s�����,�����n��4�(���T�mM�Hɔ�ђ���������v��M!��-B
��l��񔠶�m�D��U�>��9^ �
~� �[���w.oKZ*���av������� �:��r����X�l�zVj������o���O4�c��✽h��
x��z��-k�S��m��m4qV�m!����!3#�_l�{�N��Ì"]��[�f�i��ðz�S��D��BS�Z`!B�%����&�k�!P��h9x�(�P�/R�a�����ƨ�6��.�A����}��;CW�� &��d�r��9D>+pAqz~D��p�^��{2�t�tg9�C�2����AP���(��*l�����ky�ވ���4�w �`%�xӸHi/������<���b��o�I9�e~��2WK�*�?
.hwL��?�Wvr8jɾ+(�C- :4������Q/Hj`�V�ޅ�,v�8o�ݫ=m3�ם�l.l��(�	�! J�=!�V�ZʢG�⠕�$w�uC�	��x6B�� ����n-�����fp�)U��8�����UN]!K��(���7v���E���}D�'n�ͬ��w˔���6��"�I�?��Lν�ӠL�n����؋Y�������e9���}�6䎅��&�����[_ҷg��%zm�oj���j��ѥ���|��|�Sz��M���E�*<�l�;�";��=���[���'݊���=Kٸw��wf���bB�|:P3��,���^X�]��ȡ�UBv�87��[��6�UT���R:e�j)f���˟�{�&��tՈ�% `=4?b�g��da��&���>��z��z��O�*gߡ�6���t�d�̦PN:��kA���R,�ى*ҿNB�a��6�w�yS�9���v `���8�j�:�h��჻�<##���l�����C�pX`{�Mt�?'!B�NkL1�^���s&� hYZ?Au�M`�Or��W�G\��Og{(+n/z���8�l/�bW�l���@a�8p����[�'4�H�d���w+�� �=$ײ{|`g,�)�21Q�gM��\����~����o4��' mFB4RI�V��S��g�υ9�b�H��V�i�^��  T*���}q��X��s{����!Tɟ�֭D�	P�9%npm��� ���ʤ�7�����7�L *���>�s��� ݹuҘ�>� Ǧ��D+�6}�R��H*k�mH�.AM��o��:�,:/�9���V���O ��劁�.�WRF�I�שr����SP�x�5Ȯ��zM�������ӛv���4���oX�CQop��|un1
�����b��d��e��9�d;�bA��z<��jK�z����;�eϕ��g�p��@r�z�%����\���xN�t��fH�	��&�w��F�6��K��3�^io�|e%�+8�<hF�:	�R��9�9��S�#c�����p�gH7c�J�u�
:������Ax�&,��y����	^O~L��\�2봼݋6A�i�k~�%C�O���*�#�l_C�_4��;��݊K&HV�� �_�"��-��qV�zO�c����`�XU����,'����9e4b��M<��qtA±�]'��ٺK��LsQD�+�7���ib�1� ��XFM�1�o�Xl<I��X�t�ֿ��n_	�0�ͣ�
_���7��@�Kd����l�k�ϳ51�$� ��5�M*�0�R����:Q�?�������i9Ņ�oA!�f0�#�'F>�Y��{�N��KN�����%5<�3��(P>�'^�CF��kn�x���0K� �'�T�� �;� ��{�)��1����]�.4��*�U����_�%������S�4���~*���d0�2��-�f�f�\�<t�8�rh��� �F�Dj���v�˨�.ԀGf���ښ5	B��L�*�xd^:}��^�L�+�T�M�V�C�	h����jn��<��*��~�L�J`K�b����M���s@��6�g��X���ZA0�TA�򎤸v6��
�ʐ���F�_�Dn.h�l%#ę�F��y��L����$�Y�"`5:	;�|�G�o!N�Kl5���X�@0�E|2��~��(��|8�w-�Y�	��h�:���B7�#��7Do��Z��h��QS�5m�������gR��HTH��G:��#���rk�0s�d~ 6
��s�d�YVHh��-�w~ϑ@�\E�	�]E}���
��t#���Kc)�}�EW��cB��w:B���,��[0���^jJ"C�S��Jr�`b-�d��1�|@a���"��VHj��,�.���B������0
�L����7��$�V�-��̪����)�DbP���1��^"����v���Ⱥ��Vm�V	�S��׷��<.6��Zc[#�����C���N��$�No�+��هb���E�e�傯�%�D�ܑ��ϴ�q�k$����G�@�Ȑ�|�H��EB�1�Ed�j�nb�UZȯ�;�h��,bf̌�t������~'c�������f\�ZפJrg�ٴr���)��}X�v>M��~h�/�j����߹}4�����FA�{s������m�o�J2>�`|���Ԗ�V+�k�}��K44�l�2��J�#c��AA.}>[F�M�h�@�T�BP�^�?��[�۠��7�
����Vx�����|Gl��eT������.7�a�R}���$�2
?p"���d#��Ww��3d�,��@V?�Ã�৛�ʬ�iAi�x5���}���uMP��u�^�T�����,��^%K�J9�,{U����-��~�h��;�<�g�/�gx�|Z
����T��w�ڥ]�A/�OP��0�A5�f 7�(�Ƶ���C�Cf�Ɖ7�\�r\���f�x*K`-��`�uM`�Ƨ��B��W�{!���^)�2^H������_��w}��,%��(��P���>g�� 	Qs{��; �|`ܩ��4�������ȑt���*���HA�������߁*�ڝ`
�aYȳL��<3���U��y�"z� H�A~�[�1��2�Ku���;5�vw�X��?���!��x��o�r݄ɼl�;jn%��� Īڔ��8�^y�������wx惔zo��-FCI�(�h��gV�	���D�d�Q#�[C��NzN�]���N
f��͙�\���D��7BΉ�Z;F�`p��[��k�S����=xołP�R'I�FA�6Ia��xo.�>��kl*�����Vb�WS�^&��d��c��Q>&8bq�E~��#>y��6[e2�Kt;(gԧC~Ő�~�PY��((�*�`�ݳ�PyL�X���M�����=�`�7��(/kf��<�<1{ ��:jjF+I�ie:҃�M"���
	f.L��t?U8�fbj$2�(K"� U�b�5�v��QjX`{�>ހ��vA�j8*;9�X�5���ֲ���Ml.�B![�=ܡ��*�
�W��{�V$�Ϣ�����BC�A E�؉���~�E�A�)���8\@Ƕ|�8N�@�|T��{�߲Ю՚��$�UDgD�	�A�)�M�*���������>r���3�n��i��j*��F#���徲VJe�����E���8�&7���Ք-[z8���jS� ХĪ{��JS�eK6� ���7d|���z%���y�w�eX��n�R�ŰP�!��6�>=���� �5�f�����c��7��3w��}^3)��8���v�孩ߧ?���+T�R�Ijh��Kퟨ�d{ٞ��ς�b��`X�Nbe��H�1oA�.^T>��i�Lޘ�r��^gZ�/6n>tη��A�N5������
�,�i�*MS_B���9��wQEhS�h�oO`|��8���:Gw�15�w�Ҙ/$	�U���f�p���h�?�J����LlI����&���Y���u}g\�_��	$2��\/sMO��+iE�zU�Q8�
��,%ů��aŎ�p8p$��"<����H��ϻ/��5t����$Hi|����$��1��	MOu8��',ڔ�:�ԟ�4-F='��=�R����_��n�{��k��5�9tHI���Ͽ^)
� ���e��ID�N����K�Td]֨uz	�3�%)�[�Z��DH����3���{u��H�*�S���~s�۷�_Nu�I�y�� b���?�Q6ؓ�����k�Cǩ����#�u�&,��>�4�᱊��
4�1�����T�2Y/�@+��D���G�ZP��3;�PG֚�M��	���1��hSv{$J���*kdCl�Ɵ*�nu��3NbN��W���Y����vdV\2b��z�C4�Vm6�!ً�f���Lf�u��p��%r5�^%ˍ�LjtЫ��N��G�M��Ĥ=AF�w�1�Fwjr��dI��]�^d�5��8í�v!<�\5:��jR���tr�c�<r�/�p��HRd�JU�����C��͸�܎�&3�1Ѐf�O��$O����C�\�li�W_�6�vi��*���y�&�T��*{-�l���_Ϥ~;�aJ���{Hz �!�"}	�BIq@�h�wb�^;��
�X�~'ya�d��4�q}���e���A�e]���R��+]�N\�DȑC7�ӊ�m�b%2O k"��s������3"�IƋ5XV�ֺc�n�4�0�w>��x�� �(��%{Od��j�g?L&�5���9y��L��('��T�������:���̟���/�� ��f&}!T0�� ���F�F�|��{�}kא]Ҧr�`��<"x$�#(-�5�����1����&��;���}���;��6���6Ԫ$��]��@���T�Ն������=�<S�$��(�~r�N^�ˁ��f���L���t�Rr�:���́����4d�����w���b,��ld�5���чzr�HԦ^��n���|�+�Շ��lV���DGM�{�0n�d����9��L8�J�job���������bs;���p��"N�XlZ��D/���-�C���6zE�e�!����_p�\.CQ�lB%��4'tF��ryW�c�t$���"�5�:�J+|%So���Kg�\�q�X�?�0ԍ�2�����ے�������d~h���֩7 ���8DH���Nc��Q��[m�+��	����3��	ST��-G�K�#���r�%0.��)�
tݽ�SY�>�h�[��G~k �@���$�Fؼޠ`�V Ot��m�Fȗ)�eE�>�~!���2����,�>��$b���J}�?����e�U��o��?t�1OS@�����Vz�����I��痚��[���km�L�t��2��t8S/�����
)`���W�����0"<�&�Y���:/��Km��	��}x���3y.���pB�cv��_��`~̉�$hZ��&S�����Z $����*P5����>��O!ƫfn��D���o��ɮ�×E�	���3��n]1���[�j8L;�N��/G�f�5����'�H�U~"C��Y��ͬ�S\��ZR
�rB�ѴJ"���tz��(���H���}h�<YjC���� ���*Ȗ�mF	���֨��loP�e3oF�>�e|ݲ��1h�V&���g`��d4�O�2��Jm9�����u�[Rd����hW��@�"+B�+	�����p�/0h����s.xvv�,wG�����T��"�G.2p�a_�}h�C?d�
��p"��d^��W�^3z�-����@ק��[�ͥn�i|fx�>��x�Y�<��P� ��y1όK�y/�,Q�q�n�F�9�}Uҏ&��������S�<�z�/c�/�Q#Zn�r�0O�ڤo���ݥ8spAj�uPy��<��f{�(�������!�d�&���\
_�a���.�-D"���sԺA�����"U�}��YX�2]l%�\��p+ʒ8}�SO`�0(*&4��B>��� ĵCs+w�϶u�W
���4%,���\@�#� ��6�E����u�h�Q�77�'?��-
T�e�nǭ����:�<Uv���]�0 �.1~ܶ��1���K�`᧶�vRU|�:��6l����g��}0�?Z7l�j鶆�����P��vΓYj��R��H4hx�z�E-!	��cP�أevV����g֟�O#�;s���NU��U��Nb�f�W?�y]���/�D�1BI=Z9��ۏ�k�(�Yk"x*��P!dR��a�u�q��lb�.�[F��(L�Y�J�q�}W��(&`U,d��@�o��>! q0-؍[����X���2y8�tY�gog�CyxG�h�PI(C�:*bݎN�y�C&�=���՞-{�`��Z��(�/�i��r�/<lI�����e��I�Me�E��h�� fn
�uL��?�8jz�jŜ(!� p��*�
�Qc6Q���`�{|Hv�e�8��X�sjF�
֍eK��Al�x��=�!��9=��p�E�lʘ���V��$���y�BKB���  �6ؤ;E��[f��)ˊ�8���w7�N��7.�� ���-ᔮ��_�aD7��Ò��,�A༤*�=���^x�����	���djwſI�d��=��ѥse�h���a��{�{ك&�b9�`�[�{��]���En���C��`���[�J��Z�|�gz���TZԠ�Ǣ1ߣ����2���&:���*�=ʉh�.�p�дrf��R�������32{.���^�z�sMX�U�vĲ��:�Ŭ�T��R0�j߉���q"�C�E{�6��*�k`s�b��Y��^�l�1���Q>�2֧���\�+הpg�Rz6I��t	+j����N0M��!�~�n�U,	�*�\Br9�txw�OS�8�i�`7 y8Ȁ�:�EA��>����Խ��>�pΝ��`�?�z� �L���5�&��Y�eu8�ѕh���G\j�O�h�+d��z���8Y��%���Ŋ��a 9�p�a���G��ݜ�HH�	�8vm`���v�$M�j|� ��1��M
P8�Z'�I���_4h�'V��8��R���ŵ�Ϩ�l<���9V�vH�7�U�^�O' �늓�m���Ob�)Q���!ET��#֣�	��%�Gδ/M|�����Zнn���~��d�*V�贅���B u����> �m��:�,63Z�SL�k�߅�$�8��G=԰�o,p���/���|��� L�LB��w7���{-���嬳��@�l>��k慚�_�M�[����vvl��T���\C�cş��hn��l�nڔ�j��j4�̖կrgdq�:b7�z�k.���u������D��ꖘ0��p�X�r�!�%�`������F�LN��l��;�x0\�w�ߝFR�>�4���i��^_7��2,���<���:���R�+f��H���g#c�{����[pz�eHm�SJ��=���Ι���w�F& ��oz�!tp�8TOtK���\�۴� �6��iQ4ׅ���6σ�*VW.l��r_j��;�S�E�H̐* ��"�.��q{����-�Ypu�>�]X�(��K�'��,�?�4�츌�����Ax|S]�.����)�MDx7S!P�nKb�R� &N���lv�'����GI>X���ֵ/In��0}.S�
��{F����d��b�N���5�T�T�R�:�S�9_�DO7��Z:���l��+W2�_���A��!�ȿ0:㝮��F��7�{�̱���M�䛏�<��� ���,��뭜�kP�n���R�v[��<ӷ��]��%��񃈨�[Ӫ���]|���$�L��ǆ�[M�%3���S�4���~�����<�f'����/�ҋt��r^�A���̼��=Ev�6�,ݨc,
�}���F5�����nn��O!^�����P����+�	�C�;V{+��F��pNn���c�.���LSt�JV��b�N��
ӏ�F=_s6	>��8����X2�Z7%+
�d�h���DϮ6uc��+���O8K_���.��l}E;��N�F��!y�m1�GV$�3"VV:�z�|`~�oWS�Kbሚr�X_�V0��b2�_;�\Z|��������5妿N�hn�	�")7�p5Ɍ�D��c��[^y�Q	�!mP�N�$��]5L�:T�>.Gp�#�0&r!L�0�{��RN
�T�����Y̕�hX��u~�QP@P6Գ?	0ST(�{����tY.��A�H)hV2E�Ftԙ ��m߯��&�,$�$�9��юmJ�q{X�����V���Q�1��]@����p1V�̙:M�d���L�6~����L*_��-��������~�������j�^?��9 ���"�����Uڵ����m��	PfO9!���.�WM�+rc�/���Dd�����ĳ�$��!��=?��JƄ��t������������r�a���]����Dh�25��>��E�w�������nXfV�]�%��;ƥp���|fĿ��c���:Z~C���X�g�e\(�Z͏r�����#L������,sG�`��hj�j�X�sy������12�F$�1��'p~�o�a�>���|�����V!{��3脥�4�R 2�U�JHoy�!d�[~ߪI�h�@�BF�������ѐ��ʳ���p�`I�x1!	�GPGb|Cr�TN�#����.-2�a��}#��Z(j
5�8"{�d���W�Y3us���@̎���P֬�̀Pi���xkd�sn��lPCCfÔ�Jjq�T��,�򄄶�]A �9I�U�]�����tÖ����</�T/�|��?�Z�DS��E��1�m_ͥVNA�;P���7�f��(]n���B��9Ý�?3;�F+\�z��\}�1�-��Y���p�����K�v�WY�T��2����W���������}�7B�P�(�lo���>+� :VsF���1<�2����4����A��~z�y�s�`�֒�4�C��r�g߷C2���q
����)bp�����UQ���Z� ~��~�1yl��ب?�K�=�1v-��u6v�^w�����%�N��
ls�jd�Ԃ�(�� ��� ԏ�T{��p�x��ze��-���ɞ�y�>.�V�����1���{#ڲ9@N0P���f��`f�����a����D�*B��Z�t��־����k����x�^TP9�R����������li.�� �!n�U��� �WI5&;�Jd9z1�
�>(xq�4R���r,V>2TuCt��+g
GzCtK�����P�Ɗ(^�*��V�i6
y�&H��2�������`V���	I�/a�	�MB <�7��3�3`�IJ�e����+��
��LLZ�^?�Y�
j�xE(�?~ ����n�,LoQ��O`��3�v{0v�Cz8�n<��K����h�`�	ldo~��!\=R���`^6�֋�1�@$(��r���B��� �atؿ�:�t����F)�8���r��Nn߀�x���ߨ�������D�n����߶r����E~����պ������(u�_` u"ؼ�������L!�e�SW4�8{�;�v�E&�B3�KL[�ޓ�������� �+��[C#Ѷ�`��n|2.z�y�/_������=����N�_�� �As�,��=�u��iM��k$f�.�s,���&3M�ˏ�6^�6񜮿��&v�������g��T'�CR��Bj��ج��k��Ͼ{��ʅ�r�حV`��fb���˥��_V�d]>��|��M���yJgPې6$N�tD�D�w�N+�l�|	՝)\m,$��*C�DBM|����w��.S�$�Ŀm`�c�8�;�:d�r�؉��e����h���p�l��A?��Xg�]L⑞��'�&�͉Yk��u���)b��R���\���O8*+_czN�8��@w��
9�es/a;pns��Ռr�8��HTH�S�'��U$�Ҁ|1}����1b��M�J\�5��ڊީ�	 4��'���3e\RZ�>K����Lٝ`��9���H_k��`^ߴ� �������?{����5T�x�֞7�	a4�%��ĴJ`F�:��5Y������{���*����o�_������ucI�a �z�5�C6�@����k��ǟ!�_�&����30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�&ڜ4�z^�27лXo��R�|n�?S4��{2�в��3�i��R����@��r����>x�<%Vֱ)#�׳��'Z[�Ϲ,@"����4����Z��mg�U�f��Go�����X"�q���D4�y���O|�:�G��oT.�t�U���8 N+[II��
U�v|#r!��HQ�I1���7 �dI -/�,.y��1#r�.$�����S�����ڮ 0����o}�#��o��O\u�s�4p����O�>Ԣp0ut�U`��D�i!C����k�z��( ����x��R�׈ӞX����jI�����q#;r���Y�t�����ه)�9IhnB�v��r/�#�6�ˉ�7vCl�Uɽ>^M����5���Ve�)[�����R��O�>Zp�#�؆P�(o�\����9T�͋�k��Gt�_ÜH�e���ʽ_�	��k�ڪG�;3x��4a6��y]��
�5�l[�s@�5��R	3�	_�8�u�D���PsxN4:�@���e�O��jn�1+m��;�{B���b�d��e(އm��Dch~9Ԛd����I[����K�zV�v��8K��S)9�ӰV9���x����D�|����mG��-��'�e0�Nx�R�dǺ�+?����b����a�*�w��N��J3H�`�p%eWI�PjJIH��j�� �;|�@�ɬ��zu����&��!���:$�ٙ^��F��bs�u�V�:��G��TF��\O`���L� |OgY7̟賴mr\�J�}4�gO�u�T��١0��� x)B\R�iA�\������
{t�ΰy����=jL)�(n!����o�zp9���������X������`<��4t���S#�J��/��U|� m͏�J�_�'\Ə5�喢M�9h;�j�ΤK��F�uuR�4���$Ώ� g��qq�8��jd�{�|Q�C�,����xU��0���(	$x
HQϑ���R���'�i#�V��5�Q������БN�#w�c��\⬕bk�q�l���TmE0��O�S6xO��!��k]u��~��'f]|��EpV�[A!x��t���	
�i.Hp�6tO��WFE��<
���,_p��a�9�҆�7d��F<����g,��0M}lW@sp$G8wq�g$��,'����I,�5���R��=�G�[r��
��=�A���>� N˹9�JYE�ӽ��ZKۆ�-pk�Dn�K���$����@���Y�~��X\^�%CPF�-���!��h�t���r�"�d$�::��d�� ��r<���L~yn_��c#X=�:r_˟��/L�(��ƔT�^��s8�dr�MD��Z�eT�a���"	#�FN�9t�&�J����!�Of�ZaIݦx�x3�6[�u�7;g<1'w�q��Ӳop i�D��KHҟ�p�;��>���'�L���VP�UHt�<m ���i�'9p����[�D����ڳD��<�M2�EIp�\t��p+�瑴���S���#-��.��bv�ß�A��Հ�fɗfF�s���۹����0�jm��?V������~�˹ʛ��a��%[�w2�V���;3f1h�R$�)�$��q�Q.��m(I��Ɍ�n�~}�n4�r�ʰ�I�\�qBSlw�!��
�U
�d]}Kn5B���O�RN��W{����
���o�?(�]���7dcs��<�WJ�\�ꖩQf:���1��s�M>�d%�	�������v��E}T.1L$v�)���1����
Ϟ.��*Σ#ȋ������%��Z�5��N5��{�]5�Gڦ�eIX&�iê�=)`����/	�Ֆr�GSU*F��6�8���yl�F�q�Xx@S��r�{�eS��|�#s�P��7�N>@�Es� ��u�P}��b��Z��2̼׳qY,'^���=�n�&�k�;��"޿�-k��j��s�ttTW&����58a'W�l~��0"!g�psd���������5OM��"��څ�ey9v�.q�/~ڧI���kMV�#�c��k�s'
���18���?~�8ڋE!�42pQU[Ӈ'ߵ�,��\yμ�}c�p�.�R�4ą�M�[�d+��cl����g^ �WFbOD�b�RGw��l�;�갴�_EvsTN7�>?�x�D�ː��+۵c�`t7-\L��G�r��[��y(r�Ѯ��0z���yBۿH#&i���z}q���Ƕ����+S��@B�<n�-.T7���On��f�כ�荂������' �c�i�Z*}b��;);A���.V�t��{����W�\�i�kƮtE�;fۺ�;�CF�D�T�2o۔���+z'sq5Pƹ�_��Cw��btܕ'1Tp����^\��P�u.F��X2=A�QY�~�Y�6��!���GL�.��������x>�F�&�P�2_�<�[:�����%�7��a�����I+"��o��ڏa��#bD��ɖ���u�^Z����ѹ��Rh�5�8"P�ɫ�C֬g�^vִCEHpIq��nR��pvY�L��>0�p��B�)�lՅ[YƮۃ���*ݺ9|Jr�ɩ!Zr�ē�����J�4�W'��Vx$C_��}�lnA"��wgt�$�'��\�l0d� G�_K�6d�H�b�2�'�981��!��lz��<����D�bZ�%�|'�k9�Z~��u;$�|~!It'NZ�)�eݰ�v�����^ �0���J�֘�̣eބ�$���p��.qȾ �M�E�`%�����1z��[�R���,Q�����\��/��H*�z����?�G����+�q��|��iǤ��@P��~�X�)���b�i��Ay�mf�O�E}�.a��i�����V�K4's$���=�{rd|�1�.Mݾ��@��_�܈��B)�ԟ{[�� �'z��G����U�p���쳈/�\�#[���Ey�xx��]��U	G$'��l&�I/�>���h߿G�)������re<_��])@1/n��47��y�o��	C@5ʆ��<y����w�{49�[�Ֆ�^��h@	��xNH��Cr>Z%������j8���{���!��Ǽ��q��� ��܉�h|"�5e���qy�����E�E�h. ��^3��
Jl�:+�R���$ւ� ��]a��uaߗb�����J�I(�@�)\��+�c������iQ���������i(��q�� 2�'� �3I8}�6�JU�rt�'��_
�qo��`�CӅ¡�K��L���Y��f����Q/�.�X2����bK�E�К\�P�\ʴ�%Qt fX[X~=.}LJ��7�}I�ժ�?�ۓ�Y%D����:���B����#�Ā�d�o�iLc����cF�hN Y-��P�atÕQPX��6�5���3�8 3�<���.2F}hL�f����S��t*`�]�Ҿ�*�m,��E��GT�fWT�KG<�x��痁1[�a�␳/��8)v��a�Ēk��&B����M�nR���+��F�Ȁ%�R6�_\{S^N�8gUK&�����%�,�˘��t�<��~7�gj��l���c��@��A��W��Vt��Z���0���őή��/kѼA�u��5��B����9ox�,^���:L	��0+��iW��{�(G����rq�'�mw`,�=��k�6�'�(��SM5��:f�o��6�Bc阝�.-|�0�ǃX�b=G��P�k��6Y��	�˔��3[8����z����p�!�qU`1�y���j�_�ܶ���<3n��`M5~�6k{�C+��
B���{{!!���t��v̈́䭄6��EXp�H��g�X�tD1�RۃB"q�Ǎղ��s�]!`Ξ/���<^&�т�"d�ND��Y�U�y�]���"[�X/�1.�"�7�_���\�A� O�>0�'5����:D|�fe��C7��<����:�ȑjV��Ҫ�>D->��-�ւH�C������ �%�-V�
��p�~b���qQ����Q�����"��2<��e8�EJ�����cVpt?=^TI�����Fl�R��[	�ޑ������H�R�p�3z���Ѧ�jy�"�l��}���� ���R���j��do�0'�k3����1�V-��-5;�=h0b��y��s:5)�����Q��>�~~�-�A gD�)yꐓ�<�K0��ʟ��S�-WTAEE�d�(R>���7KF`�5{|P�S�_��S�y|d�t-���nDz�`�9�ZԼ��QKD�𪝛�e[-W���?B_����?�9{�B��򣺨�M�S�̂�kB��%5<�05�48{Ye����*�0v\�/��=6���ZѦ���d�n� ��l���&cӳ_�2�m9�}K=��n(��S94����t����:i�����@��������`����G��n�F�8Z�Y��]"dB��돕DܸZ���g�#+fhoܐ��L	�"�/��G4X_����|�(��-4oy^�t����T� S�I�u�
��9|��!��r�͓�[��'��7�iIżɎq���&��H�0#�j"$^x�;ݦ���z�L?�P��0������#�љ��c�u  4u�t�V��>�0Z��U�s:�iO!���G�Rk���7���D��˛�X�׭��XK�b������V��U+;���ٺ]�r�2I�ܐ��)��hs�>�o�rt������vh�/Uݰ�>������� ��3�Ӄ�E|� +��>��#���PJvvo������9�Fs��N��ki�Mke<�⦫�J�9,νo�*�Dԉ����	��ۙ�eoL'*_7	7�I�6R5?﹵��Tu�
cKWl!�Suz��>L���m��o?\��D睛�+���{��Aھ�iL�������y╽Ȧ���F�`�Y^f�����j��O�-$�:-���K#�
���&���I �:Z�-����x\��EG�*�}�͑VZ��� ���%�`������TZ^y�;ͬ�m�Im��<��1�.��X�(��-Z�s��GYlx^H�ʴ�e�աw����Ϭ������8�g���6By����`Y^rF�F�%���Jz�on ЁU�����S}tHҍ��[�>\�}�C��� ��?���h���	�a[Lܽ���q��DplN��5W;�v �hH�U�X
�ŵY�B������5Z"g���CE���a�(q�杞��ѝ'iP��#s.�8��=w9�ѓ�na�q��t~^�Cs��8�2�-�x�ޮ�y��.'v52����Q��.��܃�:��`�\uQ��}�v��[
2��s9�����	~lq&����H��.N���v�ȝ�I�����wOi�t��bo0����*5����w#�bn��o��n�JywS�x��q�*]�&�<[���2�7&Y�
J�wx{|����5�UAzQ1��>5��TE)M4�N��vB�ސ��?�EQ�O���3#��m����+��<,N���,�����P�9(8���Խ+?声'�}yU�<��2!nFU�:8��]�ʈ��)�Hy*s=��^�ʨ{����>���Tݯ`�䳒X�[�mӤ��C8�^�g���a���^1�p����ʡzHy��p~���9~]4]u�5F\�Ƨ�R���"Z��ږ��R8
Ä��_C��4�F�	�+�VX�&�w�ԋ���A��w��c��<B�P��mGb_�T�&� ��#	2�������-U�mr2S�? �>#��G���q�=���_F�naث�cZT��|u3�$G���L'���l���eiK!\���¤nT8�n�E�=�`Ƕ������pZ*!��f�m��R1r_z�������ڼ����|`��j���(8��cȩc0��񳮀4�}M �����̬�J�Q���-jUښ)����b�!`C��l�o�.�mJ�|���wb���f0�)Jb�кǎAtÙ{��d�՟��o�˯�\v�J:0�I@�����J�WW�o�maj�Nú-���CX~w��Q������I[�7O�k�c"�dQ�]�YD�|��(x?�G�ip��_X�Xcsu���]����tx�= �~�p�J�F��uia{l��""��^��=M����/T��<�W��#��:���_/G�9܈[5{
�V$�� EX&�����ic�f�6?��FL��2`$����Ƕ3�~���~^S�U�E$6��I�HB���+� ̇�%~��c�ݷ���y��'����y���dH�P�4�����)�'�?���C��v�����jN+sɁiN2����2���j�6�w�;�vp�$�� �k�2�`�o��D�F�����vG�8�>g�?�ZT-��G��Yd*>���.ű1�����Λ���;?G	/YKN=��t�+I2���O�3�pp4.�������Z��|�N�@�I����3�̣�����:�D�k���N�>@Ĩ)eOWҗ1����9��{O_AX���\(��RZ��y����hK\{��\�TV�c��K?<<�c�œ�瀃��P�9�6x��}��A�ݜ���c�w	ۆ�^e��N��qK���0ܥ퓸�h1S߯�D.�N�me3�`@�B��=,KI����� �R�������uB�'�s�&��)�{�Q:Q�S���?�S�o.�u�s�:7A�Gz�mF)2�O����Mm�.g��y<�5\s�}���O
�4TW͡��6�U�)�2'��\��\���7��͛�P�PU>J\)�\hnnNl��B�z�i�����)��D�Л����:�,��q�����i��� U�g�z9	��������%5�Ѣz��5�vj�$K )��"����!�x)��Nη�Jn8X�?jx�jψ�|�@b45 ����-������}W	�meH�\�}Rѥ9�יi��V65�Jn,���Α�q��p�c�F�94|k���l�t���b�0KʒO�ax<u��k��=��p��|��NE2 ���xҞ�$֠
��i��/ң��� �E0F�
<i+�^�n� i�����7q=Z��h��$�,��M
�mWK$��q�
I��=��9!��[��,��
�t"\�j���(Y�w���J�����>�˦h|J�Q��?�'�>�;@k��9���9�q?���Sk�B-�ӫL�X)?�%�J��u���>���q�a&��OJrjZ�1�:��q *����rf����c~2W��%�:ߓ���lHLY,���A/ߵVt͇Fv������E()Ӧa�^W"V�K�3��9���&,�f�2�Os��a����T%3���c�;��p<�x����ӿh� ��<^)H�K+�F(�;=�m���;�BL��T>V�HHa�em��ږT�9ػ��]��Q]��~�� ��w�O��8��rzp�%Q�:S��Ĵ.0Sk
)�~ �8w���fA�	��S��D�w���~��ɉ�Md��]�mut&V^)˷�8ɛjz��u���4����Dr�V�1;@�/h���v�X���KQ�&ǣ>u�(z��6�S�{F}-྿���Eu��\B� ���"
��8�EZ}�p�B�Oϴ�N#�WD��ر��
��o���t���]@7dPr��?�WI�Z\w������_�1r���d	bڠ��L��C�A��PlZ1�e�v�x8�����:7�l�:�uǣ0��Рi�� r~z�"��Ȇ�S���&�]�#yTl�W&RC��=�0��m�	u�]rQ��Sbyv��q��������Ӑ��ф@ _'rA�>�r_�)t�#��$�����ۈ2�r������P������Z��̩!1q�M^W�=��&���'�6jK��k�����-s0�t!s_&iNy�x�8��W;�\���!���s����²��}1��5�Mh2�TY|���2���ܧqkE����#M"�p���Ӝ�!�'7�'��� ��e?�<�N���R�4��U苖'��,���yu�=���n�"4�}��ڐ,Ƒ҄�0����E
�tR[,�F�z���aRԩۙ
�ܷ��̈�sa�w��>��#v����v1��ċ`A��-ɬZ�T&�-����M��}���z�o��|�BH=l#3C��� �zʓ��u3��v!�Xn&M��B׺�T�ݖ��n蜮o̽d�b���ʥ��x�j �1i�N(*�~:�(ϵA?h.�_0O$��k��W;oi����^�;S]_� ��Cs��D����`�ۡ�Q9,R'��P �����1C����/�@��5$T}� c0^���P�E�u�`�⅞NA�C����v�C[θ��/�H�.$��&�xa����d�����S[��C�9�%Q�����F�p�I���ۂ�ч�d��{����u�.�^�0q�����f�DZ��"�G"�����#e�4�^�u|CR�p��;�*s%����Y�2���c0�����k�������܈�����G��J�1e��9���~�úZ�[��J�2�W�3V�_�P��9�e��Jwt8�$_meé�l�|�HCh�������4���6r�E�p��$��7e>�u�tZYJt}��8R �5�2�	4�k=\�F���]��3́�[��W�X7��%~a��eI� AL�����/��/זrk�7�?%�:u����k��rt2�^��~�gA�_�D3��:����W�NL�
���3����W#��˹�(��ٕ&%��?aժ"db�&�97C�&zА%� � _O��aD� ��X+3��\���e;��<���̡�M�� d�J��Hɿ���
;�Gx���y�	{rL��7�V���H/5�m8)��a9�rX���<���邑�=��E��h�>����p�
���8 xL�|��Sy�K�޻�����ݟx����A�2�gb�ɒ�H���k�����	���k�m��uV,���n\��&3śC�1[ߣ�䠤R��V���;�7Vh�W㇄*İP�QI(����($Z�"c�	7=}{>���j
��;��w�B��
����
����/�}F	B��O��NN���W��]ؿ�
Ԛ�oXR���ڻk�dD���$�W�5B\�E���p臂�1�����d��	��L8��Q����<�1�G�v�4Sh��G��P	�C�C�棾���G�.̴Hx$�-޻�c��׾]p�_���`�=&`�~�a=D�'�3	��r��S�S��I ���!�d!�a���tm@.l$ri�� 肄w�#α���j�i����,u��!��=P�c�]��Z��2�wu�qt��^^��=�v�&�nQ�������N�k�7���s~��t/
�&7��8\�-WIV����!���s�>z��w��K�τ*v8M�a�b�р�<�����oqy8���m�� ��MQ��~���ߕ���'������ں�{?���"ҋ�J�4���Uv�l'Z%0,�--yC���/k�­�`4e��hr�����>vs�Nd��K�z"�F������~Rb9���k��e厚��s�h�9�C�ӥ*膆U�F��0�`O�-�����nc�{q������/�-~�z*j]�߃�B&g#�ET��tz�q�C�Æ���9[˛B֭@���NT2����z�|�ܽ�	��c�Q����FJ� �g(i�~*ظ���J&A��.��]��9��W[��i߭���ƞ;!�=��lC���D�p.�m(�/� �8�'�uP����z�C���=ր�R�aT#���^�]HP��uI`i�ӏ[A�^C��[���/9���!��Z|���&�7��x��adR�M��7'G[��|[�%�'H�ܚx�~S�I��Ԉi����ȼ�r@^��Q��ނ�2٤u�ӵ^�wF�#�Ѵ"R�>����"kyN�
��B�u^��ZC�]�pD@z�88���Y�W�#v0��0�}���2��V���	�s�[�����J���hͮ��Q嶅��J�8�W�zeV���_9D��G(�]��w�$�W�÷!l�~��;��_�Wd��f����.�93,��|sl5v ������qV�`��'\�]9� E~D��0lۊ�ƾĿm).�d1� ���qA��D6 ����3�z�<�j2Be�N$�=��k�.̣� k�E�~M�v��B�zP��[B��EԲ�WU��nƾw
Ǫ$H��z���گ���Ѯ+J������^�������XXz�� I�b������y���fE�EX/z.�@���f��Hh榻is�Vg�3�{��|�.�5��CR@�`_]2�D�)���{�7� ����$�?�$�U�ݖ�ɗ�ꀼ�>�Dp��yًq�C-yâ2�U����'A��&�ԏ/��`��{�XG#����4�L��<��]D��/��~4V��8���#	>�U��<4��:9���&�6�s�GY��߲	�9:Ny�y��&zZ@�4�i��E�{�W&{���������K�U��7�W��hW��5�=��ƨ�歗��Ǖ��2z븂�t��o�J���+s
����,+�����nƗ�fjs��J�߯���\�!~��+���ɓ��a�"�xX���Y(Kq�.�2<ii���IS`�6�-��U�b��_�}qj�I��~tC�|�¼�K�`bL|϶�6��W;�]l/B�mXó ��KI"<�uȸ����\e�%L�f�<X9J2}g�s��Iv�)�z�=��-�%?[k�& ��_Ky�ċ��* �a��������7�c��	C-��˙�O0�Q�`Q�[F��82�����߱W�ў�:�}Cd�f�ǝͿ�o��nc|����*��#�	�q�"�f�r{K�!�x��������K&a����Q'8�	��-��!ha�5ɖ�g��#� R�o۱�C���}�c<C��?�R���_U0^ḭg���ָ�%��=�,�*����t����3�g�l�7_��P��8A�ziA*�tz���u'�U��q�����N/�5A���t�7����29n��u��2�8�����5�(��)�H|҆�Ym��O,f��fCN6((H),MP������ӊӂqc�ք�)K�k@��>tU�}�y�q�P�1ӂq�d礅���`�3�H1ܷ�0���I�nC��K�!"��`̖&����j����q�N���&n��M�g6U1�ީY��\��"S�{�ݎ��m��LNĄ�tV6ɃP�YYH��Jgai�ɻ�1ޑ{��Dq9:��G� �]Hi������0��y"�pu�)a�ꔬ���]Ǖx"���/�H�.87�^��̋/�||LOi��"�'���D7��e��7h�G<rT5�	��, �,S�	�D٠����_õ4��0�!�&f �QV%�}�+��b�^��ʮ�����#����K$�� Ԙ����nH]pO��=�C��&�y�A�];��_�=;�x#i��fR(kF3-��F͊p~n��r����(� {�`R�����*d�A�f�&^p������?��6�x�0��y�ڢ:����|Q�o�>O���Mh|'Hg�sUy�f/���K��nʺ�SO��T�����?$�^r7�4`�����S�}�؝����F�d��O-�M$n�e�`����uy�w_Q&<ĺ+�!��)g-R�w�Xj�T�{�Z�c���������^�u�}��k�X����5+@������YL�[�=uH�+C-����-ʹ�I��ׅ��Cn7~�����Zb&z���p+2�G��hμ��nc�KSԣÀ�D��p�<ȿ�i��ͻ!��@\e=@7�̧�,�܎��Q��ȥ(��a�}Z���̀N"���f1��?�fZ5�9g<G;f/oW�0�'�J"?3ч&��4S#��b�|Ȗ���o��up�295������=��w^��{P��ub����A���2���jFoՊ��{B��S�[�7�H�p�1xr�n���k3���[n�Su��%������ׁYI3�O��юܒK�d��.����kI�uDK^�{��x��m+RS�齃"�Oq�Cfq����^*v�Cy�
p��#�b�~�UY8w�\�10��d���Ƽ<������θT����J&���U��FL��1��b�VJ�,W�,tV��o_rX9��l֮0w��>$f��Ð��l��T�-_��d�����R��9�]��Ux�l.�=����<co�B���٭�'��Y9���~�u)�����&�N������r&��+��*�X��>� �B��L�U��?���6e�P�$E7��$F�.�g	 d�aE뜔��`�K0z��[ۈ�_��`�j�Җ���E���UH?7zA�S�s���KP\+#.\���� ���X�`�tQrj��XHM��p�b��b����y�Bf~nJE�.����΀�h����s�9|�LIy{&�x|��.�B*�@�U|_6�|�=p�)���{�� A͝�'���U��O��CN��5B�WO��`qy2J⼶R�;�U��{`l':��&�1/ŔðM�>�K;G������%�<�]]h/"�4k`s�-���C��	��aʺإ<-g��ש�/��E$�����2�	� NRo��ZYS3��s������?{*t(�������D�ʑŸ1�H�h��5Ԓ��+c��ƞ�y���]�4u�B���XaJ �b+�������$���ݎ��]��\�Jhm�tw�\f�)���Ф����	�e�[6Q��^p�`_B(�q�B^2�.���8IlO6Q����&����_>��q#Q���ҟC�K`�Ր�K�ѧL�g����"�ivS�	/�X�k��)@dK���Ω�
�\��%%�f�"AX2�}�����BI�����LRQ%����΁�XՁ��T2��S��N��#����ě��cz����-&�������Q�ߐ�|J��Ap��ր�)ǱpĤ��x}�i�fg���6�L�(�	��=����Z��Ia���W�Dk������0�p������j2��Vw�}�?�b��'�R�а�H�������rϝ�F��������]p��=+e���7�S�	��N���S�*Ê����A�9R��I3�2�����@}�o��Aџ�� � �R��{��?�d*a��Zz��ܛͰ���]E�Zw��
��0�~%y�~�:�#�Bm�Q�r�>a���Lt�g��^y��[����K}<ʌ��Sa�`TnA�R�7�-��7���`:�oi�rS�����ﭥF2d�q�-��n�!�`8��G�<Qx�G��&�W[%-d=���F|��J��,|�(Ј�ݺu��0f�̏R�k�x��A5������a�wY��2��=�[��W���̹�x^�"��ݱ�n�����w�,��&�~���~2�(Ȼ
d��DBn�LS��Ā�x��fc�Qe�iml{�3q@���Ұ��y�+��u֣�4�7��3߱Z쳹B�"1�e8�#�Q��Z���gΫ{f�foi`�yʰ"ѐ����4e-g�q��|�\�okbt�(��!js ��VI� �
G}�|A��!t��T��;�?���7r�1I�����L���5D#$�8$�r_�;y�&���YD~���0�I'���#5�`�ܘku�ڤ4���cKM>��0�$U�����!5�/�k�n���� ��%B��E[��:�Xx����U�0�����;d�O�&.�OG׿�\ܽ��)��fh����(h~r!�S�h�����v���U
Z�>���zPƱ�ֻ��/�[S�2�7�� �Ar>�1�#��PW��o�赘�#I9��u���`{|r�82���MeI+d�X�񘆓[�\a�*P�X�����gOY�H��e|9**�i7�h6�?�?|eR��q���%�W�=�`l���eL���m�6 ?�}2D�z�����p���h��k�cL #��g�*�H�ছ���0m�o^]^��%�j��j󦏗�gᑦ���w�"��;��� 8�"�W}�Sx�?�EW�Q͞�H[�o ��%�_��y��phZ+�L;y��͹l��)�$���HZ�-ry(��Z�$޿��l�v�������Վ����9���A���@8q�ρӢ�B&Z�OY4*F��6%���%^o�$+�b7�Ƶ�Sʽ0�zK�[�]\�_"�֙�G� �?5?LSh8�	ߖ�[��7��-�_�l��5dGJv͐�h�!9�E�U�R �Y߇�^�Y�Q�5g��P�J̅g��O�f�Ep'z�y�7|s��x��l=^�����a��t��|�P�ԪP�s��e+s�y���b�v�N�3�0��m.��)��:�����q���v���[�ٞ��0@�F#��V�qZ�Ú�H��F���【���vޯ�W�Āu�a�b�����u*�*��Z�bo�1�n�B�w���9**���rLu< �ۍ����Q0���Bw5�|�2	���!Q>C(�9�f|�):f-�S���� �]>?�f{Q���J΃#��â�Q�+3��,{������8�r�{���O8�ٷ@�+�Ύ�Ta}F�G<|s�?	�F�F8d�C]�δ��)5
%�w�s��3��U�j3-�+uI��@N` ��%q!���G��tC����wT�Y��ͯ�1��Jp����Dz�y��/e�~�~�::]�d�F)��4a�����<8��8fC
�&��]��axPF���+Y��Xڿw��Р5��A��Փm��#����p%��aImT�K��ˠs�Z��ڤ2�^��H��
ۚ�m�K2 ��?b*>K�GSӅȞ�H��e�_�tl{1��B5]T��u �"GH��LT�ؙ9�����!iI��o��T��P�2&`��+�E�dB��!�i:f����SErL�e�u���t�Ђ!��9J�w�W�� ��a��P�/�~yZ�a�M�����=��p����~0-W�8��+�sQb��UC���|���J�ɶn�dd��4�0�Z�bl' ��qt�בE�B�"�m�\�(��f�JX:��K@\2��TJZ�ܼ���aW�mN�|�-���Iw�'������q��['��X�:c��ld~�d'��p�(���G�dp�q�E	tc � �&.�h�t�P=��<~���p�3��3{ڢa��s���ǫ˄�=Z������x.)as����+�sʷV/��Uܕ�{���$��3E	��K����Ei0`Ĩ�:��S�c����$d�e��s��̕=��~+�7�}42�R;�6�$ÖjB�F0˸G̴� ~g�?cZ)������Kwy������P.��TQ��=P��4~\櫡��AN��s6j�	�ɮ�2�u��2��c�j�5�w��v]�xG3k ��2s�D��^�D�`��N#�Hc�%�������-�ӵ��D�Yqw�_�{�|1�_R�����_�h2Gv܇YX⮞f��+�������32Cw4[h��H��:����U��@3��}�$3S�渼ú��a�Dl{
�N.ѩ@ne<���$[m1%���?7{�|'e�B�	U�ߟ�����xK�hxO��}]�t��p�}K�ţ�����<P�J�����9�(Hx4�������Õ��y�dO��Sbxe*��N�� �޿B��2��鄓A�6f� �q�oN��3��`M�-_�U����I&�$ $ ����z�v�>��uO1�� �!�P3��h�:�m(��������Fu��Q:�G�>9F��O���F��:��g}�2�P����\���}��O�2?T���jY��$[!)��"�c�\�ųI�$��Q���^�^��~�)�̸n������z��{u~���	�`j�K����L�ن\R�ñv�<fU�)_�U�j�畞�yG��> >I5[i��Zb�,j�	�Km���/g��.��^̮��ķ+�18�pjEڝ��Q|�G���?����G��\g��KK	^�zH��M�i��R~���aoAi��gV��$5�9��2����P���c4�s�&s\k>��l�"���8|OP0Xe O��x����q�k����a�M|��wE*�J�U,�x.U�O�
�W#i( �pK^�m0E=[^
�"fC,��*�<Q�3/�����7ށ� �r��8E,/o�M���gZ$Ağq�r^�U���F�̺k,9N��ar���O�UXD���]��\*{��8R��[�~j���>SV[D�##ȥ���d�A^-���n%Ϙ`�*ޅ{��G��Q��+�q4����-��� ������`:�����?�)<_d?�C�k#���x51o�q����Y��H�C�����Ţ�>z��V��%���Zn}}�����B�& ��`��2��L��D��x9,n���S�1����ߟ��G��i��@��ŋ@����_̭'���C0��A��&��galZ����R!"�qEl���Z�M�g�+of5p�o����"��I�,x{4��ӥ�:|��p��Ƌo�0t�+��p ���I���
{�a|��!� ^<��o��֨��7��.I�c9�R1^ ��i��#؉�$�!�ּ�b�ZE��$1�0����((#�X�<eu���4I���$>�1�0[��U�P�ª�v!iY��Ȭ_k��]�bq=������y)�y�����uX�:�Pƨ�d�^��;������5r��s,S���)�<�h�W��
"rU�k������v��WU>ͽ>D�M��`	���`��v��f�/�ap��u�/>@V#K�Pt�o��ᘄ+�9���Z�)��S����E�e�)���Ƶ�:���S�*�$��@8���|��e0�*@�y7��q6.&?0V�� ��bW����uL�b�m��?���DH�͑��MФ�z�Fڟ�'L��D�@��޺�8�|¦O>�'e	!�a^G��q�j�w�Z�y�� ��3����N��xJ���mY �R]�N�;.=x�R�E��7���R�I�r� �;�%�	���i���w+Zߚp;�S��m@B�*����6��R�ڧ��(��Z7��%��l9�͐{������BF�6:��t�?��8�:{����BZ�״���Y5�hF<'F%+��nso���I���yS~�{Ү�i[ġx\27���g�{�R V:i?�Yhï�	�[���;Mέ^l�Q�5�Wv�VhI]�y����YL�
��4�M��5����������i��ېG�]�R�B'�1��΍�s`9�9=?�z@'�ElXaC,�X%������~3F���iˮ-���I�Lv����g�$�{D�.�0��v�:�&�Ý,�8�vj;R[����㘧z,+�
�fqG�K�N �H*g��rr��6�M�����x$���b�Ii�"T*���^2�8�bbO��o�I�n�Pw������*�{���T�<����E�8�ץ+��w�}�|��ɶ�#��Q����߄|)n\������8��-?0W�QQ�˖~�:#�1T��;P+��-,�R�ޭG�lr#�`�W��8���++�s���@}�w�<�KT��F6C98!�]"�)���#)i9�Ɍ�sނn�Ujʉk��!�_;�ߕ�t`4������դI;RC�x짻���tߢ�1��`1��?pFU��O$pz)}�q�I��2~`�+]�oFݐۧh	V���B�p����n
䣶��Fa��w�Fa�+�j�X��w����F^A �/�!KWy���;���*mO_���Q�'���e{2S/�����L����>�mÏ24�?�A>D��G}��u(�D�b_��/�s�v�_T��&uTMG�n$L�����B��u!<i��T9(��f���?]�D{�7�w!L�[f�6��7[r��7����+ٮ� *��f�+x��	RC�����F�2������M�
~13�Ս�1+r�J�-����L���E�b@�+C/��0CP�NQ�}�7������0���b !*�/�ft�y����H�ݐ�6��I:�~�{���@7��Z�J��6�p�8a�	MNSa�-#`�ĊXw)@r�q��Υ��[��ڌ�cc�Rd��}��}�(9GG��p���yc�u^�C�%�؜t��=��9~�f}p��U�g�la�Eeʣ'��xq=��nFUp�]O�:a>�_��k�/�r��I�H{��$�7fE=�5���Gi����m��u$�R�J��t�o�q�~�+5߱��o6�I�J�EB	v�lX����~�Ec����ѯ��>y�{�˥nPb���>�q���<F��6�����%j���(32wkn@7D�[��jӾ�w���v��-��� N�P2'����DZ�����k �YA��	���>ч�����Y%����/+1$�ٍ�/ξ�j�nG�dNYqF���+J	q��3��4�����n=+��Y��@���+E3��хc��D:ܓ���Nb�@�a�ep�r���1Y[����{���v��=���S�>�5��,p�h���R�����?�$�K ���d�J掣���@��U9���xhf��Y���r������t�o�e^$�Nf�� o��yz���Rp_�Ϡ#���Nr��3�N�`MG����>UI�� ��D ���.�f�r˶u`f�T�:�߽͜r:��{�?}lnK��$uFO�:�G{^mFJ�O�qE�z�g�ɲ:&ҳ���\t$�}�hOK��T�I>����X_�)�p���0\��x}���x����Ŷ�S�v�)g��nO���eDz�F)��,�Y�ŕě�O��A�P�x鱪� g�]�?Uj�v�ݸ_������m595��'�.}j�'�K�v&��� �b[1��"�΄���D�8�=Nj�kA�)Hg|�s�Z����Nd��De���jk	�H�c�R����/�i�n�VZok5/O�63iz����Q;Lc�˙�ZIk��Bl"*������.0��O�e�x=K���kˀ��;���+|3|E�(����x�I��E�5
U0�i\4�$!����E�mX
�^���
&a���gw�tք7�jރ��!,�r*M+,��(�$u�qu0ɰ�e���ݺ<g�,��3ѕा���#`���:��v����>Ę�˧�?J���+�ԈJ ��5kP�Ϙ�׎�R����3��c���0FX��%1C`�}ޭs[���&�bwH��Or^�ђ�C:(ؑ:խn�rG����<~'4H�R�$�&�:`n�j�?L����⃔Bbֵw���m7�{{�H��kaH�"74�42�9�ս&m�>x7��L�O@�a��M��M�3�(m�#�;�Ba<_���_���`ƌ ׸���H����gnF;~�?�H_.��n�L�Dy��V~�XHbʠm�s����99����Ѓ���\���ᚴ�x���G��pW���e3�����SLG��WC4����Ӵ��GA�/�z���˓������n�,���m�
#VߋZ��d��\ql���v_�"�����PVs��;᐀hd�X�W鰃��Q��"���(w����'2���}�|a��w������
�hB�B�O�
���B+�}�
	B�"O��@N@��W�?����
���okԝ5��>cedQ��`x�W���\�� �?+��g[13���{wd�	����?A<դ=:�zX��c1r��v�=�����`qx�s\���
��ƅ�a���{�Z��ڸ���E�]#\��S�ӫ�&3�|�`8=��<�u�	���rҭ�Sœ��7�f�+��=k���H�Ɖ7@�1r������d�#���� ����M]���2�.x{c��P+;���qZ�G�̪�hq
x^Qq?=�o�&���-@���U��k���rXsq�<t���&�� 278�4�W���,E!&�s�_��#�������=ֲM)��5�d� �$����	�q�/ڕ��3JM��Q]��-���'xe��_qb�m�?,�V���sA4 �rU	��'M�,�U�y�:��+n��Y|�4��9��Li��Y��A����7��}F�(����R��Y���n��V�M�\s��������w��T|�#g2`��w-J�2�� ��e���t�0�*z`0�28�B�d�#�Zĵq,{z�هv3�v~��r#�"�B��	��=@T��CG�����SʏV;@�+@��� �BNi[��*����)�LA`3�.���Rv���Wn	�iR�E����;T�4�A�@C��(D�D� L�B-����'�O�Pj���C�_�Ȑ�/��T'$1�^���P�z�u�5���eA	�}�l���.��,�u�������*Q�xlӪ��0�@��3	[h}��P+%rÝ�Ϩ����Im@Y�|"��H���E��>��4]��%*�u>CE^H�ÿ6WF�'�<%�ˣ#�"�ږ��`H���\^d$C�P�p���!6��h�Y�����0�b�0�y���-��Ŵ���U���<�h��J��t�O�����d�]��<J���W��V&�=_,����#'7w-$ ��Ê�l��ΦR_���d�K*�P�9�̭�9��y�O��lh Syj������<�0�A'o��9mE�~P�cy�*z���l|���|� 	��(���J �|c��u���u���"e�@$����ë.��, ���Ee�X�i+>myz4}[U,��ٲZs�ݾ
{�ǝ9H9�az{����.��+.�� �������R�n'��;�X��L�s<�b�'#�/��y-�f8��E�B�.O�	��I�"���y@�sv���}{���|Ҥ�.;����e@�U�_0�G�wF)KrJ{�2� ��B��.f�7ޡUd˳�є5����ƀc�_y,�����uõ�4U���u*'t�1&_��/"�G"m�V�<G6���Z�ȓ�]<M��]�GK/ܹ�4eRρg���F�	�D�ʴ7><g�0�Q�=�鿹���g���/�/e5	H�NL(��1XAZ�2��y���ݖ��{��Ψ��d��r�~e��?r��J1wh��U5S�����Y|��sdS�j��Q��D8�²�JZ1c+��ѽda4��긏Kq��#o���y��J��ɯ��\ v~��ä�ŃEd�m��l�,�(^�mq^F�2oǤ��I�&�6*��?�a�_���q�nR����C��s�O�aK�<iL�)���������/1�X�y���K<A��ŭ�>�,\x!7%�v�f��(Xl�i}�]��C�IɌ$�-L���.%�~��������Wެ������]lPUV�U�ct�@<�.-�6	���[��Q>�n%�{᜚�mA&����瞜e�}��f�ƃǰ���d�A^���L*<�E��ӴuC<fE)�K���x��i����#�ax�Y���8W�]�D��@����Z��
�;�D�f�R�cH�?��q���v��o��Rd �_J3�^�p+göo��n��w��l,�����cyt�|�,�gؗ�l�ﲹQ���Q/A	����t���_���)��:�Μ��/J�AX��c��0�/��Y�沚�l��(uR�Ew��W����%�(5Pɼ�Xo��U 8meQ,yR�����6�D({��M��^��E�&��$�kc�{���e
�>vO�qd���dϵP�x�$��緍t�k�3��������(s��aO;Ԟ��!��`�g�dj�A�ܤ�E�Cb�n�NMcǞ6�M��w�=�k����{W��d'�?�ބE�6|^W�;H%sg4+K����1qf��TĬ�ՠk��!�n]�^�]���*���;"҈c�|wJ�G�o�'�i]:o�"���/	K*.���7v��E��/`O0�g��O&��fDj�e���7[HU<Ű�����?�ft���V�D���'2��@=�q3[��Ǘ�9!����V���^�b�ty�/~�mL�?��6���b�E��z�3⧙����a�hp��v=L3�9qŴ��0��I�f��4�k͙�BOIR�]I3(v}�G�W�CXF��ז�=>��� �gR��t�4d���^c�Y���q�(��"t�[���+
�0$�yQ̃:c����Q\��>B���/#�g��/yXX�j�SKw��M/�SB?To�s�#�����7yl&`�!�*�S�v��@�gHd�)�-J�nr��`�3؅��t�~Qy�ʺ������-����m���b��/����2���q�����kp'��;95�i�~�b�~Y���P����٢]�+Z����H��.��){nꋶ�f�፠�&MճM=2j�V���E+'n8S��1�-N1�C�����i.RO�e@�N��J�̺}�O[��$"H���w���kZ�ڰ�B"R�Yy���dlZX�go�f�A�oJ���zc"�L�9H�4�u���E|����z�4o���t��R�B�s t`I\E
���|�4!5L�5�n�<����7�A5I3���2�˚��#$q$���)���gL���f~˼0za,Ѣ��#
�ݘEu�ھ4#����>G-�0HM|UQS����!63�5��k�#�����H��{-��R��Xyp̊����q+=���;�6��x����נ:�ܾ��)���h!����g�r��I�	᫉I_ v�n�U�>�P��Y�H���a픃���󓆋�8/�B�>�#X9�P���o(��q�Y9�,���4�|"f�Y���wye��~�ٯZ�'"ܽ�X*1n7����F�Ӊt#e�|�*�ue7�M�6�ә?]q���� ���KWʹ�3��G�ULw��mC�Y?���D�X��0б��'N���o�L�������絷�IG$��V�4���h�^��X�{�:j_����h�������1��%�;�BH# �vb�ۮ��hx��sE5#�D^���L�I� w�M%Z�����-"ZL
>;���?)�wI�Ŕ?����d~(�BSZ��2��l�p�bD��˦�O���c|Ǭ�e���Gb8�!�4nB��O��=mY�OFin}%��85�o9ȁ����6�MSk���;�][���\���x���� �w?�!�h��	��[���t@��l�_.5Ņ�vN��h6|H�`P�3�"YB����Zx�5����Ѱ�m�st�g0�<���¿ľ'����{Ms\�e&m�=�n�m��
�a�r>�"���g��ѺA ���&m.�Z8v#A8�t�H�(��.I���Y�:�g:��~]��v���[���P����n��a!q��U�{/AH�{_<!�$/�����0D�eA�"�Bb�Ub���"*#�Ukk��O0b��2o�NnxH�w�}��Ғ[*Kd���J<�ǭ��܄%4D���w�Ca|���#��4�Q��}l�A�p�)��d��������~�?=ǲQ�%7��B#��b�D�0+Y$,|ط�_��y�����2+�8����x
d+���UC#}g�Q<�5�F��	8�q]�ɧ��%g)6���6�s�)�s����	��kd��g���1`�v�F�}�(�� �C1����0D�ϩ���@�1��pSvw��f<zv���^�1�?[~���]�fiFJal�u� �CMI��Rk��Л
q�����ٔb� F��i+��X;��w����"A���N�q$j���1��I�m���E?�Nū�	2����[x���Y��S�mpF2�q?�>ќ<G4]�ȟ`z����_��'����Tt�lu�]G)��LU�Z�U��!ʬV��4T&x����{��>���ڮ����!���f ���${r�U���������� �*�0�آ	�VҳnC���_Gb�b��M��>���:G�x���q-��yJ��n�b�V�C<�p��'����J�j�`�%���0��xb���<�Wt1P�*ڼé��?���F�K5@D}u�L�J�)m�]�=a��N���-�2x1�T*�şg<!��g@U8��2�G�c0 F�b?��.�tc�8 �u�����$´���"@6s؉9 �JMde�e=a
d�N��-bV�Hmw(��P~"�d�j[Zx��X�c��d��C7����(x�G�O<p'f���1c���F�;��tPD=by�~�<p5������a�y�����+=���YH�������X��zʊ��/�0��(t�{��$5�E�,O^;`$`i�&��cr������=$�J)ɞ�J���p���~��߰����m)6��O��B��P�ˋA�'b{~:c�Bo������J؞=}y\N-��P�M'	��p̥�v"枬yؔ���2*j�1�!f�2�P�?�^�:?bj���w;�vxRZ�w �t2F� �+D^T��M�d�߭�@������MѦ����Y��r`9���1���e�+�nx扬�G���Y�fZ�Y��+��Y�t$3E٨4�^�歯��m���v�H}@����0X�3fՊ�/�݅��_D90��]N!n@d��e�2*�7�61�r�����{��������4�����޴-�
?h�(�qMk��Xͬ�>K���+:e�� l��@M�9�Fxgg��zB��)��U�
��]�f��e���N�⁯���`	�|�=�X����.`��jiN�>�3�m`�KR�U��L�IuEћ7k% ./��M;��qyTu�͹�����@���$:���~n�d>�Su%,�:��G�nFɦ�O-��йȪW/g��r+���\��}aûO��_T��L�=��W��)�+��V�b\M�������(�;���E��`])F�4n���7�z������k&E��j�~$�ȭ������ͱ)��y򐈜��U��a~
ݗg0v�ES(5�$$��n���j�Z�K����8��!�֯��r�M�;�>�8���jN��(n�|�Yi�a
Ē�,��qͷ�"��ԃ	1~�H�ʑ�U�RqrVĴ7PiP�OV�5Jg`�vC2�����;�{�c�#��H�kQ��la1�ԃ���0�O���xܱNJ7k*L�z�Ž4�E|2�oE��A�H�xr���*�
��i��i�Cnv���LE�~

ܵR��oBc��񺠦�!ғ�}7�0���vZ,�frM�����$�ލq����"��ٙ{��1�,���W�
`���5�����`)'>���F)aJ�&�ӊW��+C���kO�O�������ց⡵�KU�X�[8%P�	�9��R�|���'?Adr�o��>�:G?��5�M�r�=0��~��Ç���t�:���iq>L����8���o����t��^9���]�g���w'a'��"�؇��n�9I�t&̕��#8���O8sa���eA�3v�����;4 <��
�~���_M! ���H�l���\�;�pk���э�@�L�0�Xm/V=u%H��m-q��6��9x8L��m����;7�ڠ{Z�p�z�����pSBm��A2�Y�Έ[SwB��~g��_�/_��0��A� �y�����d�`��j���}��\�m�'V������;���^���/\0�M��n[V���;�q�hC���1��"z�Q[�����(�%����c�}��h�_㎰pƖՉ�gB I,��A+
��i�A*�}��uB�y+Oo�`N�W�W�u��Q�I
��ojb}���l`d�2D����W� \\�ة^$�虄l1>��:]Cd�{�	O"��U2�����$�0�1Q��vz�f%�	�+��ןk���b��W�@b���~}�?}�P�x�T��]B��p�岵�&���P^�=V�_�yV	�Vr�bS��eU�%_�6j%�s�H�%Z/@��"r����c��L�#`��̟,k�{ٿD(�m#)��P*| ��'�Z�z��IBNq��^��="�k&�T��,F��ւ&ެ:�k����_�s�x�t��"&	_�1�08�i
W�s̀�R!�"�s1�l�b���"�<��Mhj��ſ���㥒�[C��q�ڴi��2��M��̴nt��'��	��'Lڌ��?+A���5�2�\4��U��<'�h,4ۉyh��*?n�J�?��4Q^��z���1[$�Е%� v������cFOg�ӓw�Rt>�930�W�>�lYIs�l���Ͽe�6�X��X�Gۂ�h`�r-i������ͣ�fz�^>�?g�z|uZ�q�B�M�#�gf�P�^zj`2��D�,�L��v���B������"T�6D�t�@�Np2�׈��.ϔjb��� �m�i:Gt*j���o�A��(.#��r�ŘWmùi1��a�;���0�CoD^�.�?�/�Av&�d�'`ԝP��.�CD *�υf�$f�T�	�^I��P���u[�L�%ǱAH�`���F���$n1��4���,i��0c����Qx�=��3j��1���['�N��%��.6'�YI����{��'�����p��Ik����u}Ke^g��5k��I���#���b"}�1�\�B�Դ�^��fC��7p������W��Y1��uD00.01�O\���>��7�ƛ�{�-4��J?���69�.6�c_��»Jo,W���V��J_��|��g /�Xw}l$�E��Iڀl�Ir�M��_kd'_Ǳojy�ˌ9�L��:l����U���{���2k�'n.�9Ls ~�9����Ͻ�M���6y���;��Ł��R0 ��E�2����9�e�R$�q�π.^$� ='3E�k���dE�[z"k�[T,���-�J�}������ԿHx��z�wH���O���+�<bԜ��/��q��̭���X����R�Ib����ΤCy���f�7�E��F.n�����ǆ�8Xs���E�j{?k�|0�.Z���1�@a��_�절��)�03{(�� ;CU���Ì6ĳUCq���X��?��P��D<yk�:�gôPUf|4��'i�&�_�/ށY����u� G5��9{��޶�<��]V3�/;�4���tU���y	�7��s��<�v�ЩH�H
$��'�GV�.�'	'�CNƸ�Э�ZR<���@���f���n{�1F�n��ǩ��ꭑ��s�Yh��5r�W�R��8��2���-0{�+\���Jy��+����C��uȏ�S������/�H�`J�����o�\����P蔤����tb��
���(]�1q=�72Η:���Ie{�6j��_�4�+_�\�q�jƶM�C`/����K�&Li���)��A�e;/��X���"�K���s�]{�\w��%�P�fE��Xa}y�����Ij��Lћ��W%�����1/��n���oK�����|�&��4�c3q�۽/-�/�V�Q]��mT}�Z���p����i������}�7�f�X�ǯ�7���\ ���_�P*�v�[t洴\�fdj�K�xٸ"�n���|ܺa����^#8����4A�?�ݍs�g���i�ک��5BbRN�p�~m��C`�uq�NؾR#?�_�I�^{[g"���Qr�3!�@,��˅�XtzHM����g7� l'E�p ���wA�vLӰ�tLB���%�*��_Dλe�/z{A74�"��B>�q|E���_ �G�7�D6*�6%7�x��(�՛�;��(���!m�[$,x�%��կ6��(�;Mb���+Le`G�C�	c�XD�{�����O��Əp�ãGP yD�C���ٔ�V�3H	@܉X���
������i!��h`�����Qj}���C���Ąnn��M���6'�ؗ��������{����~����3�Q�6��Y��HK�g�F����1𔉃��I�տ�D� \L]n��1w��ˈ����"1������f`�&��]�w"H�`/��;.$7�'~�^K�N��O/���t��zX�D	�e��7���<���� ��>�S��җ�D�Q]����O�µ������8�r#�V��G���b @��gj��Gs�^�5��A�a�������`�����p�n�=kqH�8s�œ 1�oY��������達|R�J�3'��&c��%���Һ�d�z�f����~�(��+��Uq��}Ō$�W���hD�Ձ.�B%'����
�S��9#�}��B���Og�>N��W��%�Ib�
�"�ob��f���d�ԅ�qW��\浩V�8�m�1
F��2d=d�a	�������۠������1I>vrd��#@�[�2,��ݣ�ڕ�8Z�uxS]�7H�=�L6�]:&�����%�&�7sH�=N���q�	%�r���S���]=+�F��.0��k
v�~@���r���
�:���]#X�̗j��sؿ
��e>�z1	P"5����!Z}Qj�A��q~]�^�3�=}%&�F��$w����ޤ��k���L3s�st���&Ɇ)FX8�1'W�:��y��!���s)��ZR����4�M ���i������P;,q�!ڬ�7�*�8M��v�If
@�+�'��r����ڄdr?#R���g�*.�4�QU��|'��=,,��y�ϸ"�;���7��4I�Q�rʆ�)?&���c�8�����'FG�Ӌu�Rl�|�1���O�L�d�s�\]��"Ͽ]G)�PY(�P�;�za�`��G-a�����ųC�^���V,?7zt���iĳB�w#��Y�Ha�zb磇��$<��:���#B�)Χ���T|6��l�e�FN���s鏭jC�b��� ��fi2�*b֜���A���.\��W�We��i)�ӮY�>;�k亸��C��DVYq�7���9����}'X;�P��*񄼌C<�O�Ǩ@��T���^AebP���uSr#��WA@ʪ����6af���,�$���(X����px�P��+���������[�]F��%�i�&B���vI���s��������<F��.�|*�uuNM^_CͿ-~��k܅ģ�g"u3��TȚ��/�^{��C�Zp��a�¶�O�Y)���m��0&#��G����K����%Ɠ8�%�}��c.J7����W��!�[hi����Jg��W���V��{_�=���J�'�w��$���Ay�l��d�E_��d���g$��Å�9}d�Q�l���ek�MJ��sh��*�`'f�|9D<~�ȴ����
�@��_�.#��
��ػ�i��Y w��=y�Ԙ��he��N$�Ҝ�O.V�� 5��E܈Ȳ�ʟ=�z�[LM��%�A6���ľ�����Hp��z��y�����[�+ԫ�ԔLY�<��i5̥?��ZKX��,�J}�b����j�y� �f�[�E�X.fC��&U�0c�s���=�{7|	K�.R#���`@YdD_��F�g�)¥�{ �* 3�}�����.�LU;����E��mv�H�<�Вyc�b�o�ì��U^ڧ,��'�&�ĉ/օ��~���m�G-�!�1����J<��]N�/3�4��~�C��r3	��w�k=~<�aq�����@������&��	�N��Ȼ�ZJ	���X	   Z   Ĵ���	��Z�RvI�+�� 3��H��R�
O�ظ2�>��j& ��ش�?A��[$���(�E�r�c2��&��s�}m���?	CY���'��6O.���.n_8d1�I�TT��k���A�p�ش)iqO�a��d��Móg�$4�H5Ѷ���=�
��F@yB�@A���#^��$��yލve��=�(�*�E�a2����Ȍ��X���=3��<�A�B=Z�'�+G��� (���p��n3ll{��lV��
��ۼ
���.	X�|�T���I&c��8�DʣWP0{Ŋ�- �� u'�i���K1/Cc�	3i|��c֒|�g� W|�Z\E�zͫ����	$�ɠ<]�Dd�I�(@���Q#����I����q���DJ��O�I�OZ�q`T>��5�B;02R5���>�W�5��➔
C��#/�u2L�?J!&���z�u�����"�O�x�#�] E5N� *N="�`��o\�a5�O����$A7��dD�)KNiұ�%߸���T��	=[��������`dH�i�Ĭ�G�Ëm��Ȑ��dĝ�OH�@��E���l�/��=ha@ĘL,�T�<�f�;�x��O �(��C�rR&�!���#�^6)��((���8�'v���>����sM-MT�逬��\[l�D�Py�0�pi���i���������� ��%�"?�$T�tCJ�s%�$ w��<q�M ���$�@F��#��O�<�'�Q����34Í6~-��H�_�x��?o ���p�_]H��O�#�(�ñ�3D��u�   �                                                                                                                                                                                                                                                                                                                                                                                                                                                      P   b
  	  �      �(  �0  7  [=  �C  �I  =P  �V  �\  !c  di  �o  �u  ,|  ��   `� u�	����Zv)C�'ll\�0"Ez+⟈mZ�YL�I07)��Dw�����c]f^�aPnӗ[��9� l��t�(�iҢJ�1��ݱ��׏X<X�;t���'L0+��PD4��gŃ\�^r�e������٬8R������.^�Y[�&���hq��|I:Wj��|�D�LE��H��������N^lq���ɷg�*ٯ(�>�ش'�����?���?!��L��m����3@m� �p)eY����?I��iU�ۂX�p�I*rY������SP�[��6v�PU�?ȵ���(�'��'�BcB<�M;7O��T,2kB|���U�"� �@B�<ғڈO�7mI�e�T�"'����.Ы?��p�'Y��?�I"-�����xҨ�~C|]�3���p�f��)��?A��?I���?���?I���m�1���N1�0ّPK0Zt۶o�On)��ڦar��M��xΛ6�kӶ!o��M[�}M��1c�����9��V+Hv���d��ȟ�m�bn2l��h��M	?Z}�yC�ڤ*.& �����ЫUy��Uo���M��'��G'E j�PqІ�PՔ���G̋�&}�)�n��kJ�tG�uzq"�O��x �����@��%�p7�Y��۴Pi�Q3 �2Ɏ()�A��W#�A"I� ({P�ʒ.�v�d��Tn��U��#eI%��.�����*!��nP5k��ٹ$��$dd܅b�Cx�p��ΟKz�7�O���شs)�]Ce�%Y�%�E�z����'����hhz�$�X�E[�j��U��� �D9�"#�V���eDן0�?I��-��H�/ƦJ��L#J�?����'�2ðE�:7�,��`Ѩ�p0�Fa�'u\�+�OS��Ȗ'�2�'e"JoA�d��E��'i�&M��d�H�޵e� !
y���7�/)]ax43k�Ѱ``Y,)`�I���'*�0҆ �:�x��T��dUn��
Ó4������'� yC&*�)Q����ەW84d����?A�����(�����
L�"� 9�������DA�'�p��L,X7j��	��h���1�r��A&'O>��;Zǀ�%P�Ve;���z���ĭ� N�Z��v-��9��@���ʵ��j��:�P�g�G�lײ����a�Ӥ��#�6`Ss�W�4����ȓMp�paF+.�&Et �ȓL|�9��!޲^��*s�G�|� �I�&�"<E���{���@^�26}b�W�Z"!�?eǸ�f��9 Э��@��*s!�$W=E�� pBb��s:~y�O)W!��϶F�����Y#څ�c�Ӑ5V!�d"0T���㬁�K	ڀJa#�M�!򤏯m�F]#���V)��M:b��Ii����s>|Qr���(�hħҠ<�!�D�& �YHW�B2i�,�ۂL�!�!�$S�_�na�@!Q|���7�!�Ċ�Rv��i&뙛qc`h�@&T!��VC�<�;�H�}H���fd�l��yb��7yJ�7�(?�TE�`����^1��`�`��t�'3b�'�Ҭ��yBv������t��XBaƅ)���qk!��ǅ�<$�0���� ��)�1L�8)9�����$=C�Q#L�~d�(�Düv$�@*T�,2�DH��D�DW��'B�'�P X`J4=���&"��
vX��^�(��L�S�Or\�	w��$����ا4,������ D՜��7H� 8�v��B#��?�/O�\�q�̦1�I�P�Oq���'�̘�f�[#���adf�'%H���q�'��@�wN�Ñ$�.+`���FW#6�PX����i�it�=��,��Nf.�#S�\l�ɤ��+d���'6��4�á*��"���L�j;B�Q����*Ȯ�h�Ò���D߃a2�'��OW1���SӈSʜ$i6E� 22�s�|2�'"az��0�~�&�M�����[���O>AE������Hq0I�r�xQ!��8}��V�'I剾WM����ȟ �I៬�'3x-�"�Ձn4rh����v����c٢3�����O��2�
$=Q1�1O�+�J��KC�m�X% &L:-}�!r�G��~U��Y�R�t�����y"F�,NXB��Ȩk�^�3 *B<�?��O*��W�'1��'���2�b%��T3`��e��F4a�!�$�^��}�0�
,x����%��	�HO�)�O���<�ڒ��;��}��l%5���ǃ�,h���'9�8�ag�^	��բ�M`�J�ȡ�x��lѾP�gG-�P���� q���	�'ֶP��	�t<4z�,pI�4��D�?�	�'6@!E�2J�S�ą�g�:EA�'�R��� �*S@d�xRc!p��XJ>���i��'�1i#k9�ɋy�l��S!4�BѳТw�V��	˟|�	xL���I�cԾ ��E�'�� �ᙳ�
2h�	�jR�q*��Rb�'V�9���a�
�rB♏?�6�Ț��0�A�g��X"��4ax���?����䕀C��Hѵ�C��9� 
�,��'�R�'��
F͕�~����V/	1d.!X�l�I�
֪�˃GU�U���g�?a*O�H2�����&?��O�BA��2�C5һr�x�Y�n�8��'�1�4
�������]%��uBE�ޢbΦp�J?�s�/ݨi�t�z�ύk��e�ՙ>��d�-� 5��Z&O *��S�dKb����8�t,G���]��nE<>*���M���$�
y��'��>A���(�Z��1T �I7I�4b��a��|�hb����P��郮ܴ�8DFRf2ڧ%�f����38Lj��@�	j���I�'@��'���� Kv%� OR:f�5�AIÇ8�$�Q$�Y�>�����?��b>)���U�	��$N�[ɾ�2�_
e�JPbRLX*M L���1S� !��k����������l%J�'��e�anG�l��8s�����`h�i8�7m�O�����O���䟎��O����OR�Z���a�nY��"Z=-�j���a'T���c/�XrT��͊e"`��]�4���D�ϦE��Iy���~X�`�A�\����@��%׀�:����'@r�'xP֝����	�|���HM��u�[;���F��"�h���B�H�d�Cn��XĆyX1�ɯ.t�E�S#�6X�IH��`�4���IS�	G��GF�D 
�KJC���O�E8"h�!���D�B��h�����'��'���'��O��h�cǀ!Fؠ�MȻ9et(D�$D�$��I���K��^���a6#%�$���-��[y��[~��7�O �dW%9ՈXg�*��a&(^T����?9�CL�?����?)I��O��h���<�w}�q�Gj���:P����+�TzÓ{wDm9�c�%\����3�� �jPJ�̐�D�^�Z���lz*%��,~�,����O����ͦ����-�R�G].8A��b��
,��ؗ'�r�4�Xb�@+�%Cr@F`ڱl1a( �4,;�OLoZ"�Dq�GS�(ԫ�Dǅob@[ٴ��DuK*xo�����	y�t C���Eō��!���t�nX��A�H-R�'�.m94i�=l���Ot�'���F�P���P�jM�J��0aP�x��	
�`�2��(n�,u��\++Ô#|�ң1I^�t�0FR�I�}(��|~�A�$�?	�_�f�'�O��ɀ+z����ď��3����t�'��\~r�ёX��0��I�9IT��*����M�³i�1���Y���ZdL���+������'b������Q��u�O_늅(��P�SV:A�բ*D�����2�
�E	o��8�+D��Z���>��~�0�3*D��:���$p0iP��߃8��0���2D��{��D	�аb�^���p)2D�����ߦ!bh:�B�<b��s�<qV�t8��`��"gJv��eA����-D���Rn�;Ni�7��un��{�?D��`3�Y9KAx�[�ܳk���{G�>D���Q�ǟ��9	�����F&;D��0Tŗ 1<i�	ˎG:t�
�,=�O�	�E�O0 �0����ce�$V$�})1"O$i���-i�@�x�e��>�!!"O�]�a�N����t�Y�e��ѓB"OB�r%�Ǡs��Ҍ���4a��"O�0#	�'�Z �FP�B��I�"O��a�G�:\s���4&�+����L�f�~��g�@x]Y.ЋK�̰��La�<����bS"�hv��/�dta��YQ�<I�c~, �
50��R�<�VgF�XaZ����CFڶ� ��K�<�ТY��AraQb����3��C�<iKQ��ah�-��[�b=�PAٟ��N"�S�O����/ �F�Zmؓ��Sg��H�"O����(� Ht���1DLt�{"O����sS��	�B:�c�"Ox�Isb�~��m�e,ΉJ�L1��"OP�acC��2����.4�:���"O$5�e�#� ���H�>'��6U�Ly�	9�O6!x��4W�e��	ŏD��T"O� <Bub�c �$���� /����f"O&���8i��ũ��9��1{�"OI��_�Xo'b�	9�9"O
1��EF;x��×Y���`��'$��'k�PG�4Q�Px���syt���'),��Sa�Z갼���	5gy����'�Nr��	3�	�@Տi��p�'�0��ƥ�I�|�^�t���
�'o�����;k\ à@D�6(3	�'q���$�Lv���2#�4S�p�ʈ�Ĝ#FQ?�[ꗸw��a��䎪pmFU�Bd3D�X2c��H_F��䍶@��
A1D� ��H'4�����/ǔ<����4D�XR@�߻v|�0�,Y�_伈���3D��qSco�%�U�Y�_n� bW	?D����P�K?��U��>nE�`��O��C�)�'C�hBc�^�q��tB��ڌ@����'����@˲��$�Oś3j���'��R$dѪ_���!�v�lU��'y�] J��o��dX�M��j��A�'�lM�k°W���Sw�Q9a��)�'i��j���)�x�%,�|-O�}��'O��ViTM���Ql�}k����C�S�#�l����+d����_�ҕ��E�(("�S%=� t��J?ʝz�H�@��%3�

v��ȓ����a��&%�>�bsL�8�p����9Gp����W�^���@�o����. �sm�B�I4�u+���>��M���^;ĀB�ɻ?�!��j\�P�ĝ*��Q"A"C�I�y �Q�Nt
�ՐFN/D�FC�I&��5a��Y�NCn5e�̪\u�B䉈!0�#&�pcP��w�挻W�*ړU�x=G���]�an`Q����+�ܙ!%��y�DP_���%L�(�.-P�(ʁ�y�'�3�H�h׊�B�Q�L��y�h��W���:h�5`.�A���
�Py"�
1M��eq�NB�C�d 0D��<i�d\�� #�<R�1�d����ʗ�1�S�OQ(�HU����<�~���"O,tvA�#9h���V�?��="A"O@���W�s���Sw���h�θZc"O`͛�I��#:��1��\�z�s"O����Gq��X���*}b�Ҥ"O�8����j�,�����k�CRy�a��p>��ǸN�ՠ��7�L@#�o�H�<a�힗R�
��g�3_��h����H�<��Ɯ4aLZ��"��9x�AAD�<�S�Y8^��%���-I�*XR�$�A�<1���jU��L�x6ԅ��@ASx�x(#���T��C�U�4eaC�o������'D�HM�K60��OG9a�	�w�2D��
�&T�~"�Q�cÄ:y�Ԥ!�n/D����I�#���f�ƅw֢<��N/D��@���_��Z���	"H��a:D���PǚS:ֈ{�Fj�4�ۃ.ړG��)F�D�
�q�t ���L�n��Pqt����y"��LyԦ�m���*c!��y����]�aDB�^��A��]��yR��4�y'_�1��A�a�/�yR�P'M�j$K�
��k�� ���,�y���`��\C��gS���r� �?�1�J�����mY��X�A!x�sJ�`Zƈ���#D�\��Ei�ܬ�u"D�s�+�.D�� �A�EֱU��D`ƘQ[0$Å"O, )�瑍b㦍�@qX��!�"Ol�W�Ca��(Ɖ[�g��4)�"O|�!C��|XX[�)�#[�	 �^����>�O��A�됨4�Ҩ���a�-�c"Ox�+��P-vZp�0g�w�L�w"O틓b��?H�̘��X�>��B�"O@���"g X�%���e&�H��"O�1+�.��1pv���ݙbsƱё�'�8L*�'KT��n�*@c�"Ї,�@�
�'���e��FY3�Ƞscl4
�'І�8����*�χ�E�l�x�D(D��-C*^eh�Aa
�hȄ�s2�9D�`�N�6B�\�&���!�"=D������A�Rp��L� Ύ-�D%ړj��YF����/Rj�a-1��H��I-�yr��4M� 9�#��)��V��y�J�U���q!P�N�uK� ?�y�bO3�� Q�-?G�ĕ�)O �y"��q�!��S�<u�a���y�Z8:Z�A���1e���擌�?YT*�[�������v" �Q^
��g�L2��,*D��Ń��&�x�3�	-Cb$��qk&D�ڷ@H����RmȘ��u�%D� ��K1�� �i�Ym�-#��?D�4����䦰r�i՞Eˬ�B��"D� ��%\�S�uY�cѹ%D�� '�<�!��q8�4Ȥ" NGH5ѷ��+V��@�8D����)O�����:W���0h7D��8aF
��]�Rhˏ��pR#D���c�.D��@9�(^aj��!D�$pGi��O��n:�F���� �O�H�O�T��%�Q�n�Kw�	?n\�"ObX�r�	 ��8
�`١sH� ��"O��I���V�А��3>3|���"OZ��&ꈇ��t��x|�!*A"O���oK3=*�X�5v��"O�Lۢ*�#�̥�4C�J[�I��I�B,H�~���C
q����5FG*b�U!��}�<�$����]s��Y�U*�!KFx�<����;/�	;5%��/�|�Fz�<��cӇaT��b��!+J�#Ou�<����Bn���R!֞E�f�;��r�<`�����@e�Ș�дf�d��g1�S�O�Hz��U���2�D�gEPHXG"O���C��$�}K��>�l�Z�"O��A��)%(�U`�-��B��w!�D�{�����f�24��Pj����!�8���Q#�+�����x!���_b4M�v&
J�D�엗E�	&W������<9܌��T�ӱ������!�$�{W��Z��d,�+��":!�@$l�L˶wa%&�&x���3�"O^|�"*K��$X �Õ8��Tː"Od���`Y�Qqڙu#U[�Ȁ�`�'c6}I�':���S@B�Zm ��/�90w�Y��'��8A��P�(t�JW \��Y9�'릹��+ѥ��	��)M�!�'�:`Ra�!ҹ�	�Bά5Q�'�"̈% ϐ�|9*t�.� �s�'���C��� ���۳�ݡr��mS����ZZQ?ѡ叉(=YL<��p��!Kb'D�h0��9w#��&�	�gL\�IU�2D�� �Mꕻ�NȊ3�DM��k0D�� .��ք۩_� ��\4c�� "Ofȫ�,�~Hd!�'F���f"O�԰ fی7�-��o0Lߊ��1�'�H0�����]��|�CN��1q��;���*|�0 ��M�H���
��	��Ề @�j�Y��:�����%� r
�"�-�f�p��ȓ#x��!N�'��: �W(y�E�ȓ�.�����O�*&��%�n�<9�bY�I4�`F�}�(�C�-�ly2mƖ�p>�r�'M��b lG�DHE;s Tf�<�� �%��Pçj��2��'�X�<aq�L-%�q��@�ov�z��W�<u�ĺ[ٖi�v���K ]R��O�<��(ȫ1A��+��,� ��b�fx�D!���� 0q���qQ��#D C�{W���r�1D��� �QW-J�sJ�2�`�0g0D�<���^[̸!Wf���..D����F�;�h��`hA�d"��*D��)D��a|2��_�]Tr|Ҳ+)D�T��.��S(���F���7�(�]jPD���R�,�����#T)2�X�'�!�y�b[9~�T�V S+V�b��C��y��5U�8Ao��R���!��yB�^�	z�I�ŋ,C�$!� AŲ�y"�O���	�><Y�7�y&�HQ6�rBA�:L�S����?y�L@���� 1�
�� ؀�)�h��l\���6D�4K��>m;b8[�ݗj��3w�2D�8ڀ�@���1��ݤ}��E�2),D���Q�ҁs"h+W�׭"��k�*D��z5/Ӷ �i�V�Ӽd�X��&4�t��FJiy,	A��#���2�G�ǟ��O��'S2�9viX�<9��OL��]NH\�fJA�$ZrQ��	�ln���Ob����6<FP��$�Z^�ŋ�ߟ���Ɖ2PN��	�0-��x��#>a�D#gj�500�ӻqpt���|Dיm|t����Q�$���a~�'$��2��?��4Hȶ_����U��8DC���*���O����I�"a��]�!�|8
��Bt�}rL�<)r�/R�n�#2�:?%����@fy��D���'�Y>3��Oϟ|�ɷ(rr���G�|A��"��	hl�I�F� ��bD"�4�E�@r��uџ�c>���M��ag@pp��*&T��4�b��b5!�P�t9c�͢}����JX��H��H�];<¢�s�KB<��A�?O޹�S�'�Ҝ�����=���
�h�:��y�aHн�H��ȓt�$�(�61�<A�Wa]�R�
 E{��"�'qVL��������×l�pڦ����?���;eXq&�U8�?���?9�����vqj\3d�
�]�Lh93D�G��9���5tq� ���,���ې���XR�0�p�4 N�%*�� $_2&m��p lA�k
4��!L�<,��R�DR��.��d?������s�����R-���䬁�I� G{�<OZ��hؔ�(��9D6-Ab"O|q*g� � AubY�g��e�!�'��#=�'�?�)O|�c���L9�)؛x$n�y��9&ڢPR���O��$�O��$�N���O2��� ɒ(�I�&��B�S����፞^����UKޤ/*�@p��OTHWC	�J�|� �����Jc���f�`�B�&��iЭ��&�G~�g���?'I	��pu �	#���K��L��?I���!�Y��t�ӫٰ@��K�"`��ȓ3U��0ʌ�b�8L��Y�~��d�'qt6M�O�ʓǺ1��S?!���|�I�9��t{�iƾ^��Lz��ퟠYƥ�������E�C R2��J�ˏ�i��tB�\3F��.E7V洌�%T�
Ā�iW�a��䑅�Q�F�Kdf� t�q+sk���u�Y6t"�S��B0}��5)�o��шO8���'���)�����W Q!n� ��B�*���@��dJ��#=S*@��M��I��2�ON�':F<ZƪH�P�a#Pǝ�'$`��)O����Obm{2��<-�����OV���`��Emp���
:r�b��/�O�8"�!Z��p�1{P�����O?�#s�!�Π p�\�Ak-���a��`���7w�e"]):��hF�� ޴ �PD{�iE?Z�Cd,��y"kE4�?1�����䘟� �8����PD��f�ݓP_	�"O\	��� L�\��N�<�"�I��ȟ�HW�� ;g^<@h�?#�VE�@�I;�����3�ـh`�҅\�
�C0B��:e��%4�hQ`�h�F����ѧw�h��ȓr��$�����d��rNN/xi��6(l�;�̓3j(����Q�Bܚ���+���UMZ������%}��d����3TP�3l̟F̅��.N����$^IJ�H҇NXiI�v!�]U�4(���%$Юpj�f�2d�!�$�.Z��bB	ù0��5��eak!�RxS����[��	"X!�D���BK�{hT`"�џ��g'���MKK>�ǫ�'1A����� 0�<�c������O����O��#�� 	Ip�)e.H9|����KW�p�@�kW?z*P��4-6<�P蔻^�Q���&�&C*�i���O/8���sآl��y�V�A�l1�H�!�r��3!P,\�Q�����O��Op��p>�:�FY�T`QN=;�"���e�O��D'�)�'e4��9��J�*J����sP)��k��	$.@��N�G���b�Nª<kx��?����?i��4��LR0k";����S�I.W"�����2O�=q5 �`U*'��*gdT�C)A`��M�O<	�,5�ӕjf 0��R\pTU�`�6n��8�D��6��S��'h�T�ҷ1�`�!T$��f�)�&�x=I�O�OL�ƙ>q���%�ԒfE_ I�xTs�)��<�Oz���h�󤈩 ����ga��R9��4$�$	�Ќ��>��>qb�_z��RK�4�U�{Z�]PT*��i)��C�$Z��?���z��I7>K�?ݣG+֎6n�:r.[�h��qd�ԟ�(s )}rC5}rˉ���I?�M˵�P=Zȃ�}&|�iGnky�OW���ɬ�ȟ\%�@��'�=��IǊ/�\����I?Q�͙i�T>�	'+��:����U�@6/�h�(��@|P놫K���dРIl���Of��=O c>�R��Z�A�F�
��̆()�D�O��A�'��p�O�s�0)B����C2�3�Xa����*Pyp#�O� [	��2xp�&"԰ �<d�FC��~]�����|�1��n���;fV"¾hlK�.��|��=��B�
$�Cო"��K�ꓑ?�)O����S�DNG�؀�MC�L���1�ē�hO���$���>2�]Yh�:X���"O��z$g\�N�!�a&�2RB�;�"OvU�T�-n�0豤Q�b�EPS"O��и�M{wᗑ�P�*�����y�oņG:X
���-�j���yB
��X���0va�. :�p�	U<�yr�\�=��E-sD2�i��	�y�@@��se͌�eL`"�Q��yrΆ$>N�((�O�N�X�l���y��6S��q�2"�4>l30�
�y"+��z,�ނ��r<k���y�P!x]"��~�lpH��+��'h�QuD��V�ڔ�81툕@��[[�}����9�0�3����9��Dv6Q8S��>]v�z�,��)'�@ "����r&��!���92C,��y�n &�uA��C5+����� C�@&���"a\Ju$��Oc예w��g*�`� �,�P�OB��JU�8���4N�7,>�	Cv"O�\ ��7�m�sB�/>�=�"O�! �F8�4bڴm��4��"OLm
u�+��r�C1+�>4Q"O$ՁpO�$!�R!xT�Gk��P�"O�� ץ�
�"|�3o z}R��2"O��3��x&B����&j��`P"OZ  ��A��P!M5U$Y��"O����L,�h�D*�1��8�s"O	k���]�����ߵ"��`��"O���+ГI���AE���v"O�;��L�P%��hM�>���)S"O���a�ܬ5��@e�:?k�	��"O� �����54�@�����|�"O�uc�g�;��8"fe��Yc
��"O��I�$F>l_���1�TI��B"Ot�B�iM�4B�E��#7���5"O D2�#��no�يQ�E�"L�"�"O|h�F
�E|Q+�A��2� {�"O�@��Ӫm�H����!^���"O��+��4%G�р�X�$Ĺ��"OV�i��	�
N���O�1o숝Ó"OZ0���*v����NU�V�8&"Ol����	o�,`SO�jCf	�#"O��!�	�|�.���V�/3��C"O*�P0���G"jc�R$v$v��7"O ]�#Z-[��4JT�'G�p�6"O<�At�+�\	A�a �y:b"O�	S��Ї4	R�i"�ҏY��T��"O��%�њ`H�1�.�05����d"O���l͵Y���t-��M�QӦ"O�8�p������+�$y&0�1E"O$ ����$?���&���h2���"O�IQ���YDNu�f�Y�T0D�8"O� bt�D?sL<I"����q�"O�����/dkn�{e	܅D�t��"O6��ҮX�7	��J��#��U�c"O��5��*�Z��be�(��&"O�x��+s�&e1�Ę.���Hu"O�� 钑uZ�e*�"ݝ���R�"OF��+��<�0���cW}��x�"O�D(ef�))< Ib݇
l\�k�"O� c�F���TA�
J
5c��"O�
OZ�+nT1�o�of����"OH[�A?2��"eOt!�"O��3s�߇/V\�k#m�/N|���"OlDQ�l��W:4]��k�j[���"O��	q��7��x�#ʁ�=@`���"Ov,`1I�)%�j�9vf�)g/�q�t"O��ap�9���X�b��_%���"O����H�/�� r�!@0�}�W"O$��Rh�+{vD�p��O�l��Lj "O$L���;eAf0kR�F*o�h:�"O���!W�Z���Cƙ_�d�V"OH
���b���{�"ӥP��aa�"O ��5(�aH2D9�At*��"O~�c7}�0����5Pm@R"Om�l�Y!|J�����	�"Oଚ7�؄n�~|��a�`��kB"O$h)��7����P��m�u�"O0�s��ZEƺP���S&��(8�"O�p�D�	D~H��3��%����"O�%�!�b��h�b6q�Ƀ�"O,|��H߼
2QKJUt.�s�*Op�����9}pB�� ��BP�y	֚OK�<�m�&[��٩A�ˑ�y��8^+^E���U�F(:�o���y"HC����J�0M=ļ�0 ?�y��!'�%�u���@=�$�(֯�yR�A�pd͢�lռ4>�l�G�	)�y"�(C���Cߙ(U�� Ĭ��yR/�
c�4E9�� di���y��>w�}q։�
�c�L��y+����d5e߲5�@	 s��yr��Fl�ڵB5 ڒ���1�y�$U�><��/æaqb�S��S �y��-.��\a�D��\�v\����y
� ���$n��Bh�Z�	H~��w"O�dxң�29.�LY���ߪ9�"O
���G�)�`��@K�8��0�6"O
!�)ŅF�ș#�i�a�VH�"O4D�7T�({R�Wnܲ�H�S"O*��"˖�~@$ ���V��a��"OHm�p(ڟ'ݢX�����F$ZE"O���G��3=��!�%K��)�"O���s�˶3�� 
�#� ���a�"O9w� 	�����/��-�"O�H��B��P�P��3m�jE#�"O,�#)b�2���b��a�Q"O��(���>qD��*��K�/�2`yS"O��Co_�]8J-����"���Ag"O%ѧʊ���"XY��h`"OD�ɴǍ�p�&;u����P��"O��ې���0Cj�Jp��=���E"O���Q�� ������;g �-�`"O��`�Ò�+���5�Y(���9%"O\��P�14���L�,E9�"O�l�$b�=F�@�`�ڬ(٤�Q"Ohr�kD4aF��j��"O�izF�G�uH�E� <96�0 "Ob���Z0Nq��cCǣz�I�"O�P��<1�" �5+��9p"O�b#BJ0R�{ӡ��F��y�"O�Qh3�Q�J�D1�7�����	G"O@����V*"��9��)�}q�c�"O&�ۆ��?'x8`���fcH�7"O�ڶ���8xR�@��I �Q"O�ظ!J	r�|mZŋ�2���Qb"O4��S�L�! ! ��M>��"O�!���s 5
�,mV�9��"Opq�
Pa2����J�W�dxq2"ON��T*�#q�&ph'Iۇa"�K"O�L %.��,"�i��IZ�g.$x��"O.A�e ���^5y⑈���"O�-X���.�A��_�J�|yD"O(��$�8x;���l1x׊Y�"O���O	��Iх��Պ�+�"O☠�D���
D�Gj9Ϝ��&"O�(��C�B��bʆ����"OT�;4��~����h����Q�"Ob���+q:m�����:D�a�"Op%҅*�?mJ�	�!D�I7"Ov��􇈌�ddaD�G�f'��!"Ov8�+I�=��x �gي?�X	`"O��aNQ;@��F�? ��C�"O����f_�
�;&'N�45�"O�]j H�(;�V�i%%q@�5"Ot��0+�w��"��WiaK�"O���+�L�z<:�`�4	��m3�"OX8���VN@b��:>�<}��"O
�I�f[ /���4d�(�h��"O���"����mseɝ�Mrf�
"O
E���W'�Q1�U�en�	�r"O4�B蝬2��YA��`fp3�"O� �G9Yz�� Oy-B�;�"Oʅ�i�~<L8@�@�5*t�*�"Oĩ*���/9�DP���-'N�c�"O`QB,
�˞�SG ٛ�L;5"O@uB��ʧ#�`��o(Z�p��f"O艂�ǁs���0��v�ڜAw"On����HtTLq+l�+�Y��"O� ���Cm��S�R����Tk���0v"O�<PnG$��s�ɒ$�r)�$"Oh��Չ́\��c闫#�P髕"O��� C�67�U����:��A�"OZj��B�fb��4L<$r4ѰB"O��r����x��b��ݸEc8�"O"�y!�,reXq��h�<'���J""OĀh�
O�A��	Y��E�o�4��"O�u@c-�Kju�F���V��"O�Yx�%N�Sf��ɦ�!-f8���"O<�X��+m\��� ЖD��$��"O��	�B6y@��T���u"O�ȳ���}R���p������w"O��3dO��j��:"��{~ iaE"O���a�'[���[ �Qc�9iF"O���1MFe�4����f����"O(�X`FO�`�t�J@�N`���"O�%H���	�tq���&.8�1"O�sW�V-$vͨ�i�J*ъ�"OrD�Q�P�O���(B9Phy��"ON�H�@�P���
J���1w"O��T�M��j�be��x�h�u"O�"�ZIN�$�O�`��KC"O��s� 0֢�sh@�*L�8"Ox������o�#�][j�Z$"O�9B�G � �ZMJ�n�-%U���D"O�Q����
��a��ЅDv�*p"O2IJr���k@�Kv�Cg����"O.!pA[�P�V��u�Y}�\jG"O4�j�#��^X�Y��"|�yp"O\z�kAZR%��C��xNA��"Ol ��it�V��V@����"O0)��(�rzD�p �5`�ir"O�5���;-J���͓#N��"O�!	�� .��SE��;�i�c"O(�J X/`�
Q� �I�p&�� "O�`j�OҠ#�(8%�ʌ[r���"O�A����a�L݈uiˣ?S��0""O�@T�Ĝ�kp��j@8$Ӈ"O���'�=4�`�;���!J;F;�"O~]rd�npI%O�t6��@"O8�!���`���3s@#`���"O@�3�^8<t�����P�f��p�"O�X���S�!�% �._�
�P7"O	s�Ҙ���I ���(L��"O������P�V� 0��Gf� ��"O��`bѧ(rn�Su�¼(Z&\@B"O!jv��CL1s1��IEÆ"Oj0W�B�#0����V�v"�ac"O�Y�MмT�(�j4KQ�'jy��"O�)!�C�9e�(��$�.X�Q"O���k��AR�RB-��Tf�р"O@�d!Xo� 	:� /`� �"Oܥ��#(KW��!���.T���p"OzI����=£�ߣY��i)�"O�-�H����@�����,��"OĤ���Ԇ��Q���܅J������J5A�ph�%"�,�t���-M��'#�Tx�˕hUڗG31sJ)
�'�pq9eZj>�Y�&�(	�P��'A�y"��H!x�y��
�w��@�'hP�Ól�.��-��⍿pn����'J�lp3�
�7f�#��S�t�r��'��xQg������A)؅��'�@����&�`ti�6XL{��� �a�+8�F�`��9W�~�d"O|���� �cg؜����%��ʗ"O����͗{�h�3፷Y�j�"O��arØ�2��6�J��6�{"O���a6�)���s�t�A"Or�
��ٵ'��G�;JҸ�e"OZ-p$c
�X��a�f�.]*��hR"O���nQWo��ZD�;y�Z��S"OH��ℙRl��s�d^+���(�"O��Sb$�o�*Й2�Z�3��!۰"Otĸ��E(���q��y�l�*�"O@@�T�%iظ˶��$�J���"O~����ZTز1c���$pP-kB"ON��@��)�����Jy&��E"O�t��Ɏy��+��L(!��"O��SÆ�k��9�-�;L�fm��"O��v��y��I$��	��qh�"O��"R"KvVF���DP�T�yg"OL�K���n�ec��N�a���"O��٤���②�*�l(�"OT��� 8�հD�,���Җ"O�'��GL��ه�d�$Xp"O�$�P$�}TJ�J�dȰ7�����"O,PE�ҡS2&P J��6�|�X"O:tZ@�µ:�D���7�� �"O8�#&.ەc�P1��]����@"O8���W1@����ڣR/�]�"O3b�<u&����J�;�P��"O*Uö$P�,>�	#i�fGX��"O���STA�H�h�NF�80"O� 24f@�k(�ےA
I���Z�"O�I��"<�	���V��[�"O�7�=�8$��!A\P���"OXsv9�P�j��zN��"O�q+�!�9��V</��q��ME�<��.�Tbz5�!苭q� y!be�<��ň	�Juʁ�Єy#@�2���{�<�v"��;��\�4�E�(�WgEz�<1����u�B�ӓ��@_�[�!^�<Y��(���#���a�2у��TW�<$�,%��Ub�εe0D��S�<���Z�1�|I�G�k�AE��m�<Y�(��5�<=)S@נ�q�ek�f�<!G�3aQg�H �^�T�\�<	T�	FHJ���Q�xū�e~�<��-��@S�ѡ��ĵ]$�;e
�@�<�g"R�2����$EJ�Uk~�g�]�<�0�&eP�b�,O�B};ᅌp�<i3@�]�B���I4���`�Hw�<i���-j&�7�  E�y	U�g�<A���1G8��@'����%�R��e�<���0a��īS��"-��%Ib�`�<a�Y������ό�jѮ ��C�	+`Sqx��
�J�N� Qy"O���c�D�ށ�t$ɠ(��1�"Otݳ4iK�3�<耓�JX�萃p"O�,���X��b4	^=u��͈�"O�y)����6ܓE��g��"O�D���]�a-��AA�A9'���g"O��臬ċ2��a��b�0ez!"Ol�xD�
�L �O?fĞ�v"O�"��$�2�JQf]�1���W"Oz��	H�oF4
 Ý8.q	6"Oz$A�Kծm���
EG�2my�xk�"O� d���	��9x��G]=�t"OT�7ƔL��`e��E�!2�"O^����M
h���Kc�D�$T���"Oj�r�hĊM�H�;E!��MX�"O�lb���7�ް V�֣d�0�X"O^xF@XN��e�^�(�j�"O���j�-d9���TE&�J�"O"d�
NM,���E�
L��"O�\���+I�pҵ	�I���r"O�u:�*�fR��'�Կc��I��"O��2U
#Q�� G�ՓІ02"O�I��$��0oT����Ʃ�]1"Ojt�e2�/V8k$���"O�h
6Á�jJ� ��
�\�Z���"O4mӢ�Ͳ l��ǒ�DѮ���"O�q��NLU�Pa��H�w�����"O���.L j��D� !�|�g"O������7�\��s�\����P�"OXY��G�,�Hp	@7`����t"O��cPfҪC�P�h��z|Ҧ"O�!Y�e�65���YV�4�yE"O�yy�ܼP. 9�ُG�\�"�"O��D*i�"�X4��2h��m3�"O��jI��Gb���@�b$b��g"O�a!Γ(�PR��\z���"O4��- +%�|����w��\i�"Ov�pC�';��(W�J7:``�"O������2�� F�SU�M b"Oʘ�RH�q���(��l^��"O\p�4)H�2��a*��Q%$�8�"OF�O��o�}��aZ�gon�I'"O���$�
i�d Ȃ���uj��"�"O�A��ȁ�A�թ6$C'�6�Q�"O��S�Z08O��1Yc�d���"O��K�L�\:.@WJ��_܎��"O&�z���R�T�*�IG�]1HԨ�"OF���_GƦ=K�JH5����#"O�A�M�3wo���^�Y���7"On�q�\�
�<a2D����!�"O�L���M�,$�d�׫��*���4"O�a�s�T�C/l����Q�j��xc"O�ԩ�`Eg3Fyj@���PqH�"OD����!EС�E�$��v"O(�� ͼi(�`� n�&��X�"O�(�' ��C�ވ<�H@$"O*q+��?)�;�x��	Y"O"�xP"�2��U���Y���A��"O�Lr��"~*���	ٲm���"O�	ᯐ$\B�X"�i�"+�ʬ)g"O,�3�7x�^�����;a�j0hE"O�����(/�*�h��D�6�"O� ARJ�0If���΁nؖ��"O�}��$m�:�y��Ws��Q"Oh�������'c�� w��5"OB<��{��3��kH��"Oz��b�/�	(� �N��k�"O��J��H&p��P��m�q�@��"O��#�(�8-nā��&�X�\t�"O�<�Dnݼ)hL	A�%�>1Ŕ�`�"O����d�dڢ
� �Pݪ�"O��j���>@4<cf�1Y'.�J�"Oh�@��p̚&i����+�"OҠ�H�?4��I��Z�vxp�"Oj-C� �yW.!�'/� 
<��"O� Dl�gK; ^�s�CJ=e �$�"O�$��钹DlV�s��� Vf |�"O���ц��P	r'I�-� "O�+�(�r�a0 U����ڣ"OT�[��۬v8�吧��w*H�=v!�ē�C۸�pB���>cm�7�Y;�!�$O�a�$�� K�UU6UI��W�!�!�̟lU�t`�1&q��r��$#�!�D�~M4�a��7	Z�I(���!�ą88d5z0F"i���z��ٞA1!��J�h��C_5�J��c! 	!��@���
�c, �T�27+!�DM��quBμ8{�ܻ�k�&j !�ĝ*El� 9��[�0Y��ʞ(c!��1-V���Oz�h#JF�B"O�y�)��|unPI�ׯP�q��"O�ų��͌6��i��G"��"O@	0@h�$�z�Ś!��s"OZ4"O!bM&�*�eD�gdv�P�"O�|z���'S�ĉS�	�yL$9�V"O�e��c�*[DJ!PǇIE�hٓW"O��vB�>.�5 ��<����"O��p�"H�kڀ"V�J�o"n��"O6;1�L��hP�t��Y� ��"O��%Mؖ�b��beX.yn"=YQ"O~��v+\�]�q���dUh���"O���m0q����S�h��"Op(1�I�t�8y@"�I1E)���"OJ���˗a�����#��/��c�"O��rA�][��sA���+�"O��2�]!A����ˉ0M8Pi�p"O~��jB=g ��h� ]�)�	�B"O�eRk�=V�$�ՄQ��"OH8���Q�]V0��F�y	hr"O������(b����'���o��2�"O�MBSJ��)�ݡ�Ăxj�Q�"O��&�G�N]*`5he*�"O�i��JL0� @�π�8�>m)�"O���D-2 ~1�g!(Y�V��"O05��Fڋ}��m����v��hQ!"O>$�oI�Q�jS���.*��@�"O`m#��Ϟd%T���۝a��
U"O����>�rѹ'��?)��e�g"Ob����/$��E��ON�i��d�r"OBة�2B*� Wn�9d�dE�p"OV��D��2��\��'�&pJ�"O̅i�(z���e�d�\�H�"O��NW�6����e+b�5��"Oj��=K2��E��F՜]��"O�)��ñ#$\X��
u_�s�"Ot5`qC�9}q��&�&{|��B"O��AA k�ik���?$:Q�d"O�D�%��|8"�X%	T�}i:A"O45�EiM�G��I�^:F$�"OV�x��'pH^ٳ��@'H<�XQ"O�IY6!Q��4 �DW� ����t"O�q����ʴI�,%��=��"OV-#4ڗU6�)�	��T��u�Q"O�k壖hƌ�`�)l}n���"OF<#B�À\�>�qǪ˅A���"O������
!��;���:���O(���D�>���ђ�_Y��'ʘ�◂�^q�=�4j��D16t��'������T�Sܦ<;$e�8���'5��"��mx���B`ᴥ���� �TїL��] N���Dɲ5O���"O<I�c��b�4�Ȅa
?7t`+""Ox����wo��&�3��$"OV0���}�Hr�N���>!0q"O�I���C|}�0����q��p�"O�q9�g��`wR�jg�Cg~���"O F�C�)�荂�M%7|����"O�h�İt嘒��5c\��k�"O� a�Aڏ;k��Ihh���"O:E#PGޑl��ȣ`/g"�CU"O�a�%�j��
P.�XM�4��"O�%��C�42��JO�Z��{f"Of��L?A|Y����O��0�1"O���]��F]ibjq|z�C"O��d���;�ʱi�b�Yi�P8�"O��B�ŋ2K�6��p�=I0j�
�"O ��V/[�H�I�0L~���"OD����O�g����V ��D~HK"O���׍
�~��]�����4Q`�Ȳ"O�"�D�u��(�a��>N�	��"O�|
v�Y1�,��艹eX���f"O�t��H�R��&'�C@���&"O$�3w� 8S���i��(��=9w"O��g΀.`��� p��:6"ORU0S`�N�(�h0%α=\�$y�"O(��T-vglc䙀 O�Q�c"O�����/%j]#�$<2Bc"O�� �	͖pM���R��B�4&"OhMP��J=�*��@�
�;�"O*0�4+H4��R�b�0K�Q��"O�-�@��3^�Z� %@N�n���"O,Y G�W�1
�K�E]1)�`�"O�1��u�eX�d�{�XH�"O>���c�����%�����"O���
�,8�B�A��ݷnV����"OT�xw�E�3*���k8!Eh�#R"O%S �YN�@�S�ʔ�x6�倳"Od��	��3W�:��Z�[.�b�"O0���F)e�H$R�kԋ ����"Od�p�+!�:�d��� �Q�C"O�x�ԉ		O�i�E*�
X��Q�"OP��p��(2d]P�b	�w�x�e"O�t��%�0d2� ��[�����"O6a�a �-t���
�HE|�Z�"O�q��bՔ 
4f�'rRx�0�"O^벅ҙ6�m;A�*."�8�"O��3c�F�OW �W"O�
A�����c1-��l�����"OV�@��R$���k� �a�"OL��,��*���JD�R����#"O�B����W��9�B�N /�2qI�"Ob�aM�B�hXQ	��>���"O��uჅ*�1;��W�A��%"O�YI5S}��dLQ B�:L[F"O��C�ѹ.u�0
��{�x�K�"O���@cǐ:�Y���g�<"�"Oz��1KN�N=�1qê��]&<��q"O�5"a�C6j`И�&���'.H�"O<)�3�S!1�5��@�06$ ��f"O��zD �u}��k�`β]�"�8""Od���FJO���w/N�a 4az�"O����YT��Xs
�^�.�p�"O:m�d�'c�Y�q��
��"O��ju�˘5��X�b*_�	���"O� ��Ņ�6�*��i�2d��"O ��AȊ*��̠�HPD�sD"O(a�G�4��e)D�O�7��(��"O��M�����d��m��D�e"O�ЂF)N�eBZ)S���;j��W"Ozrf)�Yr�e�@�L[�@�"O��:+N$��u�H������1D�0`�c+Hp��� 9�b郐a1D� ��S=i�9�#d�z���y�g;D�\� �J�1R2@�dMQ2(W�4�3�&D�,ȢKR�}Z�(��Hю:~bP85� D� ��2xnbT�����j�$D��qB+�e��@�^;4z�ڠO!D����L�+tY
�x�F�Z�P�c�>D��	��H46�حI�D? 
l(Ą)D��Rl��,%>��nVz�ҝ0QF(D�|ؔM��~I�F�Ek�m�!H"D�,A���<p����鐅'8�aX&� D�����ҳ"x�!!�&J4֢Y�A=D�����~����,��^@t�%�%D��i�/�A�j4����1�1Pb�$D�0�d��I��ق�cңp���Z�&/D�Awj�0l����
W@���.D�� n�&m����D�;Zr: ;��7D�%�ԭz~��s����}^�͑�*8D��W��8_�0D��Z�
4���1D����J^:�ڜ?�� ��]�<!c�^�'��8���4&󴥫BDBp�<)�F�E?�DѢ
ǭf�rY3��Gh�<)Ua�� [�Z�J�K��1� c�<y�n�:(X�A�cY�e��P���a�<	&&@�TV�}駥��#j �K���_�<�s땓QP^�A-Q��E�AG�<�ceW�:_քR��6��Z�n�j�<�$� q���C��L����jm�<Ip�S,�| ��fʹ�R,�]�<��N�V5Y�Eq���� �E@�<�ѩ_�K��y�Ĺ.ZQ3�{�<���+�*��ͽ�
L��fVu�<�W(M:m_ ]�`�W7tB��j�f�G�<Q2g�*(>L�+g�^�z���p��Y�<!��� 7V=I�፤RP�p�F��X�<A�oӊh+�Xs�JWMP���	EO�<�G��(XG�P�� ���{6jGK�<��ӭL�V�W��7��ˤ�I�<��.��0��İPX�Q4�g��G�<�gk� 86�a$̄0	�,��k�<�E�[N���ܒT6BY���Gc�<�c·�]|�X���4c�zPej�c�<A���:A֒�� �Fr|��$�e�<)B�J�OJ�u(��
����Z�<�ehȞ)�
E���ҍ9ɒ��L�<Q@$�/��L{2��	%���A5��D�<���ͫZ���q�P4�|1)�Ni�<��Fֱ�:}���9c<�p`��c�<��&�$�������2I� +D��_�<��m#se6=�Dc��DA�A�<)v*A�:�R�	6�d��
^@<!�9�2`(K�a�P��� Aڽ�ȓ�x�tB�?"�ơd���ȓ}~u��fP�1,,��"]�T�z����Ժ���݊�c�8^&���sX�@�1�� �ڤ���)�bt��@��T��/��){(�i�ܦ��)��S�? ��P¥���n�#���
��$f"O�D�#i6.��xJlA�E�tT��"Oe��J7a����%��-�����"O�t���כ5��!��̂x��e��"O���E-_;6�F���
ܞ�ҩ	�"O���@��>]9+/S<����"On��B�P$C���jS/T�
����4"O�1����b�U� ��
7� ��"Of�ꅯګ.�x��A␗S�:�"�"O>(���JT�\	��ʜ>v���"Ǒ�����F8�Q�^1�ް�D"O<�A�G۸PW@��� ގt0���"Oΰ�p��n�^�8���~L� b"Otɘ��;c唕9&��v���c"O"0b���;b$F�R�ɂC�-��"O��tBN�N��,����4I�nQ�B"O�!�M�E�pͳR�	�w�`��"Oд�ңOJީ��P?dq01K""Oʡ��
N@��['��,Slf��"O���k�?s��-k��26�U�R"O�  F�
 @l�'ƕ�j��r"O��Bs�ջ|�b�[��յ,���ۂ"O�թ���`�`<iE��6qptk�"O��vGJ2.S~e�N��EWH<2�"O؀C�	P����NK��T"O,Գ��޴ZT��M�V2$I�&"O���&G�"4�p�f��t"O�I�"G�R��-��`J2P�T�t"O�@�ԯN���!�)�5{�RT��"O��rU(S�r�B��S�
=+�if"Ox�0	�#RذSg�R@����"O��pQ�{� ��fD�d���$/D���R��G-d ��IV2�T �W�.D��0�f��(�,�cIJ*%�PT�b�,D����l�	Kn)�ôlB���o+D������\ څ��d˅8Ҝ�ȷ�(D���QD�#�4��g`�h���9'D�Ћ�aHs�DlC�a��"�z�9�C&D�$,�?-}0��gE�)sF�� �#D�`H�no���#��f^T���?D���%*�Q-BHq��K�E�Jx:��"D�<���Ҿ1�L��Ń� 6��,4D�|���LT�H"�aATr�Iu%.D���qZX=�!�g�X���*��-D���o�tKZ�c�c-pq��h D�x��A�7B&a�P(��1��	=D�����^�Paʂ�0��EK��;D����� hPp�7�$N\����%D��K�^�\����#,�B@�$D�,��U���ل�mL���#"D����I2$���"�U-F3֥1��!D�<� �cŲ4Q��W$
X�]1��>D��XsQ�p�� @g��l���A;D��6�AoY�p$$ٵz����g�+D����@C�'�H{��յ]�9q�i4D���F��~]��!����|d90�1D��F@���&-���>I�G+"D�T EBV�9���k��@4e��m��/ D�́ҵ����	ƻN	̡�Ə�U�!�]�v>`������L��ů�3�!�C6�((kpg�l�"y�t���f�!�$٣?"R���I��;�5�� �!�Đ$LtTkN� '�(���!�dT�*�B�Y#T(��ƣ[�o�!�� ,Q�1Á#��q�AQ�M9v@I`"OZ���i�Z���ۤo�<P:���"Oj is�ƕ�F�
H�-�a�"O8�rP�	YxL�a��h��IPE"OD���I&U�:��S�E s��B`"O*l
$��y�xr���n7V"On ؑ-	��ΐ
ԀX$ ��"Oέ��O��Q�"��u��"6�ɳ"O�xc��ɕy�]�vE�?� r "O�䊲�غh���򊒅0B���"O>�U�0ܺ�i �"���u�<�WhͭM$�A�H�<A?FX���Ax�<93B�*z���G!�D���y�<)U�鶱��D:C�����p�<	d�Z�8����HI�6J�Ġ6k�<��\+ �Z۫V�D����.D�\Y�D�_$�a�Y���4�2D��c��ŗ��f� �k3`,D�D�a���o4���R0bu�l+"�*D�'��(:�!x��\vi|@��e%D��	U�ս^����u��
G�h8�'�$D��DB�ళ�/DS�0�{c%D����,J ���!H�*���;��!D�$�T�֋4c����
�1��T�*O����4(���K��Z,Gp�pV"O���$���Ơ@/\e����"OE�#GG�ʤ)[c��@�л"O�L���dY(l�1m�\6v��"O���ܪlȚa��%�5.+x4J�"O( ��+>f������UV}2"O>� ���`����ϛ�&�З"O~TYp�U+5���"��"JϦ�{"O�4��Ú���,�>�t"O:�H��=4ON��fßJ޸��T"O�E1� By�u�Q!2!8�7"O
��A^�n��B#�nP0"O�� ሜW��sr�<��u�"O�,���r%,(�$d	&u�PH"Ot���/��cW �͝�xt¹��"O ��g�!m�<��S�X*+d�D�"O.��"W�^���X�j��9X�S�"O�@�"bF>**@`2p�A�qB�b"Oq:��$���S�S�~RX��r"O�4��D,l��#c�N�4t"OF�BsF��j�0@K�k#�=�v"O� s�Ȱwֹ#��ںzLkG"O��(BCE�b�<9{�nސs�T9@�"O��y�,�:w9�ݳW����2�"Ov����Рsn��@f�/����"O�1�&'�"|XS(ö/>F�"Oh�%/t8p��-��Y(���3"O���CK��	v�����Rs"OhA��X�����K���i�"O���йB�e2�	K�(�Q!"O�8�l�%�B$���yӮ��"O~@C�&[Yl�X�9��ӄ"O�mS��g�P�ҕVB����"OVP�@��8:u�icP%��2�$L��"OL��6)�6��GV�/!���"O 	��l��(�8�juBN�垜�"O�,�aX���l�%��(��d`P"O@-��#��;xj� ��XK��@�"OX�ȒO�Tc�e��N�R4&��y��ä.�NP�$���7KP�/AM�4��S�? xպs,B���lyuC�2w@`��"O�|J���-7kX�U���w�.t{�"O�|��DO�%��Ћ�
��G�=k"O���� �6C�I�NZ�Y�Z�J3"OX���Mͪ'����O:��$�"O yY0$J%*�d�K�ݦ{ٌ��"OvY(7*ߍz�
����
�u���k�"O�t;$ي�0������;v"O��!��h0�\PA,�>N���HT"Oڼ�s�$�昡1�[38�rp�"Oz�B*�,j������u��XP�"O^H�Fሹy~�*@Eљo7 �)�"Or$jF-�J�0d��G�cU"O�]KS�ߎ��3%�O!J�b��"OlR5�%c��~}Рj�"O,<�#�U�/���x��4Nr�DY�"O�d�0��64tN��R�{��c�"O� �'��q/���GU�n��1R�"O����Ń!��-�L�V��J�"O4t����p`d0�	� a�� � "O��6F�RUV� �JˣF�LѸ�"O��1q�D�gh1y�
Xz�� �"O��d"K)'�I(a��&hpU� "O�Ճ�jZ�q^~�1���7Iإ�E"O��a
^�:�b�ZD��2�q�T"Op�����#�y� �M�J�sD"O�[w�E>w��J��@3%�F���"O�q1Ń�d���ǦҹnDNma"Of<A��Z�LQG�/�eb�"O���ʇ�D�LA�OQ��pE�"Od�5�0$^�@04A��1n
\Pw"O�y��Wx2&��EEH^ܕ`"O�1#F���P{��#bBUTP��z"O�e�@�! ��0��7k8:[4"O��Y,P�B�@!#oV�����D"O:�� Gsy�ȃ�mз.��Q�"O�`�th�"N�f	i�L�6!��U�"O(��ئ(|*U��Q���"O��3���Z�ʝjBB�C�d�3�"O�p�O��yBtP�+�%I��a!"O<ěp*^����G7.���f"O޼@�"Y�xyx��ŁӨ=��"Od�ihg���cF2Ȭ���"O��s��E03�}�4�T [��As�"O�)���+B��耳J�w� �)�"O�-ӐG*aj �dD� c{jq!�"O�Ŋ��ڝ+�dR�S,7��r""O(IY�)�2�6xI����"O8X5��u�򰲠��8j||��"Op����ӿm$�� ��8k�n�)U"O^��睄0P�x�@��d�f ؕ"O�T��a�q�L9;�[�n�Pb"O�`	��X�B<c����^$Y"O �V��7Zs�=+S�L$���C"OF�1Uc[p�R%iQC�2f��)Q�"O.�j썪}=���ʝ?+�+�"O¹#�n�#3�0YzЂ��C"4��T"Oȉ�F�^��QfAO�,��@�"OnY���C./',q��&�0j�""O�ݪT�P��$,������"O�\��'I�`�Dҋ+tt��"O�xx#�C, &z3U"уAo8��C"OV$�r@L5�"�jW�� T[xӐ"O�����)g$@"��ΧiS����"O� }kR�K�y&^5�GA��X�"O�Ȳn�b�*T,G2K����7"O��I�X�����^�:�Li9g"O`��B͈+5���@1�!~�-+�"O2�	�=[-�S�ց#q�]b#"O��Z -g4������cl4�g"Oܭ���
`k�	u���W5`�b�"O��ypJ�1E��S��H8p!��
�"OƜp��|f0���%�>�Ji�"O�]C�T-~"�|�2��x bl1v"Od�a�@7p�c��P��"Oz�
��>=�Q�D�4^Ҳd�5"O�����W�h���H#$H�F�VAP�"Oz@&�7B̲���ߐR���f"O�e���? 馩�W��tQG"O6�[�ü ��!�gcǅ&�z�&"Ob��ua��i�t�q��)D�*i�$"O*Z�	�n���K"gmF��"O\��b��Sa�`��]�rWF�pa"O��ғ��#�vT!פ�@8�=�"Oz����G�NT�D��$98,���"O�$�W��>LR�]�7D/	:�a"OA)0�W<�RI*�D��� @BV"O��q%�����Ѳ�&?���
G"O����eE	�&�
��-K�����"Or��4���{H���bZ�}
�"O�,Ya�"J�<m��nA�|JV11"O����.��]J�`�2��s�6\�B"O�@d�D9	L�)�K��Gw�ɲD"OR�(s��8rlP��c��f��9�"O�<��&�7��tH��2�l���"O���MK6_��T�m���tI�"Ob�����|����l��d�f"O������;Uj��K��B�Iv�s`"O0�;2�9D�� ʚ�|�~�$"O �ۧԆQ�89���M�g����"O$]����"M*���2mZ�{���v"O���ShR���p�L��6Μ]��"Or�U��5y��PkW:���"O��P{��S������"O�����B��|)�
�5� л3"O�I�&!H4`�0��2�r���1�"O��8�*�#���K�T�y��`�"O�`h�g�/J� x�N4���"O8T1ȓ�^����1X���"O��dO?���`�T�|���S�"O���p�A�#@hb��O�jdƌ)"O`��N���a#�!u�yK"O��µOZ���
?d���"O���iN:���F暁'Zz!y�"O*$��mA�����=!����"O,:�.�#�ڑ8���5
��`F"O2m�'�Q��yP�,W%����"O�T�]�ej�x��k�5��͑R"OT�ca�ZH�։b�� ^�!#"O�S�פke�q�i��{����"O<Y � ��n$�&�Ee$hqa"Oh���e+��pu^�%[� Z&"O�t���ăD-*�s��X�r?��B�"Oh��D��%i�j��Q��t"F���"O��Q(��Jn`Y���e l��"O&��5ꄄSذ��m�c��"O"��#�Yt(iӳ.�<q��-��+9D�́�N�,.h)�������R�3D�� ��TI\������O�=d��P�"O�m�g	+H�����)6��qё"O�2�*�*m`2%S��B�~��}�r"Oܰ�p��o\����FF�JIJ�"O�]0u쑒Fl�%J�@־a�`HDxR�'蚸h�(I�5�~��)��#lt0@D!��*�b�˳�}��?Q�@�(})X���8(d�(f�^Q'0�?N]�4�O�&�Вd`�Z��#=�i���Ѻ�!ܕ!(���3�@-w��$HŤ蹥�+�J�0ǆ�~ؑ���F
�O���ͦ���L��*�;�~��@
n���X��� U���d5�)Z�}bNN#<����oݷ6����Y��p>�4�i��6nӪ��U���}�A���B4ʁ1��Ot�a0 ������� �Ok����'��i��4� ��Dj򮁃�j �d :s� ���*D���8X�L˛Nr�<��OR��?e�1&�8yHV��Y�"!�E��/"��n�76���+7����B=�t�Ӏt;p���\�r�hc>�X�s� ¥��$�zsǕ�s�7-�@��u���mZ��pD�ܴ;( �C�E�D�s�/̨Y�L���?�/ON���&OM��I>�N��f)Ɇ9��8o�ԟD&�<��1��p�P��7!
��˃� Ah<ҥ��uyR�ۛk7�1,O�k"�ua�:rv,�' �*���P��M A�w���+��(^�"<�t�N��d:b���o����L^�Q@��&���U��
F���O�#<I�'^�&k�٠)�B�&�A #��d2���2Ob�\P����I����'ʊ!�O	���	��Fۗzx�����Vh�@3*9w>��N�=8��S�JbӚllO��4�	�<1�#K)<TТ7 �'r�`uزO(1�x��v�-�?I���?���~/�ъ���?���1��	����YoHmJ�ן1S>���CҸa�,:g�H�D�Yh@��8S�#?2�\"+*�k�V�i+��L��i�A�ٱlV�Ha&֮$g@	��͗�-�j�<��V���n�Zz$��1�)[�[J�x�a�i�RV� �IIy"�	%�2E{u	6;P �i������hO�:TYd�G�a;� PS�/$Ξ�yq��՟��ߴ^h���'b.I	d�7M�O@�$�O�EP�7G��@�weVp�p���2[T%�td�O��D�Ot#��YYtp��+EAJ��0�M����ə-C��bD��n7nP��K��HOl���Ď���0c`.*_(q���@N�����L&0�VD�A�G�S�5���s��r��O���N�ܦ��ĝ^��M�"�Z�&�4хMH��?����i�>��+�`F\���CV�Ns��!�J8����4TE�ֻi]c��%���F�>���'�$ ���y�N��OX˧:~ҥ����?�4v	�UɦHs^b(xFi�n�Aa�a��U�(�G�W�}��LpB�������2֘.] 8�����f�쪰�'�z6�I&޸�h�nXo5�E�GgP�o���q���
<�1�k\$!�̙�ƌۿD�$�RB�ǧ$1�6D���?���i�6��O6����u�C>Z�R0&���G�RQs���p��{X���
��tXp���p�D1&�nƛ6�u�֓Or�'R���'f��y%,�k�b֭)R�p U�|��'�N`X� ��   Z   Ĵ���	��Z�RvI�+�� 3��H��R�
O�ظ2�>��j& ��ش�?A��[$���(�E�r�c2��&��s�}m���?	CY���'��6O.���.n_8d1�I�TT��k���A�p�ش)iqO�a��d��Móg�$4�H5Ѷ���=�
��F@yB�@A���#^��$��yލve��=�(�*�E�a2����Ȍ��X���=3��<�A�B=Z�'�+G��� (���p��n3ll{��lV��
��ۼ
���.	X�|�T���I&c��8�DʣWP0{Ŋ�- �� u'�i���K1/Cc�	3i|��c֒|�g� W|�Z\E�zͫ����	$�ɠ<]�Dd�I�(@���Q#����I����q���DJ��O�I�OZ�q`T>��5�B;02R5���>�W�5��➔
C��#/�u2L�?J!&���z�u�����"�O�x�#�] E5N� *N="�`��o\�a5�O����$A7��dD�)KNiұ�%߸���T��	=[��������`dH�i�Ĭ�G�Ëm��Ȑ��dĝ�OH�@��E���l�/��=ha@ĘL,�T�<�f�;�x��O �(��C�rR&�!���#�^6)��((���8�'v���>����sM-MT�逬��\[l�D�Py�0�pi���i���������� ��%�"?�$T�tCJ�s%�$ w��<q�M ���$�@F��#��O�<�'�Q����34Í6~-��H�_�x��?o ���p�_]H��O�#�(�ñ�3D��u�   �R]3dcct���*��C����n�>����?	���d�9T8�(�O�rcմ?�Ei$�[��x�fZ_|"7M�O�˓�?����?�4���<qK������&��R�"|�ūgJk����O�˓gBܐ�\?1��������f�B�Q���'u���//l�aӮO��O|�$[;��|�������:��=sdl<`��M����M�*Otq�5�U�e�	ן8���?U�O�.�J�ā��j^�T�Uc�W���V�'���yR�'�"�'�q���`)��Q���)�>�jtyַii���Jj�|���O��$런D�'�	K�`<�En�ikŚ��:��@8�4N/������O)bO�"�����7{v]���N�6��O��D�O"\A&��U}U���Ii?9@�Є=S�dh#�    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �T   �
  ~    �   �(  �1  �8  �>  BE  �K  �Q  X  s^  �d  �j  <q  ~w  �}  }�  C�   `� u�	����Zv)C�'ll\�0"Ez+�'J�DlӤ�;�5O���'�hA$cŨOo��b.@�`u� p�v.Đ1eʉ%��Hj���%��¯lݱ��.��?����?�YA�)Qf�)��gU"%�E��:2�⁃tC�*N����*�M��ү �u��Ⱥ+����'�6�p�a�+f��i��eX.~�Q�`Йn�J剒��Oz���
u��`�Aަ�*�$�ݟ��͟p�����Q��S2 �\�#�Kľd[��	��M��f�����O��⟀���O,����3Bv4@�B��r..X{�/�O��d�O^�d�OD���O�"��i�X�����ѿR�}����9������Z�'=��mګ@��ɱDU�=�ll�D��J��O2�	g�=�xlyV�5��3��@j�"J�N\�%2c
@�O2�'8B�'�"�'�R�'E�SӼV��7�$IriO5�}kNߟ�����M�7�'~�f�'��6�ia�G�ئU�ڴ�?Y�!�`v��c���r|�k�+�hO2d@��	Y�\a���c��Z��]	0#�a��u���j���U�� k&6͊��eq۴�*�����7���bZsտ9����؀.�^m[֣�aèU.na�!��
�%v?x�x���{�X�#�f��M{3�iM 7H�#�����&/��!�g�Y�"���R�_�"^��q����գ�4V$�v�/�b,Y�L������H�;)ϒ����q�J���!G�/q���f,�Ft��`ӫT��M��iɺ7*4��%	E���8��$˛j��ѰՇ����'²8��x;���ΦQ�V����$��R#�2t��ǟ�?A aŲ}J=��.�	%n�����?%D(�Q�#�6Gd�h���6����ɑ�b5���d�$p��S0�C��,��P�t����<1���?��"��� i��t` ��&�<n���PHM�р<����G%!�Q��Y�';R]�S�����Ф!4r��Ďا hZ���(f�f<;W�	�@�r X`�'�����?A�O�h����>���h%˘�f���a��'���'��OQ>}����zni��H�k#p�E:�OZ��I@��*5�L�6�h�A��yC�$9�	$G�"|z�w��]�-�(X	05FE&�1�
�'|vd�����$PCDkD��
�'
d�PA�+�0� 
R�8P�ِ	�'ZM�CF�� %ۻ~Tjh;	�'w��Ӏ�*|�k�f׸v�4� 	�'YpQ�s�6�Q�&�U��,<���@H��Fx���O��Fy�֦�f���5À�:$B�I:	$$�S�N(����h#BB�5L���"V�5�X$����a�lC�ɺ<:}�[n8X &�R=��B�	.P��f̋n2T+��	V��C�:J4�Q2)�1c.���i�+�p�S9rD��I�����˧C��I�g��'�C䉆,�M����>����#]+��B�I�+��T/)Rr� �E1R�B�ɭd��h@�;��!�O�O��C�Ɇ8����g$r�Tkɺ#̎���m{�l�R~���ߒYqD'i|)5O2�?�)O����OX��&T��� ��Ń�uڃL��fF�P�AU�c���Fb�,�"����Q�1��Yu�e��01E�Q5o��-����X�ن!8$�]�'cZ"<.,R'�N�_8�<"�剣o����OV���O�HJ���3s��"�E٨]H�j�H�<�����(�N52�-�J�]t��|��:��'���D �L��I�#L@#z]��� ,��	e2]�5\�unZX�W���'� II��%l��+���~�HTk��'���"6z�KH=`I��Hvn%.@e*�ၣ��S+(��0�&�3C��,QgV�(,�F�̕8w���q�����5_Hx&�rN�Oyx�e�O����1i	�(j,��O�=YS�'Ob��D��=>���B�-�J�*h��\Bt�'���'�l=��H 7hܐlBfC�.s��Í�D�\�O�h���*f��L{E%�Mv�1�$�i�X�(٠{>I���<��Vy��5hqJ����� ��LR$�)}���aY3|12Q����5bL5���	�, ���'�P��� ��u{uf<b�6��rmE&)�(��-f$L�WH�	��O$�
���T?�,Ӎ,^���P�ò3�E�+_ҟ��'d�}�����?9���?١��"`�1牞_ȴ��SC�5�y��&f��9�!	��B�|�Ӄ�X���dY[���D�'L�I� WYбa��V�d{f�A�&�(Uct���M��e8p�1@A�*S���'��776^�f�Dt<	���c�N8�bmC�]e�ғC[7P�Ȇ�`�N(����[W,�$�sXbQS���ӟL���:�٪��Q�E�
e 1Jڳ[����(����V	^�K�VZ���Q�5�$�ަ'�8{��b�<�'��$)#ǖ�<s�b�a�1Y[�taÓ�z-8��=�BI���;@v� ��C ˟(�:��#/�W�V�jP	'�"9c��D����Yja��d��$kaH?-�����R2����0.�J��U��Ԧ:�������ng��o��`X�	�WYx�,�~�`�7�Eß�������ayʟZb���dj��}�&��G��%������ �O�a��B����Da�	m輨��ʒh�<���<���T+_�V��O>�	 fy@�@��ҿ;�J��qJ�a8�V�]9䁞����z�*�$)6��4��NR��O܆����]�`��v6��HUɉ���d�%^�hӍ
H[f����ܣA�zij�&�%���7r���ь'wxY�A��4K#�O1�D�ɳ�MĽi�����O���u.�SB	�Ē8�n��W���	֟��	�XS�5*2�����H��?� 퓙O\�U�s��M�1☜��Py#�i�2^�0K��b��G|bJH�Hq�'ȜsD��&\�H̋�A�Q�18R��y!��b��B	�XN.%�����^��`P�R�\��C��&}�Xݡ���nR�e�)�ģ\6�mj���L����/���C��/$��9S1"7�S�)�	^5H\�I�?���|������j}`��ԥa���ic�M�%�V��ᒄbLW9��=�H��`�'�#=)��iN�V��y�)Xe0bJ�<M$Hc�[��@�
�� ӟ�I͟��I��u�'HR5���&�Һ���kX�f�^1�!�n`�`x���{�eC%j[)fay�'٣����ǘ4,�`U�)��֎d)��R�m��[�����$�*-0�����WJ�X��N�, �ae�'{��'��O\"|�����&8��ſ\��Q	'&o�<�SiB����ہ�I?ve�))�c�t򉀉M[���$�	.< HlP���+0Ѫ�9ՃՁ/ܜ=������?�+O����O�瓠�%aD�D/T):�	!DҀd�Hk��V� �j�X��_�]�e'ڭ���j�I���Y�+?il��f��5'�.=ؐ�'Yd�Q#��a�U�*ۃ?���6�ɼos��$�O&Po���"A�G���aFa��(>�ם�Z��ߟ �?ͧ��'���)R�L��s'���d¢X)�}��VK�S%� �,@��֨g&�9G��6��<bǑ$2`�f�''�	{��'&@̈�c� B�z����2Me�XS��'Y˝�&�K�,fϞT��a�{װy�3	�)���W �5�vM:j�A�6�ثD��� ������G�<պ��)6�<,�A	��.�OD�=@u�У	��8��ډl�d���O੡�'�b�h�T�$!��u>)�s/θ'˘}�׮�tLj�h3-7�$�O\�=a�O��#��U�-~��4.�?�&y(#�	��M��i�1�|��Q�(CĈu`���g�	b��'�@}�c�4�Q���4LI�)>�cpcR�>�̠�.D����Cߴ�~ա�,�7�pʴ?D�Dنm�0p� \y��<eBJEQ�9D����L�b͒49��M�H$�5oq�<uf�e�R�JG]�f��y�b�n�<1�"�._Z��g���L"�.�iy��@��p>�v&�p�TYh�K�����g�<�J��P�<*3��\��ѱ���_�<i�!ڸC ��gg�Aw��T�	]�<��G�ji����/�&,���PO�<D�'<�f��/�$[frHyt�Nx���������2}�<�r�"KHh��H0D����σ�N0d�y�AZ�j���� 3D��+A��m�N�`�a ����6D�\sÕ(����ĥY�s9D�Ʀ3D��X %��E�v���Ĉ^%,a��1D�HP�LB�=�@Tke杤
!���a0�>��D��ő���e��Q&�JHu��y�m� �\���M�*HJdi���y2�ٙ��\
#�!=�(�S��y"` 0��A���ل~5ȹs��y�H�T:Z%�FD3 S\Mʢ'6�y����2�,`r#��c��P�e���?��#�Y������4.��?.�P �.���.�r�<D�|`���:��5Q��2�,��1�-D�L�F�P�3�lM��L��[N�� �*D����U -�d�H5��^�����J#D��5�T�p���Ҁ`˰+���@�!D� ��OF�n�$�"fʎ$�8x��΢<i�eGV8����E�C)���E�KE�$����>D�� ����
j�
!AB	+��{2"O  )�a9{�����:;�yQ0"O��y�?��Q�C-�=���"O�P��c]�7L͸r��(8� H ��'-����'7J��BNבj�pA��.�}1�'\�9����*���{ ��+^G�l��'�����i	�fh!��T1�m��'��L"p�ܥ��#�%��H%�a�'Z�ŧ�/��%CDќD�(��'��	 �Ǆ7KДS댷@�����D �Q?Y��
̈́P����ӥ�1)�6�:D������7K&\�Td�{�q�'�4D�@�� T�j ǌk���
0D��5jQ1O<��5):-�¥#�D;D�t��ˠ
�Np�
�5��)p!-D�P�E��,G@�T�	M�Q�|Ԁ�O�0���)�_?����T�@�T�bwl
�' DX���.�< `B�X�4��';� ��M(M�,�:��ȣ�nU�'ڴ@���(7��ұd�*���'��ؑ	͋|�u�t�v�t"	�'1�*@($�b��d� �,BAyb�U�p>�tH=�AH�=�^Y�ԏ�C�<)c�*Si:��Ћ��-P0���}�<�M�Z)r��d	X��IR��	~�<� 
Z#`�mcS·��\�5�]c�<9�È��*("��aCP�i"N[`x�x�ա���*��9^w�i���G�B�T�e�+D��cD�'j�yq脎Y�t�VN*D����^�h� ,�F�H�.��xP,D�H�暘1x	�v�Q�fn<hU"+D�t�͐|1�� _״\A��(D�x�0A4�����.N�X�L��(ړ_!�1E�$ȗ)�`<Y�Y/�x�`.Z��yP-D=�qH�-S�1�g��y�Eh�:�#�1�L�P����y"`S p`���7 ��q�Z��A�?�yү��� T�ۧu�$%؆.��y�Z�@�2�� �"�!�ҫ�?��+�^����xx�U��^���G��J��-D�d�2)��6}��RB�J[����*D�Z1��)Q�.�J��N��ga��y�Hl��@��Ǉ*��4Cco��y��T��Z�:T��M0��O=�y���&6��r�ٗuкD� /��$����|����/hzћP�nq�p�$�yb"�#F����"�.��Q@���yGE�CNPE��+�@���Ŝ�y�ŽTY�OҘvҼ°[��y"LJ�-��a���'��$���\��>Iwj�o?��J��U��}9�d+r�]��B�\�<�C��#�h��X?BH��0���s�<�R�UY����y����t�f�<1��Z�\��aLU�Fw�}�p�f�<�v��[�H(�6���+ON�e�!�D���l�K^?L��H@�<Oў�*� �Nk}��"�0�,���G�L�Ʉȓ5�8�'�]�2��Z��ȓt�iRꐌA��50%΄9U������(�!��؈�F�s6�׽>N��M���9`�9͔$����tJ6�ȓjT����i��d����N�N|���ɣfx#<E�g
��00���3�V�"u!�D� ��)3dS�F�p� ΍2_�!�� B=+��+V����jG1q�Y:&"O��i�b	5!���t	ɼO1UIU"O�E)�&��o��8:��ɂXtd�"Ov��I�8�Ga� }	Z$W�d� �O��1@�ߕ��y
��;��؛�"Oh�'!D�3�@e�2Ň�p43e"Or�jS��W3p	�$O�^�<`��"O5�&	?	�Д���ȳ~]�q
E"O�m\/�2�[�tp�����'�hDA�'l������4cL��p1AybIZ�'ڔ�S�I�eQX�ˠ/�ug����'w(�ZD=Ir48 
R?t�]K�'��Q�m�+Q㪵(�I]�!N�-	�';$�3��9�̰Θ	E���'�0�֪اnR�)jQM�}��)����x�Q?)���WYL,�QF��7j�&$�g.D�0���V-���R���53��1D�Ĉ�nN 6H�5�Aᖗ#��!�3D�(�3 I4YIH�
�Ĉ�B^p Y��2D�t���j�N9���� <���<D�����Č(��!O$��(Ä�OB��)�'/#��v��@ȣD�,�$�r
�'qth�q`((F�U"#��3 i�i�	�'�X`�� V?&��yX���tt��'δh���[_�����[>@�x�'𤽠f���"���X3ਛ
�' �}�2IC�lj�S�kċYhp:)O�MRB�'�F�!�a��"B	�e�0��x�'Ot@aPjTY`f$��T���`�'�h��1ܼU��&��_RL��'/ <�V�Ĕk@�P�$ [�� S�'"Xz���,�����ěN	5r�1����p�>�Bǝ�e�&	��È$z9
Յȓ���y��(i�P�96 U���i��9���`b܈.�YWh�4oPՇ�J5>��
��������z0��ȓ)&ʜ��#ǖ,�H�]�]�܆�9��l�B�uHE��@ד|[6�D{R��¨�H�R!N�	\�$y6��MM�({�"O�p��~N���eÙg(8��t"O#a*��$����ꁹR�[�0�!� ;X$hRo*��� #��*l7!�� J�X���&VTt�B��`5!��3A�t�R�Ll��!�9R�k�8�O?QV��G�U�&�G�.Ƽ*c��I�<�UE�%l��S�R����]I�<�"G�&q�%�
=N�P��E�<1����/B�@���G;O@�]*'��C�<A�f�x��H�fD7M>��5���<�K�D�T�j��%��S0��yyBD�p>)���_vLE� ��t��<�HY&{�<�Ҁ�Q�\��%[�+�T�<a�U�j�ZոT��8ZK��b�T�<�@��<S>R�˵�^625{%�l�<A����I�QNO�����\|x�lBi��4�4�]ސm�'�?Z�.�(C�&D�,p!΋�`���R�wS P�	8D�\����8��٩t�.R��T�8D�xI����}[���#��B4l�K@C8D������6p�!�'.E��!D�8�����)�2Ę6̇��D�ɣ� ړ}���G�T��48"<�D�̋"6��![�y�95�z�y��L�n�DtKG���y�l\�y��A:Uh݋gu,��6����y
� j�0h́	Z}�n��F��"O2,����Ab������QB"O�Q[�
ס/*���6�۸)���D�'V�����S*p�0H�B�/�J5"�oQ�[��ф�	t�p��,��t�
��$�,y��,���#�	5�|Eۆf�B	��ȓf+J��a]�w(�"/�Y����Ĝ�Q�&ޯ�� ��L?D�`���Q��1!�;Lh�BkN�']65�'��Z�)$2t��Má<�8���c�0FȨ��R��ui&ӫT覵�h�)a��ȓW�J!T)KM'FT��Ό��t��ȓ:��E é\�@��%fȐ��zs��^/>��ŢN�����7l��I3MF��K���R_	$0Ĵ{�#7D����;�<���������5D�,��l"X�P�h�)�p��O9D�㲡߷K4l[�ߍx��9QS6D��Cu�_��!��\�f0�
��!D���a��m����Z�"b)ӵ/ ���E����|�d�2D�fBhx�d �yR'��]F-i�N�.b��l�&�y+��i�t�oY$Ҵ�1�C�y��Gxp|K	ȉp��D:D!�:�y�nÕ#vz���T5��8��'Ş�y"��2se�)���E�(ڰ�@����?ɠIFM��������G�[ȪuՅ��s�|�&�)D�`b�%��S�.yz�ę�)Fv��w&D���Nd4�Blͭ3����ҁ"D�����>M�!�Ԣ����k!!D��ѐ��t���e���~КW);D��ѓ�W&��%�"\�_&^8��7��$>�Y������a�B��BH�r�xd�rg��˓�?����?�>g�� �X9,8|xh��B�}�N���_�N�R����6.�	�$�G	\'$EyB'�yϊ%�u�Ԥe~��W��m'������(t��M)}F���֥1`�`�Dy"k�?q��O��Ls�
[�0�И� ΁�S�d��(O��$"�O@]Y&��_�b 6�>���'�ʓO�"-G&J��$ؗ��Z�dI�'v`����'?RP���O/B�'�pɛd��uT����ϋ�*��;��'V�q��C֤o�p��D��C2��#�edEZ��4�̓e7�Ih E�v|�1��K��yr�2�D�!\�:Զ�AōT7&�x�Haܧ6NE�%��&m�T��;o��Γ[����������'����i�R��V�U�,�9�+L�!�ItL�q�đ
}φ}��o�,tў,Z���Ρ[{D��E@��x� <�C�>�����O:��q6Pl�OV�D�O��d_�����]��Q����0�c�h�7N֖�e ��M	�EĬ2���k�)����?ᨥ@�	Аin، u�;m�M,3� Mॡ e�����b7Fx"g:wxn���Y�w���Ŝ���������F{�:O�QB� �o ��j��3�@c"Oh��!˝k���[�/Q�L�̝:`�'�L#=�'�?y-O���3�C	�0��2K�-V}� �M4	{��c��^�QL@���O��$�����O��S�>p)���� �j&&U�8���qS���e�P�	3D�7ְ=�D�V��4�6��|��Y �%�'q���hD�_3Fź���E?���ቢ[0.�d��j���N=8r��Ŋ���,�$0ړÈO�� ���y-��#t�O-pH�+�"OB�# MT>�����MW�080R�x�۴�?q.O:��D��ܦ́�(
��p�'h���B�څ|F�d J,G!���	+Y���ݟD��@�p��q��O?�`�&�wO��'8��+�@
f��$�u�Z:yx�E|�U��ș�j�	>�V�#5��{��"��Hy�"#N�	~�
$�W�'^\�	�l�|rqi9Qέ#e	"'g hJ�CKy��'���2�'\�h&RUC��B	����=��I��B���_� �a�O�X^� �@������H�5��ꙡN" 9���ȇȓc|���
I;��� ׍�6Cn��ȓz����M�$��)H�nЈ�����S�? r��G�8c�q1�aO�6�5H3"O�Q�����5:�W�,��m��"OZd��-��~����� 7@=�dJ��O��}�@׼̘`�C�X�$E)V�^�~̅ȓS�dL���*u����A[sh�� *�QB���&�
ő�N�$Y���dٌ�CVɗ�\5�𡑮��c�"=�ȓq,ja
�g�i�,s@^�1 "�ȓNE��Vm�>40g����"��	 *���dE�ED���e��h�������z�!�$7b�xq�V�ۜ>˚��c4@!�$D�,�����W�n�(xҵO�g4!�P?�t�����!�N�����k!���w�����'٢$�z\��O֯(�џ�A��Mˌ�d�������n�H��չ�W��O�(�u�өe�lj�p&��r��&�4">G��L�OA�ɒ0L����#3$7w��K���5Y����2Ȑ���4UХ�v��
c�C�	�:HI{�u�h]x���_��� wyҎДT���B$�#/r��`"]0��$�O��D#��?A�'������?b�`4��Kہy��1�Ó�hOv��D��?3atd�G Kcպ}���Z7/�'걟������ѱ���ME#������'ˈE�J���<iW��6� `S�!P�P���[FJ��e��T��O���Oxq�p�>9��tf���|�U� -WS%�5ȒLc&��O�x��h��.R"䠀��v�Tq�#��4E�(�*�>�f�>����M��Zm�d��'Ř�E&�!P
X��.�?Y"��S��]��?=��[�IE�y�ǡ��sE��I�/F�H�TD&}J"}�-^���M+�HP�-d�}�EN�G�ТIdyR�W����3�ȟ*%��WI���j���_��4��I?�tĕ\�T>�I.Y|�<��q��*Y��Х��-FcT���!}���1��D��H��uR���	*� +bh��H�KD�'��0�@bm��9O�ڇ�O��c��$�)�&�%�T�C�'�0T��� H���B��H�Xy���%2ظB�I"� �!��X�W`�i�bȝ�}�6-�OؓO(���D�|n:z���闌ȗܦ����Y�:��hO��<q�i��n�VX��_��As�{�	~���O���Ӂ�30�	�UΏg)FIh�'�x�2� D�D���ʓO���A�'���[��b����]����!��}�<�çηZܔ�`*\_�~t�e�{�<!@c�>,�AC��UG� k&N�w�<Y@nڍ>�\��e.ËG��rR�Cq�<�lB�ڤ������SDn�<��JS�@uJd��k��n���#Sn�_�<i�Ț Wl��e�=I2|��l�Y�<	f�R{>�R�\
[�s�Q|�'�l�S�'UE:$:�VOܕk@M�*#$����>�����:D����()J��>9
ʄ��)��*�Y�,���4���q����ڨ�3l��=���x靂~�z)�4#��3�I:cJH���y��-�9wGj�ڰj��	�ld��Bˊɓ�%���V  �)�e��q�c&�z�"h�� Z�����
6r*E����Y�|�o��W�tс�`]L����e��Ԧ-�s���ܸ��/�$i�� ����?������e�*g��	� b!�.6]>��Oꬠk!��=6�rIXR��*`��N<	���	8��!�o��FC�܋T�S� �!H�L
i�(]zt��4w�RO�]���'�R�զE"�$O P���ݰ@%�UQC'T��x�"M��HG`��&%��V��p<���'^S&D��OW7�6�@2�Y׸��%�i���'R�O$�����'L��'���<��0�
�4+BЅ ^�3�����&��'�j�a�ߦ�2W�!.yb>O�{RU 9���;�$H1]�Dj��J�5�@�F�@1��N^�Db?O�ɔ�^���*��F�m�8 zW�Zȟ��'��q��|"����'g�p���n��Q�TgUp��'Ir9�1d�?Dv�!b��R_` J�T���4�*�$�>��@f����M��O�6���jT��h�H^��' B�'�ם����	�|z ��r���$%���qj*q��x����:	�S��S�/�T9��\A� f������&�L��1A�.L�	�5/H#=d:�XQ익-}�M��'}�4s!�I�2���gF����4���Z��?	���?�"��^����R�_�FFdx�b#S�!�$�1}z�4��숕w�d�+�T1qO:�oџ|�'��-��'O�ihJ���T_�5���
�23�f�Oj�DJˀ���O��k��@����9�h������Y���)���`3,�q�mP���#�,��Q��+�ja��4��a׮߆�,��i��7P��*�H+� ��󧅫I�d@��$�D��a�۴�M+�� ,ҍr�ގ2O��ĭБb<B�'�'��)�J<Y2C,��,��L��]z�-J(<�u��/yn�e�QE�=z������/_������$UF�xQoZ���	i�䩊�_����<=1��_�0���"ȭi����O ň6��O�b��gy�ع2���0dm��U:օ!FP�ē
Ĭ<Fx��4�?B��x�g͆z+��T�����Vt�Ir�S��:m�­�JMԹCb���o��Շ�������A+괣`fߎC�@��I��(O�P���_q�� `7��b)<��c�O0���I;�i�P�׽��4���]��!�$*
,CCb�όT�N�;O!�Ğ�gi8i�RFՏ$O2̀�Õ�u*!�D���`О<Z�1U#Ѻ2!�d_�R�₣�2�i�+�����'D��"@O�>#KT#�i���T�<٠ [֒��6��c��`aGMS�<q$��7��� g�M;�d���J�L�<��B<y���lӳ]����C�E�<�S�#7���SfӲ
���["NX�<���@6#5B�P墝�ͬ8��E�S�<9�IZ�@kv�B �V#9�E���N�<��fu�q�d�#t*Q3�`B�IP:!��UT��Hb��ʹ}dC�	�\��B�B��J��4� I�Pv�B�	��=�,V S��@ t`9R�0C�ɹ�J!��S�]�p��M-��B�	�S�}���ʫ�d�I R�`C��$��aD��z*t�yg�HT�"C�	a����*A�o�(S%��D�B䉥':f��j�
E���*�-����B�I�H�65��	�Y���cKJ�KEvB�*a�T�7�G)9D~��*S�`B�I�:�@�ꔪՐ`^r�i��O�5�6B�%x��AS���9$��q$A8�dB䉟tmԕ�(P�86:�&i˫F��C��0hV4q F�ӓ"3"���^�C��C�I&��
�T;NB���j@^��C䉨�DŨS*Xl�"
�'�f��C�%X��a�MȰB���%J��C�I6���k 	Q�����N�C�I/[�ܩ	�Ņ�5�Ja�$A k�rC�I�)@ەl�r� 	*���Y#~B�I0b:(Bt�JhB�� ���ovB��-ik�)k��ڬG��`pƆ߹4lHB�	�_�z�a�F�T��Kb��i�LC�	=W�h�a�C�G�KH�^�L V"O� ����@��b�,���� �"O��#��K�"��q靈�nT
t"O\+��6t���%y\T,{2"O*p�N�5It��`,G[�d�"O>�	2�K$$�2ab��z��j�"O6�"��عew�]K�/@6M6	3�"O�H%gJ����P�V/d��"O���(
3C1�L�A@��4c"Ol�g�Uՠ<�  ԎB���"O��G��-	��I�$��/�Q�*Oi*A!0Y���r �Ƿ>vD`��� �}�EΆ�c4p��/B�e ���&"O(0�b�R�-����S�?T�9�4"O���g�i�u9�ƙ�u9�8��"O�e!�h��k!�i���>��첃"O|A�eė�g��̢RřM�	�C"O­Kq��>��]�&Í �n�H�"O�y
���S|��I6b��,*s"Oĸ���4�@|!� �<����"O���䁙�J�½�`�1���$"Ot��kR�EL\i�Q%6m4q��"O}�Qk�g���r���w����"O�i�����\9!뙼-�!���0�����݁l��k��z:!��Л0tع󆋠��Y ���4�!��Yղy����H�a��3J��D F�U��σ/k!�A�`E�y�X�W=�p��J'q<p�U��y"^����ɡ@�����ϔ �y�+#F��S
�6��Zw����yg�_:vPK0J/`�XY��]�yr�֨q�0'��#�>{�ȋ��yB���T(��r���M�\��N���y��ɏOǤ��#.�����y�$N�`���dM�4�TI�-�y�i
�'
���À{�"����:�yh]�@� �7F܊@.8�T	!�yr��3����A���?�H��Ҫ�y���J�{��9�����;�y���A��҄@E�Du�]�%�8�y" ��&� x�*L�9�q�J���y��VxQ��H�"�D������y�l�=P�4z��(81��	%���yR��#R�L��b�M�.���%E��y�DӔ�` S�ՁY�)X�� �y�)H�{��s%�B�R��4��=�y�T�[�P
,MBHթ�(٠�yǒ=����f(1������T%�yb��.��Y�GG7�nI��y"��
*�J���AT�M�F��y����n]K0m<.�TH����y2��4t�ڀ�XR��R��y"�	o��=x'*��PI@�RR���yT�`�&l0���I5�U)�'�+�y�l�'j4&�0D��k<HyjDD��y�E(�8 Ѥcם^N�%त���y���k�b ��Y�W���p���yB���rIIbn�9[\����yb.���c��L�\P�*��y���zrpP@r��9S���(�X��y�m·k�p���Ô~��y�2H]��yң#]HL�����7p3v�Q���y�D�	-��S4e�4p�E�0�yBΕ7+�T@��JzZ�ճ���y�@�0銸�PeөxG����(��y���9J(Lqz��+R��yt���yr�+]�l�a��+V��)C�<�y"���.�*�C_��B�ۂ��y��4;_�<�C�A�ZN���S�y�NQ>�� fɘ�bxTe˚�y"A� ��0� �\h����	�y�T�J����r��X��͓ulH'�y�g� ��I��L�<Ke��ĩ��y2KJ������>k�y`�	��y∓�2:�"`V�c�00�b	�y
� �h���?m�̘ҷٍ�8�kF"O���6iR��Ѐ��b�2}�"O��;��3K`�P̖S�25�0"O��c�o�.yX����(0ӄ���"O)1�Ӯ�l���	�)v�P�"O��Rg�M�opj�g��4�$�F"O�Гb��8��e�sPI� ((�"O�puѡ.W"M�"d>\�IW"O�E���[G�h�'�S%9;N!�q"O� ��*�}�����@5�xt"OL�X��]�]X^y��g|ʨ�5"OH��Ř~��Q䌽0��h �"OIJ��@w_�h��I5K��݊�"OnXy��}&xt��@��9%"Oh�)4���kz6�{Q�ܚo�81"O�i�f&V�V�*Ոa��%ӐU`�"Oh�����,����G�%�&t"O�B��B�râ(���7R
b���"OB��Rh�a�a��F��+RdJ�"O"Agf�9g�� �Ơ-F�,�4"OH��c!Θ8&x����\:K�-�@"O�pi�E�X֚����=AnuY�"O:E�&��
ܨ�R���B��p��"O�2��G4n�ڜxpeN5 &,Q�"O�a:��%w�8�CK!&�~��"Oԛ��x~ɣS���I�-"O��[�'C�j� A����7Y�-0�!�݌+v�r���F�j$��y�!��t@H�h_5��@�uQ<o�!��_C@h ��ˏ&Xt�g��|�!�$T丩R�j�,nР+��%O!�dT�ax��Pԥ2Bt.M22#F�Qp!�d�{�Ii��ťX:H2q��0t�!�D�.��e�SI�>Z/�#1�Q�[�!�H:8��I7(,,���Uq�!�$G	?F�	a���A>�����!�d��.f��r�nM'4d�ə&Cr!�dӜ/��욁��B2���A�w!�$�	j�>؈��ę���E ãnS!�$Ƴz�f��E�N-	Ui���hB!�Q������P���&,�5M�!��f��kS`�9:l-!f�Q7/S!��ɱwO����Fdoʵ��If'!���gQ���决i���:�W)7�!��>A֣X�\٬!�/؟`�!�d��� ����Ie�0��-d�!�$֪S�^l8�l��TN8X�ꅺh�!�C�TF�3��x:Ag>/�!��K�,�0��)�� L0�0F�"h!�D9y&�0ǈ�o�T�Y�E* *!�R$$�(Ƞu������2E�<F/!�D��G� d
 ��K6��k���!y!�$ʂbWx�Q�"� �f�yeʴY!�D��dH��D�G*L���I�Ȑ�!�$��m�r-��pS$eQS�(w!��M'wA�)���:{;Ji���!��[�'&�Xeꍟ'И�C��V�!�$���(�B#A���2�R5
�!�D�/W$*��F��:���i��G�V�!��Щ��p���l�L��v$W�}�!�DC�"��bf`<pH!�0�
�@0!�d�5a%41�Z6���g��
�!�d�
C�6����☁�p�Хf�!� !)�j���y��u���@Q�!�� ؄�p�H�"��X�rB�AYtuAU"Ol�`�x�됡^g��h��"O�1(�@˥}���bE`9��Z�"O��k�$�;4��+G(��e� :�"O��j�#��!��] 	Ӫ(��"OV�����5fI���dҦ"O��{��ε	n0��^��["O ��1���T�
�Q#K:h]"[t"Oژ3���
%}x��&tF��h�"O��/̇h���CcնA+�;'"O�h���' QiӔ���!Z���"OLL�uY�W�ԁ.&Vs����"OȨY�jލB����/�DfT���"O���+��s�� �mN)K]lY�1"O���DL�8=����4!�N0��"Oj ��.K�TP����<�4�B`"O ���[�?�X���N�>�<�b�"O�;3K�%a�� .��%��͑�"O��c 
(t��/Y%P�
,R�"OН���T�*�#���6��e�"O
PC�LY2l����N{�ABq"O���*ߎ�BM�5�C-(nD`1�B,�r�i�)ܤ|�ԃ�B,<O@��Rd�8,<���Ҧ��Y[5"Ol=�Vn��0��|��g�E�L}��"O|��/�����/R��^��"O��1/+v*� �P�W��|B�"O�H����	6 �"�N��B"O^�M��7­�%-:�� j�"Ox��@�53��#�ݒ6�n[�"O���n�?0�����Bc�	[v"O:(#�#D�U��L8&ʟ:Ak�X�7"O>���Ƞ<YZ�[�
�eH �t"OƘ�"�>L
4
��V|� v"O���7C������$D�q��"O�!���X7G�3Ǎ�\����"O���7��4��q�ƒ�����*O:�a _�>��\y#aѣP�*	�'��h$,ڢ*ȱ R	Q8<r�A	�'�\�q0i��Q h Ұ?����'�R�(V�B��`Jfe@�]��'��{��O�O2�XX�͐S���r�'��I�0�J*7�� ��>�`��
�'U���@������ 2$t���'�8 "��y���WR���'J�ԁUn֢c�vA�Rl�%.�M��'�2�h��J�$<�C�6(W(D��'�����iy�@"R�ܟZ�z]*�'Ϥ@���$a�>D��j��Q䌉�	�'ĀX�Ӌń�\sCEG�[�\�	�'Sf��p�,:��bT�Ν<�J��	�' L`�$%V�p��M�%���x	�'�=Y�@�3"�s�">��	�'S�|�2�Z�7�|��RMƭ.f�]��'��Q��+C� ���P%G�%�X���'0\�"��)Xd^���U3 ����'�
#����4���D-Rh��z�'VD��OBL����L�At���'/��y���j��%�� �.�����'�p�a�L	L&T�O��1�]�	�'�^UӁ�������"�*t���'K��C��
�s�.�S�/4Ӛ���'(�y$�C�?Q�(��,�5*����	�'D��;�!b���#UfPA�\1�'8�{ś�5R �S4뒒{3���� �Q�N��*���3� ~� -j#"ON��oU�(�6����	qD��@"O"�(�O�4���z�EKe�\��"OʔYb�L�j
^h�ꙴpM�m�"OL��1�G2R����ӥ���"Olh�V�g�6-D�ĬE"q�"O&/>Ԉ�Mȝo��y1 �/n�!�D�".x>�	���� A��
���<�!�D�8/�4�&M�.:Bv��w�ږ^�!��L.����eũf��-�Gʄ7~�!�ӝh���nW��9B����7!�d��q6-h@���;����b�q�!�$�'����R���¯]X�!�dȐE�4T���-b�D)x���<�!�$#��sFg�#T�"�*�e%�!�dNA���IM�L�L��$&@�!�܃#��U����Y��Ū���{�!�D
 ��y��ǃ踀`�_U!�Ӹ-�F��,�|X�H�B	!�N�zg�ɑw"H�m�*� ��w�!�D��
�P9�IP2Ǌ5R�a�/�!�O&ḁq�s���qoN"!�$/SZ����O P7�({s�
�G�!�dP=I�S��K:/����	�!�䙧|�	HT�=&��2�V-v;!��
����B)N�@E4�#�Jܬ6.!�H32v(�
�O�Q�f����.!��8�PL')�7m0����+��m	!�٥~&�!WcE8.,n@��̦_!��I:���E���~�x�ˤ��ai!�-}4�ҥ�U�x�Dh�A"��oZ!�DԺ9�4k�`�J4�EF�	}�!�$Հ.~�� ���(?�� ���o�!� �T�D�-��Ӏ'� yz!��X��0��hF��_|��Z�'��ܨ2�D�#��a�Fɭ�rUq
�'*P�֣�3��\��Q
l�\r�'��e؃�#$t0&��1Z�'���*I�mfb��-I��Jy�'�\�wNY<?�Ĥ
�%� u$�'����礜�3���#0'hjH���''�e���	�`�{#�H���Q�'��)��M;:-���#s|��	�',E��?D��(���,7]	�'`�Y�B��;["v0��9��HA�'����GJ
�x&x�!Åa��c�'�~P�F�5&n5���$6��'�` �-��|^Q0kD�3@��
�'��x ��<$\�F	Z+� �
�'�raC���-+T�Bӎ_ c��@
�'x�(H1EZ�X��u�b���`�J�'��Uʔ�ɻT NdX�	�=�fT��';�0S!b��M������9:����
�''��@�
L��$:/
2�Z X�'&`9Ȥ �1a:��D�(ϢAH�'�~�X��֔gF�AqTLM�%�ʴ;�'��M�wDT���5�t��5xT%��'
����@����5ä�ي�l��'����&�aQ:��jZu�LC�'����c���w��2i�Q*�'%b�/Ś+�p]��v��'�L��3V�b� ���\ ����'��| 
��b5c��°(N���'�FH�Nݖ|Զ��R�N�XU, ���� \�HV\��
��y�f<� "O���_|�Bh��iC�,U��"OL��u'�I	Mi�E�w�XD�e"O��QG�:�X��E�.�V=qA"Ot���Y1TQ	�ր�0�c�"O��6�\5W��y��V02X�4�"OB�`��ڠξ�P��G�l���"O^� E�?*[dy��*����M��"Oji���.���)2jr�zuJF"Oj�YŊ�ue2���
<�4��"O`ps�FT������.��#�"Oni�� ^�.�K���8����e"O�5�ٰ��m�9s��l+ "O�mCjʟ�֨��LQ��2�"�"O"�b���7g�6�C ��/G0<��"O��A����pRB�E(j�A"ON�[bo8T�!�M\�,��"O�`���B���V���3�|���"O�� ��́[|�z��(G�-:b"O��A+ĹD�P�sF׸O� ""O�ؘ�%�Є�f�rGи:�"O*@�E��G����̆?Fv��0"O`����n���ڗ�<L�tx�"O��Jc�S8F����
���"Ox�0lR����d��.$� Iv"O�h�#�0'0f!C��4a����"O����� "��"�'c�V$�1"OB�I���*+b�E��M�@����"O&@@`ŏW���]"I@0��"O�U���	(�ٰrC�<��	a�"O�h���T��Qs��4�Ш�W"Ojx{D�0y<hY����R����"O��	�^J` �efM�o|��PP"O��s��ْ5�a A�+<i{C"OvA
$��*W�x��bċ"&�<��"OX��D(N�Q�j����A	"O�H	cȍ
r(x���֪{� y��"O�Lٗ��� qIR�Y'~�\���"O�,y�T�%.�A9� �(di���"On0�/ϑF�~U��$C-T�4�!"O�u`� I�x8��$��\Ш�5"Of�z�)�.@�PĆQH��A�"O��u�ȳuV�QpDkS �2��%"O�A��-���ғ�ʁ)�(���"OL8�q!��-�8�1	���p+P"O�k����M\X}�r����"O�m�G���{&��#&����2��"O(ɐ&-��+�t��C��܄��@"O:|r�ˊ_h�U��eD.D��\8�"O���i�'z��Acqe�3|��ȁ"On��F��XS|0�p�Y}޾�Y�"O�Xa� �ty�`j� afj�D"O��!��H�WK���F�5QH�k�"O������xM,	A!C�4I��M��"Or���ҳ+�z$�s"��z�~Փ�"O�tpVO�k����CgO��b���"OF=1�)ֻMm�EK��>J����r"O��cGOƥ���s%��8>�g"O��iɋq�tњGDX�NdЊ4"Op<RG�|����3F�A1"O8��A�����ˊ���T�"Oh�9��ߝDlX�БHj��IX3"O��:'��_��DKU��(���"�"OH���K��R��Q��ٲf�@@�"O� :e	u��h���b
��܈"O�la6� !ZXV�@�;V޲�Ʌ"O�ehE*݅R�!�3)���a��"O�M{�ł,X<��(��B�i�C"Opp�C"�]OL���<٤К�"O���1FY�fL�(���&H����"Ox�{�N�n�����u���aR"O옰��K'^߾Dv�?T�ڍr"O�2Ӏ�(lZ�1R5B<>�ґ"O�݀��E6N���l�* ,Z�"O��I�+C���L��!W�i�11A"O�ABw%A�R�@A��G�,mx�4"O��(po��!��pA�F(S�<!�"O$�ڗ(V&%��8� j�V8NL�e"O��s.�kk:��r���HF��Z�"O8��� Hn���'�]D�k�"O\�U�U~�L�G,XUହT"O�h# Ô1cF5����=B�l��"OPl��+ĮW���Q6x�6�)�"O�H*�-�SL����s�(,9"O�L1�bو#�H�ے�R�Q��U�"O����DD'&&���\b�a	�7�Py�L��Dn�;"e�|F�R�}�<��F�$Kt����F���ТRz�<!����a%KƢ�u�D��@�<1Q ��W�АB!ʂf�{G��3E��{�)	T",��e���<ɕO�e�Vu{�II��*T����O�<�V�螵9  U4�X��l�A�<�1�-w.�Q�G/�L��0� T�<��&�PII��Y.ް�b6�v�<	�d��.�&%`pM�)hH�c W�<s�өG��q�i"�
Q�LW�<�W�6P>�!�A�P�D��Ra�S�<�#`�,c4�@�-~o�LSs��P�<Y׊�&uM�I��J|�p �5�]K�<��LK+A{��ӡ�9.z�tOXD�<��bɆ�8)�&�/;X�5Q�LRB�<��C8l���E�
#��<��a��0���c�~�#a]x�<�i3�h�#!�"��ERF�v�<1���,�k�M�4�e� -Rv�<�A����V���3������Ss�<i���:H�-���)0HN@+��
m�<	Qج@���u"N'�R-k��@a�<9eDĈG�vԲ��%A6bt`5��u�<�Q�-Z�0�k��$1 ���PZ�<��I�k��DR`+��$*&Ģ�C�X�<)Ì�K����2�y�.Ͱ��z�<�c'݃z�W�)Ru,�(3�Rp�<sAV'	�X݂&Q&:>%�7��m�<��*\G����@*]�^bd��k@�<Y��:=�P����M"�� /Mx�<��\�z�����C�f僱*t�<� �Ě_P��b�>���3��h�<Q�	��t:*�5��[��Ma�<qƘ�-�������#��@8� Z�<w���\N��pc��=���!%�W�<Yw�*$#l�b�1
�X���Io�<�%]17J*���N�Ŗ$�� i�<y��=2@H�ᄁ3V������J�<鵈D�d;�ʃf�q��1G�a�<�3
��TH�ԥ�Ɖ9pN_V�<��ў1h��!"-W�3a���T�<�f+�7�R�Yt ^2{�pK�M�I�<� Z��be͒A�X=��d�0"O\��)�)n)��
Ai��t�
T"O��x�F�0�ε��M�g܎���"O�]�C� N�̺�ၙ�8I�"O��8ċ�'(�"�Z�4(�hL�v"O�|�S��H"좶�خa8b!��"OH��	^�K�DXQ�-�$�б"O����S�!	|DӔDPe���"OH� Wg��)Bv͊�8X�4"O��Q�@�3WJ��ɔ-.U�LQu"O�q�bF�%�P]�+�7%V��"OZyt�v���I�~p�-r�"O�����]�F3�Г���s`|3D"Ob�8�y�`$��fD�H�zYD"O|�a/�v�/C_� 9�"O̸{�,�B�0ę���P[����"O����@�b�M��ęV�bt�"O� ��H�8	��P0jJ=<�h�y "O�h�f�j���kq���&ضX[�"O�hX檟; �U��G�1%xde��"OD �
)!�0�*%�)Bi��!"OHI��ʍAò��&_�=]P��c"Ov��KΛG\�T�Y��T#��yr�-[����u%�lB�S����y��9��U�aCҖ'�YE��yȅ�\o:�he�=�^��w��	�yRN�АA��"�X�h��:�y��U�e�&͙'��~VV��!�C��y¦��j��DbT*1�0����yB#� s﮼��M�/��p$-��y���'v��h����]@S�Ȉ�y�����h��
ג}��r*H��yB�Sb�p��gH4r�0QC��yb���#��i�RE�F�1P��)�yr@� ��-C3����r11�8�y���[��p�W��$ِ���y�c��s8pR��E'D;"<�l���y�;v��Y0 ��S�V��V�
�y�5����'e�HB�P�'!Q*�yb-(G� p��	AIX��l�*�y�AXL��j�JG�9�0�+e���y2e�0/���1|Z�����yrC]�O/lA�rl�?D$�P�m���y��љ(F��C�o�/:��ɣ1n��y�'F@�"�aӅ�4��{"a��y�⃗*��S(�/;�A��ݱ�y�ő+<�Hs�U�Z�􍺡��	�y"!�%S�-��hM {�~y�q�I��y���$F�̓"-Y=*L��c֌���y&V-Bd�E��`�'�#��_��yB	B\J����mStu�u-�	�yE[��,M#1��{u������yB����Sw挏@�BhBԃ�y����?<,YI�ȏj���fi��y�o�/r4P`r�M24	<H�@��y��s5�` �рY[±{���yB�Y3'��j���5&(��@�H��y��)@{�u�G���NQ��Q��yR�ڷ@�\,��lS��rЩް�y�ٞm���ǮȬ-b�a ���y�E�' e@�K*�$8 
]�yJ�k h�B?�,Z'Fϲ�y��H�Ix"�qG����q(��Y�y�+:���`�}�z��C�y
� ��&.]6�
�cUoJ��65�3"Oԥ�⧖�$�v��A�^�7H��"O��P!�-M�NQ
���tt "Or��cA�'���e�:8~�i��"OKU�H��&C,wgaRr���y2j49�J�`w/շh<�#"�Ҽ�yB@A
R�. ���#]
tY�ś�yҥ	&g8��:�cU:R���bW郎�y���/F�1ɤ]�!8d y��S7�y­̀�q&�[��|
�jM��y�!N�z��1�	j {ԭ���y�hՁ|u��jd-��x�i�ś	�y��8_�x�����b�@BE���y2��0�D��Ks�l���˒��y�kٙ\�("$�n��9����2�y��ևU�Z���l�#Q��FK��y���qў� q�T�1�g[��y��`Ҵ��f���:��l���4�y��^��*a@�#� LK���yr����-"r*�!k�؊���<�yJP9n��Q��l���	��K��x�'j����nƟ~/��A쌞n8Y��'�\�:I���h��n�g�ܰ��'�Z�7�"P
�kZ����Qd<D�h!k^�j��S��,&R�IL:D��r�V�S���Ӆ!�1P��q
8D�D�T�X�,�f����ϵL�E��o4D�P�R(�CX�0 ��J���1�/D�liEJ֖3S�T�QE��
��j�9D�02�2%�2e+GX�=d�$�)D��#������kץ�:�	P�:D�����$�yr��4q�Y8�9D� V@E�HP}��oS���F%D�<���0X%.}Ra�ҳ<�.��Э#D����n�f��CV�E�IIV�r�N"D�Ο]:L z��޺i	b�� �2D�8�bCH�%����)��z`Z3$>D��w ��{l��Rƛ�Lظl �;D�lk"�9s���[U�Z�Z����P&=D�d��B[\@XЋ�@�ֈ�"#;D��C��J)Pjz�c"Q6g v܃4F-D���b�(�2��B�xC�mJ!�D�2*������)�!��\�.B䉋B�,�r�ۏ>l�p�M2PB�I/(�p�h�h��o�+�Ά'��B�	Q��ʲ��`tv�ST�CD��B�I��,�a��%M�<��¯��,G�B�ɶY�Ӥ��*xW���q͉#z�C�	Re��0,�4?ڛ%�K��*M��N�D���Q)!��bu�0cJ��ȓ ����#��;�,��+A�l��Wm���RGz�X(�aQ�m�b܇�5h��h��F��LX�C!oA��ȓw�D�SC��:�T��rdH)�ȓW>�cahV�a�f��C(���P�ȓ6|�;�nH�0�&���V�I�ȓ6$�(��̡e�ĹQÏ*l�����U�`Yd��Z��5	�ѡkLe�ȓ��3��l��r�W�i܆�W����'����h� �?!�D��B��u(!ò>E ���f������O�Ep@"/9x��Rb'��Q�l��ȓ� Eyd�W�4?iʄ��!�f���,P����8.mf�XQ��;?%��S�? 8���X�z�.ѓ�!�:O��[b"O`�K�%��+�z�86&˒o+bE b"O������* �.����tȉ"O\Ec�^X�ҩK��D�r�@��"O �Rp��#|	\�g� .Eq�y� "O�;n�7r܎�����"b���"O(�J1xv�C�ʅr���"O�\c��]#��({��G$5Դg"O\��v���WՄ0��O�Iz91�"O��1���'~��U[t�%��<�"Od0��e�
^PE�W��򂤹R"ORd3W	S�<M�̣�m�W�f�"�"Onu[��(x�d�m�:[���p"OڐQ�ν}Ȁ\�T�B� KW"OlȐD��7=��Bd�� ���Rd"O���⩑����!�#��Bt��"O���(�'G��]Id�-+N�""O����+Du:az�+�F���"O^���i�!3Ȝ *O�4�"O��p�F�wNn���k]�B��u��"O�+�ˣKYn��a���v"O���.�:Fo������,5wD�'"O����*�r�V]2��.�yҩ�OP �DH/������y�K�qFM{4�D#����� R<�y&�{�z��e �e���*A!�y2�(~��p�&K�U��A�yBJw���"4HA�
l�M�C�[��yB�!5L� 	"�@ᅀ�y�b�Hv�y&C�Sj�Bn@��yb�:))d�e�ڰxzQ���ʏ�y��&� �R�]>N�U*6���y� �&6�,1c�i�]��3ԧ^+�yR�^�Qh
؁6��^������P��y���C�\�c�9Xڱ�����y2bO#K�|��aN�23��-�*��yR���o��iQ��ðf����L�y��3%����/k�Z�ۧƮ�y�+��v��s��M�z�&�N�y2������\,	����!b���y�(F���I�2�+p)�C&D�2	�'�ՉT��3yn�A��C6C�Q��'������,o�܃�J	=5�v���'����ą	LН+F�.Ѭ�z�'�
U"�M�����;�(P{�'_��
�|̲t��Ȗ5CRQ(�'W��/�CTU+�H[�0�����'�	���2��˄���$�mi�'���12	˂f��PS.��|;
�'��AgB@6�e���R� +�'��e�AE�3W���R��}��ܻ	�'�29�VKO�o.02"��|��A��'SV���h }Kv9Qh7JE�=k�'�m�è�1k,>�cAǁ<=�x�'�&���ܒ(��݂0C�*:T\L9�'�,ZqeP� ��T8p�ͫe���a�'���i�ղr�l�vfٕP�z��'�NtH�C�#2�H����Iq�H�
�'�H�U�K��(1JVW;G��1
�'�j��b��L��U�E>>#p2
�' �8�����ո���+़�'I)Aq(ڷe��-z�)�#V�`�	�' ��2�	 *���F�/��		�'�@���eV1(��	�'�u�`���� �q����.c�Ƚ���(L�p"O�e1��'xL���D=N01"O") ���O2<��#/҆� "O�����*�(�a��͚]T��C&"O&p��Wwx����;@04"Of�9�!�8�Ⱥ�gJ
Lq�"O��ҳ��c7d	�"F�2��H(�"O�9:�JÇ8�j��֥
�S���
p"O`��"�DyJF�	���je"O.qJ"��p�h}�@�WNڌ���"O>9�OT�?�2zQj�(ؐ]K'"O6��g��P���8�)ߙ,��p�"O@\���B�n(�| VN�/��56"OV�1�dɜ�HPJ1o^�,�	z$"O��)�*�s`�a�Ô� ;vݙs"O��J�)��ܥZ��	�]$6�w"O�L�7C�N��yp3��k���X�"Oh]˵�/xeZ�����	M�L�Q'"O� Е�� 2U2�z7��)w��Q"OT�jW�t��蛐n�UN���&"O>lF���h1���b�O�\�fx��"Ohl�5�@�pu
٫NM�J�v���"O�!֮E�J�n���,B(H&��b0"O΁�@���tӕ래'�#1"Ov0���ߴ-��{��T9%�Di�"Ov ���'K�!��_)Z�@�e"O�§�V�/
Nȡ��W."��H�"O���#f�)�p�-�S�,�"OH\�0��q�� �ȣRt"�q�"O����� "����eUN9��"O������~�̍3�,�>��P��"OPh�U�U5M�L<���S����"O�}��R�BV�s�j]���Qu"O�]�@.ZW��{ CU��%��"Ovx�mW��ƥ����N�*\��"O �z3Ν5:r�0�P���j��!�"O昪�!�4P��#-��ޝ"�"O�)�4�D��!���zs"O�Hp���Щ����lcU"O���SK!�����Y;�� ʷ"O��pUŏ�\嬁�V�
�K���E"O6�8�}׶<�
�Z�\Ʌ�=�v� ��_���rg��7���z��p���ql��ȝ�)ϔq

�'`�L�痔T�Pl����"(K��
�'>���i�\�Ui��wX ���'�B��u�1���%��p�����'6��ran��f�Nt��� m��{�'��|B�nY�%�8AY�
�x?��0�'�d�Ċ��%Q,t��m�k��h��'͞r%`�7V<�l`b��"I:�'��=�7O94R��8�_����'����k�E�z$ʶ�� w,f1��'0�9B1_�@ $��,Y/]O�=b�'�@q���0Q_nQ�W��RԀ��'e�q�fH�.�ha�艣NҤ�
�'�q���R�D�aF� �Ig6}�	�'�Lz!���n�δQw�TA��U�	�'9�BB	�X"TD�,4=B���'o:pJ�J�~'~p�b'

p\�'����NO
hŮmh��Rb���'�Vqp��!p��m(��V���'�tչb�*Y�H���L)w���'Rq��!X%��;Q�Ҝh`����� �����K&6�3]�R�2��"O����h��)z�q#Pk�>+ ���"O$mzu�]�K4-��I�2`X�"O��� +�	�-zt�U6.f��;�"O8�۲�qj@���E!
y�A9"Oh�؀��6d�Eё���{Z�ts"O�Q�.�)���w.Q~evU�"OR��a���8�bqjgO�'.^��#"O�`��(�N�|ء���	X|��"O��cj£��\�f���iRΙ�7"O�A���E�nM{���dQ�!;5"O<aSk�*T����㎿=�v"O���Rg��UGW�O�PL���l�<�!):w����O���\PDk�<	��C.oRu��&ͥ\��A�a"j�<9����_���bkּ$�{d(�e�<�Ecú}�Ҥ���N=Y5D��`�K�<!U��:B��L`"i��=�2��ep�<y��jK��V��<dN�k�<�SK̪.2U����$ �l� rϖ\�<!f�I;f!`�:���: ���"V~�<�C�;H*p b�}9�|@��^�<ubP�[Խ@��@aRE��^�<9�~� ���r4�`Pw�s]!��=9��P����,�H�8Vǀ�<G!���O��Y��J�T����6��%[�!򤄢,���KD���Y� ����-5f!�Z7��TRa�R �b5*C�_#>F!�D^,��9�A-�q�� G&Ч!�dA#=0���-�*���ҍ!�䑫uP�SeA7x��A ��B�8�!�$�4Y�L�*��%~���W�qY!�D�(P���{g*�=�~��E/� e�!��(��sF�V=v�.�G�x�!��F��Ae�
4^yr�c�2d!�ܤb�~a�AǇ	��Q�#dמ9I!��2qy>�cBG9_����!"!��D� �TԨq�ڄoST�I1o[?!���>	$b�.1AH��P���Q�D���D,���@H�U���`bm.�!��� ��	+�䔆�Z)p��ڝ c�	Y��H�*�K��I"YO>u����; ���s"OT]�0��D#PYӧ�<�։y2�>AA�'����A��*p�\�Y��'�h(C��>$�r������j/�|2�'�ʆ*��%xƀ#�[
k^:@��'n\�(@ U,3�u�ˆG���'<ִ��j�o4�dR��ޫ1�(8�'��X	�F�/_�񙵇�5x!�|��'y��3W�ȝ����e�2f/�1J�'Htг��$s�P�	�F�X����'�8lb��&ъH�g�$O7���'�0�t��²`�w s�Ÿ�'�<���%�(��GG��A�3�'{z���jH�f`I#V����6�'D �s����E�y�Zd��'W�4�1��!�=���$�c�"�c�<	��N�S�M�3m%cX�,C��Sa�<�����,�4x���*L�|����_F�<p-�JG�Б��''8��v�@�<y���|xf甚j4�ɐEB�}�<I5/�#R{�0r��#�N�C�w�<�v��# ti�%LL�*S
����s�<�C�n��R���W�n���r�<� �(Т� �G�� hI4�@���"OL��&��7R�Z;_�YI "O<p �G�iL�K��|�(�P"O���g��}0��`&��_y�92"O�T��݇}w801Q=Ds�e�!"O�I�a��}���bD�D�;�x��"OT�%�o>�x�"��r�@�P�"O�0ce�
�H��%�DlP>�޼S�"O�Ғ�ӚT�P����9�re"OL`Bi�&E���IU��/xYD�K�"Ovtˢ͖�G&��
W措P����"O�$�gR����@f�0Ie2i��"O|@�r�׻SpA�0Ñ���x�"O�	 ��vr���$'��5#�"O�Y�eƛ:$�x�eO���"O�{� {�2���NU.J�A$"O:X�1M�
��0��_xa#"O�0�
S2.�j����]F�4a�"O^ʂG�'�p���j�EYQ�"O�U�E��~�%C����y��Z�$���v���EJ��yreP/$� ��I��")�Ժ�d��yBmE$*��ʒ(�����Ϯ�yRJM�8U�%����5���iG��yL��}�(em\<'2|A�j� �yC�	T08Qs�U����X��S�yB!��oB�U)�+�%'b�,
4�V�y��T��,\�BȑQdx D���yrOˏ�\�D��/+��X \��yҭ#&�^����1!tPoּ�y�̌mO��3�"����h��D��y��]'��H����\��b���y�� ��99��Y�N��r'�3�y��gOb$�F�̶z^θ)s"�6��ޔ��LoX}��9O(h3����$h��'�A�(�*� ���z�,H;jz�@M�eP��������L?nbD@�!�.cHh�h�g��Ms�
B?T`H�f͖,���t�Ԅ~�� ��,�s�x�LN�^�<��+�5����uӚ��b�'���<��o�D�~nZ7{�u� �I~pH#F��fbt3��?�L>q����=�^�0u�\ _/��@���.Q���۴�?���:���R>�m7���"AZ�p8|A��$^�X"P�*O�0�!
VЦ9��I!'��Y�@��9"7H��
S�Y���S�-�(:��z�%Ȣo�ԥ�iA���`#�rI��;�Q�h;N�{���7@
}B�Ѻ���s;.A�g�L<��i[\^�-zJ>� (�pTry���̢gu�t��+}}��Ӭ�?Y��_؉':��'���v>�����L���r�T� ���h����O��ل�Jm�z��c��z�<��l�&�Mk�����|"���䝐9��L�䣆���H��h����#`Ga>b��D�O���p'Kqm�ԉ�-��g�Dl�b�@�O?��Ar���X�� ҥ�H-��Ȉ���	avx�&޳P���hua��b��E�TAG�#���,j���5�яMw�$���
�X��i� ��ǎ.���"�C�Xw|�q� �O���<Q�����4LvD0���C:�Qj�	5���hO����%A�k�IP�"Z�y�V9���OP�o����'H����j|Ӹ�d8�II1x��j��ƇVƘS iDE�qO���C2|:@�#�H��^S>��C�xW蔻�O��
,J�_h!�T��(=i��$ �m�H90'����C�ؕ$Z�[k]yDdx��#��i�mM���1��PC�R�'��OG��h�Wƌ��0A�'d�3.����-�)�����%#"���4����A �q�'����}J6�i¿iK�h`�@R�#"Ҡ�I�Y���*�'��l2��qӔ�D�<�OL�'ق��AـU�0�*�l�8`ٖؤ?~^X�靵�&�Y�]�P�����Ͽ��I?p8�V�ފy3N����殮�����N��eJbiBԦ(iLS~$̳D���Hm�aj8:��`"A�y-rh���i0HmJ��?�B_���<��5:�Kń<;nI�qa@�)�\#��@#�?	����D�O��'���5H@�lv��A�>~DT������I��,�ߴ��}�:1֠�G' p��ك5ז���Smy2b�l	�6�8,Oڈj!J	�k�������0�����i��!�|PXW�ŕZ ؘ"�
�^�ڌ�SB��� LU��� L�Y�"��,X(�kv��k��	�`X�e'*Ȉу�$S��S�1Î�Z�|�"@�)�P��
HSp�H�j�G)�$�x���O*(z���͟4�'��*��U�_�6D0�[UD�($��<���?	�S��R"ذ��Bŀ\>_�:P �N�8%|`oڜ�MO>�'��L>��4GpM � @�?   N   Ĵ���	��Z�JvI�*�� 3��H��R�
O�ظ2�>��j& ���OP�se��c�T|h�L���$�6���ْش�/�Oe�'������͓oO�:�W8K8��s-��]�ڠ���N�P��6��{�/�#<���g��A�Ƽ/�"$�!�π(��-5_�H��gP�=E@�#�`�<qdi��gߒ A�F}R��z
��C�X0`�����`��G����%���u��Ӿ�yB�X��4�S�`�l�I^�"ɣ���xӊ-8��&X�j���<&��NY��~��αN���� V|~�3	� m�w!@�˧�YJ���[�K�-�!z���A�I��tJҝ|�c�9���.��!�
1Æ���yb#t�'�l8Dxr��r����� dK�� n�1m��#<���)�8J���Ċ�ab�x�YV[	�O:�	��G'ȸ' �۲.J�q����3ț=}�\�ݴ[("<y�4w�ܑ�3�1P�����zi�ة� 
f�KvT#<�d)1?�g��k�6h"�"~�~	�C�DbyR�L�'��l�?���֒c�IF�ԞU�)݈g�"<���"��`���*��P��,8Z6%���ө�1O�$P����<orѪq�L7�49waAu���,g�#<Q�3�D��%�b}�����t m�>�W�
�Hھc��!U��H���"v&v����Y��x̰�������%!CN	������	6?��`S�O>R�n�!F�,�L�]}"<��K0�n���I��x��]�򠗬�\@��TS~	  @�?8���5�͕
��lARC$�x�U�<���	�O�``гm�2�f%Q#�"�[.9bN�zrF�
*���{Ȝ�"V�"�B�Pj��
�'��|���T8kɔ���2��=����5\����?p�ê�":��`�@ U;nΞ��O�N�E��m�f.�*pC�f�9e�a��&��}i��RCN����pԸ�pNB�2�&�8�Ũ,�8(G��F�&�ɈA@���O �bL��:���H����/ ܽ�B�?�A�hz`NY�$�*p!�N�`�dh���?��<�R@B�lJ���<\�<�ci�O")D�''>2���S�? �ș!IӾwt�͂��XB��ۦ^���S/�*ɖ�PF_6tk�Ę��_�9�hY�r蟛���8=�d�j�%[�D��D�F�8�ΓcH<�c
����D%�~
zQ���=����)� �S��%4)d�]?9��G�6� ��Im��]�n98��6(WX��Ys�r�����3D��Ͱ��ܰ)�p�C��ݤX�����I� f�-�k׹|�Q�����Z���00��Ot��,W�X��'�62�ˊ�r�H15`�:+딜���$��`���K��R�6M�R��qH��țA;@� �c��`פ_�t���IģTϟ�0Љ�sG�}h��'�^�H�IE�d	���H�7��y�'(�9Po�<A����+r+R���b]��L�C��O��b7D?E�5[�Ⴠ��9��S6I�#��s<��_J�)��@�A�24���"sz�݈��!:Ĭ��^8�G�O�$y�� �D�*�@����������0�,�?�Tl����f~"�'�p�S�A�G\J���"طF�ڝ;� _�15؜ 4%�.(-�q�i]�s� #C��BVZ���bضE�εk�����D��7հu �+�BO����MYlQ�,j͛�s����+zܚM�� 4��Jul��a�&\k%J3�Lx�E�,W�x�(�,B�4W�� �Z��=ͧW%��˒B��~�����I!��'P��>6,�I
�����UQ�U:�N�٥�MK%�ؿDږpX��V�4�`D�u�Q) �D�{�-I�hO?m�`C_'����)i ��ehf�h;BkE�S�<�#`⌣�����0"�D0y�8*�Z!��̼+sf�,?޼K�D�>9����v~��'#H$0��C1��D{' ��/Q���ŀ <>��H�s
`��e����^B��C�x�_h(��͈�h�`r��>�0D����8ʐ됼8FY�7k�W�H�aWC�0b`�����6{��i���Q��͹�	�#D;���AY{o��=!��Ի|v�erfHP�s~U`���~
�h֛-��TCR�]&�Z!h�d�<iw/�{�4ـ�Ǘs����C�<�'j��
|h	�ʛz<Pxg�S�e�h�'�5n�0�c���B�	�3p�!��Ő1+|&�u_�Zw�C�^B�Ĝ� ���~&���C��{P�1g"��J�8	�B�74�|)�a_`�����뛹t*^�p��ؤS�����|}��)��W����&Ϥ`���2d��pr!��G 9��yđ�~�%n
xqOց�H��0<1f��(�P��H�.x�ЩK�AZ<9F,��2�����r��j�2���s�<��?9�h
ps4ȁ��H�-/��Z�WA�'���P�; Ȳ�$>�����`� pѡ�W?B��1E�5D�$A��B1����C��M�9�2ð<�O�Z*ZI�$*}���%K��ŀ��1qM���,�:M�!�ę�l�����@2-d��q锘���O^�Xuc�*7+��qOf�'b��{�t��v�ǛS�z$qp�'Ul���"	b@Z�r�O:e�	�⥊Z2l�pvUi؟�bR���u|З�̕J�l���%�?#�i0�޼0R.���Xw�N���D�L?~̀��"O$�X���k�術�����*�]�����<?�2��S�>E��%�(�Lb�B�.r�60�E*���yBB ^�z(��fjyt�{�ƃ�^&�'���J�DM$��ϸ'����4i�%���G�!
�]��'����E#$_JX����5g�^�J��SX~!R��'�:�J#�X/���[V/O�CY9!�b7����N9�=)b�1��lL�T� 1�N}'\B�I�g6Lpr��îs�����L�0B�$E&ґ*0*ɲ��0
�=Q�B�	}2uis+˩E�h�$��]�B䉒$���'$����JL�B�ɗ ���Q��li1Q��ON�B䉂LX�C1�$��c�푰%��C��:iNq�aOU�E�x�5@��|B�ɢC�	"Ƅ�?�v$�E�4B�Ij���鱣��'�F$X��� A�"C�I�&*����¸&a�R3$�+enB�Ʌ9�ɹA�	#j�UY�
[,B�	+u��4��T���8�r�
HU&C�	�TA��c��4��`�
[C�	� �I�a�71`�(+򀛈9�0B�I�7�|��o�#$m��C�lB�I�q�J����0S�x$�Zd��B�)� ��CQ�̮0����P-GѶ�r�"O,"@�<y �ᡄNKo�y�"O^e�J^f�n�A�T+;6�"O�}���'��E	�ٷkɎ�K�"O|��D� 7��̓�
4 �NB�"ONM�� ��q�쐉�`��L����"O������6p�r��
a�}	�"O怚��G;�6	&ș�V�fh{R"O�p�a��\�f�Q��C�|/~ub@"O<%�&c<{�T��fv��Pa"O��Ф<���`����PH�5"O���䖞3�-!4�5[B��"O"Aٵg�<�Z���ɳI6 a��"On���8~�6PQ���+$/0�;�"OZ��u��r�jT6'C0���"O��z�k�5n8��B� ��e"O�i�U����C���{.�#"O"�@�\ �����Zu�%�"O�9�Kߙw�<���d�?'$Q#�"O6yk��4AW
��1I�On�"O��0�#@?����[�i�T�"O����� I堰8a���%&T�3"O�7DM-�r���j��0?j!�d�/O��<)�jF)zÁG��!�+P��+��g��HB���!�E>'e���˃$�P��@K3�!�� nj�h����]�N��S!�!��U7`W8Y�]6v��yb�Exf!�$*8:\�[�ċ'Y92���=4�!� �.��e�ٹ"�Vm��9z�!��@zx�i�6�A/`��D��,��!��2%0��*��%�(i3�E7�!��-0$��Q P-Gt��ڃk��!��֡�	�g��`!��(��!�DK�!0nY	�PjD��(ػq�!��
/�bM���� |�4t�A�Ӡ	�!��}��� @灴=�BH"�I̓:�!�d��qb��ՄS7 �jP��+T�!�� 'n� \����Gɢ������F�!�$���ip�$"j� �;B��8
�!��O!܅���B
VU��Q!�ȵy��$H���\̼J�LSz!�D�<��k�CQv��ŀ�=x!�dF�H1�(�T�`�"D�T/!�$� �e��(a�M
���Ga!���,��$
2��7b�V�k�̎6�!�䜣 ~��ӂ�<2�0@BaKQe!��;Ll@#B'��1�$|��AȪ�!���$y=��#ק�@�tpk3�=�!�J?v��yL��9�6<��@W�5e!�Ƞ����D��4F�l��<2�!�ѲjWnhF�@=G��A�t���O�!�+.��s@ÇY��:b�*:!��O���\��cƙ*n ���;{�!�DV�U�H���J�/�\�qsKπl�!�D_�6xP�k6{�����V�&�!�D��<"���Ց$��EcNߧm�!�䉌�Z��+�@<mSW�ۨ"q!�Ę6x��;+����o fk!�d�5}��Ά(>L�DS� 4Z!���ODV�V*�% [�%��ŐT!��E�t����2`GZ�ˏ!��P�<�z���	`:(��W͌�h[!�dW����[��/���ѐ�W�^_!�� �a�2L��+Ԕ��EK�;�REy�"O�XXƇϒ?�p��E
�+���B�"O�qr��6lI!�	�*���W"O��	��@�s�ڭs�JR�`�6@R�"O�%b�ϝ/q(�9ؑ��\�X=�"O�,r��_���R"o�"UpQiD"O����`�,����@٥X�!k�"O����f�n��1�V/G�7��m��"OD�YrI��@�^�8��/]�x��"O��� �@ u�,�g��D�<*�"O� P�W�+tPBd��	lBLZ�"Oz���aM|���9�nU�_�x�$"On ��
��E�Bq��O��v��"O�HbwGW,h�P�d-��|�j)R"O4(&���S[4Q7L �o�v�jf"O�`�@k��A`p٪���+$��S�"O�\ �+��@�Hae�9Q�eJ�"O�9���M"<R�Q�h �X�X`�"O��f�kh��H ���^���I�"O.qB��ŜĒ�F��R�.���"O2eR�&�5��cgNاRwX�X�"O*z��܁���"�֦F��h�"O���O*n�<Pj�l��A��!�"O��ߒJFar��Λ'�:�#"O����ɛ1�f��¨э
�y�g"OT��f'[yܺt�b�ą!G\���"OLa����X��hf�`�!�I21�Hi���	�O> +f��l(֔#Џ���iKcØ0�~�朁f9���:d�,I9�@]�S��@�#�3sy,�S�o�
б$���?JV,x������l�	���h�d�ұ�wdL�,q����>B�I�,��\¡DU}	������*�(��O%NPaЇ��|+T�B)�7/��L�ᄕ�~���BA%����k�8k�ă�k<d�ƅ@�F��{��V�oV�*tΌi��9z��J(&\t��1h��6l� 0�n�#ϸ�2bEF�FP9c�q��1r����(�y��!5ڙ1$ʎ�2<��i���'52ѳ��Gf���dd�)Hx � 0��6J\yk���9|����Ф�s���z���6�@��g/ݟ�0=y�&�_7��Շ�;�>(B��5nf���#M�[w���1i����x��ǬZ;�(��'
;�4�$�j�q���R� ��!�)A�~�So�1DB�I�H8���
&a'~ArRh�]_��$��Y.�x��"�ʀ���ȃN4�!��B%g-pi���^Z��Pst����M�,�.�˰���v����c��YA�V|l�K��?��<Y��!
��1��B>vL���Αw�1@��0�(�s���?�C��D�z;��C�֐	���3�D$�OD�`��C��x�{6�/"��%8Ř�^-ǚ��Ð�.�ڰB@$�q�b�	�4 Eh�+�*azB�[+��i�HY����u�%��ʚ'	8h���1�yZwL�����D
"maT,�=Z����J��[uo�1�,�T����"OX3���@��߯y�`����O$��;�r�%K�$q���W�A G����=Q��hB�ODV]K�.�<X��mS���z=��gҀ��Ƭ��5��ŏ%L\K�$(Ѹ��aA�gV�Ty�T�L˂O-�g?�녹w�d RC�l|���Ǡ�D�'�ڱs��M�'`7�<��Y>���K�D�R��8�I#h9�e�)ʸ1I�ȇ�	�F��@�l�!F6�q���e����D]����;ȉE��gl�=b�PY��a��Y�rh'D�p��@"�v�jP�Ҕ%�F���������ԃk�
]�{,a  P�];�)��A�EfAh��	�;�b)@�+L�0>Y5�A�\dJ���H/.����?2����\P�
$LĪI*"�#�)>1����\n\n�j�S4��'��@���@��)M7��@Y��^+�>��tGBH�S)�:��d�_+|nP�&)�J>��%^�c���n�+�.����Ɇt��z�B�iC�l{$�%M�`-rN�%_-�<���̴D&8�'�P�B��n�Np�ܴXI��V�׊�5,3}<���L�67�|��`Ϝ �y�g\#pmL�Ӫͽ����@M�1�?���<��ܳ!̚M��,qB��烘t�Sf��g%�)�^�iC&�y����8*{J����7���+0�󦝣_/�ұ��	;����I>?qw͓p$",1��3OR�;��»k0H��2d$���\���`�!ϔ�p`�����О����6c%�-��ܒ)�ě�+�2*��顁���J�%�IZ��ҤG�h�Z5A�
�<W:���E^(HP`,�v�Փ�Kş(JD��/�%+4X�>�{�? D�A-]\Ox\��G <�S��'�Z��#n��Ȩ��h�$	�veD6E�&p ��*X��y�Pʆ!SFPhCdKb������
�| E�>Qn���I���@	�%SS��[�'�p�O�"$Z���X��,w*<k.JQ[�Õ�?~^(�%T33Bxԛ��T����'E#yWN!#3�'���r�	',��1�i%H��ݱ�O$,Y�.O�J�&U�ů�c�d���B����$��M�,�.��� �O:yP@���N��ԛ!�9$� ba�P
j!:��'ȑy�\�F���~�i�>9N�D�c哵Y-��H`Z�o �@�D=O�����$�7BE�Eɐ`�~���^BP��E��`�t)#�@Z�>ͳ£�^RT`)��3��� �?-0^-��'��iĆz���@�H�� Ŗ4r�ZĘ��C�J�G}R)�
\tyC������©t� �h��5��ᆬشn~�J��B�i'�u[a��O�]�fg��aa$�0<ɖ��;� ��U0`i�Ph�gDs?yF敍c��=+�e2=#�m�&.�ekH�8F�X���cBٴj��WF��o �s�N��*7|봩V�r``C��/uAv�0���Ѽ-It-S"zx�B$G
���mڒG�&�Q"G�/tDx�Pa�Ѷ)��R$pv�]5Y�>u���߿_ļ9�R퓁w�b������p��T���u*2���� =v9Ī� ���Hx����@��dA0@��_V,�s���N���1��D~�(�>E�bްt�H���*��O.ȩ��(a�c��KV���ÅÝ*��)r�ʕR�f����4��o[��R��/�:b�n	s����0<�ԆF�h����%���^�NH�2HA[}�L�C���7
�A�D:�C[7B���B�ɭ{/�D	�4HjfHs��U�݃ŉ�'�x�����4,h,��#���B,�����*���l��3�֠���Ĝ�%*E�п	B4 c�L;�\�!��[�T�әw$� L����s̝�36�y"	�'x����"/���A�0d^rai  9O()��N
+�{F�֕��I�wPdP٠�x�����j�C4`�-���!�Cy�a}��fȦ���� TMzE`LI&h슶䙥�h$"$V��*e��M1T��RF�(2xR��G�W�G���D{B#S�W1@���-����a�s��	$U�
oK/:	��1�=�yBG�4���Oſ1�|�闏Ο�y� ]��P�33-}���1dg>�X7�=�3�;uвu��/;8��хȓ:��L�gN �8р��1��@��/K$��ɳb"V����L<)T�.2P0�m�3�B|bc��mh<ɕV8|�4�bt���;��c��Td������0?9�	�Fa0�o��`�詑uF�y�<��
H�ĩp���;N\i!e�Lܓ'����'D&O<L���0b­a��;NQJ�8�O>D(�R?>�%���ս{�3�ʽ5M*����:�Or̡�a�:���� �Սg^��W�I�I��*�cñW6�OE�����C8:uj�ƅ�M�je�'A.`+P&��
�2FM�-F8���.O�D��7X��N��|��$*A����� 0Ō���Cq�<Ѷ�2*c ��菪;�����o9�Tr���ጠ��g�A0Ṯ!�ԧ4*P�T%�}�da����C7@��!6q�e�F�M�ح��ɍ"fv|;��'9��懖U2�*�fEW�a�����PNA�DKȚ��'i�>}�ceE��8Bm�m����I�$�WᎿ,v�x1O�\�'��|�ѢD8#nT�OQ>U�"e��̔�D��)r��I@"O"D�(��Q�6SuB%E.x�բ�
���	�]���5#T�3�	�{@N	��G/J�pT	ǀS
�B�I�zDD�qԣ��F�a�R?Cz>�'��E9�}���R�썡@E�8=V��׬�M\���G��P�y��o�
�@���43�F`h�S�yB���Rt�e{5��.q�y��B��y�+׏lf�9P���ht�A[Ҡ��y�f�&'��Ggɤk��(�A��y­@�fR�9�!� u�K�
���y2,:��M�g����@l��yb��1�.D2GB>a���yR��&&0�r؅����>�yrD��~P�T)T �#_��鎥�yri !3�bX[5C(@����kڏ�ybn��r�����q�TrN��y2��yzi{(�/wux�8r���y��?lL���R"2@�	�.���y
� Fhr֥�'M\��!�%41l�3"Oļ!�D��-�tq�m޴,x��"O�}ʓ"[�$0��D]8��"O�(b(6��!I��V*����w"OvA	�O�&%ׄ4Yd�7D��Ep�"O�)n��[0�131�����"ON�!���:E�H�*da��{�"O�ds�'�� aF�Pd@�8�̠�"O��Y���wؾ�A�@'w�Nt�"O�#բ 6�x0C��F~�@�"O.��F�%��\{��<[����"O"���_3������M@��"OB���
'X��d!1h�6xOT���"O$��s��R�(y!g@�M=� *F"O|t���L=}��,y��H�}8$�d"O��C#��lD^%+���hK�"O`�ȥ�kؒq{�ƆV�l$�6"O��ґ��3Y��X $�(H��xc"O
p���(w�0�0��<7 	Z���,���O�ax,�W ǧF��I?g�D�0L\�	�|8��Ƞig�C�I�g�.$Ӓ���j��1��q*xC�	;�)��b��%nۘwΘC�Ict*$P���n��d���"�fC�	�n�P��"�J���-)>C�$���*��>?�Ub��;x�2C�I%ӈظ�+����"���72C�������=-a��93M�)q(��HOQ>��%/
*<�������ovZ��"*�Wt�4��#\:
�h�ɨ*�]xU�~:����O��8c��G�Q���a�`��L�aY�m̳Y|���6$L�фX��I4�'w,rA�W�V�g�U�a��* ty{�w��s�.�:��b�w��S/:F|cf]"B�x��0C�:r�^�Oz�� c��r�1Oq�,6h�)3�2�P�,@�Ml���Q�¤b�3 �4c��|��c���1�*N�Z��<!��D�(i .^�p�qOQ?-RE��5$,$�ҍ� >0pɒ�U�XK�{rY?��'�O���3��� �1�dN"�>e��O�3Z���鱟<P�	[x�S� r�OM���V�HA|VY�'����{Ǥ�o� m��k�&��1�Qp���`�O2�A�6O�dJ�� ڼM4lx6YԦ�a��	7�D������?A���#8V0j�m�*�)z�-���M�p$��Fl�IGcE�EN�Aۊ��'JR䋆:�!�Cܾ|��ꂚ|�c�>�Oq�bL��O&,dR�qU"�u�\	cQT��Au�5�Iֺ�?��ٕ;a���)W�`����`�v�<�p'��n7$p��(D)Aܐ��c�t�<�q���M)�a��	�y7��brFI[�<c��,P��$h��(T��B��|�<�e�T�?�Ę��� �"�p"���v�<1!��o�~�2`�S��Zt�EI�<i������7�M�mw
�+�`�<Y��}�4��UJW	 P���wdIr�<I����z����l�![x�#u�Mb�<�,X�q����c!���.�cr?T�0�� �<%����U�9r�)q��6D���f�#'
r3)�c��[El1D��@�G �(�`3F/7F����3D�pc��M�yX[�V�E�3��$o4D���e-�3ԠD��L�R`�1� D��Жo�"=��4c�#�;�b[e!"D� q��4B��H�󥄤Rg~���5D��
N�*:A8��R �5l�E�� 4D�hk�1���� /H�҈���7D�ԋ�^�%&xY�D�Sڍ��e8D�����7<�	a�I\���-qU�7D������P>�]�ժY����r�9D��ɐC�[K����
T�w���f9D�`�$� ��z"mR8>�J@z��� >@ڇg��J�J���[i<���"O�x�FE�\��0d�M�H+�"O�9�G
�� ��Q��ˑ?4Vջ�"Ob �)�zp��〤�� :d"O��b��P���Mz��I[�ԁ�"Odܻ��S���U�ӣL��h�PA"O�l�AR�q�S*c2���"O���qc��*�`�W��%)@�q�"O԰6�ʴ�x���� �Q�"O��"2��X"}Z�J�#�r)�1"O8�;v��by92Z�&�`!���y�/��Eg�aQv	D9�^�aG�-�y��ƑE���V�� ��@ 2�y�%F{�`��B�fa�U�^��,��`���
�*�	���� ϯUXJ��ȓ^��x�
�#����.}��ȓ"P��0D�@~NM�cl�EK���ȓ[��e�F]�6$��bFF!���/&����Ll1�	b� ��x=��84��8E�ڰ0`�A�.�(6���J�} ��sK�a�(E�@��'~>��Z#�L��G�3NP1�'���r�m-$�t���/͍/���
�'�ĭ���!E!�Mi&�3*��C�'�F�%N� �S�K).T�z�'j:�9@`�3Q��l@A��i��}i�'%ܸ�ug�=��:6��L��,��'��M�L	�g��ʥ�!=nʱ��'��؈�m	�_�8i��ě�2�Zh��'I�0�Ķm�r�t�	q:y1�'�B8x�*t�0����?R8��'�~�)� %������3aF}H�'�J�10�<c�����N4-��Ё�'�4���mF(�zup �Y�%n�e��'�rX�bBԬ|�"�j0�F-�Z��
�'��]��K��D�k���!�V��
�'C�TE��d(؃'摧�0a�'$�UG�=Y�]��B����'oB9��*�v)�+�	�9�����'�����O����V�,[�\��'� ˶�Ϳk���2��U."`�h(�'�n}���ȴ�pX)����4D�LA��0s@E$���]����Ï<D�hʰ�"(^��Ê�p���*O��)��ץ�ʝ+��#D����"O�-3�i�`��㯓�H&�Y��"O�@�A(�=,Kj� �m�!Ć	�"O�Y�d,��9�V-��-̥
�hs�"O�q�e��/߄=I�U4SZ�*F"O�m�b|n|��+����5"O�!����'���� � [vH�qw"O&�[W+��8
���F�:sR�I@�"O6�"U#۽Ƃ��s]�<$�DB�"OV��s�P?,��"��A�ld�D�#D�X�� T��p[��z#�+Cm<D�ذc�y?B%�t�Y� �,�F�:D��t+O?.bz��-�3j�A�#8D���b#Rk�� K�k�!�� S�a5D�܉f�݆Z�r�����^(J�ktc>T�T�����@�X�:�BM'k��x�"O�����$H2�;#B���H���"O�� �-�1I[F)X6���<�"*�"O������ 34(h�p�Q�"O(=K�䝵hW�q#��Q�/��\B"O� ެ��Ϛd����݋N�.�$"O$tg'�$/K\� �J\�$� a"O.�!v�Y9)z0H����!���"O��4��o7x�h	�f!�|*�"O���t��Es��+wf�
"O��`A0��Ł���+"<T�s"O��*Ů�&�,�CeJ�I��� "O��JseX�zU�!뀁Л5ʾ���"OH��+ҤO�����/$�h���"O�=�b�K�G�sa��;���)�"OZ!R!h��.���ZR"՗mX���"O�	��GZ��.Ÿ"�& [�"O��;�n$mk�\��H��"O�	I�d�:D"V�B"KH9.�ъ�"O��b�Z�6N&09t�ҪF�d�e"O*5uB�<�*4C�55��mx'"O��J�N�5٤���M��Y�%"Ode1-͘*��K��8�zh"O�5��Cԫ=+d���'[D��V"On�)2�G�5y6)��R�8�"O������F������?vcj��"O؝I �� q۬��B/ߪ%Rֹ�A"O�$��bROU���C�Y2�p�"Ola����N�䑱���:!�,��"O:�R ��u����u
�4o��m�q"O�� BJ�L�|M`��զ?Զ�"O\T��(���T�#p	����H�"O�@F��6Et���"�({r��"Oܔ�����,(��̲A_PDp"O�0h7�F����ID�,�`l�T"O����%��f��ߑB� ��"O���s&ȣ%�Lа��=
�mJ�"O%�#<i�ppׁ]�S�|��B"O��3C�q�@Mc�b\ *�����"O�|A2FL�-⊭*cl����i*�"Oz����*3.i�I��v���"Of��pFY"dL�b5���U�V�f"O�Ȋ�%J�E�d`"�J�b���"O0Q�"ʐ�WHViy�CI
K�P(c3"O�@��b.m��Pk��8q��tY"O�����X_v`AZ�e��M��y�!��͛ � �%Ұ���Sf�D��!�$֌v4ʡ��o 7�6(�F��lv!�d�7������=q���g"NWd!����q�	L2!ɠM���F1`{!��4n=Rm`%���	�����@߲]!��g0���#�_�	
�$F� S!�D��&l`�eBt#�{D#��$A!�D�v&���l��XAzQ�D��~!��H$2t��T&�Eˊ5�r.K�7a!�$[�57 �	���=z��(T,�
0w!򄁇{��u��o�y���1f��k�!�<r��]i�G �R�@A��H E�!�䆔%І Kg�>i��ᵁ��k`!�$��(Ƣb7AP�W��]9ԭ[�^!�Շ_�QǤݹP�`��vl�%!��B^���$�$���t�F��!��E.4�~9�����3�=��I9�!�Bop����Q0Bn��r.M*d�!�(�⣕75�a[��|���'�h�v�<t"2�*�`r
v�*�'����n���ܱZP����H�'����Sf����f���q��'h.��׀
4K60�qt�ق}�t@
��� R�Q��<��3aA&(��IS7"Ox��Pf>*^�����a�"Q�"O4�9�lز����h 5rL�"O�����֦O�A�G�#L�n�aS"O���ReU7*���@�26��-Ä"OT):e�Φc��(�#`�5sX> {�"O&�dn��]���'.k�~q��"O�Ȱ�ӎj'2�+%h�i��8��"O���� �7L��1'���)K"O��i�����\����"Ohhad��.���A ДJ5"O���M"k��C� \�@�f�@�"Oցc&�Bj�"�.D��pf"O�H2�A� ��1p�Κ�J��F�V�<iC ח<�R��s��>~�,=��CEP�<��I Fp��zW�>09���E��O�<I���=��\���S�^�FT`�<�'-ã+�\�H�MLj�xf��_�<A6$�?,�j� "��D�5:��X�<)�ғh�t�b���X�%���H�<Y��&SN�RУdֹ���{�<qTJ12P��Ė4�Lp�6DG^�<Y��P����ꃈW�d �6��R�<�0�3q�F�@�^i��d�c��L�<�D�p���p5��Al�1����K�<A��N1NG$M�A��Q` �c��b�<��J1��<B��9�i`��B�<q��[�
�du
�JI�]yQ�S�OU�<��m)h9�)�@H#vLd$9ҦDR�<yUL��b5�cR \O�A(��r�<ѣ�q[p���MRżu��p�<y�Fܳv��qɤ"��F�KDoZG�<AeIBr�<p�]�t�y�@B�<	Ң�@� ���YN�q'�T�<1� -$�EB���-AwV}��H�i�<1%�1>�|x�ñf6@P��b�<I�H����ѥϒ2Z���My�<�r؈Z;���a�H6t��+@LMt�<A��	;as��"��c��S�̘J�<aiJ���Y��:�^��� r�<14膢6���F�\l��"��j�<��IX��5�����~Cp(�ld�<��C�h-Ii���b� 5\.B�	� hl���L����r�`�=)TB�	�X�r�����7}Ϭ�B6hī��C�I9y�L�%k�{޵�E&k2�C�	�C��u�hQ Yd��3����+,C��/�*��2$$��%�r%�f�`B�	�U��@  �P   /
  T  �  j  �'  �0  �6  
=  eC  �I  �O  EV  �\  �b  i  Po  �u  �{  g�   `� u�	����Zv)C�'ll\�0"Ez+⟈mZB%8牶7Zn�D7sF��aH�-똅�#��n^P�Ĉ.~�� ���DV����	��o&U{��	 ���'o¬�a dW�~����
��V�
�[���F��vp2E!B��a8��4��R�rԁ�&��*U�0��I�u�݋3���m�Z0#n	%ye��IG�Fh QCڿLh���4/�����?����?�� &�-�ᬌ�\��e�)���j��?�'�i�7��<�����C�'�?��>E"U�v-�J�5!�A�=\E��	���?!,O~���<�CĎ�a��'CBk��"�@�3��@�8�I��#h@��DG|2�ieʅ�Ԋ�W�:9`@`@�r.�x@Ǥ>9�'�'U�� !��)a���r��w*D�)�����'���'��'��ٟ̖O��X�;��p���޹G�l�C P-%��h�^�o�1�M#2�i�"Fi���o�!�MKV�i�2Գ]sj���Ɏh���e L-�ў,
��)��<dY�q�I,IV<UoO4>�ֹ�C�����Ȣ�Q-�6-P��q�ݴ�R�O5L��T*[B���Ǎ�j'x5 �j��f	�D��'��� �eH|@��)RN�]�$�{�ː0� �i=�7m�����%P7>_�u�WMV�D�PQ�@hJ�M uP�D^��f�R�4V��f��|S"�`�}S]w@�]�uI��F66�!a�El.M���%*V	��H�*����Զiw�7M�ʦ���5Z~r���H� �(�*�K@�n
x�����=�te�FA9;�T�޴!$`02��Ю J6, G��>L
�Z����E�Q*�aVM�%��P�"�?q�B�'�ҏ$rM&7��O(��V�	�j�!q�%^��\5aH"G����O�ZR�O��Du>�(r�=��X��'���=;$�7���6�Q*f���U��Q�|��&Y�R�rb��3�P@o�<��\ѷ�D��,c���
U[.Yʀ�C�J���0�e�OH�$3?�oI�o��\�S"m�)Z`�W����	��?E�TCX?��x�0��:�D��o����?���'��-�G�%�F����YW"�S����'t�ܠ��iq�Q���0��l��!��#a�k"D�!��(o�J9qN�z
�Jk D��%�����g�S�|�ȑ!1� D�X9�)�0#��,ڱI�7S~��S>D�(:�j�]b5iw�� o�H��`C/D�,�0"�8I���wAǙ}nX�� �O�phC�)�D��d�D�/' `�({q�E��'(�|*�ߍ��1����)y�`[�'���cW4Th���ϑ�?6>��	�'ˎ�iσA#ʨS��;�@�	�',�2q/(s��l(q��.@���'p�����z�*� 2%�2E�(Oҙ�'��:��a,�BVOȖI�83�'cf��lP*+��B�
��|	��'����I��L�!&�%:d��1�'��${ ��p�$��%���0��M��'3Z��"eB�C�`5�ul��.���ϓe�Tݠ5�i^�'aH���jK���p��X!pn��x5�'�"o�6G�2�'�	A#���c�lV�V@yeF��f�Z��E	&��q�dL�!�4%H!EXA�'k ��7�_<J8�DM
�
$맊���]���� H ,*�╝.Ť#?���R��I��p�I�c�`%p�(��nn��Xr��� n��'��S38n���P��Ē�{揍#�t����̟�H�'_Τ�Cj�,\���e�O4�3f�.�'�y7�
1H�(�;��J�y��{E�>�y�c	~dMA���x��������y2��P�&��#�	u'68I1���Py2e�
o!��D!K�'�^-��MNt�<A�ۓ`'������I׶��E_n�<Q�i�2Xx<�
T\V���(�Mc���?��xӂ����̀�?��?�ӿ[�EJ��Hɡ �+.�p9� ::�� ����8�rm#�a�� ;���F �C�hج��#��d�BŚ������ׅ^N��%����(����It�2\�^u�r��6&�A���%�'��ɴ ��D>��O����OF�����~t�<8uD��<�8�&�=D��X�		�PY��ԼY^�wB�<���i>��IFy)4i�pİ����c�,=p!��l�@S�+�1;���'B��'�r������|���ܸa"I����&�L@�%%N�����.��{��9�zȩb�&iwdH�!�[<AU���d�r,�C?��℆��3��	J<�����UB؀����'oIv�h�EP�<	q��Q5�x+�o�p!Th�WJ�I��M�N>�(Оs�ߟ�1fi� ^��u����**�F�s�ǟH�I%iyΜ��ܟ�ͧw���U�H2��]0���P�6�� ¼i��c�a�uǍ�s��'���6��&����2,4*�B�rӼ���@/�2��VO��0<������	m~�ȓwPZ�j��° �&�RU�����?yӓK� :U�ƍ_l�(�a�T�Z0���	 �?9��QrWj�ۑ��氹@����Д'�6x��'��>�ϓi"��k$��M�A��k�a�,�'����8��+ËȽ_�f8J��2)Ӣ����J���&�^P���ɽR����w����MO�k��}����b�1�G�������~�nG-�����*G���}*��Z~�U�?�t�i`x6��Oʒ���iե+ʉQ�j�>B�,���Q}����O����O.��D�	�1��Y.$�ʅ���n�џ<�����Xlh�+ǏI'zc��(��9���?���*�1G�,�?����?��{��,�Y��qkf$:UƂD���C��œƌ�>�?M&��|�<Q4��^b1#�d* 20r�Ovc�5�6P�@�gݲE��b>c�4Xt���)�� ���q@��"$�O��d�O"��O�c>˓�?�"���Zt!@w��*}�iY7�^:�y�J����11�)]*}`��&f�0��$WX���\�M+-O�qP,8G+�-)s/̠���K1�Ȁrꐬɳ"�O����O��H������?y�OPazQ��;ZU"q0'��$�*�p�b�hi�<�6#�5���=,Ot��Eˏ�mϾ�kpj�N��=b  �X�$��*W5"ü�J7.�}X�T�/T�vƎi)�� �!B�Ae���X��d�O���:��X�O� ���/���B�jRh*���'0*��i�j��t��J7`��(M>7�i��_�a�-�8��I�O��0�OC(�D����@�� ��O���c/V���O�擼)wF�P����P��uQE� ��M��M\ 9\���A&U:��i5gX����&h(�1�����`"ݴ
�r� @�^�_A�
aNA!�x��Ɂs���O��E��Z󪉿HKm3�%[�kD�M'�8�	[���a���@�44��.V�]p��f9�Oh�	�J�5)D�>�6��Ҧ͑5ھ����'gFA���	s�1��Y�>�(�;u�����s�&D�@i1��[���)f�Ķ`S:Z�'!D��2����	�0��j��E�`���;D��*3(���r$��z(����7D���e���x����B�X�g��x�;D�����@Ÿ���D�mT�โ�O^T��)�'h�L 1�%�LH�d�����'>b1�E�D�NV����bʺ`��1i�'x�
Q���B'z��W�,C¸�@�'��4��T�OaLm�ǀ��:�Ƹ
�'� �Ō�]��[�B[�h�	�'�`�"��"1ƍ�$)�>�L	R)O:����'��`S�� _T�t��N�1�h��'2���j	��l����=)�FpP�'4rD�T�*�PV#����'���cvGV�L�p ��L^+}l�)�'?R!�P)�,� �T>��\�
�A=(��gp�K��O�n��P��q�j��9�f|3#�		|ت�+S]�(1�ȓ=��yK�ސ$&h�L�3*��}��Ub�����^�L��	ϯAj�q��'� 5�w�\9���±?04���W�:�s��*T1���I��PE{�*
��p���?u�|���@���M��"Ov�ѥ�ȞC���P�Ղk���"O��p#["�����G+fj���"O�������Z°��e.2�<�i"O�đc��^\q��)<���a"O2�	cN�X3"����$r.�r!�'��z���&�F��t`�GR���2������ȓضȳ�dڅnHb)��KX+`����Qh��qE��5���&i, �X�ȓl�h�*BL�3$f��Y���Ipa�ȓD 
�;�JD�Iް���.#�\��e*���枃���"F'\|�&l�'��Q�SCX��ȨeS��I`�K�6�\t��S�? F�Xsiܯ:�,���F�HbZy��"O��IU�M!̩����-�
E"Or�`rLE�����R�D#	T�9�"O౐�.�,v�����M�ji�'"����'�E���[^�\@��l�X��'�����!���u��`��-�'B�jE��r �1��U��h��'���V��0�)PF��s�'�YP��_�V�Ɛ!���4���'�D�A�dN�s�� ��������b��i6���%`�8wp��7��!�������n��=8����!�$�VM0A�v͚)pLe�LY��!�d�%lk��r%�N�iT��k��!���:uj�B2x�)��U6$�!�ۉaT|�
��g�<U�#,�7Uq�*��O?Qq���B�ajUX%�I9���T�<�,F?9�hTC?L����R�<�@̧F�d�%�ҕu�<bgBJ�<y$��()|̂v�W�T���Jz�<����	#n�x3&)��VVLz��A�<���_
!#�[q�6d�j:��ɅO����+��]��)rx0l���Ķ!���$-X����E=�X-$��5�!��f�n�a�֣ln���.־:�!�%'n��B�Gq]H�Q@�)j!�?�|,ĩU1cJ���A^�WL�}���~��
'J�Q`��OVx(*�k�y���U�m���V�E*� c7���y�	6egLp��Jt�n
g�ӑ�yr���¤k�ֶj���S.�8�y��.8�$��Ӌ1�p!B���y­�i=vhB$@����)mXK�ў�!�3��lE�� �iZiP7��#7����l���A�$:b�$(Yʸ��F�J��bY�t'$�!��?v�^�ȓ-[Z�r��}o
M�aù)
f�ȓ9R���JӷS�fu��
g d��a&83�e�%�����ZێD�I���"<E���:]9(h(� W.M�^�s�+a"!�D˦��d� o�"0�\�x��9p!�D�E����҉Y 1��uC�� }!򄂌Y�V�;�i��y����l#;_!�d��S���\)4���DPZ!��-k�̕�� |�rf(\ d��	�'���$+�p�B@�����-B?o�!�$���YX!ѓ�-�j���	�'M6Uz&�E`hb�3�iUQ�� 
	�'
��
T��&����A�S- ��p��'F* k��?��	���B��"�`���B�f��"Z4�n�)�c�ai�y�ȓ{��H���:y`!c]�M�ȓ��5SF��S�x� `J�3քe��hb�U��A#	w�ha�-P9G�؇ȓ �U�,F
x����R��0�����Q��qf��s�z�R�Sf=ZG{ң�+����@x��Ⱦ����юD%\���#"O�ȁ�-��F`���� �j�P��$"Ob)��m��4B�X�# ^�"3BD�E"O�=�ЋzȌ�"4�D'p�"O:عf��N؄�Y"�%��Y�"O� ;�  ,UX���ρ�N�L�yV�'���;���w� �2��:r�R�;��U�E�V9�ȓW���+���%g��8�*OS�h��S�? �t�A(���څB�r���A"O���&f�=�P�KD,قaR��Z�"O� ���J�+2�\�B�D�l�S"O�-�$�>4Ez�*��=����X��+�.�O��rb��87�!"R�H�+���á"O
��E�Uo�u�#f�'qj�"O��pk� R���V��b%l	��"OT�@UG�W��ɹ��W�)���"O��g��=W(x �ȍ���i`�'6���',r�X#�^�!i���s�U= Px�'��:S&\�n���oJ~e)C�'��u��܃&�@z�/� r��i��'�$ s �@�R���U!b�"���'��}��G��14���%��07��Q�'&����W����*Â.�������]6G�Q?�rE ��r@����<�<,�!	"D�`ô�-RHy�T+�;G�
tZO!D�8s�A�a|Pp�d��ع��>D� vF�U�<��J�@k� ��>D� (�)A�&xLs3�	
%���T�>D���s�	6�~P���@�j�X�"�O"m�D�)�'7���B���:FdDW��|��'5���+ �f�)g�.KzHdc	�'*蘀�  !�zhVn�7G����'�p!`@%O�a1N��u�B�C��(��'QdH�f�-0$��F��B��l�
�'+F%��+�',�p��єI�v�H*O`M��'*0Y�'����,|�V���<s|��'=������&8x���ɍ�0����'E>թ�h�>�Y����.6�C�'���t`��
� E����ȣ�'�,U�Ӎ�duF�[��H(~*4�������dJЍ�F�����9UA��rT�d��EH���	B�ĉ��%^�k;�M�ȓ&����!�8 � 	� =X���*S�:�@	4�9��8|
���mz�4"�'%��鳶d8�b-D�ܹ�E�Qb���D<@�6�Rtm(�^���F���2n��(��iX0.��[@���yZY��Ȣ�K�.G��Y�IJ�Y�VC�I�=�b�a""�//���
�=�2C� 1�\��(��u��L�6L=C�	ni���L�%q��SDț8�C�	4>iT��fK�'2&h�O"����
�I�"~R�mQ�* ��B��-�d��.^��yrlR'Rt�1�ˀ�Z�2ͪƤ���y��Q$1L
��p�B�B%���L�yr^�WCL�	cd�48�v�1����y	�m�=���+@�̢%ڍ�y�E��FX(��R��y}� �`H�4��2��|bI��x���(z8x����'�ybM�]B�����q~,��7Ǘ��y�UT���PFbRmlꖅ7�y��J]���HB��Z�#6��y⇄�R(ĩC3��5��ek�^��>��*�x?�Ŋܺx$tB�j?>M:���P�<i#�
Va�L�E��[츀abL�<�$Ϝy
$�����{�z����`�<є��94��f�ق>6&�"�^�<��$@�A��+7N��|	�av��n�<Is����X�g��'HD̑baWn�'F,aJ���[Y� Q���^�<��{�+ �!��M'TB:L��gT�R�.=a�	,E�!��J<V�]��Ͽ��p��(��Py
� � �N_�#1$Qb�kF7v�Y �"Oؐ触J&}E;$�U_��P$"O��2�T:%h��0l�Y�M8��'\�X�����(c���q呇��b�Ŗ0n��@�ȓMf>q9G��GrR$
�YS��ȓ>�q�'<���/�,{  0�ȓ/s.�h!E
	T �#I$@v�t��U�i��"G!3���u�ß:�p�ȓ2�������v��"��؞s�H}�'m$\����<�wI�k�x52�dG	'�C�ɏ5���4j��A%�X��ɴh�tC�ɕ9��Q�p*;7�,i�bI�o�hC�ɳS6~��B��#�x�JCD��/�JC�IBm�Y��#�5M3�i��T��,��$�f+����{��ɈTo�2�H�鈰y!�$�T��!�WꁟM��%���=yd!��T3E_|������+D،"��\#V !�䘺E/�� ņt��Y���L�*�!��z[h��7 ��T�!�Fi{~=jcf?@YP��#u�ўhxf�%�P��c A�vH��!CL5��m��lhƀ{���*x�>�s�&@����)s��x���a��]�s�D1T,��cF���G�bg]�F@S~І�+zDj<0�$�"��`Q�X�ȓ ���RÓ�})�l��$�T9���V��"<E���ܡ0���q&���Z6<=H��Q��!��6(,~)i��/ �x�G��;y!���$�a'C�
f���&�k�!��f/R$Qw֕HR^���+cv!��T�T�P�I�C7����%a��3]�@)��5�Lp����B����_���Q��D)/�N�FT4�'v�uRGc�&��pXc:*�P��Ą�t������(
�d$>{`MC�L�b��f�K�Ye:A
��;�I`D�1s�����8#��Ĉ('r}��m�&π=��Lѯ��O]q�'���V�(Ze�"-�r2��23��ay�	u���"PG	�*�X�IG36bl�g-0�O��'� ����*F�ѱ��R4��,O��@�2OH��0�3}��ƹb#bk`+��y�����y2Ǜ,2����AZ�aV��S�O2�Z=!�0�;�F�'{�Nȝ'+��|v��h kڥs��)�8mHГ�@�M�L\��@�~��ΓJ��Iٟ��䧫�䖷sJr�B�_�~Ix4�Q�U�w�!�dծG
���`� �uR(�kF�Y/�ў����iA�M��pր���VJ�nB`m6��O����'7�2(����O����O^�$к��e�*%��	�<Rx]ْ��G����.�H�[	�(wʺ���I�n00�Ɓ��W�V@СHhUXPkr��ڟTc��+�����!)FxR�ͰR���5)0q@����d�7jS��'Sr��h>� ���� �+lN���'�!���BB9j'a�C=�A �?���+��|�����U�1��*�#I%R�q�'�����@�@W)9��D�O����Od�;�?�����f�nגe0Qh�@H�@&M+*��Qp�.]/ ��(��S��	Ó^���y��"e��@
�U��l�T�J�W1 L`-G=���2���{���A�O��P&�8lҹ��F[Y Ř��O��d=��z�O��㡠	�f��� 
n����"O � b���c�ѓ�Ȗ}�db1^��C�4�?�.OL0�nB�T�'��	�-m����q��],�QE��-���J V��'tC6W!r��ˀ{]�ק��%3�F����52A�hE��O���GR3c�Lؔ��{�SS�d�"�02�H��UPR�#>1Q*Vş��J�'b4���Kj�����M�{R��'[a~��^��\��)ݏ~ޜ@W��>��Z��b�(ܞ&.�ܠ2���,
X%	�d�<9%��&�?i��?�.�z�	���OD�$�<kk��5��6}hP��Uǘ�$T���)g��Ԣ�Ĉ2K8NAA��[bdz�O)1����DOW��}�F⊢"���V>O����S�|Kb�B ��o�n�Aש�A�Ok��렩��[�
y�3閿
uX���'�<���?9�O�O�)� ~���a�u�4�yB�/r4�7"O�����N(�Z��4)T�&�I��ȟv��b�N.�
+�$�v�P����[%V٠���O���w+Y�E�d���O��D�OR�i�O�蒱�V���s�
� u(����
�){���(տ7�2�{Qe��fj�'H�O�Q�HɉE�ly��_�E�0��5fR;�f��)чv.mZ5�O|�����'e0� ���Vؼp����8-�^���O�u��'hr�I�<��ǔ�d�@,��=$�1�+�T�<��ɻ-�؈$�%u��hAmYԟ@ ��4���D�<&�vU�I0!�A%N�ܹ��I	#`�5A�-�j=�1��?��PT��O���a>̀��Y2lQ�"��w���R�De��� H��i�m$��ٰ<��^o}����9��tp6(W�J1����.��Y_�
Î T�ay��]��?!�m�FnD�S�ԗv�&�q�c��?�����'��>���*�r�a:]��x����z�<��eٸf��4�"C4F��q�My"�uӢ�d�<��FY����ӟ4�'غh��Q/P
6�p��9���>@"���ڟ\��.�RLzǄ�0c*�-`c��$XV�c���%�T��d]���Ҩ6"z�	&tǶ-{1��[4��C�B��J_w @ q���7�pu���J�B`���� 	��'@1�r���	�y��d�j
pi��_����I�L����O�f�v���#TV���d�\yr��)4����ɐ�9j�䁂��D�O`���O��?��'�� �$Ll�x����&�2��hO"4���0AnA!��7Z�j��d \��'#��ұ�t�Ӕz���ɦA��>���摟 ��'��I���<Ѱ���Ϛ��q�S�|�Yp(�w�p@ �Op�OP0cR�>!Ԙ���?>D �#ALI�zt(DPRC�%լ�O���h��d:����p�ۢu�mq�ǉ$eê��c�>�r�>�+r��R}�dgQ�dې,޾s�7�
�?�@��I����8��?qp�ߴ	��!�K��NR�I�MH�P� A4}�&}������	�M�vj\�������6��Y��cPSy�Gٞ��	��ȟt�!� ���x�a�=0<��$Fd?u��g�T>片w?�����x!Aظ��`��{i��'*��-�I?z��ʉ���Oa��	+� Vw���M@�R�U��q�$��'i�S��'<�ȣ�'+x�	��q�����ژR6���"�������G+�H���/zh���.B!�$�7&1�)�<p9!��PV�v�'��'�(�g~P>7�����1Z�CO ���%.��?��	[�]����S�*Zr��0ꄊ�����!�䈍RXU9R�c���EA�2:�!�G&`������M��J���*+�!�ʅ2�f�Y�K��`�r�=�!�$��ܬS�!�W�C�D�/!�d��֬%����q߸Xh'N�"5$!�۶h1V�yцh��P���>#!�䛕^�Y�e�_ 3���`�-ҏo8!�Dɹ62�B�ˆ;C���C�!�Ć�X�zd��gĮuW$���L�A�!�d��I�2�ChĵV�I��)�!�dß;"�P��K� h�%#�B$n�!�H'a&��SfP�?��]�f!�� ��O.,�Q��F�d�M#yo��#Dl���i1 ��20�(Q���͟5d:M��MD��c������'�!�����$�������ʭqJK#� 9"!�S������9l&�%��ʁZT@J0�4상�P�7(�(���4|qN|��hL�%��&�(Ӗ��x�^�K�a��j��eB�4D���'�N=pg|1Ҳ��	����4D� �m:N��ۗL&K�IJuA0D�̈¢���
C"ٕ���`��.D� ��;�t)a��Vz�3�:D��Qr`�z�4��"��Ĉ��8D��:�BX�J��N�!}*��G�8D��(E�Uw^ 
pjޫ4HX���6D���BᘞQ?ƌ0�F׀@���e+4D�Hk�!
�A���b��i%��i3D�`(`W#m��s���T18�S,>D��AT�s�t �D 	!2pC�.D��B�̀�- p�a3��W'Y�L�!�� �ԂsG�4TR�|��ۀS=D��"OT�6�]M���1�Z�q$$qa�"OF<���ӃVq�ݒ��6.j��"Oȑq��=����,#?>�A�"O���#��(8�ıZ�����\z�"O΀�4��+l�X��OŜ�nȰS"O���ff�!*"(V	o��p�"O�ӒOUD�~��`�,Τͩ3"O�5�d���R�@��+���"O<er���
�J1PҀ�C���"O����Ψ	�y����~��g"O^�+��Q<y�����G�<;d"O��#��{��QQ�"08����"O~�"�nC������u+�Ȁ�"O��h�*��A�^�k櫆�>��I�"O���w��;��#'
J�Ij�a;U"OV �wJZ�[�*=a��S�<_�AJ�"ODM�Q��,��J
4Ȝ�"O�M�&	(t���!�J��B�"O:ez�A	�&}��B��C�Su"O�=;a�޷}z�y��L�>�aC"O�M��dȠh�j���^�se:���"O�D��oϠw��� �,��r"O�<AG�T�*c"����ؓ
�f�g"OF���Ff"d�a`.�	S~ʵ[b"O���#J�xO%q�
�yhx��d"O��5ܜ�x�B�C+xh�0"OT ��莎`�,a��i.���"O�S�K�,C6L����O�m`�,sE"OJq)�@�>B!Ι
���-tm�ݹ@"O6T�#�N�Jڲ��RL	yv"O���J�?� �$F�%<<���"OR 	Q+�B���E�>\�z�"O~�DQ�i��,���K	8R�Q�"O.�9��ko�x �@]��!S"OF�0S#߲x���{���:鰅��"O&����T1ZŢ�YFŗ"�P�Z�"O I�A�=4���e�^��a�"O-���c�ʔҲf˥cI�u"O�-��h��4���&��}4���"O�5 ��δ89t�K�o�R���A"O�	 �#.�r�smɇ1>��&*O�}�T�ܻoL��Ri9n��S�'3�%�c���$l"�Ӻ4[�D��'�tt*T��+I�B4�0`�B7D�|�S+R���Ŝ��$RG�5D��ó�B�@�V D�%dVt[ע2D��Z�ɶ>e��B����*Ъć%D�����ʊɤ����=P-�=�Ɗ=D�({e��"0�OZ�@I�ݫg�8D����
�!R�X�J׉
n���$�3D�4rCB$+uИ��LU;/��$Pl2D� K���0�iA)�,>�����1D�2�V;�*-cQd�
�<�)1f0D��c���=j~e�Bw}l��蟞�yr��_:z�{ �M]4<8ê���yR��2�٠u��B��p@�-���y���%�Ɖֵ2�p���6�yB�'^�d	�fI�1Lj�X�M�y�凵#sV�#�hA#+KFѨGh���y�m݈UvV��J[V2�`�M��y� QL�l۲�Дz�v��"	���y�I� j��5�%�J`h�)�-V��y�ɟu���P'N�U�̐���]��y
� j$y4��r�(�i�T% a"OaI�o�5gT�7�8t#Ҽ�D"O�:���_����0	E�>��2"OdpZB�:���c�(סD�@"O$�٧k
���a� "�m{s"O�U���C�=� �B��ۗ����"OT �ԍSE�F1�P�{0ؒ�"O�;�
C����RՀ"
��)�"Oh��ц́=!Zy��@���
AA3"O�D�q�
s�u��/�(g�X0y6"O��Is���D.A�a����"O�	8u^�]A;�,NW�> `"ON��Ɇ�F���V,�6���(�"O(yQ�-@�dY(4RǫB�0����"O0�Y#�P�,T����Z��ޤ�H�<1��҆rے0���3<�1��,N|�<�$��� ��C�č
e����NC�<Y4�џq��5+2���/��S��Vj�<�4� ��0/�?dg�a�"��d�<���)��K��g��Д+`�<�jU3J�b<1��ɱ8渹��C[�<�����.��=)Ea�8ke%���Q_�<ypc��Z-$�"��ĞI��icŇ�Z�<��͈[ڂ "jЛ7]� �m@[�<I'��	�xG�H�t��$@��GT�<�p�]Xs�U�ǡ>I��}�V��v�<��T1��)�d�:;�9ks	�I�<QQ`օ.y�0�� V�j��7ͅJ�<��$�>	��c�lG�,��2P�l�<��3'�T` �@E7�����,�]�<��/4?0�1CW ۄM.�b
�\�<���_1X�j��[�&A��� Gs�<��ӫ!��'K�r���r�n�<��B�9U�$iW��k�d3��i�<wAQ{	��BL�������b�<Y��_5E��pAR�^��##�\�<iC-�D�<+B��-$�!L
W�<��kF�Fx�`��b�0�<�˰�Yh�<I���?�M $f��$J#�a�<�/��qx6�[�#��v���9uO�_�<�4�Zs_v�Y�(W�Dg��'
P]�<�sHQ���v�x��_�<sL]<��%�3F�č��a]�<�4t��vɛ;Di"�;�ADW�<	Q�K7Ͳ�e�40��2S.�x�<ic �kj2,
RH�� #"��3�L�<���'S�^�iA��* 〉�D"N�<!�N�r��h	){�pA�Q�AG�<D�ҳ	�֘z"C�;/�x�ƌZ@�<Y#�:O4hA��݆O�u����<Q�!�)@D>��5S��B���
S�<ѳn��_�@E{p%_9r��-�Hg�<�M�� % a6aɩ2XT�Y��~�<�ǁ�=g� s%�p�f���}�<�v��1�M�6dR�8����&	|�<���C�z��Y���>Ⱦ�Y�z�<��O2!�0p �D�0*��|�A�L�<�2	Э7cb��Q+�0L	8�0�h�G�<#�A�^N�9fd��HC�bOJ�<�ւ�2i��
Q��G(���Ԩ�H�<dm�3n	��'��RnJxX� �B�<��%#̠��uCԝ6��/aeFB��5/�]A#"��d�<C�(6f�^C�*8$"X�f�Q
s����,X�6C�)� (l	�Uqʦ�K�%_�1	�A"O�塢���9n��1��(��K�"O�Ȋ�g�7I�̡�×N��pڄ"Ov0*�ˏ1|���7��F�����"O� BK)5Lt�J�]�y"OV�2ĉ�]-u	��*'N`�%"Ol)CeE��D+1�'4=.�j"O|ha ��_�V�3]��ۢ�Њ?!�dϭ%e�0�*��:��aܬ}!�$=Pڊ�3iD7!ܰ*`�W�k�!�$�%��	�F��I�ިx�dD&o!�dPhݰɸ�#� =�Ȅ��$!�D��hq�K��y���e�!�$1,���*S���t���¦�B3h�!�;kr����X(^��k��U��!���
W^��[`·�`\�2r"��!�DC���X��G�Y�P�`�`�!��/u4EY߈Omn��S�7ZC�	��,l��*�����5m�Au`B�7��l��U<EZ���d�YbB�	�N-�����:c��HÂK[7)`B��Q���1��	:�ȓW)�c>NB䉝�޹h�d�7}�p��R��^��C�	<p�:�)�(�@�j +Ցlu�B�ɻ0|��g�ѭ,	(�!�aN:k�
C�ɏd���0�Єe���9qB�A��B�	3^�
��F�Y�{�{�L���B�I8{�� t�W'h�����A Al~B�5}�T��ɝJ2�J� ��-,`B�	.g'�1��cJ�j1�TK4�?V\nB�	f�v�1��ވK����SeA��TB�I9q�8�e�!h�lp��oDn<B�8�Y�E�G-�h,��i�5�B�I�r�U��m��e�u�O��C��?WѴ���=0���h���;Yn^C�#;��b/�?8�Q�Q�^�I|C�ɡ@�����4fUЁ�rVC�	>:��0;�j��G�"����;�C�I�VnjT��%ΏQ�P�+q,L �C䉹 ��I�Y�)�$�ۓA��d��B�ɂO͐xk��s
�Q;�*Jk�B�ɧ�Ψ�So�:"�`�� ��B䉿�r���=:��́we5�B�Ia�j� ����t���H!+�
��B�ɀq��Ȑ�'�'ʜ���FS�B�)Nl<sE����@%j�X��B�ɮ,�8LzsF�O�\�)E/��B�I8(�")���:u�.!a�0&|B�I;3w~�  Ȑ�=0�کiKzB�	)���2��4(%ܸ��G�B\tB�I%Y��R���V/�U81��kcB�I:8�H8c��/�����˂�mc�B�ɫ]�L�9U�F�8Ĵȡ�
�Gq�B�)|��WǊ��B4�0�V")��B䉅$�p1rK�����d��/&JB�	X�l��iW� 
�J�	�B�IEJ�=�U��'FL�� �$�"$EV�u�B(S��I�2����0���\N�ZQoB�v�D82�B�/4d!� �8LRp'�]?R�ʔސ1D!򤘂M�bL�� U�]h0;@��>`�!�/[oDH�b�<O~9��a�=�!�D�_�X �q�]M�bA!��`�!��J$kr
���	�&�r�&�G��!�$�E�
�	�cѢq�$D����c�!�� PL*GY�(h����ɖnu��`6"O�!���&�h��R�XU���"Ot�f-��~=�4��.Tm+X�@�"Oh�aTB
J�����8$��4"O�p�˫hh�`� �֯)-�i�"O�ZUAw�ڼYS�,(|�"�"O4[��QqsD��؂>w� �"O8h6G�?d��(���mj�i��"O:�{�AP2NHbL���F0fPBHrs"O�(�S�J���a�� '��+�"O<�3���?c��,#��"Nih���"O����dɺ<�8�H�LZ�=�%"OZ��AU�N�ll�HJ�zH0��"O�!�R$B!B:� �3�����E"O�̰2�A�w��X 
W �d�+%"O�P�G��Y9�i�2�Z}"O�с�/�?��3�n�q*��B�"O6�X�kZ�n3�Y�����z&����"O4`[wD<C�D}��m�&K�y�1"O ��։�.{���gG��t%8"O�M�ckN�9Xv)��%D'6e�M��"Or�[�O߻NÒ��5EV�3ü ��"O� ��IU4nQ)���X7��u"Ot���_rU�yBd�^�&�(�p"O�(#�U 63�$���	,x.�o.D��@�fN�#�r���y��*v	:D� !�c, l��%,�2C�Ь�f5D����M�cCt9ç'u��*�>D��e杉
��!��ݨ4�R�!D�D`���C[�`�7�O^ʵ뤇2D������o�tx�lDo���x&D��sS.�?@
9կOe)�dE/D�4��i�s3ʐ����=���4�+D����B� ��D�ƻ~[i"+D����j�D{�ȟ7}�$k��*D����R�/,�R�(ޓK����H)D��ɷ��7|f�Ia���[+D�$)T�5Ri�u�ņ��}�f5� -3D�����"w�(�`0�G� �����A?D��j3����,��*�#)��Dr#�=D��9"�4k�<�Y��IY�p�A:D�$��߽-��0[O�%R_l��6D������P�Z�1r��#{4�w(8D�̒�(K�WK� D�ڡa��9ħ%D��@ �G;�՘�
Y'ь! ($D��J悃l2Phu(��|�R��%�-D�p)ǅ��`1��a�L��4�RPA)D�0�$F|��NӀ8t`:D�(D�pf�,k�tT�Ф!z 0�D�(D�@q� %*a�I�q�&��0���:D��3� ��?������^�I2�P+e=D��q@%�H�\��G܈Qä���:D���ݜ:-����^=�����$�y�$�3�r� An�n����Be
��y�c�'lu
�;�E��p�N`�RMӘ�y��^�T��uP�A�'h����u+�y2c�=�� (��_/uL�Z����y�L4`LI��ř-ZdrdO��y���3��`���:�bm�Wg�o�<�1+�>z��RrI4,�^����J�<���e�L��LY,h�K1BN}�<yBeec��� Kh�ň��X$�y�� 5�CHO�D�<h��c��y��РRtp��@�>{r��2i]=�y
� 5XGB$v�4�:@�O�OF�=&"O8
eL�.:�������p���!"O 8+e
�WDҝ­�!�J�ʲ"OΥ� ���#R<躓���4�
�3"OPm{���t%B��囹C����"O� �$�ڤ:;�5�.�J@V"O�52Pj��@Xj�'P!�D܀V"O@(q�f���0�ݠ8���g"On(8���)>�X8	2얙l�"��"Of�Q��$⚱x0#�p��P�"O��9�h	<Khx*�a�&G� �k�"O2!��;|�(�0�ֻF��ɰ"O��z�F�6.�����2��lk�"O��Ǝ	 m�|XT���A���V"OB���Ha����L]Cq���"OL(�Ȟ�U`��"邔g�(h%"O\z�@45!֕��#:�j�Q�"O`�@��1�yC���O3̱�"O��	,I=��Rs��0'�A"O�,"SoO�sC�\���*Ƅ��"Ol��CE\8��=*ѩd�D�z�E2D��k�9^b^:@�
6,
y��`>D�h�'N�;i��M�7 �<yR�A�?D��aɌ@*��6�I�S\"� 2
8D��@q��'>3tP!U�Q�`!����L�<���\�V�DYJ�b̰<F�:A��@�<�����L����0j,��q�Y�<���_�E��!��w&���@��M�<!"Z�Bf��af�0
V	xEI�q�<��E !;uJ� �垉���iǬ�r�<�QR�5̸Ro�ǆ\	�-�O�<ץ�'JB�*F7Np-�tHN�<�kE�%��YPpꏰ@�T���G�<a���#���5��	<��P-H{�<Q�)Q: �i�f���Б��g�R�<���5�
�8'�Z^K ��3�VH�<Q��N�\��� b-��%>��3�G�<y�G���-IG�P�#�hdS���i�<�IW8Ҥl۲�UIɈu#Ai�<���
X���PoN�mcx �n�<I�e0 �{�*��j�42�LE�<�S�V���ԢcA. � %"fƗ_�<� ���J�D`[A�8� ZӁ�D�<)��D�w�pɣ��]
d�!��@�<� ����Z��s�ę2u�a�<��S�S�H�12�Y�D/V"b�E�<Y�mܚ~�<���H�Tcv�+2)^�<�p��egR�C�I��� ��\�<�G��'|��T��<H}�ɻ���o�<���H�b\���'�Y kd�+U�f�<�FjT	~�h%���>#`5����~�<)�o�3z6j"�B��S�b�p`B�z�<	"烀5�X���Q�L���'��u�<��%ī(��ѡǷQ��):7�Vp�<�25r���Ve³g<8�K�<9gG�f��`��(��>	��E&Gp�<	����͊b��kD��Y�
�Q�<9 �<A}�qh�a�d��qGH�<�f��,yr�0�f�Uy���n�<� $�'�����ϼ{@��"�g�<)����x��gR�4"�4�K�<�1(�~�htjB�"�:!����J�<��F��5��
�x s��TH�<���^�S�q��1`�ebMH�<� C�K��m?�1��C�z�|��"O��xuG�1B���7H�#r��ؖ"O���ŏ�X`8 2�':���8"O��+�.QށF-R�X�p8�"O�p�@��->=��Ð�gV�t��"Oha$lT3��iY1�K�B@���"O�x2�V��������u�"Oh$�f�Y��4h
��]�&����"O,X��X4h��]�EB݄}�ʨ�c"O�Q	�`ۨm�x1��Q/-��x "ON�2AL��q��D��'P�y
"�`q"O�5i�F�/a���Y"xޔ��"O� wi
�(���;��7kor���"O�4���_-ae�M%�\ 8��"O�m���	�e� ��\���"O�H���]�����Vp�b1"Of9�CG�{���y�ܲzO�1�6"O@e�0���Y��Y�fg[��r,��"Onݸ�Jֳ�b0�D�,t�`�b"O�L��iS	Wx��㡤�!L����"Op���� beV��k��64r"O������v�=���R)����U"OB0z��<71��a�(;���7"O�E�À{;���0O��v����P"O����SN��]��L&�$<¥"O�����2\7P�p̈́-P3��S�"Ov���FW&~ߤ��C�#Ӕ��v"OZ�j�'�T���¤ǒ/7~-�"Oj��D�6窐�qğ\ūv"O�m�G*ԿR%���v =��iU"Oj��:~�n�2a ԯ^V��"O�]��
�;7�����S�-I�iۤ"O�P�lU�!I�4x�"C�̠��"O����8.�C�@H��ZUs�"O=K4iM�	�zG.�&���P�"Oxa��̓���s��k�r�q"O*�x'�`)v�v�!Zܲ���"O���j��q���5�A��H��"O��ՄK�[Р�������P"O�K@���ұcŁ�`�L�hc"O05��Ax2H13�R��0m@�"OJءqc�(�m���$��ӡ"O@�Ռ�
J��ad�/���Q�"O҉A*¦A���(��A��E��"O,�A��r(}ؐ�׋� �;�"O�91�߹4!4yK�b�*:Y�=��"O�q3Δ"�ʑ`f�����;r"O�=RSIΕRB#�CR��Lir"Od��l�Y�3�hU�]Ĵ�+t"O,�i���Uw�s`�Ȓ/�l�"O�M�6���S�L��󋅪|��	0"O�M�F)z!�M̓D�:�qT!�2d�!��ν.�(����ڟ2��I+4A϶]�!�ܶ2y�Ǐ�iZ9S�B�;�!�d?c��	�q��9:�6 ����&�!�˞)�d� ��G�4r(-`E{+!�D@�G��(��	�L����]�!���C�$L�a,öbM�(�a�BT�!�)��`B��O��M!0�̥`!�DY�k�"تǎ�r��)Xj�F�!�D��:&�:E��5�r'�>�qO����
@r��1��9r��S�|�hݲ1����i�7�"8x ����y��	̩�	�2px��L;�y"�g��1��Z2#���;��R5�y
� �bS�jXĐ�#�׹�(@!"O��)�@�9?"!ZB�ӭ!�l�!"O���Db8
���ѫ��ͤ�"OP��w�F�VX4��C�O�!Tj�8�"O,:��<$����		_^�0�"O�\;�J["`�>]�6
vJ�}:v"O�$B��-:� 	��O�Y�@�ys"ORUPH9Z,�"��"8�0"O(���Z�A�!��8Q�j��"OX��G��83��1/}6��`"O|�swƜ�>��	���!_ԍy�"Oj�qMG >�	�q-Ө}X����"OR��P��@*���
I�YF"O��ڦ��	2<2��ߚS,�2F"O��p�_v�V]�OA�N�v��"O��"UA�(g�1�����aL��Y�"OB�J�jN[�j�x��SQ�i�G"O)�t�(�l��/ڥ>L�Ыc"Oʌxଋ�t�4���.V�&L�"O*TS��țs�P���M�N8Ep"O�U��/ҡDX����!�4�RK.D�D�"H3o�݉c�^�0�\�$�9D���c΍*O񒬐��Bpp*�N,D��(�
Ų�xё��<U�,l��*0D� ��P3{�2��G�G)x�0D���ƇU�G���6`ō\���C�N,D�D�s�/2v��U��2:5�E�%D�H��bY�#n���&P>h�1��b#D�`q�űp����K�!s�(#D�tB�BC(&�5�3ę�}G~�`� D���d�����3|�d�P$=D�٠ڵO� �Ã��c*2�5.D�����,+��%;d%ϟj�QC,D�8sdă�){@�$O�8J��cS$=D�`��%S�Ej���3�X��h*;D��Qd�xY;�`I}���/#D�X��ߎ;ͨѤ�J�iߢ�"S�?D������&��˄�2JԵ���)D�X0e�C�2F�0�8-E^���N5D���afߨAP|x B�4k�dujF	(D�@0@�V(E혠�V�V/=����!%T�d�WȞ,β]aj�;<攱C"O��XdAӸf���;ↂ��T��e"O��
�=�Mib�ؙ<��A U"O�Ը.�		YVeȻeQn�z�"O�1���	P�6|9r�{=� �'"OH����2e�&����.%��W"O-�6%]���D�Y$B<�Y@$��X�<9�D[���ׯ�#?~q �n�V�<ɦ�A�ΐ �iC�_>�pd�w�<�t�/8�da�"&JD�>��Ƭ�s�<�sC�>SVa��ț^גI����U�<���>]>�ӑ��azT�UD�N�<9�NAu�BIy�.ӕD�0�d�K�<�hɂVx&p� ��K��+��O�<iR Uyd�С
� �f��P�L�<��ъ�D�1 �<�R=���F�<�v����ɗ�ߍiv��w �@�<��AO�sh|��� w�p\�ƦYb�<qV�`M�d� ���>S"ng�<)Vfʁ0p!C�D�Gq��2�l^�<!���:LG�xeGA�o;ڼ��ƎX�<�R������u���r������kM����KӚ �Ti`���;H��=��S�? jX�e�f��H�`�Fr�K�"O:�J'�z�-*e�L5s0<��"Or�˖ ��vT`�9 ��:$:4(:�"O�z1e�(cȰ8�� �*?��"O.Y��F�Z�\��һ%v���"O�u#�"]$rxd0	N�U<(��"O�	�dmM.~4��:\hT�r"O�hB��D5��	 F�|
Z���'���r@L�`L꼐�F�Oa��'����L�\��D#L�l��	�'�p:D�[���j�*��1)���	�'a`i�c͍�Ed@$;�e��~ۜ���'Q��ٶn� j�@�-�z�ܸ�'̰(��FA�k�8D�䊈�s�i��'L�0�f��g�J(p�'��:����'����W��J��+�@ 0z�4�
�'�, ����X^�9�P�č#lq9
�'�h�b�
�D��((㉜"�t��'��mr�C�y�6U�f��=0y ��'BΉ��@+ux6�*&뇯�6IK�'�F�ekS9?wĭ��H[�aSl���'�Tm!s�W�Y'vmPF�>U�M!�'Dq)��2Y�\�%�H�LLd���'ٴ��W�S��0��+�71/��Q�'�X(��f �r�#W�˒(�V��'�Z���.I P>�(dX=!�ЕB
�'�p���/	�d.6���ӟc���	�'�b��U��"���/ܾ#��t9	�'VDrǂ��6���Y��sȘ�r�'�P�	"��|)4ِ$�=��]�'�� ����1*�t��c ������'��ĎݖM�lĪ'L$u2��q�'BrĈ�-A)hfy�#���3�'�X�Q�+K��C�J_�j��'Ȣ����HS2I�陒R�Е��'z���}d&�R��	b�0 ��'���7`ՠeǼ��g�9*�ظ��'��p �C�k�*���Q5 $B�'�2Ũ� F�=�(��elCk��Y	�'<�-ɦ~�Phu�M�z�~ur�'�b�@��) x�<�3�ǎgF���'�`��M���q��_��a��'�R���瑜\Q���)M�dm�D�'�4��|�t�XB�����.O�!�B.Q�F�a�+ߏ]C�uY��Tm!�$W���(`�F��3�.�RC	�!��ӻ>����W G�A���	B�bt!��M�@�㠀B9֬I�N,a!�$�Vef���D��M�d+n��B�ɚ�H,��@#�2����G�i�`B�I�GX���Q^
K@�ƻd:^B�ImV�`t4r��E#
(B䉢L�>��r�Y�JBB�B���)ݰB�ɏ'��I�H�v�ĉ��LW&��B䉩k���ˆn�%�1��픪QF�B�X�&,
х��so�Z�R?�B�	�k �� ΐ>��у��T)aN�C�N�jq% 1q�v :�'��P�C�I�b$���S�r�R���"~H�C�	_�%��,Y>ej�� 4鉮	���)ړ�v��w-S�����G��޽��k3`(�ᇀj�r�q���� L�ȓ^���l� B4�Q�D�U��lvXC���,h�T�c��LɆ�S�? 84(��Wv�l`�#��1�I�"ORQ��.�w>����T�"Op��Q�b���8�^s�6ls�"O��R�/ŧ-˒��/X;D�6���"O���*�nh�h"�G�{`���"OTT#1�YT��,
� L��"O&m" �i�)����_�
؊�"Ob�2�C�X� '�;D9T��"On5Z1��#M^���MFnJ�!�"Odm�e�O 7����4��3&1�"O�9���r)TC���<c���#&"O����f�;,,"�D+?v��!4"OLu���֯>�8Q �T*����"O����H�K�D�7_��js��`�<���N=O�x4eT�B��Q�TG`�<	�bYC�����	��%'�b2�X�<��Ɏ�g�j0 G�Y�#5�8q5� T��x��U$Xb�  a�do�ᢂ�(D���DXU�i�èՠab��+(D�,�uf�
o��@�ҽ(��es�
(D�h�2/�T_0�ui�9Cy�M�q�9D�0�#斲��Q�MJX\1�D�"D�x�'x��i�A��3,�(��"D���s�p��P���TE�\�!�5D���'ϊ$�
�$�k1��8q�4D�䒁�u���HE��mhZ<�C�6D���7��$��Z$h	9n?�Y"s�9D�ZgL��T�� �-����}���5D��zc���1lZ0�dA47�ba2D�4BѬ�%INJ�I�e]�q�L���1D�Hb�j�(*e�d%�"g,a1D���!j�&*dD��j�T.��pF0D���c���%E>��1!����E�dB/D���Iɢ1��F�	�<}"�D�!D���T+��e����Eۗ_�ͺ D�|p%١M�JpY�3�N���#9D����C�5<-is��Ԉ�Ä2D�0�W[ 9#�9����c0D�x�e�#~�!�	��W$�� $#D� ���?�^��FŔ��br�<D��V�&Oʥ`�lP���<D�����W	��B`�nY)rG;D�`Bp�M+JN��§Ĝ�L��)Ua:D�x��)��43�5�c�� h 9��(+D�	�㑺�v�Qun_%1�&XCGk4D��CR<�1��>����1D��7M��_���v��7���k��<D��r��ݯ<cL��!ZbI�3�;D�����_�U=<����Ҕ'�|<�f>D���c`مY$�r����-Jhb�k'D��{��
cZL	rcLZ�#�PK�&D��Ư,�LU����(B��!k��*D��@oT'6`�������w�%ᓠ'D���@ߏ.@��4Km�f��&D�L�u��7p%@]âI��D7�Ҥ�.D��r�ND3w=6p�L<g���Va,D��N-C�2X�A2N��EK��)D��@���/���%�9[�\���3D�\��C���p`��ilVx�0�6D����ʬv4z�A�$�(8	8��6D��S7"�/8߾�K�ϲT�`��Um4D���2aX�@I��/�U�$lj�.3D��� q/ �8�
��AI��i�+3D��5
�"##>��@�
=��U�6�>D�� ��X���GL�{g�P4�TxI"OhABC!ʬ4�0+6I�%�X�9E"O�����sR,I���Q�S��\�"O�X���NJ�ԡ�H܂]�P��"O���hӹ'ٜ��&^��P�R"O�([�J��hY�ާ2�HRC"O�13�ݑ$w�ܺ�%O�cz���"O�l���Рis<Tcu��1.���"O�,js�Blr��c��
[ifd��"O�-Y��#'("�b�E[��N�a"O�q�� �7ufp�$��>dQUi&"O�$��c�l�r�Ň�J+�ɸ"OʰJP���0r�Z�$��D"O^8(h8(�H-�d
y����"O�s�N�L���0L�oF��Ф"OX85'%����*F�h��"O�{�'A�T�a)� d���"O�y�Q)[3;dIS��-xr�`�"O�E��DK��2m��I�I\�в"OD��*E)<���B�$�]7�!�"O�T�SD u��)Kp���A4x�#�"O���f��A�!
Y��u"O����c��+��(H6˃A�6���"OD�Q 
�.A�b��%c��P�"O
1y$F؅TY֘栆a���%"O�P����J*�Q�5>�8���"O��#f\튣'��"�D<�NC�<�옆3����G�$
��)eNW�<Q�,��5�t �"H�h	%�R�<�&�]�)Ef����w�6���@V�<��-�s���¤��L���r���O�<�Q�;"��0����=��$��R�<�����YF��E/	_9�13��d�<��␁�.E�i�	�2��4AY�<�ߋ{���`0�c�a�cNK�<����
���+u��Jt�}��'�B�<��CO)SU�y�'?�襹���@�<y2��>��hd��<H!\����}�<���]�]j�iJ���[�:���HR�<�BR�8�
t���n[L����U�<�!�?p�QXDCx�ХQ�<9R@M�v=r	r��#IrT�DKMJ�<�d�:%a�1 sH�:��-����D�<��lH$nejl���-�j S���}�<q�Gӓ]��A��eߊw;�+��OR�<y�ş{�x�Ǡσ@����Ys�<Y�Ø,��XS@�� t`�-�$
{�<108��TJ�ۤc'F�ÒM�u�<9&ƅ��x�$gZ�a]� �Bu�<�a�d��'T�"�����u�<�qi��G���S�Y�9�<x���Y�<qv�L%d��;"���P)�f�S�<Y6�D p[0�Z�s_� 5)�C�<�Ħ#3�n]�֫C�[��0�΋~�<)$jՅkRdr3��� ����2`�A�<!qI ��R�����(c����i�<y� �S� �X��*,��1�o�a�<�n���=�0�$jbh)�Pa�<��[;U��YY1 l��MIE�<��[7u������:<��A	6��F�<�æ4JS*MK1Hĳ�lԸ��IC�<a�/�Z�
P�S@�V�4�H�JQA�<A'D�
`��h{�i0Wy�&g�z�<�Z�C ����a�)C�YX L_�<� <șԂM&@����!�	�E���3"O�ͩ��+w/脒2��V�pYC"OtU0��rg2h4�^*�eX4"O�-hQ��u�l���ՐY�-�@"O��#b��j�^�B�-Пn���A�"OT8#��s��ZM��n���`"O�����7����+��lv:TC"O6Pb� ��F�jأ K�`,�R "OȤ{��h �(�$Ɉc'�0��"O�y℄�3Vb�����<���F"O�uX�-X?<�e:D��4����"O�v�϶;��,���]&�<�RG"Opi��fYNR��;��ҥ%�\t20"O�,	�cD�Pr
C�g�J�ف"O���&�-{�j�\6u�h��"O�(�S��!(�J��)�t� 6"O�0�E
@����C;�R,q�"O�\I�Ė}��8��X�"��f"OP�!S��{�X�����dS2"O�j�l�Fn �"���[o���s"O���Ű�$-�e U��Ad�u�"One�b�Rc�b}	 �ܖ*R|��T"O��#$��2�50ÅG� +Zݳ�"O��xT��$s�T��@$�6-h\ȵ"O(Q��j3�+��^
��d"O�h���^!��A6�<�F���"O�����84�PbT\T��4�"OD�ri*mc��i���p�
"O�X�ΛsR��p,�&Lf�}�Q"O�X/ݷlӊL�a)I+l�`)�"OR()��P<Hi~a���;�
Lҳ"O,���K�+��I�DZ�>ɒ���"ONPR��"	�
�h@l���B���"O(��c#�;Q#�XQ2��~�v�`�"O��a��$
�B��� ?�A�"O��$Oa���SiN� $ڡ�4"O$�"%i�����F�?�-�#"O���G!R4j�!��4�T���"OB� 2�F1�811��IC�"OK�����H!*������Ȩ�y�L��7&F=3 ��4-�Փ`Iډ�yb�$)U����G�	��#����y�(JBI&��-��jn�2�̈��y"!�)�di�I2s�5���yrIȨƜ���F

&j�p���yR �L�������"}�(e���yb ��+���/��FD `� ��y"g�{�X����1*#����y�䌀X��a+sF5`����!�y"`ԶH����ك,8� 2� �y⪈�m<D�r�GG�?B2�+�%Ϋ�yb�B8g�Z�;Сǘ:��!m@��yB�ƐZ\8TЃ��4V.�p$��yb�?{�4Q��F�0��ѹ����y"iV�	&��Uo�9t�LH�#bC<�yR�4lO.��c���mߊ��h��y"K,�|�PiލRJ�,�	���yb�A
[���� _L�(�2���y�GW��d!���.~�Hg��y�KUb��L�B�ԏH���Ԡ�yB�X��P=���KX�pc$n"�yŭ}f��c�CV�8�b�'�yRŊ%���7&W<q��x��jZ��yR��&�(��W�dz��CL�4�y
� pQ!P(�Y�$%Z�l�"O*�zF@S�"��炚?9w��!"O蝛�� x�HdPV!	/��� D"O���)H��
$"���@l�رu"O �z�� f����({]��@"O��A�T���⠓�0O��b6"O���Ç�z����W�R�10*G"O��r���s@�R��u���"O�y�#�V	o�XIX�E�2=����G"O0��C!�ws�p��V'l�c2"O�)i3i��!kȂ¡�q��LP"OFWJG��ڸ�+�) ʊ��"O:@ O�5Wh���H�V��i��"O��ӀK�p�0�ԻqAZU"O���`�7�°��ؚ.�F(9�"OFY��,X ���e�-��À"Oh�pӠ�Dm�aب���IR"O����B6W>���%�u�vP;%"O II�$G4f8<	Z��S.aܤ;e"OJM���ބ<���wĆlX�s�"O��(F�U�=�0a��c�-R_4�#g"O�`�l
�u:Y[�(�")>�� �"O���E��2� �AW�O���"Ov`��l�!m��=��!^J����"OH%c��ґE5�9B��P1?�.�xT"O�`�@Ԛ"(��Z��6j��5h"O�	�Vd�)#W��9"�ӑJ��y�"O�сv�DCҌ�U.�<�E�5"OZ�آ��D��­�Cx36"OZ�X��G97�d��6͑'�9Z5"O<Y���;es&E��	�(�ZA��"O�ؕ���M���ËR�5���%D��w�.@D5@O�pu�i9��!D���"鄈G𩻶A��:�p���3D�,j �N=X�J���<IL�d�dl.D���GR&��\��7km>�V�0D�,��-O"f��d
�4k� �E-D��Q!� �uw������X�cF,D�Hѕ�o�R��������n+D���G������bUH{%�6(_��yҧO47�� B�"G�w���⠃ؖ�y҅�z�:����9XN��a�=�y2��)���p*ƬG���#��[��yr��>�D}�oJE�h);��R��y�%U)F=����N�F:������y"G�U�&�Z��̑=�
��Bٖ�y���D@�ѣ22���bl_�y��QA3|�r���-�n��G
9�y�ȞH����*,���9E�Ǐ�y�ڡg ��
�Ň�(d��C�yb�Ku�m`�� z	Qt�S��yb��q� �Ȟ���L�Cb���y���n�4`eN���5�_��y�選w��{th�}!�,�5@Ʒ�y�g��&�����#L��$����y��p���c��)B	<��dž�y��z���c	�9�2����5�y2�ۨI���au�*��Ha��yBbȫj�P�"Ą�8���Hq��y2 �����f �>GV � ���y�B�09����G;#�ؤYS˒��y�lVL�⸳���!*X����@��y�ˇ= 1eh����.�%�d�ʛ�y�_��j�c����!�BA�y
� �L颮�<���;��ÜN���c"O|i���j���s#2S�pt��"O�����+�J4slƦQ{�a�E"O~�ZՄb^�mS#�&_L �b�"OL�n؏2�t�0�A�A<��b#��ҟ���d2m���)I�2�ܘ�S�@�86-�`�aqO�dB�9+V ��$��ZV �i�Ν�[���Op&�زؽ*b�I�f�Ôi��]���%	��c�Z���آV焪P��m�'-���!��X-�]y4*ɵhT��Fz�m���?���Q՛&�'\�e�<у�@��`B�ܣ����q9������I8�	<&�����8-���!���>����dKǦ�`�4�MS#
�\��T��
<"Ւx�E]?�	�X�F�'+�i>=����!A�� �&IE�eKbo�>��1 �M |s�УW&���� j^�/q�J��w���ð��A�[#L(H�6B�⦭��fH2���j�Os��������H�k��������˕�n�)��Ħꛆb��?q�e���'�?7�� q���W)�#m̱�����J�$�O<��5�S�S&g�Pp�#����� �hxv�<q�i���ig��]�-(5�`�V�����F;�LʓyTFX�c�i2ayb!$TD�&�ج��ӈ���H#0��y�b�nڴZ�+�D���Z�I7�/��H�	O5U�E`���<i�X1���ԋn��T(��f��D��h��c/��ZP��Z8�ze��%�v)LM��J���t������8�ɬk���<q����Ĉ~����f��-��ʴ@F�%�$$��bV�� �:Y��_�!h�		6)n��6R��$�p�O��	�7�9��f�&g�� p!,(��d�/$��M��ԟ��I⟐�Re��x���`r�D0/ud�[��U��zW�ـ:ԑ۔�Ǽ>k�xXvm�;D�p�AB�I�eS:p�g�*Z����W���@�6�I�@�B��r�L�5N��tO��">!D��Hn��F��$��gĬY�,\Y����K�i��[��IJy���*7
��T�N'6m���t�!�D��B�b�b�.C>Ah*0P�3��D��5ܴ���o�Bmn�$>X�d�#;=����J��<�6B �!�	ޟ$&�*\e�f�4`?qx�G^�7b�i��	�ډ��-T� � ���+� �HO�H
�%�\����e��xd.XP���|
 O�h�Zš6��GX hdnx�' �8���?���T�i���(�պ�(X;]$Y����/�?)��O����0�B51��%#P�Һ9J�A2�"�O=l�M#ڴ���2H���!� m����l?ц+ cԛ��'0RX>iSvGG؟�����鉂�l�={W�qerh�Ƙ {<T�5�ݻVI�G�ʌ�9@q�?��Oa���j<��-܇It9:!F�w-f�{a�i|lQ��7WV.,Bb(�{ZNe1�dT���k�ѻ,�!���B�Q�� �/X��E\3�?���3�6�'�?7M�.1�̨#Lɍv��wNǍ18���OF��$a�\-bm�+t��Իq�I�v��g��'�M{�����I܊[��-�3n�|S�)%�Y�Guĵ&�Ѕ��9� p   �    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   `
  
  �  "   �(  �0  7  V=  �C  �I  6P  �V  �\  c  Xi  �o  �u  !|  �   `� u�	����Zv)C�'ll\�0"Ez+⟈mZ�YL�I07)��Dw�����c]f^�aPnӗ[��9� l��t�(�iҢJ�1��ݱ��׏X<X�;t���'L0+��PD4��gŃ\�^r�e������٬8R������.^�Y[�&���hq��|I:Wj��|�D�LE��H��������N^lq���ɷg�*ٯ(�>�ش'�����?���?!��L��m����3@m� �p)eY����?I��iU�ۂX�p�I*rY�������Rk� CC�N�L�l5Q�l�;UѠ���� �'�"�'�bÌ��Mc�1OX���)��( \0�x J`
�'b��"=!���n��S��/ #���f�}�5���YX}�7O*⟴����!�':z��t�ݬ-�$@�'�Wat�1��?y��?1���?���?�(���]�>7.�8'e�$G����M��x����ʟ<n��?y�4�?��i�v7��ȦQ۴�?���+VJ�+3hȽ�*�A��]��hOD8��iT��нp#jM�~td����#�6�2�ډ7��$�Gg@X�6mW���4�b��\� �bBˉ4���� `�{�޽I ΂�G��H�i1�
�7!�[t	A���)��b±P��mp�m~��%lZ�M� K��((��e_�6����∊�gK���3��1_��Ѫ#�i{7�Ӧ ���z�h�9��E���n3#)����?�!�B�� X�3�ǀK����np��el��M+!Bϥk"��1q�RN�� Dƚ�`���JT*���J�2jp��icn�b� O7C�t���.�\2��'l�O�x�oފTdR)i����d��9O�����ğ`Z�i�&�M�͟Č�S�V�%.�ɨ��v�@I��'������	ǟ�og��R'v�xb�@�Dr
��`��s�������B�C>0Խ{�:��H�Zy>h`��]�?�GGڢ FR0���b�a"�H�� �_��'$���!�����Ϻz�>ճ��D�j��O��2�)�'Dz�,co_	8�:��vė�Ml���ɇ�?�D+ܪ{�"!9'���Q�v|S��[�l�?�1f�G�O����J�ν��$Htdj0jF��!��7��e#�+#1�D�յ�!�)2%Hd��&Fe�UƉE	!��I>)�N,�/�Bͪ�Q�i�;a�!�Ĕ�<��T���:&+RF���PE"O��ׯ8[ <�q����'}H���S?w;��ծÁf��)�#��ц���l(D/K�o�t�aV�	eV2U��O����&+M�X�����K�5^��ȓ'�^=Ȱ�FE�m���4�ȓscx,bgAӴ,e�I1��Y����Cl�a��@+���z͕�l\��'R��	�����%�8h���D�#b�J8�ȓ ��vGT�kBd{*_Q���ȓC��q��nA�Q��3W�������3�b ���x�nY��L���A��BJ^���Bp���B��)�^X�牮_���ڴ��D@�w}숃�M	B4!�Ӫtx�V�d�	̟`�	�����DB +�A��,�5h:m�u+ݦE�lH#�ė<���oӒe#�$�P���a ��
n�pb�ʯ[�v�ǥ�n\:�1����� %lrq;��K�Y0ң<�#�֟���ϟt�I�@T\Ѡh^�@���Hd�F�6h��'����g��=kt,ۼ}�>�F��Oں��D�쟄+�B�q�9⠆�eԤ�"��Of���x���i���'���`���4>�N�(U"S���P��F�Hf&��	՟D�*��9��E�%>�N�V�.?���(�'�(o�<��aL19�Gr~��?hPcr�G�_4$Hb���l
c?A[��_@X�r+�!U���:�6?)%�ԟl��k��@�'jb�P�#eA�-\,��腈q��&�P��L�����e�ڸQcVX1	�tEb��4�F��>��U�ȅf�qk@M�^4�̓����oy�L�o��d�'���'��~+�4h@I�U���C'�)�x�[�B�1��ah��s1̏c�g�,*`��IG�\�w���`�Axa K{�TYI��\f�<��_�g̓d
�h �t��S2�L$]�	d~�$Z�?y�����?I�Kly�,	eH(�V�ڴO��)�'a�I1��	�$e�J�:D�.O�MEz�O�"Z��c�O�`��}٤.�c�hZ�Ŭ@�� �4�0>1������C_Q�� �%ښ	L±��%k:p��쎶.�B�qOJ�n`�D�Bj<���79���脩u�a�@�]=_<��B<I��Y�A66���I����� d�<ɤm���u���2L�j���a�ɍ�MO>�1�ҡf�O�jPJ��?�x���ڐQ|~9���$�OD��O���S�85~�h���X�h�ҕb�t�? ���g|��b[E9�y��'��-Ҵ��'�R��.¾r.7M/U�kd���M+�K�Gax"�X��?������E,B��5a%:���4ȶ^��'�b�'�
�
�K�$q.,)bE�N�"y��� !���
�9k6M��j�Ѥ���?�+O�MӐe���'?5�O�B���8� �H��r��E�#Q�R�'�*�X��
6^5x�Zw��E��p!qiD���`CO?�A؀=F%h�+�{5�8�cm-?�⢙5Z�*@%�Ӄr�ʬ*�16)>�)(���I��ፀ�@�]�E���$�;�b�'1�>�ɥu6`Q��螡+�`4�CC(odT��j�D�z�M�T4��Jc�
'ML�DR:�'r\^uCg�F�p�@��QBN9;v�L������'��R�'��l���;9t�99уV�F��@r ���?.�@e�	#O�m$+�"!�b>�*'i9�����֜�p�ͭ,Ǫ`��5||�飌@ �
X[j�w��`���� �g��[�'9��*���˶�ũZಐ���i��6��O�)Iq
�O��I��f��O���Ox1���L9��d�Uwv%�s�.D�2eh+mM>Y3'kд8�h1�T��<���'�M����D_�b��a�ӆ�"���ա6I3�HI�J9@m2���OF���O�q�;�?i�������L��2��YY |9x �r#�r�5�9)���0�`�iĄ2��j5����&њ ��$[ ��`A�N	��Ph3IďX/��9э�S���t�U��5$�h��l��Lr�A������O|�O����O\�\���W�",YKV��th����{�<�Aˀx�@EX�!�/}LΰA�/�a�I��Mk���ė]��l�ٟ���d6�a�b)�*K��@�6GU!/���	��r��� ��ǟd"��	�gZ��U�y�x̻[��<CV��>-~�)g�ܚ
OLц�ɦ`8���FA�5��aa*�5FXY� �6<Ӯ$��#�p����'O�噦�'���|�~�D��5���x V���Q�H#Ֆ��?)��O�1O�!3���+�́󲇚(d ��w�'H�7m��tK@9@dl�E. �)g��k`-oLy�jM�3"�6-�O6�D�|�Q	�?y5(�1{Ev�Z���%��Hb��X�?��}5ȱHM�Li@��'��S{�d�=��E	���*K�)3"�ɰ����.ePZ<+B�Q�>cq�-�>!�����Ⱦ��+_�8�n8`V�/?r�埤�ɬ�M;����'��D��!O��{���[~��b�b5���?����&?���'s],9!�D�`���$��^�'a�7�[Ѧ��|j�!]�2�y�++c�dp� �՟����N��Fy��xP��렦�!� u:1lԃ�ybj  #�.�S�,íI���π�y"Ǵ$
��Q'�M>M��x�d�C*�yn9n,V9�W &O$	�����yR�5E��)�ϔ#xU�귢�)�y�T#!T�¶k��j|��I������|�C�3QG&��aT�J28<b+���yMNe�XF�?�(���C��yr.W*#O<1��O�Rj�y����y"h�e�,y�����}aԄ��[��yb,�*QV�I�'.�t�4P8jм��>��C?���D
��f*߶Y}�<�g Lb�<���"���Y��,Ѱ� �c]�<yq�)AH���p�-/��y`��\�<�����V|���]!?kt���� t�<��A;Z=\�UKÝ���z��o�<1Q��m��q��˕ �f�;U�d�'o�����˿ss�����RXK����r�!�ߗ�cA(W�C��k�\�p�!�dD��t���?"�(�ReI�q�<��l�&���� �3�d��'�h�<�U�L�=�ؙF�,-���O�}�<9��օ%��-�RYae�W�L��-p��"~��F�}�
xy� A9]���P0�yB�_�A�rIr�!%�����GB��y2�MZ�x��쎢z�J��/���y�H5o�� s�D�'s�����\��y�I%]�dj@�kj�V/J��yb��1t$�ckʽm�Ј���:��$QV�|�P<S�"�	��u�ڌ��D��y
� ��t�HXu��BM�0����"Oʅ0��B��rt�T�#!X�K"O��S�ˆ8D"`�92i�p"O�I;��T�`*.X�RB��e�b�BU�'�Y��'�B�AtGݪ�����.m��K�'<E`�L0?�H1rp��
t�'B9�"�	+��M�'�^+���'O� ��N/Cᮜ�1�$^�he��'Z"([6�->&p�!��'[O�5J
�'��EP��P:5p1���V9j��I���V��Q?��p*S�(Pʌ�� �)l�hAY�L,D�@G�vtE�`Ē�^Ϡ�� �(D�XzujQ�hag�ޤnID0�dH:D����ߧL �E�e�H ��t�R#D�JFi\������v���&�+D� ۲�W�f~�R��C t��A{��O�h���)�^��) æ�b��ԛp�ʃe��h�'3 a'n�:|�x;��(_��m)�'h��h�I�+oӺ�(UG�#S(�)�'w�|"'���Z=K$��
D*�4R�'u�h���t{L����g�Zu8	�'�~	�!G�B�X=�� K�/�l8�(O�l��'*(18�G��.���˘Q��'���jq��'?�a��ΘkT�xP�'�nq�DN?���p��i�lR�'���k�Y�V��X+ʨq�'��b��x���Y�O�d@��0K���_���ʖe�'v�
��F�xF�e���x�"��7�B���/��`�ȓC�d��2ł1_�F�b׃Jt�܆�RkfXXKK�@�̭����5Ai@��ȓ~�V�1a�κ,|n���02����0Y��*�N�&)�:�#�$��DF��F{R�)ƨ�v�a���1�)�d@|�$�[�"O
�P�!�#r��"r�F�>a,�*D"O�D�%��˶���O�LC��8�"O����=�����U0.y#0"OlS�i�(W�yb	O�|v4��"O����)�
d\Yj��ӡ��(9��'`�Z���ӧx{��S�	 ��i�!�7{L*Q�ȓuو9;b$U T7"4aN������P���8pl�'K1���荻g.�5��m*�e@��Q&"�ũ�AT��,�ȓr���*��8`�l�h�9_�^���n~*�AWm�9mP��8��6+oN�'J��	�)�B�AE�ޑg���!EC��$�P,�ȓR����b�̃
�}Q�IƮ0��L�ȓyu&t�G�Y$f�*S�)>6�Y��%��;��3e�6�3h�0b.b	��`�pT����#�IB�Z/y�(�����I����nT��áă-��ݢ"�U� �HB�	$�D��J%��`��N׹<>B�Ɇ)iR��fAɂ��,+��WH�B�ɝJ1�E P ����`��f��C��1.V�0�	�-��}�7�P9=>�B�	�C9�� F/�#ת��%�8c��=yt�q�O���C*׎g�¨�%�J=/���1�'��1阩Wb��إ��%��,(�'�X����4XqJ�B6�0[�C���y�mO^�`ܓQ��`�����c��yb*ޖ,4Bp;b��XG�љ�燭�y�D
t	0hpMWL@h1d��?�`��|����Ѝ8ӌ��T�Z\z"�4*�@��%D��qԥ��v��0�(WxD`��L#D�� F��l�B5�B�"�B��e"O�XB����~���y֡�(&�����"O�A��M��[� �Z4â:@R{d"O�0�p��=v�Rۓ1H���\�$���4�O �:��}F�1�#���N ���"OR�AْN���ba�}r��[�"O�$�t�]�af:���oâ"ͺ�ȣ"Ob���J�WF|���&����"O�в�����B��	�t	�'%�O��Q�O����M�{uRq�5��9���`"Of	�vGԧ\Ob�Da��O(�#A"O�U�A�{v֨��
K[���Q"O��SnF�^�t0ip\�-�ٙ�"O0�#1+��0��0S�TI�6xc0"O�(y���F���5�Ή�,y�/A��~R��̓2S�H�"l��L���q�I�<1��CIX��#�2`��mq�f�C�<��f�X�1AW�T�!GH����<!�T�*����X `<��H��Iy�<�Eh�gq��A'�8����_�<���W<T�L0�ؙ�F��s$X�8H�
3�S�O��)�
s��p�F&M��xa�"O�41ăGfl<<A��L5?��L0�"O�*�L[�bw\�%[\��"O��iB�OMl�ɖK1|Q^	�"O���2��-L �C�ˢ2��Pd"O�8� �	+7# ��N�!H��#Z�p{Å;�OhY�1�5gp��"k��I�n��B"O��Qf+!�Z�j̎=�Hy�"O,�AcK�(g�&I �	Q�&���"Ob�v�'a|�Ԡ3�mk�V�C"Of	r�Ҵ$yL���ԎL�ftk��',����'l���wcN����	�
Y�k���'9bA��KQ� �t ���q״��'ڠp�cc��,z���[�hܨ��'��!8&�B��Ђ#xhB�q�'��cυ�i��8 �\�E�>`�'�R��ơެ"��!��f��k��DVk�Q?=�G��b|$8 �[�^**�P�(D�jG͎�4m�\P��/i&�J�'#D����S�S����fE��H�މ8bC D��ƅʖ'̝����搽��9D���d���,���Y%B��d����C7D�,��I�5kA��ȇ���So6\���?)�"�o������&�ֈz�.m{�K��C��M��2D� )v��1B�LQRk#�Xb��=D�\H	E���(cgH
��ti�E>D��Hv�I3�D0x����:8¨���0D��C3OQr�~�A���0`���b.D��paԳALj�ᣇ�	^H�Ja��<Q�hPa8���H
0iE�-�����o9>�)�`,D���hV�4�LT'!��2I8d��(D�F��+�誢��*qH򐠡-)D�B���X��Ȑ��_�	�ִ*��;D��Zw@!!+�݁�K�QP�䉔�8�O
rc�O��"$�)RL0Գ�$ʕ,��qR"O�����+y&��0��b��ɓ5"O��c��	�	|�� [<a�h��"O�-���W�}+�&)ֱO%��x"O:�Ie��&��G� �@���"O�˙��ĭA��U�����I|Ɯ�~
�/L )n�}�`�X �\ĩ���d�<y �E^P!�U�D=�%���2T�k3@	sEbC�A��G��i�0D�� �m���ӺB�T�Yr�U�N��M`E"O:,��*�nV|QE�/rDXkG"O��x"�
�l���Ϝ3`�R�@d�'=�]����2$L���ˎ[SL����ǰ!�jh�ȓg�¬jA�J$��B�#n��ȓDs�3�?P�J��F�Sb���#	d!H�);2��am �01�ȓ"���
�3̚l�m�QK��ȓX���,��(�zD�	�b��͕'�\}�q#&�K!�#�dk�_��R%��9�<l�Pc=]���Z P�v�T��&�` �'�B H�Jð�����J�{�������ܮB�\��ȓQRF��
�,��U:���?m�҈��	�,��U[L-( �� ����ۃ1uhB��n��p�Ɉl�(�@��'m(C��52
�B��&k�h��jGzA\B�ɼ+$I�/�%g왠'��gZ,B�I��b�1C�J�-.�UBE
]�H� B䉹{���!S���{�ق�l5B) �=��X�OϾ��Q��0\� Ӆ�ј<V̔j�'U���)�zT�bb��'6p�Y��'a0��ܣ^^��pc?,����ʓEt�X�A�Y�q�Cab��pD�S�<������8Dt��_�D`C�Gj�<����'���rT.�'wjv��V
矀��#4�S�O����GT#��%[RF�Yr�a�"O��aII�w@�"¤N�8P���"O�%�5��A����1T.�r"O8��R�
W��S!O+��Q`"O^p:��͍v]d�:���2�$x�Oz�� �YtAсA�.X*�P�A�O��'�N˓��1h�+r��"��'��T
9}�x9��ɗ %a@ �T�]RBhB`���'"d�!D��T�Lş$M��	�&�O�I�Ad�D�#żJ��1��䔻6�d;o��>�<�֍%0F s�j>Y:���TM��B�L�^�l�i%*�HDY��ݟ��|��X���׉	.n�v%�Sy��'�a|B��0�-Po�=SD������>YfV�`� r{R�xW.��S��]n�dyEGy���'��[>e�����T�I<\����G+�*1��X��{�|-�	U�*	k�
>#=���T�W�o�04��ݟ.c>���oW�+��U����K����gm�T�AO�.y����n�}p��h���H��Y;P��V83o�&s�X� �'�(�����?9�O�O��I�_�1�s���F�B6B��7u0��ȕ?Ƣ�y��*=$�=i�ӻj� y�'D�f��P�����������ɶZ�hi	4Ğ��\�Iܟ,���?�ݱi?4т*�2)�0��\[�|�
��M��*%��76���gK'F��� ��'��`�1$��<��hH��խ�V%ږ�&.$�X��#�]n1���]F�U�س`L�6A(�)�iK��'j���?Ɍ��s�tzǔ:Y[4�з��:�p-Z�2D��.)r.�*%���&�nA�d �r��=��|�����2J��� �[�Ei���@Pz`x�͉s����Ot���O����O��Dk>!��A�:�����Y��0�w�$Rd��>���F��0�� ��$[96�L`�"�
M��0�#
�k3$�rP"́qD�)��"�3Wl`5�Ou�'f��.8��B�o�PI�,{������hO@#>aB� P4T�QSZ(ċ���_�<�妆1�@�j 4�`����\y2Dr���$�<��o��"��S��xͧvuFa��Ҟdm��KZ�NsB5�	�#�.���ҟd�I�^�eA1��W9��ئM�-}s�������k�)2 �q6���H���2g�ɪ+B�QH����$�I)�-n��P�Zw�-9�'D3�0�QؔX�FX��d��%���'1�rT�"G�3*����Œl�W�̇�	:4�݉h<���G�К=��#��'�b���4bTAY�8`$�&oZ�z�`0�'^�A@��'[XxVQ��O��D�'�D�����z�� (Ι�i��Dac�'�,�L��"�P��T� 68���F-��c� ,�割��\�b�5򜼃��Շ8V�)���KO�O&�����:� � rf�"O��y�'}n����?a�O�O��)� ��{6o���QB�8@��}�a"O��C��)u�`������T`C�퉨�ȟ
Xs�H�H@��ӋI�F8��V�x!��(�3�����u�Or8�D�/¬\��G3��S1��{�(�aV#̀J��t��	��P�2Î
�$Q���TT*���sۚ0�Ub`E����xQ�ȓ_��1y��I-h�d�{�������ȓ��-@P.��h�|Ż�
T�K;��	�{���C-^V�r��U��t�	��0D�!��#t�,E��皩~0n�x3�Q+�!�$V�&T��@'�7i&`QfC�z!��5 l�{�+"h�Hm�¡�7`!��T�Ppn�[\1?@�� �@�)Tџ�c�@���MJ>��E�k�jI2�!�/.�ր���;��d�O��D�O|�H�V�c�>�9��ϵ�"���)&Y*���(مY��< �哃0�8�8��[�Q���ɕ�`�|�1��W�Ҿ1�`K�i����O7ð<	�R�#�*d����Q�֔��?!��?�������N�]�tm�
(��p@��&�?��������:�dFд�vLg'uV�K�&�O�E�'u�3�H�F.}K�d[�_lT��*O@���Oh�%��o~rȕ"a*քQg�@�B�z���=�0<Y����>=�1Z�������]8(�Oj7�5񤉿��O�Ը���$�v�2rg�L���O���Hh�O�s�l��&���i�rM��;���@��!Dt0��'uH�'`T��K���K|���6T��8+ ��!pD<<r�'�����yr�}r��b�::c�m�4�!5��(H��J��Vj>}!�~���_��̀g��6���ñ������!}��X1��T|K,�X���@���!���Ѩ�O�a��>A��>9���R��Z٦a��g2}x|K��)U���#�<�QY�DZ�O�Ȑ%/�w��	Q.�8d<2�������2}*��DD�M��,]^�������z�=�,�9������
kyҀ29"�'�8 )�'1�dx����Jب�3�����'+`t�{fڔ��9O$����O�p��\�.,@���N�#�'��)��I�I��|���҂���a
'/�B�	�^tcD��=y�ҝ@s'� [{66!�	���Oy�s�
����D�w�>�s-�]jI�r^���	QybU��'��S�iB��F6r��J�
8A�1'��D{��4�N�W,�%�t�6��Cfe:�y퍩[܊! �eQ�[Y�,7h�!�y�� ^��E Mx����Ē�y�BÚN�vY"%i��F�mYc���yb�,8��#��WD�Xa����y�h�@�ڤ �S�V,�b��y��͵_���x��R
���
:�y$T>z���j�+;Hl|�sE���y�!�=BF��N600I��y�E(qF<�A��Ԗ+��<��	[��y��^wJY���L@�h����y�"ߤ+at��")����k*��'�r�aUo��M^��@'�Mvx�7�X�n�{���2��a��B�"�VA$���Ӡ1�M�G1<Yr��v� �(s�����WD�8!���ɧ���<�p�ːkJ(	Īd�&oD���$؀��iU�42 -H��-�;ai��;� AE��?9�n��u���-�
�OP���׊P閴[f�p�ĥ#"OB|T� MՖ%�C��)zV���"Ov��!��Av���ʑtoN�R"O8�Ys��c��uр��9l��P"OZ�QM '��d�q/�R�"O�����L�GT�(t���]9����"O�D�4&�4=��J0�F�:<DLڤ"O`�S��TM��d :%�|iR"O�)��9[ab��^y�'"O����DڿqU�,z���hr� �$"O�ev�	�ZӘ��Sb�-Xt=&"OvȘ+«:�R!@B(�M0�P��"O�A�Ri�b�nq��^3k,����"O� ڤ0���8��G]M(��3v"O��aU�C37'�P��&�g	�R"OP��v�
�,e6�"���8Uh-�"OT����@���W$X�BG~ś�"O���LU	I6���fڜ<N��"O-���X	]�t��&D!di�"O<0P��r�^-��Z�~�@���"O�|��$��*��x��`�����"Oș������[���p��1q�"O�Up%�<�H���M�E��	(�"O�����T$7���Ō	O�x���"O���a?!};��Y�(���"Ox0b��T�E�̄��"��R�0k�"O��@g#L4Rh��r��E�x�"O������?!7��E#Λ�v<�'"Oh��⩇*u����5�޽���"O����N�,�����bMk&"OL\;�CT#�Ɯ:ń q�q6"O��Z6���X���Z#N7}ߤ�k�"O.���E�dI2���Z{���#"OH$�H�
E�Mr r:!s"O��
V ]I,0�!�V�]Bܲ�"O2�z���<o�dIPlǑG�\:�"O` �K	/`S�p�®yE
|p�"O�0��)2@ %1���`>���"Ov���㍭C��ј�ES.)2<�B%"O�@�F�v'VQ���%9����"O�y{RO@�W$�1�J!+iD��"O�H[ej<T��ى�b�
FPx]HU"O��SCI)
�͒�G�@�D�"O�9#�KU)���Q(�b��,1q"O��[��C�G�("�Ӑ,y��(�"O��2���%A!�D2@�Zj�}��"O�5xG�ʺ�|i�H[�xZFXI�"O��@����r����"��&Cl�	�"Or9t��P��6 F�=	�#g"O�DC+�%M�t��ªr��3"O����ؚNDV�R�L�k|���"O4� vG�
a��C��(�-8�"O*����J�(�tK��Q�Pxa"O�E��ö*�$�b�ͳpU�q"O���V��/o��#Dm	C9\i��"OZ`���U���XIa��q8d���"O�XKD� �|E���G9@`��"O:Ј�ٷҽ��I����"Ou8 )�9�I �T�6�
���"O~�JE��6\��5�R'D
j��"On�ʤ�28~��k��J��Q:`"O�A�7�ΛU�:4�9r�N�+�"OfQq K�=,`��e�nLE��"OPIڗ�6�" ���?OҸ��"O쩉�KB�uJ�FCR�*�z���"O����"֛l�yb�AA?C����'"O*,����S���0�e�&.����"O��i6Iɓ\�J����	�w�9E"O(U�7"XNqE�@�«Igt��*O���P��ky�0�Pc	.*�j)��'��](p�Y�E>���!��&Q��'�������Ph�a(	T��'�,2�+�U��{VD5��A�
�'0^�o�KJ*�臷Z:t��'S�-K�\���2��%)d@lP�'+μP�h��q�Z���	c�8	�'��,c0&O���b��Ǯx>����� ^�2�d@�l.:,+1��L�@�s"Od���Q�Y�E�AB�
' ��a&"O��J0l�L�6�G �NJn䃅"O��-�)�"3��"Or0H#����`�@!��jdc�"OJ����D5��I��#m09!"OҬ�T�n�ȉ{Seߎzl��*"Ottx��̢^�:U䐧kK��i@"O��S�:w���EDZ&��"ODYV�ǳwF�̪��טLD��P"O�9Y���y�r�"#M�qH���r"O:	1�ʊ2H�>P!�@
&|�p�0�"O�)p���J(RR�Ӆq�Z���"O4�Ƞ�>#��cEȁ�(��-y�"Oܔ�M�Y�41�FîF�D��W"O���1[� ���G�o]~q��"O��k��z<��b`
%_R�0+�"O<�:+�+tYX�@`߭OFaH"On��9e�>� ��N7.*��p"O��R�R�K��t×�"jN��"O�y�A/[����y��Чs��1��"O2l� @UWҾ����r�n�W"Ot�Ң'�!��S�/��Qs!"O�\Z�'�X^ܴA�iv��""ObŊ󎐷E�R����ǼMkRu�q"O�iR��'L��d]���4"Oz8񷮌�A ̼1�.�
�H�6"O� ���vu�����7x�e�"O�z�YH�mX%����D�*lj!���~��m��� �.��k]�!�DÌaF�`(�q�~�3g��c�!�$7� 3�̈́���xWҵ
�!���^�v8i�'_�j�n�`/ , !�6	��cfCL)>���T�Pc!���&g���2��;}�sd�]�!�D4\�����ggp<ӣ�W"A!�$�(J}��œ"INNq�.�=1�!�T�*��HXdL�X9�h�u���!��'�
,�s�ǌ_U@��A9(�!�D��X`+ā��R�d(k��	!�$N	Q��ŋa
J�;��i��/�!��|T~�c�_>�\��bc�w�!�,F�B��em\@�x����B�!���rd����9���3@��e!���"Ek
��2���;2/ӰI;!�d��B���Md�&Yh7��!��ѱi����A��8I��"n!�D²@{�9���"�\i
���6�!�.0�"%���M��R������W�!�d� ��&�.zR!zR��*\�!��ü17�4Bi�9ؾk5�	~!�D�.p�-�pE^�'2��B�DM�=j!���R���W�$��V�Uj2!�Q,�-�Ǉ�_���!�d�48��Ą��b�i��ؽtE!�䋼d\T�s"���N���,,[>!�dӷu{�����VJ��$�wiE�0^!�͗~1^����06&²�W�i�!�Ė�.nzAQp�0}�F��%=%�!�d	*0��Fx�r������!��A$h92�A�4MT�"� �N!�'i0���T��NU���ϖL!�W�=s5Aӑ#���j@�A?F��$ &R3�,�5*8}b�E��#��y
� �MА��"Ѭ�)�ޜ-o��a"O�*`޽3P]�6$�(k����"O��BRHۿ6��А�@"aX��9�"Obl�Sc�434�8�g�?W�V�҇"O.��aHP 7��e��$���IA"O���hP��H�v�dyڲ"OPI���(�\��#�	J�j8 �"O�X{�	UK2I�$�� ��ܘ�"O���Bc�w)da0�� �H�1g"O��E�q�yQ�;2���"O�����1�����-KkQ�"O`�����L�<����"Ob	����[�~$��Ā$�x	�"Op�r%�蠴���n{�@��"O���1b��#N��D�Dr|Q"%"OV�Hs�N�BĤ��Ѡ;Y���"O>��`�?K1�dfN�Yv�Q��"OԼ���׃=�"�V�}Y�	z�"O�H`Ģ@�~�y���[ N2�D"O,A�`Ԣ68��D�V,QX�"OF�b�kA;Y֘h���(s��A#"OnQڂ)Ȃ\��D@���d�b"Or=ӃF� ��X�!��|��xt"ONY��ٳ\`
��b�;
�M3&"O���� ��-1�ӕ������ �"O�L����<A�XɈ� /gz��#"O2�5M͕9��X� ��?.W��`E"O�����=h��.W|>� ��"Oڐ�6 � 	�EyBL�K���"Oz	��&��'D�Tö��b/�Dy�"O��04)��Z�� �JX�:z�&"O�虇k�-Csx"�k؂4�Z}�q"O��z�͎+y ���`�,��H
�"O\���EN!`����I*Dt�ED"O,e�Pf--�6��q��?y����b"O2=�$��ѴxF��W����d"O*�OL�b��k�JJ��>ԓ7"OP���͗M\H�pd��z;L�2"O4�����Ú��aS-R7X���"O����E68�YVGE�@L�"O�����Z �������t
�'B6���L �N(C��NުH�
�'������� 1��� 11c@��'� %9��S��&�;�NQ�*Ϭ��'�r]��$��P�����$a�S�'vȱ�*Q�#s�Q� !3gX(�
�'�>�q�Ȋ����EN��l�_�<�DJ��i��m��l��Uа�BL^S�<AR)+(�1ه�
��!����W�<�BH�z�>\)��P
W $��jJV�<i%��]5�� �`U�:�z���j�<	����CX~$h`k�>Y!Fu9��h�<�t�6� �Gn	<T)�D�j�<��ˇ�^f���ჴ5����Af�<�R�-lĲi-b_����c�<IdIX>}E@��%CV+P�H�@�I�<aЀ�R˞�k�-N�*²�`P�A��� �&���[��V#M12T$�,
��'$�"LU.M�:����0D�����T�0T �F?����a1D�Ѧ
F�_#��t,�d�v���K0D�(� &�+5�8�Ղ9����0D�	���!� yc��S:p�F�*�n=D� �-Ş�By"!��}:�4�.D�xq���kI*�V�v�����?D�� N)��d�q;���JVbS���"O���F��FX��7�HxR�m!4"Odr�;(`�i1d��8���"Or�[d%�KR�0D���./�q��"O��+(�5�vU�7�۱t�01�"O���'֑r�0�;�m)FW^�	V"O4����,�Y�Y�"TX � "O�Y�wȒ?w:��e�7�#"O>-��j��J�B�5��P�S"O�T30 ޺(0֨��� u��W��yǑG��,��͑����QL],�y҆�.P��R@jW�P"�BB��y��˰P����ٚ8�R���_��y�F��//>E�p��&^�n�a!�K�y�F��Xt�����סR�L�����y2�\�(Ј�Y5F�Cײ�+�����yB;F
ҥђ&�'4�aW���yRG3[�T�����_Qn� TB�&�y�d�?6<Jy%!� 41�6����y"�F
�����e �8��(�y¥�x�~��QM�
)����	�y	�P]�e*� т��I�y��=�4L�u@w��mU�C��y���xk��A#F�����/'�yR�Y{81��_�^������y",�+5����ǜ�u>�l�,��yb�_�q��a�����k!"�;�y"���P�f��&c*K��0����y�����`K�͛'���e !�y���o�<��h��Δ�B/�>�y"�5�[$�m� ���@��y���X���3B֋:� �H�(E�y"��?~���V��0<��q�� ې�y���MAv5ZS�E.69��!%[�yJ��a��2�(5�L��fT��y���?U]r���<�`��/��y�j�s���C!$.����HU��y��9Z��Y�hɔ{����*[��y�8I��]0�FF�Iy��{�ְ�yr�E�E��U���0I�`�h����y���)L�Ơ�'E4�.b@<y[	�'�h� ��Ո�p��K� A)H	�'l����F>\��`�c,�+�(h[�'�lɁOܼ+�T��3�+����'� �x� ���BxІ���7�l�	�'��|�g�!cz�ɥh?3��2
�'C<Ű��A�`
���Ԣ'�a��'��ѫ@W*?�B)!T��#�4:	�'ղ�!�W��n��a
�lL �'�:1��Hn�;W� ��I�'�r1���E�Q���P��\��I�	�'<"� rDU$Y}D}��ě?~(�b	�'�<<rG�� �d��e8��l;
�'Y� `a̛�^����h�Ҧ ��'��6��S��ѐD"6-�̰	�'x�K$�OQ��
�d�*)��eb	�'/�����X�F\��"T�K�X ��'�T�h077��s�A�4K�`���'�JaP-גI]���s�¾$H�'��x#�Z?] NX`Da��uU
��'0�<���HbUH�jȨ#����'�ʗf^� �Ti7�ZMm��0�'#0Yx�@ɼS��jO�s���1�'�,��Z5@p�)qD�0[�α���� z��Cχ�
-�ِ2Q9���ن"O�S��3i�V�PU� F�
��C"O�uZ�j-A#6l�f+�>,��"Oʍ�c�5k��P�kΗQ�	:2"O04�B�G�(!{1ʝ�!��h"Otd[j�7�R!�)�!+u���'"O���
9p2p��Տ?Hz��"O��pEC.:�-�/&�����"O����A�5�8BD��{��r�"O
I��d�vU����n��:ݠu"O�l��B���A�m�Ln��A%"O��E��yE,��ƕ�[_|-�"O8DZd�H=���r+ě&x��z#"O��� Տ*�x�)4.Mp<!��H�]	�@.��t[��QY!���|��y�F�|�
�2!U� C!�SSZ���@��(� F�]�!�$�`�� :�ג(���H�;Bf!�Q0@j<���T��Ab�W�cI!�Q�iRi�"�����ۊj�!�D��4D\lD�a�>���P�!�d�9C� u�f�Y�~<*Ű`H�??!�$�w߮���K��N��0h�%%!�!S~@�Z6o�p`
����7!��0��)�'Jd��C�N �$!�d��dND6g@�8c�Pt!��:sO 4#c0R� ��3O!�D܍.��ɪ�%�x��p�ӶW�!�˓|X%1R��8e�@��`���!�dR8d�B|hu^�d[ �! 
t�!���
;Qr�H�J ~+xl(���)|�!�D�=J�zX[��ɅM"��k�D�!�E'i���	�(��|�d�
ʓ!.�!�$ ��@,�T��+�d��A�_�T!�ɭOo�Y8��>PXT�T�C�.!�.5te��L*�N�(0�!#!�DP0k~ȩk�d�01���'x!򄃔T$��򇠈� ��90�Aa(B�+`Jt��%�
a�$����'�8C�+K���zvH�(l =�3�C>C�9&�F-p�߄?���0s�÷>�C�I��lżh����'/B�3ޔC�	�{�����
F�VR�5{��¹b��C�ɓ#z~m2%��">�����c�+NlB��<i����� �4c�x�p�jY�{�lC�	�d�n<2UiؿR�J� DV6C�I	>�p5�VO��%X���E�x��C�I�*r�(��HBa����՛BN�C��F���UW�L4q�`��Yf�B�	�u6r�2p$�7+��E�y�^C䉪
+�y�C0���kc��O�VC䉴w��)R!ה���KA�Ұx�bC��5NM��%��?~�h@��A�4C�ɝ6�h�K!��22xtpi�����C䉙pAB�j�ʄ$�b�&B�m~�C�	��x�t�<h#T�?f��C�	*�5�P��W�`8Q��,w�C��cFr���FG�:n)�G	P
OrB����2�, F�,���\B䉨Kv��zSɛwZ�h�ՇA�BB�	~)�xa��J9 �N���c��/�B�	�^���xJ_ @�$��#D�s�B�	�V��݊E�I�<<����(V=:��B��
0���q����f������Q��B�)� L�j#N�;��@���N�a6aa�"O���琿z�,���}?�Y�"O܉��'�9q���`���F>�:�"O�a0mΧ ������Mkt"O�ň�a��;~��v)ŕO�J�"Op���G�x�8-�ɞ G8D)X�"O0M�W��4QV�W=~��9a�"O��q�mK?j]�IRC.'2p���"O`���c�b��S�	6Xj�3T"O&�
���O
v���l�3`��}kV"O6q)�C�)*��ԉ�	U!�5�t"OH�`bsa�(��U���U,N!�Dɢr;İBrd
�%��
E֌8��'h�eʕ�,2�DHV�C�~�qQ�'��i	�#+cR̸!�zh��`�'�|��U��3�Z9$�m��)Q�'3ajC�ܗ*o�Ѐ��0���'��;S �2�Z`�*��Yl���'��L(�L�.��`�ժ�Y�1�'�J�b��H�p<��Ē82A�	�'O��J�&��G Z�1w�2�ച	�'�̨�S&�2,��A��B���J	�'w�1�dkU���.�t9����'���A��C� �n�Y�A�h�$��'\�"���
�b �� �%��'&��r���h �Y9���Xya�'��X�GnG:��yJϓ,9�n-��'�`5� �=��`IE��8���8�'�8pK��������$p^D��'�T�ؠd�E�e/J��2"O|ez왺2�&��cL(C��py�"ODy�cQ�$PF��ĢD�N�N�ٳ"OD-�%�sR�;Gd�,<Ϧ�""OmK�嘏r�x��A�//�p�@"O�9���]�6F��	6�E	 ��,i�"O�yx���> ��3�F��/m�"Oh����;e*f��S��+epM8�"Oz�['�fNJ�!97�<<2�"OXĒ������kć�/��x*#"O��U��nn�t�S��9$�p)0�"ODܫA��*N�$A6�K�3���"O�T��k��C�����1��4	0"O0ͻQ�\�J�t���7]A� �"O��
�_���y��$0U~E��"O
������<Z����^	 �"OڥK��o"q�C�#=���"Or0oQ':q��	���w=��c2"Op}�%�A�
��e0�J��0�"O�I:�K���0s*�=%�9�"O~���i��)T��5įX~d��a"OB����t^�Q��b�4o��P��"O�U�威�A�N��V�ڜ&�\��"Ob� J/rF����Ms��1�"O�t��F�\�$E)�n�<�N���"O|��e]5w'�c�֦S����"Od=���V�A?5��.	N5�%$"O��ѩ� %$��m�ֈ�$"O���
�R`p#��$dRpL�0"Ov��ڤ_�h��[�2D"��P"O���I*qK���D�r"O��u�_�t��1����y�!�PV���b���3�Z���`��,'�' ������#2��cM�			�'��ؠ5���\!���%G3j��'�h���KN/:��l��,��J~�}r��� �t� o�:W�!��OW.'���ya"O�x�c?�v�QB��/y��"OpqP&�_:ĴX�L&v8�m;`"O>�! �E� �*��D�N??4���"O����X2a�<�@A-'��"O���S�4�r,��]�G���y�"O�<�c�A:H,��6�&0s�7"O� �]d��AjA�S�	�kD[�<A�ʆ
<���"�bژz�|X)r�Q�<Yt�ϛe�N���H_qfIs�	N�<Q��̾9ʅ�BӉ)�r|���L�<��Dݗv	|1�e�ROh�q��E_L�<1 Tz���JpX��a	�J�<1a�P
y3ҋ��%�p�F�<1	�-bCh���G	�6(�\a��E�<9מ0oh�ꗬ?���ٲ�G}�<	Q슉pP�#N�;|�٘�g�v�<I��0J=i@���v�J��0�Rp�<W&܀Swxd��(\��}���@�<�DCܢx�x"�اt�f�i�`�<����lΞ�Q��]�	����f�<�C$&��u�֝'@���%��{�<� �G'dj�Re��{�N��'c�|�<1�^z�8KW�E�4O��+u�Xb�<)�A
�c"df��z����e��F�<����<: ��q
]#Y(d;�,Vm�<���J�[��i1��LV���m�<���7DdJ��5ON��ÒgTl�<�@-�+2�Ѳ-�5:�z�c@A�e�<�$��z�،J��Q4$PH{��z�<y'f�g��x�#�$f�
{!KIu�<I�ѥ&� �g�"_JD�
7 �s�<AQ��;�&B�g��1ZT�r��u�<I���<sy ��"�ʤQ�9�,^}�<���� ��%����
ID�<q��LC���EB ("0��H�~�<��n��݁R�^y�H��{�<�a�@9{�@1�H7i�-�o�<i�h�"Ş�3bc��;�r�W�Qm�<adfҼXJ,y�#�1r2�ãg�f�<��=&�l��l�	d`� �M]�<1��E�?�̜`�C��J��x�IBP�<�1��,H�R'�8tF���IL�<�А'[$!B
ZefJ�rEkZC�<Y�'J�h�����P���ř{�<i4��-h6�l��ˬb�����'�tF��f�ѣ�`�J�x���'��aVϋ�/8`���oNJ�J%2�'���G�$8<ܫ�Ayʤ��'y�(�*�5�ʠ���#��'ULervb�'gA�JDf7SZl��'�4��
j�. �dƼ���
�':� �$�V=|K�53�.k�Mx
�'7x��4$іY4��HE.D7��6"O�UJg�ئ J����.ӽ`Y�%�g"O��c�Z.L��}9��8a-V:v"O|t!�L�
2V8�CJ�*(YK�"Ol�T�D�$�ЄO/7��kd"O�A1�ŕl�"}���Y_��Ȩ�"O>�p�_+��黶a��[�Z��E"O,3�%C��>lӇn��i�Hy�"O��3����M�A��(���`b(D�4Ђ�:r�х�'͜����$D��z�J>G��z�@� �h�Q@(>D�� �ؙȅ+T�R'�\d��}��"OV�H�Z$7�I8C�AG� �CV"O�D�����3���^�LqR`O��yr�8�u��A��i��0WGU�yi^��^h�S�4�<�se"Љ�y�	L�w�v ��:(�vI��D��y��}.@�#���6c<�
t�L��y"�W�#�<����10��tx�#�?�ybc\�ږ�x�C��~rp� '�R��yR
7O! �	eh��$ܞ��㚡�yŋ\�t1U�\�mY�xhA�N.�yj�(���3R��8_�P\�0���y�m >�F�a �+(k�I��W��yb/��s���h���)w�p�B���y+eبؒ���$鎬�*��y���k)���E�A\�R⯊'�y"�Fr�+5�Ӟ#��y$�Ƒ�yB�ݵ{=d(�AN��	[`��&⇃�y2�(9{>�q�D~|��R6$���y��!l��9�'�q�~���#Q��y�J3��q�-A�t��U���y��V�{�
�ѱ튾i"���̑�yBFނX8a�6BC#W����&cC��y"LLSL�|�B٨M;���Ed��y���r<��W 	�I�!��m߶�y��
;9��Q@f�D�*b�[t�«�yR�!@�ȰP�.թxt��2�P��y£	Q��� 6���R��0�y�� 0A:���ڒxZ�q�S �y"ō-d@�%�a U(&!��W��y�e�4k�zȳ��_� �����:�yB'�\�(��F)/����䐑�yH:HD�c*[d��1+2����yr�
�,H�1-!	�B�a��]�y2�KCC|��JY��:���f��y�J+͎��Xq�٣2JE��y"���>/�IŎ͝bD0	�`��y��Z�[��c��/�fL;�,�-�y2�߽1вt)Wiѩt,Z���Ǐ�y�����D�c���n��8��͵�y�� UW����n� dҥj��y�Z�
B�ʶ��`޼�"���yr��l��HD�GJ��{B
���y�a��2RH,<_�`�T��9�y�,N�&�0���]~���4K<�y�
�"@ h�nW��`
�J�$�y"��`�T�BQ�B�����y��Njd�X�Eɯ=<�q�����ybB`��	c�J;}h�[p����y�)	�1�^`���rz���$�M��ybgq�H3�F;gM���щ��<C䉆D�g���fcĉ!@ �-P�C�	�D�,���E����->~Z�B�	����Q$j\]��oL�0r~B�	�t�y{�B׽8�t-3R)K2=�8C�	�6$�Q��N!�G�I\C�ɠ7|������7�D��A��8sL.C�X<[�!-\M�@�F�"$C��˟Á�;	���O�8�\l�0�*D���T�]�a�*y�%+Y�F|�!f(D����e��k?49��k&w�8(Б�*D����V�?�2��!S��0�Ȓj4D��8��]bE2�N\�_�H� �7D��Y�+�9�n�٦�7;���±�4D�� �����8!�B�+�D
	����"O�����53XP��B�(��Ƞ"O������XH�,XD$61��ha"O����mQ�PhY	5"]� �d�� "O�,S3B�r=Z�k�UB���"O�)
rbW�TA�<Id�Hc5"	W"Ov̫䉐��> jO����4"O��a��ŮX��	��G�4�t��2"OJ���
?a��Q�#�b�8R"Oƌ�NY�v��I��a���S2"O����K
Gxj��G�r�t�+'"O�hH��]�Sة� V�%ː���"O\"����=� ��r��ئ}!u"O�:w$��/j�l	2J�E�V���"OH�i���2�\D�������"OB�h�4 �� D(M�6q��"O\4y��D�K�^�ⴏK8T�[g"O����O��B�$�:="G"O��9��N�r޸�PcӃ}���HE"OE�B▹rcA! #ԆK�:���"OtqrL8��qb�W���"O:<�&͵�������-���8�"O�$X� �4�  ��I8����6"O�]��%�	dX|��[ah ��"O@@H�g��%��̫�M��%�<�ȣ"OpH8ƈ��F%��Ip)
�h��y�%��4��l�GO/��ѷ)Ϩ�y�F
&�ycd΃3��\t�=�y���h]0�j%�;ؐ+�O��y�/S�$��k�F�D>���$�'�yRI�"��DJ�Bɾ��J� �yb" �-�T���&V�f^x�tc���y�á$1d4�Ҭ�.a1|0�c�y2��H�ڴ�%�+Sc���eQ��yB�_�J�ޝ��OOx�U1�Ԯ�y"�ҍB��,:���R��}�a'J"�yr�hI��Pj�FD��ғ�yRk�#g�P�тų?6Z��Q���y�#�q2�7ʝ�6�z/�yŎ�l�(�6n 9P���	��y"�޺mq\Xi	�3�H�� E�yb����h����"��|RP����y���6�b�bk�!B�����8�yb�b�H9r�D��T�NC8�y���X�C��!���
q`��y�Ş0e� �h�"���F���y2gͯ.�}�BkQ�MЅ@����y'5EV�<*G�Oz��`"�<�y"Ní�
1��4D	�Ɏ�y�m�8t�8*ڔISg���y�ŉ w��冇 �Bqy� �?�yg��;�  f�G��!Z<����M>U:���<�<�������Q���!�C�Bm���0l�=ۮ�ȓ+l��Tbw{(��,��~��ه�ZC
)keGJ�j�����JWn���"'���s
C	{*j��"��^dxX�ȓm�x����0a8L��,^Z:t�ȓN���(�(�� б�l�4�<H�ȓ<]����	YBJhy2�_�2��ȓr�����B;�عi}t ���@�Բ��9f�T�ٵȎ��\�ȓCG
ɸ�FL[ZMP��X�;%���~tⱊ��_��髐���v ��S�? ��@��

�U�a��b���c"O�a�ȁ�9B.)� 럆�Dr�"O��+B*ˀs)�T����!�"O�d��M��QN !��� u@�"O~��3m0��YS�΅�u;&���"O��0��έ�ծ�� 9�"Oℳ�D��!�b�*&ĕI�0u��"OR��GB�n���C=�F�"Onl2#��U�`�t� z��z�"O��K��ƟߤY��Z�
��i�"OL1CV�I�����ؐ�2��"O� �fH���Di����hq"O��Ip$GJAQb���=�<h�"O��`1�A�4�0����*w��[�"O�X��fM�5V��RC���zu�"O|�	��I���D�B���1w"O0�s3��|�0��'����4"�"O�-���*2��'e]a���;�"O�H3�b�\PT$�WD��F�~�y""O�t2���O\�@��(/g:ez�"O"Y�� ]�"`x�2H���<<S�"O�=�H_�E_b��%b�<t�
-kF"O�ň��8	��U�w�O'?�&TI�"O�t�1BX���ihF��	 ����"OͣV�VG�БǤ{�|pE"O�]jrțP+x�s�O�4���G"OX�@�SVT(3�&�:>��0#"O�<�櫆.�Xps#T�!:�a1"O�������n6�Y�F�P�j9����"O��h�0lB2%����7� m��"O~9��k�3:$� r�% ku699V"O�|�G�ޙL����&P<>���p�"O܍x�O��h��F&eO�"O$���Y�~�ʠ��L�:��	�"Ox�أ �;��1��	z$X�"O8)���)b&ĢO�1	�%�"O��Y`�������oG4#_���"O�,��A��8n����5{�2�q5"O���Sh޷v��@�%떋nK*5#"O��	�	�>FA �1:=R���"O�A���s
�8Z��Q�����"O��a���c�`|{��q�nU�6"O� �؅��ARO��s�!�D�d*�k$o7*N��k���,d!�DІ*#np�V��(>��Z�욤~c!򤓀1�\U�Kÿ
4 �뱫��FU!�F�@�R0�SΚh�j"jL.F!������â�Ǌ9�LE�_�2���R�
4�Az�|�a�!�ine�ȓu$��ӷa�=	��šQ�˙r��\��;�`Es��V2����Id@}��Py��p%BӅ1��O	������4m���; �5�c�ta�A��=8X$�w�0��燚��j(�ȓSߌ�R��5wb����F�4���j���+�ǎ6��pE�N�n�ȓf��{��RZ2>m��$ǂ$gА�ȓ{�xH� Ɛ�X�sb�.��X��/�H��٠z�~ �I_Վ$��	��Q��
�y=��4��v�B���'�:��D��,s&�hW;Z�4��,L���")`hBE�4B����R�ةA&&b�������f����ta�����?7�����N�tB�ń�S�? 済bɌ��4d�`���R��"O���cƺO�2�e�sJ(��"O@hP#��-V$��#�'*�h	�"O���&�g�t��b䈎N�"OvUW��!YP<X���+�d@7"OY%nĞ������0�v��"O:4if -Ee\��4�ON����"O�}���̾;�l������	�"O����R�xeę&����7"OZ��n׀\ab�h2%4����"OD�X���4不k���/G#��{�"O�m�ceJ�!뮤ɢC�?0Xq�"O*�s�@ӄmZ�t�a:�����"O.t�B��: ����&[	5�d��"On����f���ʐ,�E#D�Ɇ"Oj�xo�>C) �ȁl�p�D��"ONiPι+YIs
�p�~���"OJ�rq
��t��գ��-�d�ӓ"O��#���Y27�����`��"O�MQ�n\�^�:���ƃ���"O�TS"
�	Y�^$��ߓj�r8��"O��PFY��m3����r��"O�85�,r�M�E�G$1�Lm�"O�J���|v�����q�m�"O�a�g��:}~������<J���"O�I��+�� aQsA@�1��K�"O�i#4,F<��X9���SJ���"O���b�ƭ4���cPh�J?�R�"O���KX��R�폆,7��Q�"O�u3#Dė]�����Đ;(6�a�"O�DS¤&����| �"O2H��n���ډ��蔄{�9PC"Ov���HӶ��)R#��25�DX�"O���B%<-4�Ї�k붑[a"O�}[���}���a�&Զs\dA�"O�E�ңX8�CҤ��z����"O�ɡ ��ƍ�@%�&]x
q��"O$ �t	qFu!��ru�k�"OX���GKF-� �'a��~{�@y�"OČ!��e����sfM�Lq���"O�`��n��Z81��&o�R�"Ot����'H8�8�+��Y_RTڑ"Oj�ّ��(�����ȫBSFŒ�"O���Æ/h�f�3�ꖶ��@�%"O�d��,ʱ�&(�b*�45�0��"O|!��Y�@��[��ǭx�İ��"O@(
(G#Q�Y0a�X���9�"O�(��
+.�p{Q�
E�Z"O�5R�c?Ǣu��^�2���t"Oj�k�e��d�8|��Oٮj��{"O�Xi�m�S:)i��HT[�"O `2�m�Z ��ƀ33݀uˑ"OXdx#Cܮ3ipC��d�0i�v"O6=SBo59$v��B� _���)�"O�Q���\j歫� B�J�L�8�"O��zDM>9�n��Eb\5d��{F"O�0Ad��%A����2�W�N�r���"O��j1㉕4
�L�G���LJ�"O(�ņ��5���G\��>XJc"O�D+�ȝU�43C�W��PE"OjT:�@�B�$�0�$~�����"OH�p�)N�mdF�� ��0vה]h�"OD��HQ���v�I�-��4� "Oȡʢ������	إ#�f|�w"O� �)��s�2Y�3IK /�2��p"O�����$y��CĈw��y��"Obq�@��x��hȟO��Y�R"O�;`L�?B:T��LY�$���"O�r@�7yR���!�6s�9{�"O�W���i � �,԰��"Oni�E���� J-]:�q"O�8�"-?q��P@���%����'s�i+�,F"`�r��`�W=|�q�'��pSh�-;���!m�.���'���h�<�=��&m�)��'戰e����bҊ,D$ȔdWM�<�Ţ�%_v��V��$���c��@�<� �_#	>� �O6~EN�xPL�|�<���6-�P%�R�4.�(��kP`�<a��h1��%J�@8���[�<��͓�t@i$hiE��@��
4�!�$۹� I6�
�	�Y�a�!�$ ��1E�[_��L��,S�R�!�K�&���նL�Di#Ԋׁ0�!�Č� ���A��vr�Y�JZ��!��s\0�r`L��]c�Gi�/r�!򤉦y�>E�����:��	ɥh !�DR�C����5�L�4q>���(O7�!�Ė�*NZ�XR+E Gk���� R=�!���>+�[!F��9	59�@J�2�!��P4��cbT8������$!�΄t*J�S7L��B��蟘 �!��^,W�p1 C�Z�t�B����W�!��P�u^y�O�y���4ꆞB�!��`�uY`���U��,7�!�d�d ���ǇU�fp�m)[�!���4�p0��JZ@�c�J�0�!�dՁ�Z��.�/1�dd�Q	�9
!�,O�|��G��
@�J!��� !�^�a�*�8a���Iឈ u��� !�DB���� �NR-U� ,V�|�!��sF((�u�]���ЩGD:b�!��*4�|Q ��_�~%B�#Q:!��Yr�$�TC�]}��(�"�)�!�d�$P(�q�Ԓ��`"fbH�9
!�T�)&�)p�	��-5�\�!�d��H7,päS�p�$��A��^�!���#eo��[���:0|����]�Lr!�dT�e����B�;�d˷愵SN!��T���(�;�.h�Ȟ�=!���Y$���!lɨG������Ǿ�!�\( Ε
QK^'2����CLQ�!��PU��XB���<���Ń��2�!�d��Vv�𓒡��"5��ΏL�!���
{�C�$��d����X�!��5��1��՚O(���V�_�Q�!�DV����&�h����h�!�� �Wh��C��>[Φ��Ǩ�>�!�H��܈vM*�z�b`ŌZ�!�D��G�D�V��WN�J�!�dӿw���GdY� u$�t��N�!�d��l��	�ӭSXz�!�˃�j!�$�����e�]A�h��T�!�$V�Rl�P����wS�K� �n�!���u��s���1D�#2�� !!�$�?��ē&��@� ]"�G� !�4u<B%�!���>����Z� !�0c9�K����#��3�(�J�!�� �0����7Te	��� �0t젱�"O�[���3^,3/C�0�X�"O�	��X
Kː\�M�*ݐ��"O <�2%�5�n�pAO �D�n���"O�Q��۲s�d�m"*���	V�	���s�%�6d�6�)����P���4l��]BV� �n'qO,����%�R(p�
3}ll�v(߫Bq��J�Oef�Z�&))@`8@�47HvP����
&���f�ߍ(T��K�A�;�h�'Wm���ӡ�7#�b�a� G�� Ez2%���?I��3�v�'���3~���GS�Xh�(2d$�^9\8�������I6��)ȽKF"���&��h4������9��4�M;��8;^Гp���\kAŗz?1���jM��'�V>���M�����˦�:0�X�K�0��	�in>�[��)`�'��5�t�"�f!R��A��b�?e�O��t��&��D��j��(�NXv ��XV�i?d�b��3"�<	���������#�}���\cy��!G%!?����(bX����Ħ�)G��O �n���M��∟��l�+$��ip ��m��</n����?A+O����H��xs���7a3��Ŕbב��l���p'�� F?� �B�$Z3���"U)TH�<yf�Nyi� 8@7�),O|����S�3�Lx9��;�Ȭ[e��+K��Sr��M��G�T�*�'H%2#<�+گl���3���,�ufC/[�l]kE�ĪG�X���^<UQ� �OK�#<�㎟�,�@��R�	�]KS+:���O�<'AzӶ4c����ßէ����8+�ʅy K�R�FC�B3�ONO���ʉL�|�����<:��ɣXp< ޴d����|�N�d�*OX�ca���F��Y�J�D쐹�J�YX4��`�O���O��D�.����O�����a1�����4��B�Y��DJ
�"R�)sNS8C��U�+��O���1H]�F�V@���3����Q�_�Ҩ��)�|(��*ҍS5%%��	�'�(O|b��'ɛFE�(ʠt)�΁�=ۄ�׍+T��m�ԟ �'��U�<�~ZuCъ9̶��G��.�
�F�N��0�S��-����E�������x$v��"�'M^6�٦}�	П̰)���M{��?q��߭ۡF�2��H��c�8̙�cܺ	�@����?y�1m�#�D���h ��\�8P0�q>��d�D�[�`T�P�C�3_�b��8ғu�Ȫu$�4pUj��Gȃ/o�%�Ɗ�={C><с��r�v��eoX�"F��%�_�'�`�Q��?13����i;�RU��2}9*h �d��i�p۱C�O2�"|ʨO�t�ڐ\R(� ���B��B��'j�6-æ}o�<T��0Sצ��aP=!�*���L��6t��ش�?����i�*O����O�7�Z4F�����[�Z��4k��I���_�rA1�,ï6un��g�q��	�|����5&�TPB8�KS	�h��	��M#�i~�I�M�2h�@6����bLq`@�J�����Q4� �H�nD�&��h���֦5���O��l�:�M{���i%��i���ǰI챱℁��f]A��O��(�O�m���(Uo��
1c�eb��j �	�M��i��'���2R!a�ğB��m���ŻfR�,�L>iۓ=�~9�  @�?ݬK0p *X�d2�%�%s�qO�,\ � 7�حsbJpA� �]�$��E4H�{O�H(�/��V�h���F\)n%´�|�'�T��`!�B<�S�Y�/�@�K>�ӆX�'�A�G�?^��R"�x��8u�����P�2���E�\���c�"�?)�`��є]Á�^�8��)@��@J�'`�5��;8��rNXZ(9!"���<_Α�G�	W`�T�ʀ3b�(I���l��IH'�O�``̐���$�%aWDHz%c��!FF(�t�a��	F�IA-PBlв$��8#8���$��� !�v�$�c�3�)z����y���@��% NNQ�,k�A���D��<(e��{���-i�Q�G��ݓU�^�������L��Wn���hO��É��d�a)�Ȓ�����O( �2� ����.}��s4�|��*u��s0N�" ��)��/��|�VX}����w�@�p��<T_̡�!`���?YuO4K�Z�A���]�ƨ��ȇA�'Y�p0JDu@@�3��
�_z�Z�����` �pf��I��[&�QU�ɅH~��C�߂i���rl�>G��]��o�/q��챥��۱��a@D��A�a�F�%ф&T���Naʁj�w���	�K�z�(�*��1�"�k-O2@��i�S�4�A�9-f��(
�B������|1.Kў�F� �$p�@����t�̄I�Ȣ� �#͇.ԮmQǆ�19�(f�,��3=��	yR|�E��65�=�w�"!���挳F��/{$T�˄�Y���d�+���CJU��Z@�q��(R]Q���Q 5}�r�8�T�H�Z������֩} �DPѪ�����P�ēv�`��'��8jv蝚:�ܽ�)ɼ%�b���Ǜ�&ި���**���9�!Q��ܙk�Ӏ%�x��vB�S��;,O�㷆�U���'-��3��dHE#��Ą��D�1�0Q��'��eJA��L�*�q�I�,�*hcV��(x���G��0ɰ_�H��	�J�h��(ێJZ��A��� c�Dχk�T)
���)m@����;O>]��BA�L�Nhv�^nX�0r�o�2b���WNO�h�j�"�<TR-%tU��^�6��H�Gm���O�	"a��7������I���y��xR�2iVT�� ����Z�??u� �4eMYOҍB���wFM�o��L�Viߍs&��'��1�a~r�F1��qG��B:� �"G��~Us�^�]���*���I2����_%g�`��wK��� �&O�[~Tq��Ӂ;ݜ����|Sd�R���S��y����x[�O��2)����3�S�NN�y�T���
��HsOH/{-���d�7kլ�6!��T7�1�C��Fx��'���%��::eN���$A�W��9�J>�E$@�S�qOz�`�(ԋ*p}�S�H�Q�$j����)1M��H!�.bF�iǄ��r�1�g��aК�>9�M�t?����+P!�j�r�bی��'������!���"&�C� E�5�c���Nx�mS�(��|�!�3U�褸g�X/DL����d݇�p?� ��q�D� ��ܝ4���JGT ��'���x��z`���7���w Н��n ^�	��.�T�*���N��#���bC�I��zX𨈏s�<0��P
E�亦��aG�;�h���R 0§T�
�	�fT����9y���x� τvZ�B�I�0N�}�5�ҙ�.��cE�^�	� ç:c�����;\���C�I�P�Q�@e*@7}�����,ݲ3Ox�I�&\Of!I���#z��G��`�8����1~X<�P剘�:=9��[�,��$�	g�D�rFD��P0d�c�!1)��7�p���.[(�P�1砏;�2��A�`��G��  l}�"�371!�� $m�4�V�C��1�r5�=��N�6.#�$:RL׍q�~Xb�cȳ-q����Oꄩ �(.�P�D�ŜA܈�[�
O�tЃoQ�<.��C)I�cb����5-p�d����YT��6*�
��X��ɘU]J=�viرi^�RA���%�'�>-y2�ڛ���������S�N�@Qa�ɞ'�9V&��P�B�8�lSܩ.� D��`2B���3}B��b䄅*���J�8Ӊ�(��>!�@�@�2�pI� ��u��耔�0D����[���gLm6hqǦ�y0�)�@A�F%��G7���>I�I�\��,Uy�E+4� 3��b�*$���ш��=��:�O��1��ݚ1��6mP�0g�y3�E�w��YǓO�UC`��@�ލw��<�f���ɝ�p����'<U(����]6�x�#KQ7eC���W��QH<9� ׃v�x�X�s�P@�WY�<p�50����ő�G��I�Do�@�<�L�C>4�0-�;c{�Yԧ�v�<q���3{t tn�@p��I�q�<�F$
ʁćڵ �x�yAo�j�<!c*�7 T��Q��+&@=�S �i�<���9.ڤ�ӁD)W������q�<ac(����eh$I�h5K���u�<�T�P�x`�ʢNP �'�x�<A���V��9��F	O�1��c�q�<��喞m�F��a�ĄJ�V�8`�p�<�f��6��@Í��Bۼ�j�iX�<"�TZ�@9#AWj��c���o�<�����2�ԝ;�,;.,�P�d�]W�<97�x�6$�Î0^�Xm�FE�U�<	���	#7C^51�z����S�<��E�L�"ݳa�C0;-�ə�c�N�<)�*�"��������l� K��K�<�ǋS6t�^4�&�[
b (�T��K�<Q�ܸKϐ��dǀH��'��B�<1�,ƾ
Q�x�Aj��(�U�Р�{�<@�8k޺l	&B�&1��*1�S�<	�d�	42��1�� ���1#�N�<A1��**�o�U��:7���!����@�YD/ۦkK����D!� ���0�J�?SH�%�7�\�t�!���) ��9��m�=	�<#aDP"n�!�$�Ք��G�yD�c��6=�!�䎌�$dkC�LJa�)��!�O?|�R}JL�b *a�[��!�%L�И���$C���
s.��S�!����5�ѥ�[��UZ��K�(�!�ĕ"4cb;�� �$�t!�dV�h�����0V ��%F�!���q܎��r'J�&D������,}!�
�d����$ș\���C1�q�!�
�1��aA�F�/��a�5��r�!�DS�{G.=�B�I�F�&��v��3V�!򤛖SVDȀ�+�����H�a!�d�	4����BٞfD9Ks��G�!�DI	�"��$
�|�@�= !�$�H$�`�ݶB�Z]�A�6HK!���Z�䣁L{�X�@J�BK!�E9L�L�h�'YuRd�s!�	D��`��a^!qN���=&!�dL�6 !��/�
|��E�Nf!�D�$��iЩ|�JP��_2b!��X��;Pe}aMM�*6��d"O@H RF^�V�ԼT
ڬ����"O�ph2��5�����px���t"Ox��(�'�`���[2TlJ�x1"O(�U䊐*r��K�&W0(�Z5"O� v�����1S�&Y��^�G��u
�"O��x��͠9Y�4�u'�8����"O�����\.>�p'g�<���!�"OPAr��f^D�'O�<Bn1"�"O̡�a�"�")d,6d �xF"O�3��20�&���-&�P܋%"O��P��I�p�H(#AT ��	@�"O4(��bO2&���!��V��(�v"O �If>p"u�P�ܴ"�Ի�"O�D�e��'Vg:�	�%G�Pj�BC"O�Q�f%ւh~�P[�	Ѱ�ptH�"ON౑�b�t�zʋ�C���R"O~����ɞ��T	���
�C"OF���S�z���nY�x�
��"OʘCd�F�x����-�4;lp"Ov�'. !���ŇΎ@���"O� p�'��j��Y�A��,��ش"Ox0)4F�
*.�"F� 2k���*"Otг�,^�s�������\��"O$x���P?#�*@9�n<W�"(1�"O2��P�30��Y�T���{�:��"O|`%�"v��crk^�|�4�v"O����Z �Z���Jſ6Q�%x�"O�<�����r�i&�?J��I(u"O�`�b�.�Z�F�..f� �"O��  �)wSd��%NMj�a"Oah)�$���Ӣ^�	�(w"Orĉ4@�\�A���г.�0a�"OH!�&���]�f�:�A4"�f��0"O61c@e� ,���喟@\DS�"ON�j�KŭtWl���EI"y . ҵ"O�ya�>
w��P��V�y��\��"O�EE�
G�8�׈�A�Э�"O�l�e�^�,M1�1�<y�"O��*O�\<�� �"w2-��"O@��P�F#xz 4� �V�v�1e"O�5�pL�"JNA�g�M�BZ���"O����c�Oml]C��'Z�k�"O���{!U�Q1LE
L��"O�P�wJ#{k�r�ՇB=�"OR�Xڄ
��x���D7Zt�T�'D��g��<8��'D�?����%�0D��X��G1i�^�SAK�$uv�3�+.D�xb��@�nP+�D�*(D<�7� D�(�7��$ \y��8#H���M!D��xA�_��`��ݔG��툕5D��{Bb]�K�$�cV@���w�W��yBM4lb�� � ��>��s�y����\����r��ãN՞�y¬�T�p�SC��q����"i-�yB�#_L�1sA�9c�t���ED�y�e#v�`�Q�K-:bp �hK��y�%�)Ye�<�[�8B�S	@��8	�'~2��dL�%:�����d�T��'��Y�g�>A��2���(U��i8�'� T�%� -3�]��K3KU����'
��e�ӗM4´p%"^�E�Nt��'���y��:1-��˴�Z�,�����'�B�CH u{���$攫�ޱ�
�'���7��$�z�GC=ek���	�'F��ZC&�'oJY����?X��� 
�'����Sk� ,~�-�V��'���(�'à$)ǩU�e�M����0� "�'h�CN!+��!�&��|��1��HO� �t	���:Kb�����9�F$Q�"OtpHr(C c�S���64��\��"O����	B� ���%N�v�X5S�"O�����5����Q�>>�X�"O$�f��*����NN�F(��3"O �IP"]+{8���!��a��"O���d 	*���%�	!*�,��"O��z�aT�~��0�Z�Z<������I�Eִ�RgO�"�@1(R�J��B�	�sV��6FT���!;�"9� B䉁#�P]0UM�"�(M�dѼd�C�Ni�% r# �35��8B�P��C�I�#05�AȿsF�}�%��v�C�I7Z���a������+ B�_�C�I�3�,�T�!S$zT'^[B�	�m��de	�$��)휇9B�I�-da �/
�a4�a�'�F�P�.B�I6������� �|���CY��C䉹5�2��"�l�2]��H�#q��B�	�"\�H����;��}��O��$��B��t|�ԢscI&7��@�	�Sb�B�	4��Rv��^�-8�䈢�\B��5qZX�J�ʈ�xq��:-B�ɰ3d�A���̹u&��j��""�BB�Y�$�	�o�_6�X0�	a2B�I)Uʐ�r�_�0s��"O �#%(�b��h����ѹ�"O|l��@P!ZLf�S��(��Z�@�!�S8o��Q �.��g_���D�!!��>�jp�'�ï,<��&�Z_���;�O��8�L_9��L�ĀN�|T�	&"O@;R������h�/8���[Q"Oʰ�4%��2s�0s"h@�,���"O6D�ǂP/9���5'�=fٌ�d"Ou���H!4�
V���������'�qO�֩� "���CF��dU�D�)|OZ��k[�m�0�$M!L\\K!"Ov<�A�Ʈ� Eۧ�� W8-р"ON
�%�f���vc�xn�Ye"O y� ��9y`���AB��"X`�h"O��)Dk����L��gŷbh���"Of��C�Ꚑ�fk]�e
��'��ɱ/�6Ւ�̈́�d$┢�	
�.B䉍	V!j%l����|eG;i<`C��!=#�DJ�i�b����_/O�*C�ɛQ*�P��F�dŮ�A�o^�t��B�� ��ǩ�2�0\(TL�AdC��
{ר<ـ�/L�$��Y2
��B��?7��)0��x˔L
UHSXc�C�I!	V�ֆ�eؾQ��Ǐ�Z/�C��:�uz��Hߨ�	�B��Z�xC�	�J�	`d�	�!΢IɃ�1{Z
B�	WSL�����a�tգa��F��C�I 0��-����$9�0�U�Q�`��B�I���dqb�=7���T�Ι:��C��/H���"��G�,��,��B�-�C�'NP���Vy<��amM�TK�C� cV�h������=���K+w�C�	�KS��c��$2g�5�"L4�C�	�`~9����+�F�[SaV�+Q�C�	n��A����x
��a(W�-�hC�ɒa��mvEZ�f��U䔙�LC�.ń bB*�.Q �0�ӍHC�	�h�¤�8��`��(_C�)� T�j�A�JK�;'$G?}�$ x!"O
E5)�g��IK�Ó�{�
�"O�5�Q���c�H`т�8j�59"O��y�H�F�0����^W�ղP"OԤ!% _#b�U(7FZ�O\:0��"O�5�q�����ء��1X?�L*2"O�Aa6�ås���
�Э:h`J�"Ox��Ul��8�K�$X�H��	�"O�A�U��+\dxy��I1`�6	��"ON��R@L�?����e"�3Bt�Ź"O\��U�˜u���+vf�fb��X3"O�|���VJ�(�t��"?�)B�"Or�����iJȠ��0r�_5!�d׫f���A�o3�њ�jH�G)!�䁪>���pTk�L/X����M�C!!��'��mD+�5{d١�
(�!� [޺<�3��:aĀ��)]�/�!��D�|��PɈ�eQ�! !�!�$P"xt���MWg1�TC���p�!�D 27r�(ackH(_��*/V�]�!�D.N�Q��.Ϛ:!j��5��>P!�$N%L4u 6OߘF��$��N3!�$G�4���*:l��@�,�;T�!�H�)!�� �+_�t`�q�K��f�!�DE�@�GO�JJ8��f��R�!�I����֥5xh�0��NM�C䉎C{8e�c-��VJ��'�	��C�	&�"��bR�`�ҴS'`2f�C���ِF�'���gE��{���	y�&)X�e9yC�d�u�F:�!�E	d%2��3(0�(e��a!���x�j�J��'*,%{��/U!�.�Pڲ��K;��[t�Q'T!�Ğ���Jc�I;\!���O�P!��y]3$	�*�Ȅ!5��RF!��=�b�Ѐ��:���*��I2!��ޏq�y1� ��R��L�w!�D�;Mb��qUD�l!Z�+�r!��0_�
����C�n!�d��R�:�v���D�];4CV��!�C�<�Z�-Xw�%k3��h�!�d1r'�!�% �>Y����;B�!�dU	�n�HgH�k�6�����t!�d@$U% ĸ� T� ��r�͠7Z!��L� ��PB5������CM/dO!���,Q��	@C�H���hFB�Y!�$֟d� H�-B�w����(�i�!�DL�A@P�p�W"Lzn�S���&N�!���uF��+V�N^[:1�7�)z!�d� N8�|��ʂ�G�2�ȅ$P�x!�d�#)pb�RG(�hΪ9CQ�^X!��].�!�S���p�M�#W!�$�?1�`�a���(��0H����oT!�䀩v�4Q9҇��W 
��t�HD!�7�~�qd��?m�ۓ��2!�H�<�zq�B���m�c,��w0!�$��z��	X�X��|�*� ]!��C�Zkl��!�r�X�(Q52Y!�1W�N)�5g�Sr��Z�P�wg!��}��@N�
��:�j/g�Jy

�'mz]S+__R����˵Zz�C	�'�N������/�}�f͟� ����'��A���'^ȾX�en<BQ��'b*y$	{F�H�R�ļ�N/�y
� *��'�	n�D��@���r��b"OTԊ ��=�n���U �p��t"O^E	5ʓ�C�m@L!/q�	{�"O�I	r��5C���*�3d[�4��"O����S[,$�Q
�	@Z�a�"O|ui c�Y+ƱZ�"�-a0<;p"O����o��A��{A��"O��8�ν��G�ߞQ�p%x�"O�!��){�.��`��S���Y'"Oi� Y	dP ������@�����"OF�
� *D�@��&���"O&<iG��2J\^�"FOV�k��aG"Or2� _ m���Ƨի*0훓"O�x��FW�S0�D�QF(Vq�q"O�A��N3]���qD�+��x�"O�RbU��Y�e�0u<-�7"O*}�DϞV%h��ga�u<�,""O(�;ԍ��]�ؙ�v��S*���"OZ=��i�-�eӣ��X.bț�"O$%q&Y�*����D��$"O���O_GL]pRg��xt��"O0���ᖈ?�R���凇9m���"O���&@','�Ez`�ė@O�(�"O(<�{ځ�Hܸf�|���"Ob��m�$Q@�d��)�pঈI�"OB5�&i	#O�؁v�])eü�Q"OLd`��F??Z��F.N�Z� �"Ot%jG��8q�#�e�e�.Y�"O���ѥ��2�J��pOb�9�0"Oِ2���&��ha"l��*e"OZH�5 ¸����d��Ĩr�"O�y����Gs�Y;1�2c��C6"O0�s���N���qp!�=p�H�p"O8�)�O]Wp�	ƯF�F�JqB'"O�)W�ʞvL* ���%B����"OH\��l�0��4A���?P�N8U"OɃb��7�=0���t�"l@5"O���1��.�pQ�"��=%6b�"OPp ��-u�T��P�ҸsHY�p"Op��b�?ydJle�T�{�H� "O� ���<?�^TCѯ��sֺ�CV"O�	V/�lڥ11����I��"O.!:�
�>y�b�£��\YZe"O0[P��R�$4`f�,J�P�h"O���UmS�n��a &]���S�"O�(�a&/ؽQb�ū
��ࡕ"OZ����N���*	R���q"O��E�����SI����c'"O���"�cxl������y�(��s"OM�@���L��GF�3���Ҕ"O� gP>6�ZD� �7p0< P"Oꉊ�j^�#���(6�<
�y�"O���kO!6�"�]�w�6��"OΌ 3iȂ3!��1���0?�"�*"O0�3���|��-(5�"�@"O������V�p���̦2��0`"O���$�H��:8���������<�Ǡ[I�	ٵo�)>���:%�z�< B�6�PR�!�-`8��0#IN�<)�ᙖ&NY� B*^{^ DD�A�<a�F4"��-��Ɯ:-�H�m�z�<���ϝ*�z� tj�i] `�Zp�<Yd��9�D���ұ~��Qq�<9�� kG���R`�&1�#Ώi�<� x�{"�R.���`19�Hs"OL��f$�3J`|��K�2�P���"O^-zc�S4G�X�A����L��@"O��d�@Q�t���-���҄"O0���|���#G+��Z���"O��yj����|��T�&60id"OR�8��.X��Qb$�EF"O�q�Ei�,id�
.h򊴊�"O`XR]�X��ua�ϗu�t��"OQ���B5g]� g�9Ħ��"OP�1V�&1�����g�3\��Y"O1* B�:DN,P���4M�D�D"O��:��]��lcG���q����E"O�!�R.ρd�Y��ѕ~��� 	�'Ȱ����uƄAr�b7o����'7�г�Z(f X
�C�l	B�`�'��I��Ē�c.ZkD��b\t	�
�'��aN$]���+^;Mw�9z
�'��@���=��R�^�J�$�	�'/�� �<+�t��HA�����'�"�!��=jFp���>.x�[�'�n���لX"Zْ�jѯ0�x��
�'�P]�dmo˞�
 (ɂ]e�E9
�'I�US7�M�tE+$#�Yݐ�{	�'qB��+\�0C�9}�	�'T����ֿ4(�ˡ��:��Ѐ	�'�#P�؅g�1��/xi��'f�0�N$h�*��HX%)���A�'I��Vb�%w� ��N�P  P�
�'�����zWt�%��y�����'�� 
�ː,�@�-ܐp�z�x�'4��pa2���d�T���!	�'����`���#���tݱ�'L��H��GA��[쉽r����'�H�0$S�:��a��#V 9{���
�'��0���Q���e��b�T1�'��jƊD�,�je@�,�VԮ��'z�DA��R:
\4� �ꏆG����'A�e� iͲc�h*�8KQ�8;�'h�y$�ڻ�VȨ�'/8r����'J&Ps���r�ا-��ZG��'�n(��*���₹TT�I��'^���R,dI����L*N�$���'<��K�F����C�[����p�'<FpJ&ĝ�y>��@�נA.�'�r�2�Q$����_!W�� �'���t��>iLm�W�A�w�p�[�'5��i��bL���2p��Y�'�0����/	x �懜��.Y��'� �Y�KS Ux�r��I�6����'-���o�#=;*l����50ZP9�'F�XaQʆ�:�6��BX"<���'7�YP�25�.������8KFXr�'+d���A� ��5ZR�.3��)Y�'��Qs/�$dF m�֡B�/&M��'����3��
#�~���Ŧ``	�'���J�	"z��F�E-<)���'�bs�Y�C�ГU�A�2}���'��u�3��8����98!i��'{
�
�e?UZ��i��4tl��'�`���2a���� P.4c�Ą�Y�¼����`~vz����!�t�<qE�O����4B0c�H�K6��r�<�7�Q�<���q���P��t���q�<� J}K�N!{ɚ�Sw�\�>7��C4"OD��r��*A���+Ṕ!�l�"Oʅ�T�ñB�4`Nߧ
�2d�"Ot�Q���4RZ�y�OӾV�@�"O�I f �=����.q�b��Q"O6X*a�ٗ]Jt�xC�T�����"O�u�P�O���w�Z%v�0�"O()�¨���
�KÉ^X��'
ly(�ϔnĤb��|�d�
�'�BHʃ�I]�l���0$g��#�'8��i�b�
"q��0��
�'��
���\C�-�$+��|i
�'�*����ϸj�4�PRG�(��͸	�'�*�k��:-y�u*��W��T)��'���#�4�Z{h���J���'P@89�l�)$���@���DA��'�,��Q�օX��z�끠Z����'Y�5���^3�eC�Q�)���Q���/O�r�%A^��ܣ��_�f��KR"O��(օ��x��Yp�ZK�q�"O����Z����� #V�`��"O�abȖ�y+ez�K��̚@"O@;f!V<6��D��a���Z�"Oq3��R�8Y�0q�@��P��a�!"O���cD�*1 ��1!EQ�"���r�"O���vMU�N��!J �ƀD�����"O�ы�{xDŃ�V�{ʗ����hOq�$�2d[�QLt�@s̉�h:M��"O���$��O:\5��퐄� "O���?�����VQ�"ORl�A���
���U�AK@^�{�"O ��L:t���q� IT���"Oh��� @x��\���F	��S�"O�
�fÛxz^AXX	s�-" B�Y�<qu�.e�n����<SEj�qVA�o�<I�1l�"�KB
�(��uk	j�<�d�G(#�6=�$N��*~���C_�<�% ���� �^ش�R3	V\�<��ȹ#��2'��egkW[�<a��"8&�[e��TcD��#��X�<Y���NTFE2�	�{�Q ��TR�<���Ͳ�] !�	����D��J�<Iq�Y'�l`F�S�h%
�#%��E�<�B�	�B�����3wkV"dŒ �ȓJv��aP�n��`"��˜z��ȓJ>��j�q���E�tD{��'��� VB3,J�����w��F�NL�<A�����&1�� K<
��q�<!V%	'_��1��L��*�!���n�<ag�#2�@u����� ɖ`�<��c��f�nyMK4�J�@\�<���B���(@�τ5�L�1�m�<!CD�gi��x�8=��!"VK�a�'�axr�9t~�:�HF�w?�� T����y"Dл;�h�"��lv�2��T���x�W�O&�P�wc�3�z�'�*1!�\#gEvh�VLR	{Rj	⒮F�Py��E\��f��?"�U�S ��y�/�*rV��'��'��B����yR+
��r��G&E�B-(����=	�y�D�#n��9�#�/2�	���y"#4�D���GF:[(9Ѓ���yrh�v�dJ��͢%���3G�(�y�`�>]D\�����5�q3�E�9�y
� B�j��
q�V�[G�5z^F�BP�F{��2,n�Ui �9y��cS"X�P�!��Θ8����Kx�1*��.�ў��l8�I$�Ƈ^5 M ݈m�*B䉺b�.T���Ԁ4��d�voE�C�Iu����i�)rt�xf�����C�
�лf㜹j��Z���I>fC䉜v�VB�M�~"���G�4C�	�}�Tx�!�S���0�kX"C��;R��GK�"ܼ�{gB�6��B�	 @E����!T!`��ŅP��B�ɵAU�@匜j�\���OWt� G{J?)�h�
`Ƽ����cx|m�pB"D���1�I(�a(��=q�!�3�>D��{uBR�YK��h�����:���O���>�ѥ,U�NPԳKT3�3�7D��R��	5D���%p��D"On@ZTFY+{ఠ�7��D}���#�(� �Sܧ!�N�ʇ�;6رJ�hV�aǂX���^yR�Y�%t,`�n�H�A�aD$!�d1qd���j�-$�1�nݹ<!�dX%bL��'\:u
|����53!�D:JȄ2(�'�����F
AyR�'p�|���ܲdVaAND-u"
u�����!�@[jX�bƇfvR1��"�!�
se��Ss�H���J�@�!��lW̤���p�YB��j�!�d��A$59d��.����E��]5!��ΐoQд@�DA��|]�,�"g �}���0(�&ժS�B����� y���Q*�<A.O~�OQ>Փ���U�(�h�g?u��)�k6D�{"�ŞjǮeȆGM"x㴡r�4��hO��$Ï{�HQU����c�ՂE���d3���z��z�
R�Q����VGM&}&�1�ȓN�Ω
0��C�Bd@�=K�����5��X8V��F����֥�8Ur\���IF�')���ӢPY>-˻d�0,O����OH�OQ>��C�4r�	���y�f�1�m-|O|b�l��/H4�R����410@ʶ�<�����M��d�D�Ď4ظ��AԳGU�B䉔<BD���k�`�J���7/�|B�	�vDY��V]6`!��,dB�	�S��Q�,�p�S���d��C��!�LlC��=c�<� ����O��C�IX0��F)��5\6���ڼK����"�&�
I�"Ϸ1�p|��-��7Э�ȓ~�"��eʹA1"y֣M�4��!�Ɠ `�]+��.!�,�+�b�D��8��'�*��f�lv���q��=B�,�Z�'ǶH1#e�q��Aqc؅J���(OZ�=E�d������"�:Z�����y�m���m#�D*A�}p#C���y���:٪p��µ� �9�D���y��C.i�����(=R��
���y�/U�so������$��;�i��y⦁.T�����}���LD��y�� &��ㅅ^�j��hFi��y2��.��e��%�)P�ȱ�hV��y�'��3����&�E�o����'��y��Y�pSTY�w�ڸgb@�f/̂�hO��D;�}�j��bh�,w��=x��\]��`���hO?e���JW�����3;�*�Q�op�<�@�� ���xT+Y&�*��a;D��f��8T����;4���Q�3D�� ����!`�����n�9_�T'��G{�O���:筅�b#*�Y���<�]
�'�:=)���M?��0��@�G��ٱ�'Q�A{f}�����D�%3)h�Q���1��+@�Ŝ���X�N�nQ:d�2�SV�<�@Ȃ}!>�0F����!ƁJ�<�d%I�4ԡ���Qr� �d�����#?���/>	��H'�BbY��ӥEC�<� e��衢��qb0�#Z}�<�#�(dzZ͢���\����W��Myb�)ʧ"�j�'CU��Y	`�J/1�z���nnD�ʆ ,�u
F�\(2�X�ȓMz����
{�<�{V�*1��ه��8L�`>u�hk��K?F���ȓ2��%bnK)А���ʏ�8e�?ӓB蠄x�H�%����.;6�ܴ��{	�� �*]�[T�AQhK/I]�x��j�P��% �:tI��!�ȇ�Y�(: �M�j�x�Qd��c�
@�ȓ}+.Ha�ǈ7�B��+�V���F�P�s��8�ّ�.�f�� ��v���������{����<J��8��0ړ�hO�ɾs݂��DC"v��̂��/�C䉎:�<-��Z� z�����?H���O������p@�Pc�R�x젶�дo��j��TI���=DV�4Z��a� �'�y�߲9hxK������b���y�IM.&m�#�� u@t��Q䔕��&�S�O�굃��(�������b$�i��'�J�k�Ο�Ma�����[��i�'B0!��Ș!r��!m�@�1�
�':`,JwlE9�1��IAH@
��yB)-��j��	,��fC��y���BN��fj�z��\���4�y"��¡�djp	 �!6r�����������Պ+,�)��ϖ=G�bO޸hR"��T��f���p%�"Ov��b��\Gԍ��˖L�H��'H1Oj���'H� 6̋BC;S��qK�"O� 0�DV;{n�T�C�	"1�����"O�`B��6h��� K)����"O�2�V�1�H`�%��@<��"OYj'�ǵP֊Iأ		��xy"O�xP���
aڹ��[��D�b"O�l�r)��o��#�&F�6�|"O��x�`�"�� �PºHP�"O�PX���b{�@K��J�c�0�Q"O�ѳU��S�m�v*�X� ��"O�(9Qn�	8���"D�w���2"Of41u�E$���T��t��h�"Ov�S����[$�B�LB�9@"On���HY�!���z��~>�|Pv�D&�S���,%����1�֫0��CQ�!�d�<O49��I���h��j9 �!�N)��A�G�z9���ǁ�!�ċH%W&U�g� �`�-j��� ��Y�)�'o��]+��9f�.xrW�X���$��劗�	�I��B`��h��
2P����>	t-����+(�F��''ў�|�dӏM�S�>�r	Ы�[�<YD۰e��c+�	4�dЀvJW�<��Գ@^}'�Y�@�Lå��Q�<��N̡nt } �Н2n���Bx�\�'�8I�*Abm1��[	b��`�#"O� ����[���ٛ'�0e:�"O �*�5�P�zAC7���J@"OI�/�);1����ۣN���a%"O�tz�L�+1����'��FWԑ�"OH|�5 c��dr� 0I��"O��Q��@	[����j!9Ʉt�!Z�������&��|�&[B���` A�	2�u�もb�<���ڔ<�`I�I�����᠇S�<��ϋD`�@��K9��H�1dDR�<E��)t�5۠h�L��Eb3�R�<��C�j��`����a�V��� \y�<���b�@�yw���qj֮�y�<1g�?�|�b�J�ZϘu;��Ku�<�%�FX��UP� Ø{��Q�C@��D{��)�#�<|cD)��[P\���	IzB�ɿTq(+��ĨAֆ�ZԆI�vB�I�gjh����)|�,��,^(8B�� O��2�^�(�n��Ӊ7Z�B�Is�40����0Y�P���ȈK��C䉷P��(�/uO ��#.g��C��<@� 	W.��H�ՙ�=�
ç\��D�1 تSgV�u*�%t����,��i9�"I3U�����C9��ȓT��i���y� @K�)�ڼ��B��y{����g�"E�I�F���ȓ � 쟩Q�|ք�:�:��ȓ`5���盙&�pP,4(̆ȓEo|uóbQ�=��4�w��|�
�&���I�GjZl+B�:<?Τ�
�<] C�<q($㡒�q�`۳-ȲY��B�)�jE��bʛL"ƈ��,�,>�B�	$n亙��A���L�n�=#v`B�"=i�a�f �[������̓P4B�It� ���,/�EHf��:9�B�I�(I��K��e<`kE_oHv�=��,&���$��T�Ĺ�A�
�`�ȓ�v8��6iN|��͔�|��X��L%�eKŮ�R򖥨V��8=^Y���x��6%��ӄ�����ȓNN�=���܎q�xP@շ	�H���%��|;�0�Tl�c�ٓR�Mth<�T�L��|9�+�8p�
v�>�y��8uO0�+T�M���XE�G'�y� ���&���&��d�P�CX0�yI�s�\i�ŚpP�W#I���'掭 
�O,���O9R��hƈV��-��G�.�	G���|�TyK�i�0/�|��ȓ?��tf%��D����&ʖt�ȓN(`0�#
�j�#R��[�ȓ]""l��O�9z@F٪@ ����ȓ�#0��p�"�Z����d�H����vAJ%�ٕ��¢�eqHD{"�'�B���D%u��I��;lL�!�'��W�']>8��ę%�2�'�xM/}�\ᛒ�K�KǬA�� m�<��ٹ#Q���R�ܜ�@;u��h�<)�/�*`*�b�D�-	ʤg@P�<���	YӐ9`�]6K���IN�<1��T�pY0����Ɩc�Z�Q�lDM�<��Lļy���fD�3&�+ ��S�<�@�U�O(��镫H���5!O�G�<�,Y
t��H�+ˌ	:�m���|�<�b�?4��Z�*�|6����<�F"��g����J0b#�	��O~�<� �,���F1*����HN5->]c�"OJ���hXu�	�g�cL���"O.�����TƑ�c�T	D��0"O��V	��4U"-Q� ��Wg�y� ��Hpv���ׄ50`�n��y!�Z���q�N�]̀�VO��y��DKN����2���ӄ�R�y�L%Y��Q35�R� �l�r�m@2�y�o�J2�u0�4(�.�����y��k9 i�,�v���� �y�o��<�(��IT�m`�[@�L �y�D��?�8!2��u��Ų7	�yR�ςunlyQ����f=B� �����hOq�<�n��7�R��V�@�;��a�%"O�� aL�g�R\J��Y��p&"O��2��'6~�L��hD� �F�J�"O�I[�dT0z8z�;�-$��=��"Ox�@�Ѣ/:�CDN��;sD�k�"Ozh��AZdw�!C%��V"%�3"O0U�P��U��e
]=DyRc"O�aP��Z�> ����T��"Oj���@ܽZ�|5:0 �p� �"O���i��f�R�X$5(ܩ"O�a�3��~r�3iG!֘I�"OP�AA�[�UU�5��W�,��UHV"O��P��pwy=6�@ģD�'61OX�ȱ-ɱ>B��S����k"OV0��� #r�̣1`��+`±�"Of�����j�*����nk�Q�"OҸY�b��D��`���+I�1O�!��)�Ӛ��i��g�a���ȱ��2P�C�0^8�V�d��q��Ђz��B�I�SNhz$/�T����EP�A�z��2?�5䕠r"�b�D=h*%P&J�h�<qdo�ry�$1R������${�<q�h
����(T(�94�\b��Rz�<1A�IPąP�=O��Q��m�`�'�a���!�e���V>l��� ϒ�y�A�=U	D)���ˮi���5�L	�yB�۠v���Ѝ] TVj�U����?��'ǘ�KE�HsJ��ˤ��$W����'�X5Y�IC�:i�K����'������=q�Jz0��l�h[	�'����(��Q�����2Q]Z�x�'9Vx�׃�8��a`��ъ�D���':�|[4螣<�0�"�"�<	���'��9��J�.*��C�GF>�"����?ٜ'�4�F� f^���2OH]Nٺ�"��%�	-9]tà���^�R��6^��C�	�,��h�'�Ƅp��T���C䉥p�Re(�ʒ1K=R�q�ڡB�6c��@��#�Şh\%���#Ʋ�h�叇`x4̆ȓWd�qg,~�0h��σ|���ȓZ�֡�@��Jq+�j�=|'���ȓq� }�Gt�րK���.�z����=B��=�d[��68���ȓG��l�@@�!|�J���-9o�h�� �)�&@�#��H�U
 ���'��B���Ӽj��m��-P)��p0j�Pg�B�qH��J��F9��0I�c� d�B�I5+��,��g;�ڸ*�"ѥy�B�I���@I��f�DY�UW4B�ɕ�l���P�o�L�ҡD	� B�	����Z!g03��ԒA@¥��"O� ��q��9H����Ǟ�|�ɠ�IL>�9� �P���6�˴D�޽���6D�(��iG�;D���	��i�7D�|�EĎx��a����>{t�0un4D�<C&�� rs���#[, ���3D���Q$E=��H�
 ��l2D�4�HRK�Vͨ��҉F��a��2D�h�S�оBA�aѣs�|0�l3D�8	v"G���"�`�	�lB�2D�\�S.Eo�t��Z� x֘1V-&D�t"S�@b*L� t�&���т�9D�85JU�l@Fk��k��8�$D��k�d@�E�� �r� R��&I.D���w
��C`)��!J�;�t��4d,D���tBH��(�+���<)�!J>�����1(6�3�G<���pB�r�!�D!JHh���IMj�Հ���2��\��y�n�3/�ej�m��yr!�;ux�I����P�d��*�y�	�Iּq�D'���=���?y����$AK�4��	¼_�x}��Ly
��:M�9���(JF��H������'�jqs������rp�0#]~��Ǜ*��a"O��H� ٽmq��EH=v�V9�1"OE�EF$#�>�`�#S�-:r"O�T��j����91
�6�&�"O�!���W�+�ڗ�J:<m�4"OL�r0K:WNZ`)E�ƺD#���W"O�j�IM�T1 ]�]����H�hO6��$�%,��*c�P��]Z�j;�!�$�+��k&�@\�أ�"�!�d�X�𘃷�ɶ���[�aD!�d"x��8h��UD5���>i!��S00޴� ��1�� ���h�!�$<P_zE��IP�+u^!�d�Ԋ��3�E?�����F�?!�Dt�H89�,�/@�%�'�^!�_5K�YDd�6��1��M�!��!��0�@A�P^>���=�!�jN�L@Ӥ�����ض"� so!�ɛk��RGBڜ���0'�:a!�$� oĐqS`I�3x$�%\-k=ў ��S�W���°�Y(�C�mcVB�I�%���傑��
���;�NB�I�@Nt��AB����W�_�B��!~�6q���׈Y������و4A�B�	-�ڭZ�)[�6!V<` K����C�I93�0oH:l޹zd�4p
�C�A��p#P&]мٶ��B�	�I�`4��鋾9��@ �H(m~�B�ɷ4PT1a�Hڵ��ȑD6�B�I������bO�0o�AB���G��B�I4N����L�g!�@� шg�~B�t#<��2��*/�1;�j�	ȡ�1���4�eW(��!%� =!�D�2|q���jS4��a��Y�3�!��̧6�ܙ1���<���bE!���Nu]Z
�\�Ή`� G��!�?;�@l�f���|���1�ڦ�!�݁i��Z�-J~��ic�l�05͡��Q�)p�h+vU$��U�v�ڶ�y����>��'oI/6(-��Һ�y�kݪ4��Y�6ƾB]};D 5�y������	 �F�j��q
�n��y
� ��&W�a�H��5�U�A�|1a�"O��t��1m1>ܲ�N��LiP"O��c��mlTp��(ٯU�R�"O�<#�e�ȸ�5N�7C��z�"O0T��E��B��f$� �ɿJ�!�DT$%c^a4��<�����E��x�!򤗶�0��$��Tfyq��$f�!�4g���TO�<L6]P����@}!�d�)B�5�g�(Z� `2��T!򤂶I��-a��9tVh�L�(p�!�ܟV����Bo�2}��ɻC�L3/!�6}A&u@�e�)9����Dى!!��O�g����`��0���J�$և!�$P�h��݊���V�~n㑘O!�$�=e���7ɒ�N��}��J�#E�!�$�i�z���>'�����}[!��JbX�D[7x��B�Q->!��C��ܒ�'� X���1$O&!�JnPJ�$��o�T`G�Չig�A�ȓU��1��^$x��ɱI��I�<ɇȓWr� ���9h�N`��Q(mB��ȓM�.}pc J�XwtX��v�`�ȓ|�R��D�9C!-XZ�e�R�<A�*L�e��S���1%}�T8&�v�<�j�`�؉�UD]�	�>�E	r�<	�'7�!H����,"sLq�<9􌑶dtvY�W股Xi�pP5�RA�<	t���:#��i-G�sS�{��Xz�<ѣDQ?y�5a!��t9��1�b�<��"��fb�i	��U��3�T�<)DF�i�a��v�� �ՠ%D���e�H&ġhMô��"D���ӈРm(�@蔅�%1�*l�s�?D� Z� ԫ�d@�ѭ�!�X�>D�h�`��Y>��P,��DN�K�0D� ���d���hB��,@�Ʃ:D��	d�٧Wo�����o�
����5D�`�"�q�V�*=��@@�G#�y��1S�L0���(@p�(<�!�ǆ|4��B�a2�LiE���B�!�˷wM�tB2��2<(.��W k}!�� �vL��Y
5�����C�y!�$ǆ��h��NAI�z`0�-�c�!�Ɓg9 ɒ���m�ȍ����J!�ו
$���^��h9Ԏ��'3!���^�0�� �U��(�[F@߬�!�$Xk�x��vT\͂Cm@�M�!�$U G~�Hւ�+��ղ����!��J�7�h�6�P�#iMbg���D!�ϴ$7>yCa+Z�Db0���]EJ!�$��N��P���R:�,e��	�Py�'Z�3|�@��EW�Y�e[����yR$�=8��-�7ї��}����y�7X�\,1&��#,h�ۦ�yrlˣA/U��[�v/&�J� 	1�y2f�Lj��S���n�u�r��yB��`�$y�D�i��ْ�׾�yrf�:�5͗L*R�Brj���y�+Q�{JL�KOBJ��yb*�!&�jP���=�lE2&���y�Ϸ@����qe��R�c�iK=�y�eJ�Fc��1���$@��I�`FM��y"`�l̀a��c�{��%�y"쒘RF�q��&�$��X��.��y
� T���̕e�8���� 4���:�"O@Q�$	�ld��I�\!�ܱ��"O�FҦ��s��P�(̐�"OHAɶ�M(
�"�c�+>b}� I�"O�*I4�p0�i?D}L��"O�������B�)�i�M�N��"O�Y�f�� .��*o�{Lf�0B"O��y����*kn8@�ę,Cl(�"O��	�
�
!��ːj[�,�w"O�:w&_0�< Rv��+<2"O�=���ј]8�o� RD�$"O��B�[L7��Q�;���2"O�4���4��P)� Z��x�4"Ob�)���;��GO�+G�6mI"Oa���� 0�5�? ��+U"OFY�S"%ά[��*\���0"Ox�:�/�X�hiH"��CF��CV"O�P�������&���p�"O�y��P�
8��iժA��QT"O���`�.k�8c�.7�|���"O��a,�z���U�{�HH �"O��	G*'4�ɃK�[C�!i�"O�$Fl�b��,��)Ϊ@�p�6"O±��>�\����,���"O���&զrGđ��O׳E�<Bp"O��C��}XF5 ��!���"O~a�)N q;&�2mÊx��IP�"Ot�	���^��+W��Q��s3"O�M2"(�	V��Mq
�4��i"OpX�- )#��,O�hhY��"O�-����!/o�,Ó�(f�ȃ "O�\�e�E�rp��C+D����"O
	{rB�-���A؁,;�!s6"O�Q��O#��"2c6JȀ��"O����ѱ_�����\�<�I2"OZx�".�?s����R#�/�T9�"O� !bO� ���ɗ��MH"O��PhFb4��S!,�@��"O  K���4�d�d�t�.�C"O�J�/é5�(���Zf�02�"OX].5	.��b.܍"f&l�����y���8�c%H��
�"�o���y�Ƒ�[p:}�1��,]���1�y����i�j�W*�(3�EM��yR��-N�d(E�݁K�\e!�M.�y�i �;خɱ���I_tQ�W)�9�ybؿG��!�46Ek�����V�y"��&e9FE�M�%�g�ָ�y�/{��ܞPeF�'kP=�y����pm����(���1vn��y�OZ/AEv)"pdZ��� �#�:�y⥙!s�怊I]�:������#�y"��4��hggL�GWz%#�š�y���L��{&b�27��"$�(�y
�e@X7�NZ�}y�,Z��y2�� &��mC��@%K�FT���y"�ҽ ��A��PK
�,� (���y���L�\I5cD�Nh�y8 j���yR�5x�̱"�Kلl�JG��yR�Av�<����{ify��GQ��yۀN��i��j�l�4M��H[��y�OV13q��P-h���쏹�y2c#Hr�ЁaA^�X0*|�����yB�I�Ѩ��'ծ��Fl=�y
� �8i#i�U暹c�B,��͡1"Ob����T�JzY��C��U��"O�t�rNԔ}��������p��"OB��vOתSK�+t�A�X�jE"O���$M�
�~h�����p�I�"O2�-�t9��+��1=��)�"O6ձ���_����[�#�dٲ"OĤ
7wx�� ��ƋmUZ���"O�im��d��a�N�p��"O�]`�#0D�JQ���/`K��[B"O�ԃqdZ�<��1��Ȇ`n�y"Oz}ab�ӏe�� 3A	�f��!yA"OZ�L�m��=	rV!:��,"O�L�6M	 L�RAi��4~��� t"O�m�0KF7}A��j�:�f��"O�` �^'%����	���H��"Oj�S�<��	��F�T�0�k1"OحB��x����%_�^Z4( "O��X�Ǔ�dI��D�!iJ!r�"O(0bi^c�L�҂�>8/Ԍ�@"O���R5I��JA�ۄ`;�1Xv"OVPJ������j�똦h�� ��"O�l��jY�R?@�I4��<�>�sq"O4���\bB��������D"OXd{#*P �0��7�ߢ��y{!��֓=&VZ�� �I-C3jǭJf!�d�<6��H �H�rFv�bEfT�g�!�DL��|��I&&�n iÇZ"2�!�ӵ	��@��`�)�F(�a��j!�M�B�rS���d&� ;�*1\!�Į�t� Ӈ�'1"��CJD�n*!��D�l�^�z$j�<(��K�"!�� pƠ�E�	�S:�p0���*!��F�W�$� �A0!~��*΀D�!��Y�2�0��cK�HxN%O�K�!�$լ#�`�=qvĝbPNP�>����S����E�N;k,LiuGͱ�y��'y�^]i3�V12��w��-�y�Z�N(r�Q�&->��dK2���y2)ǂsID�b\�m�Z	�Qc���yr
�	h����cݧ|6Ĥ��g���y�+ݗf(�Z�'^�G��q�L�y"N�#X�.���'*iR9�p�Ӌ�y¥��%N(j�A̠!�IТ^�y�@�p��4��fL�˦)ig���y�˓J%�}8�Γ�1�����J^�y���6�j`��N&)�V�xa�^��yҡιm�0P3C'DdZtBQo��y%H�Q�Li)1;xXZ��AG��y�ڟW�9(�D�AxN]�0F�yB��9�t�卉@N���F[��y�ʖ2w�ri�I�mRRpc �Y4�yRɕ�Q���⍘b2�Q�fL�y�uvNt�������^��yRi[���#��j��9�ã���y��9�Bq��D�\�����"!�y��ů<�F=��H&N��9�cf�%�yR�F&�骣�B�1�ְ��	�yr���(TH�JGb�<����%D��y�.J�D�4e�lH�gz�����y��V�,d��V��'g�h%2��	�yB�]�W4|iJʌa��M�����y2��G��j�N�	��%)����yB��� g֑�юŕO�"��>�y
� . ���=��%(	Y�7&f� G"O�<@�V%�]���a%B��"O�Z�� �1sp��숝C1ht�S"O��pIT,rv�5��D�9Hq �"O��Q��=l��	�� �Oh���V"OXx!��ڎJ�P�R	GO���"O�t����7[l)IW)˲@9����"O��(�F��N�� "���l+��p"O2x�`�m�T��K�~��"O���fHw��ffժ9q\8B"Oޜ붴�z�N�X�Dؼ\l"s�"O��04��
j4F�{aFA�"O>��J��6#ҹ�ɔ�R`(I2%"Ot�IȕZ���z��)<��	%"O�e�,�C���QDf�$94Tx�"OT��`'!8�Z�$(3�(6"O�M �<�%��2�iP���y�8xҴ#�D
�
��p�]��y"MP�����d���O�y��BKrI���p�1F`#�y2ψ�+�d-�� �J&4���F��yb��
W�a�>+��
F�y�΀������I3fµ:�ߨ�y�e��J�A�A��&����QLW��y��%�j�R
�� �~@�Pʑ��y�/�2r 2|1�X��� c��'�y��G��xaЁO ��(����yB���0�U�6(TCK�a��"ם�y��X�Vi�2���5oȭ3��(�yb��ېE��MǞ~{f$�@��yr��4fxv3D�D�y�N���h
�y�@X9{�0�Q��w� �YR���yB�*Xal��W�g�.xĬM�yB��:C�Yx��)d��4#WJ �yC��#|��	`CɌY_"�Z��ו�yrO�<~��Ȃ1b�>cx�Ɗ	�y"^iR, Rs#D�6<J	`�e��y��A�ZᚢA�d�z��5�:�yB��p��U���(O\�<�"���y"%W�Xft��F�!F�1����y��Ր&K@�з ȏv�����g��y2��z�(�����P�R�ϊ�yb �<&Ҝ�2��C���T:�'1�y� H ��}��Iږ7���rJ_4�y��V%^��H�!í(#�9
�e�/�y"c�p�m��H�=R� ��C�N+�y*	<('J8#��]X��5��fļ�y�B�.}+�@p �ȨZKH4h��֒�y��1b�m�-M��#CC��yR��k����c�FZ^�!r���y�$I����M�@h��h��y�o.'����"8d�$��hJ�y�cR1��@���K�gs�������yR�<d��0��R	W�F���Ϭ�y"��&�Ђ�������yR��C��@�#��|p�[�I��y��
��<�� ;{U��ÔǕ7�y��P�\Xb�o��t+��[��ּ�yR���u�x� ��>f&8	D�	�y��-4^N�2� �[g���S���yB͑:;� ��rC�	��y˃�H)�yR�ɑb�TŲ�*H;S!~�R����y�	�I�ᚵA�b��;�����yb��$pT�}��ᖃ[Q�ͻ����y
� �Ͳ���W�4��a��.���G"O,-��Ȅ�q'<�	�ڝ*��\� "O� �ݮ	�����"p���"O�qA�����r%+U�-�(D�&"O:�ؖ��J>�5u�ƂN�82P"O�X���J s/�� ��׍8����7"O�s��E+b�d	B۞.��ɹA"O�@s�l�
A�d�P�E��Q-�yR��l��%�@�t�Zyõ����y2�ˈRT��6�IhEJ�30˒��y��>B�=h�Q�[�}+@W=�y��4-���d��C7�,P�	*�y�l�z�0qVaPw����J��y"�¶2�)YN�?=��Z��ղ�y��E
9r-"�h�6W��Bk�%�y2M۴�� �Sk��]7ƭ��@��y $Y�zUC��X!V��f�]��y��>n9�5�"j6]�h1�H2�yr�W&����q �_� �:��N�y��T�@�~0r��^���������y�a\p�Ǆ�,��yh�A�y�C
-�vp������������y��۰A�ʔ�uED�T���k��ye 7�H��3柲RL8;����y�2]����a>O�Ƙ0qi���yr�3�MҦ"�	H��{�g�yb��
n���[B�Ȫ<�B���'�yB-��PPq*Ġ��5��k � �y�g\%<!2����|��"����y2�B `��(x�A ~4�P'��yR�[�(��2��]�*39�!K���y�!�"6�:E�����raK��y�E׸'�Աc1���ȑs�'���yRA!3�d���F,sF�q���y��G�=f͐2��y(v	��	!�y2G����Qi��C�o$8�	_�yr�8N����+gJ�@c�y�
$FTy��JE�-�1 vIX'�yR��c
� �0!L88Dڀb���yrX�xX���KL(��1��e���y����z4$��ـ��9����+�y"��n�d��gI��"<��eZ��y�&}"�XjBhPil�W�B��yRL�Z, R�C��z���7E[��y#J�]n�C"ph�AP��y�k��m���ч��X�4�]��yϏ�h?@��cϖ,�l��-\�y2�
0��Z�ˈ+!�|ɸ4M��y�$S�O���{��).�%��i\-�y�iR�(r� qW�HT�����y�N%2��1�`���@�H��y�fΒU�x�bg# %]�ش��3�yKC�a	
����&��E�,!�y2K��2�r�퇨� ����R�yRo��L�L��Ĕ$+�X�)��y��2�p�V	I�TtlǏn� B�ɣ;�\���+�{�T|{���&4��C䉁#�h0�F�,�I�q��8]��C�	�2w�蹅ϑe� [���^��B䉈?b�I	�"J�n��p��n�#�B�	�Qr�h9u ¤/Ȍ,9c�B���C�	�����e��&Hpd�T��90��d�+"R�{�n�<���o��J1!�ƻe�3�@
} �����P�!�� �E��>U��-S!AQ'@�X��p"O����$�	e!�=�1��_ք|Ӣ"Oj���5�D����Hb�P�e�|��' ��El�TF	'`4!�4�@��,sr��k�ɂ�	h�!@`���y"ǌ�]�]	�[L�d�ǌՆ�0<y���:h0t�֒��\b��.�!�d؍j��S#@=G�JmZ�nV�O!��2yx��#�
6�~D��G�D�!�d�{H��Z����y��S,]X!���q�L�����h��mFGE�'Aўb?	�юǉ��� E��	~3���_h<9��H�4�r���U��PkAk�G�<��d�J�:�A0�B�. p�+�,�z�	h���ĎٱE��W�fdiz�6�O���.\��ಃط<nZ��f(+A�C��㦩ɐ���4�ƴKbD�%h��(��E0D��E�4R�za��&Չp��(�p�+D�P�V�,x9I$˒�X�$�*�$q�|G{J?�PED	r�}@qn��H�De*g�'}Q���<A�}�o�%yM���i�/5F��w�ѡ�y'��A?n�J6�6� h�����0>�M>�A�um�-ۤꔘ�^��cO�<���7-j�bMM�YZp�ɡ�Q�'Y�"=�O������.Lʔ�р	��16� 
Ǔ�HOF�B��/J0���RSx�k"Oz�)q�F�tXBYcb���zm�L�AiM������N�F��!�A��
  �ō(:�!�DF�d��\��U'bP���2�-�I&�O2����5T�}�ճ��ݸ5��D8��'���fd�2!|�#�G)hyy�"Oz�dh��G����ר��\ZX�'"O�9r�>%5�]q�^8��m���>��'�0#=��t�ҵ�8��mp�)��ȅ���'\�ɏl�L �d�ʔ]@��@��RS��=�	ÓU@��n����D�*�2��� |�,����Z*�=1*�#o���	p<Yu� j���g%jvpZ��KB؞$�=�1b	�C�P��&D���:$̃|�IV���O�$�z]j�q�#�/K6��yyґ�$��|�"�_"�a� ��*��ځ�K�ð=��O�-���x��TW:�ك T�ɠ��WF��c���f��٢���g��=�ѕ�(��	U}�j�
�;5d٧[�$�J�Ș��0<14k9ʓ$��3 �?&q������4Ё��/֕*�@�>���˰�	/@ֺU�ȓP�<�i�=�$X��g�9�ȓ5 ��0���ph�iC�!Ζ �=ۓm�r�XvC���^�z�l�J̅ȓ+�~���%X�6(<2�kQT��	s?���A�
��ō�>O�9���~!�d�{�:�R2F0{�����O�V�!���!5R�̳3��4&Ղ�ꣀ&cz!�d�O`�4�Kj��m��,Ԣ1W�����.}��)�S%O���u+�8,�P}��d�?����#��6�\��o��Q���֬D۱O~��6O�����Ҽh>ha#JI#Z�~9q��!|OX&H�#5�$���~��i��i����^R�>��B'�5=�T��G��g}azB!p�@�OfT9�^�?���WIQD�D�f"OB��L�m��$����3zt��O�|��d�XIaJ�"}��E��@P�f��s0�
P�U�O8��S�p	㖋ӆ���zpd?0��'y�	u�\��؈_d��PF[/?�L�1C�"��ȟ� f��� n&��-�XA�Y�"O���Wf�F�)���ݜ5AF+��'��&��֧����/.��� 3	��ɪ�\��!�13M�,ia/J=���J6�A|t��0?�VNL�d��6W+���תY��y���%!�cr�!��Pe�y�'�95�$�W��4R܁ ,ز�?�B��<�a�
�a.�`��+K�! �]�<��!�-\̈�`�I&&��P�&e��<)M���'Ή��-�D� 0�Z25�l9z����@�ē-=��1
D<$ ���@��$wLp���Ԇ�I�2��y��]�9���4��'*$@���4�!�B�3���Ӟ�`�m�t��#�O6,��_6y�X�+͂�����|��i�)$�1�(A7$-b��� e$��*��!D�`l2�"���V�8��A!<O���x�IL���ළ�T��5��m�xɘ���O����w
�]"�aCz�<%�$#� T?!�DVu��J�"D�R�<y��;'!�D��]԰u:�mY}��ܺqBϏx!�d�3>n(#@�Ӊu�8�c��J�!�d%e�DQ�Uc�����	�a[�B�Ih���ԋ\�@j0"�)w�B�	*'���V
1x���Su�؄}|B�I�I��S6-���
�־%�"����I@�}rv K��v0'�t�B�	��(aOΤG}>m�6*�&C��~����	*� ��,?�"]�#�Z�QV����)
rH�{ ���FJ�1�C6]�nݐ"On��‖B@��� �������,�S�'t��6䛪7�(Ir��n���Ѭ�`$\Y��ɤ��t��t�ȓ`����$!p��d���F��.��ȓSh�ifiM<w�t���O&PQ�P�ȓ���0��ܒ,|fHڤ�� �F��ȓ	�xae�خg�T��ۄc�^��ȓ"��UP5T��
����ȓ;7`��V�G]�L�B��!r)�9��(�h	f�I_4�#1�� p6��ȓP�`T0ơE,�ҵ�#b��v��ȓ\��k��пN2*�ӶX&,�ȓv�
�{ā�$ ��ؑ���4�Їȓt$@��5�N�'�H�	��d	]�ȓm[�`�C�B/R���Ɗ+G^!��~f����msd����#�����/�(lZ���<�Ԭj���;\(JD��	�	YW�G�h��� j�Py����	�
�?0QҜ�q��݆��ȓ1�����Q3<(I��"�;6�l��^I.��(�h=���J9:�N���K�P���Si:R�Q�,
�,��6�v�ŌyO^,A烃��R��ȓD#�� �-[A��"s\:�ti�ȓUn��LE$ot ��3oЍI��4��,mp|��ҡ���Rŏ�Ȱ��u=��A�k��i�Z�b��L	;)f�ȓZ�<�d��Qؒ�b��S�O0��ȓ<�BdzS�ΓG��Z'L�?,Ђ���S����3�E�
[m��8�����$3d�� �Q/�1����d�"���A��d �n�/%Қ��a$�z1�)���`S��Em4��p͊Pv�х�O ��qn�^��`���ЕVjͅ�9e�I
ԉ�/j-˲G�u�����S�? ���g݌[҅P4��^>F��S"O��d���5�JU��h
�F!���"O�|�	׹H[�I��G��L�3C"O
�y��(,80P�6�;ti�"OPek�	D�6d�y)rE�8��*$"O~]�A�[ ��$aӪS�>Ͳ��V"OF��$�M ���&�8A����"OF�ӓ ��<���X
%�����"OD:t�E?^܂h��D�-��Xc�"O~��sc�'m�tL1R#$\}��r0"O*K7*��82by ��]�3xJ"Ob8:��J�W\L-��kƴ~ ��c"O�+u�L�M�ހ"D�I�0��pq"O"�d�C����*�,L�L$Z�"O`4���]>��|��jQ�p�b���"OVhroE���T"���4���r�*OЋs,ƮLT�द�7PD�A�'���*��p�p
��E�����y�HʾH��ā��G+{�d���y-H�c�4h1B@D=8?$�Q��R��yrfN:c+�`�a��0��m��*I�yB.��<��`�S�� i�DӁ�>�y��A�_��(��Hk�D4�ц�yR��%>���b��`bb��y��Uj-��2���$٫c ���y銾ٸ�C����۞4ʂLU��y"�Ԓs��*��Ƒ1!�E��y�KE耡�ك� �T��y�툋&��ijw#��
��p�Ĝ�yF��r�E�8�b8�b1�y"L�Nv:�q)�&-�ޕ��Y��y"+Fj����,;6�:tV��y��;�����3!�5�����y� މ^E�X
�lƨJL�Ks&��y����)�TN;JҠ
�	�y�M�,�~����4K��8B�F��y"cY��qhU����( ��V�"=�)����0?AuM�AZ�tK�5�mh!�f�<�b�E3���I��@�}�*9h5.If�<�C'�8ǌ�+�)s�z�@�TY�<)S�$�&d�P(W�Q7���x�<��B�;<����`�.Zќ��p�<��Ɉ_c� +#�4�b��e�o�<�qh�V�2a�!�t��I��G�<���q�z�n\
�~��]}�<i�JTGzڕ2��, �2�(c��z�<aw��D���Շ�"}�9AP.Vh�<ْ�M�7���u�HH�C5IIP�<�#�����SԤ_4PAd�9�f�<I�)݃U��f�6�Ȅ��BYh�<����_'ni���^�0��bʊo�<���E37�L�R c�.<Q��NN�<�W"��u����Z�
�o�K�<�4�*L�b�(�v������@�<)6� a2�)��*Hx6q��jU~�<9v	�D_~���Փ}|6���At�<�AF�H�`��Gg�	m���Z��V[�<�b�̋'�!���ڏ}R�rׄ�h�<1���6:��B#�G�� ��Q�<1��իY�dX�
^!v0|uGL�<�AB	�%�A(�E�� rs��H�<)�)�M�uQ�`j�V����M�<�d��&�Ќ�t���s��(�b/�a�<qǄJ�V>4� �]�4ա�QX�<� ���T���"⎵q���*i�E��"Oܪ���/�"�$U�%�����"O���'�RBi�SMۻ9� �(w"Ol���M�u����ׁ'���S�"O��3�ƎM$�,sW�Hm6���"Oư���\�4֘����L:o���"Ot��Ș
 ���&�Z 3�Х0"O�Ae�J�@�B�"%�/=吴�"O@������.��eQ�NK���"O�����F.B�nd3Bb�"�i�"O��CЉƢ԰����J���Ya"O ph�-ϼ@�r�b�`����`��"Ob\��e�u,�X��9f���;a"O-)B�H��S�� a,���"O\��A��
"�`$i4(E��(��I{^P��鞗pU�8��J@ ZX"�)ڈ^=!�G���x��g	�1�ؕ"!hO�q(�䓽>N����4��,j�� �H�<���� �B��!5���ٴ/�>a(������J�}�Z<��Ъ=;b������S�M`X�<�'hF+<;a~#���L�h'���x��eپ#�h���b�Z�D%��O�ڸ��M�'x��xб+�.!�&�F|�)�r���t��]ܧu�D�SȊ3�ڠr���$ ��Oo(��Ԃ0�(3υ, �rEΓotF�0��1�Xҧ��6�HB�FY�\5�I?.J=x7"O���ġJ�c��X��P:�j���(���Ȇ3�h���'�6�Hp�əK;6��A��Bؔ� h� RIG -b!�C!��O�X�6ǒ�Gr�D�b6�|�ʟ#>����`ញ;�R�SU�>�/^\�K��W�.�>�;C�#���Q0Ü^ f5�ã+D�8aU*	�4 y!梘z6~}���@�AhK����'��}����p��Œ���//�z�ƢA�<���)D�(Ɔ�:wEإYt�?�'t쎸C�|Ŏ�[���\��	�����ȓm|s��� =�)P�MA<6<��ȓ.��,��в�n��C(G�`�FȆȓ#v�(��-�*7�Ũ�"�*��&�D��+Bf0�qk܊&���ȓdJ2<�M�"6a�� E�X���I1ːlh�Q8�$�!'=@o �`  H&>��]
ˢQ���I�t�t���p2Q�����Z�:����~³�,�0 '�X��f8�%G�N�<���]���L�PL�G��`1v/ �<��LM��pY��/}��)μ#^�Ah�ZG�dK�ō!�DH�1�$da��2;��{ф�.L��Icf��W���_��x�逮]opx00-���fY�����~���h���X�6&���q�P��bY	AL(N�\�+2'Śh���j"CL��z�f�<"��� S%İk_:X����С� (J(%�DL���u�'Y4@�'�ک�}b &Q-h�DRD!4d�5Yv�K���i��k�L���<���K� Ę���)Q�&q�����]%ug��˰#�6,��Dܛ8$�e2׆���)�:l\�1��d�+hQ5� ��!a��cv�@���%ЁJ�<BF+�:e�����k��~rb��x�d��T�=:�H�G������
�x| ���O \JX@c�^�}����O��W�LU��Gtpn��W02�n�4^=`tw��td� ��,bl��P ���l���`pa��10w�5{ӣU�_�.aؑO�y�O�S@������S=`▣��vI�}afN�!�Э1 C!k>`�Dy�CtL�mqv����!Kv̎���&��+�+O�%Rf�Z@�P�lL�l�Z��'P4�O0�A��.B�'�v�˕�2c�$q�O�5I���.̸���3`���QMC�8̂�QSdXӦ����	�\ႃ,I0O�H��-�Z����.:�Q>�	����h4�SWV�sr��38�=��,}5�9��4��c�| u	f2p�s���.���A�R�N�XF�W�t��Z�L1O8�+��Ll���PiO3R[8���'�� �dF�
��<�O�'=�@y�4�#��0J�a@�y<��'i"~�̝c���fB቏~T�0�&��O�4,�E�4{L�ʓ64�����8��99�㟕/�A+Ac�<���>�)�H�f<��
��RT0q��'+��p��Oƀ ��x���&s���`�>�N�*�C94���"��4²ر�E�!��=���'�,�iX+�'`�Ҥ�Yk���� �3�L%��{2�A��{�'�,*� ���	YU�Es�'��C��;/�4�燓�a���		�'�:E!��Uy�h[���.	�A��� I4&y�rh�+�(�&���K�ۖLc����G	 MXb"O�$!��	˦��ELɀ8�D�Ɗ�3�@���J�_Ŗ�I8�H����N�ap��o�|����_
[��B�	- ��$@�"��T�$%R�H�7$��
��&.�-b�#w�bpK
���£Gр#,�t���C**��I�;�b�Ȱ#D	;L�2`�E�)��5��&w8dP ��+\`��vw�!�v
�)eI&�������S�J![�@4ꈀ`��?ǀl�)Բ$@S� .�&"�H*�x"��y��x�.~��[5d�u��Q;�IQ�/�`� c��e[��hEkB4af�9�B@�$:x`օ�W�&L&�R�g~��=٢9 �[���������'4��e��
9}�Y	" \wܧ=¸,c`�3>8D�gjU!#x�-q�32&�s���|�F	�'^��0<�g�(�$� �H�8j$��G��'#|֠���̐蜼���O:�'$�y�g�Pa��d�R�h��?H6�R$D��e��dD�Xf�L��ɼRNB}9sD*)22I+�f�L�d�0�\���R�$���!�N��UC^EQSh��,> q`ZMj��'l�xȪc�A,W�͉!�E>���I�x�)$@�k�l���jǲ ���©��;��A�U���[�`{ ���%�³�_#����Z>uz�HN�Tt��'���Y�$2a7̄jč�({2܍�B�F�to^�is�Ha�d��O3ؙ+C��V*�#!*C�6��H�L b�����a��&�����2� (B&��/,""?��B���%�S/���yK4
�c�>���,� ?��Q���O�K!u������U+�Z�d�:�r�E˟Gy U���E>�8{Uo�0U��Q��'�(�8&NY$B����\�����o�D���1�C�]�R��F��f�uzܴ42B`@��_h��׍X��@aa�@-s���d�¬�0>�å��)n���kƬp�����-��^%j1�Ԏҡ4>�3'j�?8���uB�L� -R���0���Y�&�����N}���D��� ˀ�H�Q3���(Oj9�����E����Ob�Z���p�v�#̱9Y���G/lOH} ���:v��%�J�t��dC�xD~�-Ľ{��ѠB�s�h�KI:͈O����OS8Z�H n\�Kx5q���y�ܠ��	�8\,���ܵ0?Ը;0jMi�2��ě�L���f���2�@"�<�~R��4~� � �I��`\�ٴm�cXY���S�՘O�.Yr W8A�0hC��	9���'7����#�C�̲6�^�y V��T
�?:�$,��o8���g��,��)��Z�r�OΩ@��?�= $&êO�d��'|��s�ū�N��Q�Q�9�~���\�%�T�X�ԛ���c��(�����-d� ��Q��g��=�C���t�>I��� �@p�'uR<�Am��?9����EL��*�nV�?R�	�.8D��@C'^��ҤI�bU��,�>�����$�"}z�"Q�T5jI���t(�4ʄi�<Y�Cϸ>
�i(/T'G
n5��X�<�R�X?E<L��a�fF���M�<)�KT7�b�+�1�(��N�<A�*�b��_�"yn4��O�<YT+�7�,yv+,��0�eFH�<��>h ���03ފ���F�<�QE��U�\"���)�{(LZ�<q���6\N,�x���&w�0=��V�<��(�Z��D�!	�533\��%QJ�<��̉=S[@���Źe�����bs�<�'�
�X� ���G#&v�li��An�<� +�008�D�@N�P�ԏg�<�A�T�M�����/EAtv�9q�]�<�#O�/6z�x%��VYf�z�jq�<f�qMd(��O��0��F*�Z�<)�ȏ
�<p�'�¦yfBi�P�<��Ij��Щ�A�:�i87m�S�<)ǬQ�>�0�$=Ŋ�#@��G�<�&�>[PHRP���8L�TgUz�<���
�r��K����J�z��"�u�<�0B��6 <9&l# {L$�HMj�<�&��&w]���U��+[���rӫWf�<� \L�'M'>���1���d���j�"O�X�%	<�*��#Ǵ�{7"O��cB�BeGr��4M\�7�yZR"O,�K5m���� uCӛ)����C"O��9�`˼���2蟕k�ȩ�u"OH���]�JS��x�����؂"O�9�8ў� � W�O�:�b7"O�����V�(����0�M�I���%"Od��V�W�v)��nK&o�H�9b"O0��B�i��9b�ą
�ZBA!��YT"d$�n���2G��!�0.�:�BH�'/�	�,�KR!�D8Ud,���U��I�I݇H!�Ӹ$|��H0g��K�-"eJ�hK!�D�.d\�B[�k�����<5!�d��8�¹��C��}��Bw$!�D�|�x�֣Ёg�\}�7�	�!�$W�C�у@�Ⱥ`�z1��R( r!�H�fv�:苄Yy���iQ+!���8� �`�\�N&�S��!c!��)#s��C8-��bE�&�!��?;��-�GϘ;l;p�4!��!�Ė�3]�!�Ë_�f��`��Ɣl�!�d�RU�@�NZ� ��؍W!���7 �nуC.��c�~�b�� }!�$ݓB��D�g�I/���J*	?K!��>�&}c=`w,"��[�(A!�D�]:z���Fɯ�܀�0BĪ6\!���b��8�'�K!�ܘQ�H.;�!��:l�d��L �ĘA�D<!�䖅52��H���S궘�"�:t�!����Vp����<Є8cs޻5�!�$Զh����CDװ4�@E0��' �!�h�z��Mרw��u�Ua�<!�d� �8|�"R$^V�A��!�x)!��
�?ڍR�B׿hL)�P �.+!�[�X����(�UBP	[��. !�D|r,e*U��h���2/��!���^a�R�v�<e���ʻi!�d�*B센A�/�:C� �H�#Y�}o!�W��9{%�T��y�Ul^[!��ގ\i�\�1aP�gߜ��L�Tg!��W�%4&��[	��9K�`S�Q����ȓUI^X�4-��tOؽ��H��!��������珌�4�θ�V�>V� ��Uڢ��0��jj�G����l��h�zG�ʌQ�����AI�|���jT� �¯Oq��ˑ_d��4T<�ç@|��I#�*k)��ȓ/����f#�/� ]���V�R6����yP�9�e
P����
@��@���:��MN�GO0�*�O�z��؇ȓ���b���G`$E�Kԗ�\��8�.�r��O�c��ju�V(����ȓu�=arh�&a�� ��ȉJ��}����5�S-N�3i�����m�]�ȓo��1,C����Td_./{T��ȓ?�@�G�I�j�T�S�ȅȓ���'�$����'��6�R	�ȓ8 ��L�0�tH����	P����yK\8���K�|7�� ���L�r��4Ұ}"Wo/"X�D��L̀n�< �ȓ_!ZDPc��Lqt�q�lI'>��ȓe����#eW
�g�c�z���S�? l�2�oӥ#
�x�(���:���"OR S�F� O|n��ǃP���8�"O�$��&?:*��,�>��XP�"O�����"$;�q@�5<�<uh�"O�袁"�|�J��eH���HBb"O�MD��N�Q[�g�)OD%�6"O4B�,`�ڰS�#���(V"O�4��]&y�XH�V7JtnT�B"O�L�'�O�:s"i��A.`S�pj�"OJ=�ƣq�n�)���r$�Q��"O<}�D�R:��R�a��9�"O601��0@�L�0U ��Y���˔*O�5
��Z�K?�]�'bË_~,���'��y��I>RZ��(�ƒM���'�����F��Ħ��\:F,x3�'��:p������T�\��xB�3D�d9�'892����h�C��g>�B�I&7�<M�e J�hxX�� ��WdVC�
>�Εs!S�-Rt WF֝W�#?AV��	���?��0�R�R�B�!�ž�r�(�D+D���Ƈ�@�0!�C�Y�R�H��m���Ʃ���^�&��}b"�C�Ġc��B�N>�xzӫ]f�<i� ǭF�-RcE�Z)y�� ^~�h��)�\ ²�Y@8����a��x���yg&�O�,��c��&�9��K�-�صҐ�3r<�������Px��V�pG2I�g�*%4.y������OZɒ�nI%/��B�����25���0Ek��t8 �͔�y˭r���s�#�*6ܪT���y��>b4̙r�@m��8�&h�2�P	%:�i@+��GˬC��&��l��▖0���0���%ɾ�,dr5C���mN�����,6�@DH�`[�<�
Dٰ$=v�a~��:u]r��%fΚV�V�zc�M{�)8��K<`d�LeBUR"�/+j,��q@6+NDD|���I�N��5�Eܧ{��A0�e�����u(�,jp%��l.p+�ȥ<�1Q&���0'���oF&�I�	���S�Oq�Ȣ��A/x�X1�ѥP��@��'����4�*�h�'5��q�K<��"�"k���D��X�D��S� Tx��R��Py���<�� 3��)J��T�����y�ۆ6L�0z��^~B5Z�ꑌ�y��^-|,�i�D��W1hY���y�/B�|�ӗ'��YC���"F�y�K�� .��acޤ[䀤�Ƈ2�?Y&�8vN��P����j��h��H��44�����&])�	�c�����$8�:/(y��B���Oܴ��#jт��3�ȏ�p}`	�'�2$��Nޱ3
��s ��~��)��'��	���>��O?M� �E�C�g�C��f-��$D����3a�j8����V�T�K!?a��XF�(�2�a6Oz)ai,Q�٠�2V���S��Ob��"��7���%<ғ)䚕�e��p{�	y�A��(V�D9#���h�0�G8\O�@S��F)X'��9v�[�ti��@�N�nw����з��C��d��wcě���O|Л�K�	a��k�Ek}�\�O�P������4/By�z��S�L�xnr�?�rU���-�q��%k�n��{���@�1�@��>�|��X�P�"�WB��2��-�&/��G�l��$�r#��x��Z�j�V 94K�` ���OZ�C���q[h� T���PŐ�؂!�K/ d�1����w��%BB�����?�����1Z���I�0|�D;���O(�)E�3�j �I�6P��#<�&��>0�4H�V��P�1ҥ���%b�C�ݢh�J�0aE�!Xp�Px�>�O��钠*s���Ru#	 D��1Be ��q�/�#S�h$剁G�ENR����vN�$�my�@Վ1dL�'�^3te� P>N���e�##㖭�é�AU�C�L�to	�.�E���1Gָ�R�H���0$1�{J?y�|G��@�˂:0F�(���-���е��D�<�#�c�fR�"1hȟ(h�峟�	ѧă&�&�h��5r�^�bh#ړfL�I1 4J3b?�ҥ�<0�p��̌�&Y<��� �O\�+i��Z���P�%C8KB��� �]0��ļ#��1�%�?xӔi04�'x@�{�h�1{]z��O�'��Y{�AP�jF��#�vն5i��v`��٦C�> C�Iu�F�	�T��[F/�4Q�vZi�C��<*�La��2Qh��pA��<I���X��O4�8 ��[x����'��h�׏�#؂}��㐳	Q��(��L�4�Ր�O����/��T��ҥ~\P�k��I�Q�����S�Q@ ��%G.wv�<���ƅ
�nC�	S��C�%B!V��ôeG]�`B䉠Y�p �5j��'X���d�&y��B�	!�&�\�(	�5�	�r >]a"Or0���X*[z�dsŃ�#21z�"O$�"�P�H���%�+7�u��"O`t�띈טIW��,?�X0�"O��CTn@:�h�ۡsj�b�"O���r�88UЩ�AθM�F2�"O8쁔`O�].��f��2��*r"O
����߼4C��΄�4�͉��O�	ҭ?t$���ea�M+3��f��P+���6;�!��	9u��A��32ĢГ�̄ �����c�F���F��Ah<��#�4h@��%�d`v	�F�c#(��%�oޘ�%�+��/)��i{-�o�PQRbݏm���9��G6A�ax2�R�yӊ�Y!�A�zIV�r�F��U"�ɗ활���$���F��J@�8���I*���S�$�q����LϞF""���_r��yw���P0�����;�'	r�f�K���Hy����8K�cd+\����'p&�Kw�܁cb�YqB��;|fe�1�'vP}��W��8�쀇��p���NH�x;q�F;�p���v]2b&��22�ӧu��6�D���^��a�熽��!٦a�&u���ҥ�8���X��,�(�}��k�]?���$؝E|b<s�cB�p4(D����

{�8�2h�|�.&ā"$J�#�#?	t�tW��%�OJ�|a��ıB�IץI#Y��HЄ�O��`bӞ<�e�+�D�>
B�	���[��� �GA�,��|��$2\[~��D�:�X2���
1'P���'��¾i���
�F
9��I�'�PRE�inN��c���s6���*�B7
�#}�Z�!`CX��s�jN�,� �B���A�:��L9��-!�]�'�ɦ��
qje�O<����ڨO�a1�]w
�P�GȻ(Ϭ����-M��i��v�	�Y�ֹ��"�+|�i˅�s�h"�@�A��rᗟ��*A+
��1H��IY��YA�E��Iz,�c��%�">�r0-� )`	/}�֠g�*1��.I�9�p� �7#׮T�!�H���O��~c�T�鍝2�(E*2
��yƈ�k���y#*�d�d��k�4��C��kR�l���0R��A�R�Hs!�䈈3jF�@b`V�
g&� pCS�Kx�I��d������x�mU� ��}�1���(��U�����0?q�J �m��X��:n��Y�aD��f��P97z>Bቍ,�y���o�pp��@_�b��>���Ѷ����O��j�`9�R���`W��yBÖ#*u脙�nݣ�X�����Lt�X�{���!E���D
P�O"����!�D(g�h1�s���2(���$7�!��U%� 0#�����Z��&��!�dޡҒ�SPI��� @��� �!򄟛Q�-k�(�/C���a��M#;�!���:[�Np� M+{�4Z�&��E�!�$�?�  ����E�U��Z����
�'����*h��u����1Pm�u�	�'�P�Chyu�tx��$�$�q	�'�> ��;I>�-т�	 ���'M�sc^*��l�!����h�'�r�3D+�2T�~�H& ��Zn�`0�'�����2�0�zfH��Wg�Ԛ
�'��{�Z�9�0E
�[�,z
�'����dh���^	?�r��bB�yB�[]�,���۪6�n�9�@ �y���f�M(��A,��@c����yr��@Z�=��A�&it$IJV\!�y",ĒG��XV�	d	xDYv�X�y
� bt���ҭi��X-XY"O0��L�?6��Q�B�v��7"Oj��7fM�j��@���r���"O���Vj8�(��I3x�<�"O�����<���6e")\q� "O�c%%��F8��:0��<$�b"O�X�N�"�����Gϼᠵx"O�q)�鎳k�`C�f�$Ѵ�ك"O~���_O�D	�0
Ȥ]�"OJ���Ɏ�J��b�	�d���"O��J�J�@����a��TWJd��"O��0��T���
)ڮW>���"O��*%@i��!�+E�HC�!�d��.���ĕ�iQ�AQ�D+0�!��VF�����L�Xs��q�(̟�!򄝄sk�1+�E_�\�H��	9u�!�dX�j� �F��FY�H-��L�!�D�<akӨ�)0Zh0���TY!��Ӂ]i��q�O��/� �"ξ:�!�$,g��!�	JՖy(s X�5!򤛥����F�H���3� �4�!�\(��9Q��� ��oɚ*�!򄓈aW^}���7�,�s��Ɓn�!�ժ�N%0A��2p	(�m݆*�!�D�N�ژ��(ݸ��ek�В !�I&"���rW�=k�Xd�G��4�!�ğ-��܊�ߟ
��f߈(�!�d�M��Xa�$l�8��GŒ+8!�J`/:�8�d[�d�u��@�J!�l� �X�.�:?[�50$���+!��&F��(�p-oT��$ˤ^�!��<_����*H�DJ(���C�-�!�Γ=w���DF�<J�	�RA�1k`!�DZ�fPD�Ae�ď���iT��;BP!�$�Al��D[)s?��@��"i!�h�ؤ�_� USɌ8nC�I�fԱa-^�`�Z�PlC�ɽlJ�l@D;I� � �i\C�	��b��ڳDj���b��-�^C�ɐ=�a1�O1-��`#���+�xC�ɉ
6���L�X�<P��d�fC�	�nS�����/O]�x�%G94�hC�I��|�KƊַi���6	�(�bC�	,�4�Xd�&��8s�e�?	�C�I�jt� ��'�+��L�r��YV:�ӶɁ^q���d34�P�e(�>��<rcj�V�!�D�7��)T��k�~Qp���)~!���L�� �قt�P�+D
`�!�D�~t<�8�RթT�V�?��M�ȓn_�ؘ�kݮx�I��-H-��ȓaQ�!�#���8Kܘ`��2td �B�Ό��O��	j����m]-������P+*����P�x�g�!VUd�á�|ʟ4�����y�Iɿ�-�5��?���LK�A�'��<3�'n�O��#T���Z����:�&TU$�5J�+�yB�XPdV�����?�����e�~�iFfT+Q8IxA�ܼ����2�\��i���?�9� Ƙfb|�zP����e�`*:�y2�(,U�!K�����	çH:t��\R:԰����;�l���HTA�kZX���}�"|J.��T"q��19Ĵ"�T9�B���`����a� #L����;+a�		3Q��T����"2j�% �7'��4�J	Oi�(�0��\�y{���t�S��,��s Yl��q��W.�q�`��9�˓_�`�çYw���t致d/���6��U5 ��egH^~�M#'�hD2K~�O|n��b[<�2�c�)z`.�����97���]�ꅱ4���ҧ(�<Y2j��pH��K!-��� �W�<�\Һ�Bh�m�)�'w�,��씖^�٩�O�c�­��S�? (1@��ו]VE�@��,Ry�\�W"O�� �%m����"�O�\��	R"O�5@6I��>����F� YC��p$"ODE)t�  �@E��$�1:ٖp�e"O ��Q/�a��U�'J����� "O���V�P�1��6�<��"O�����z�
m[�r�:&"O��8�"�R�1:�d��W���J7"O@�0��=D�v�4JZ<��$�#"O�,�w.R`{��i7�WY�.�f"O�%��\���eQ#׶A��"O&p�4��	2�N� ä��G�蕓"O��1�u�.��A�V"O9��Ȓ�X���<BQ"O|��l �P&��I�`�:~����a"O��7��X�z����Q�4M�"O�`� �:/ZQ ��W� w�T�V"OL��j��}#��2g�0�"OX��O	�%s���0 �1R2=�d"O:��q��@:mI� .@�v���"O4���D��fc��p��RO���[�"O�q����1)�Ji��XN���"O�1����|1��(��6G�pR�"O�pA�g��2��
G�?���"O��c��Ҝ>�xZ�h�K�H��"O\�V��Bh*�"���G�!�"O�y�&@Ȫr�C���"OJ���E�8�0ت�H&u>>H(�"O>��Ƃ�L^�R���\���j�"Or��$Y?j0�N[� Fd��"O�M��HY�Wr�	b���Y���P"O�LHTȍ7$U, a��ޯsB֠Z�"O��YDm���� #�0T*�t�"OH�����B�`�𠆏�<��"O2\iF��8��u��OM9,�D��"O�9��)�R���k�-��D�L9("O����|���+�!p�X�"O�hpO���R!�'h�jp"O��0&Mߵp�n]��ET�K4>Х"O�Q�J˧^v�p��E��!F`�t"O0����ܼp�
�4fêdکk�"O~�a�5�J�Pa��_n�1hc"O,�s�ۤVT����X�c�r���"OB�Ck�'JR����!T� h5�"OdX	1�Ͷ/�f�9����~�YR!*O�U�3AF���� O�=$j(-I�'�ZP9�a�+T��k��,$Q�t�	�'8��Av�{���rT�ܖq���P
�'5��rӎxe���Ȋ4H`���'��@�gR?x�b�dD��ذ�'�d�	�P�ԭ)��~.>�)�'�$��O��� Qc�S~@P|��'x��0L�ӾA�s��}���'z�]�a����0�lS�n�@��
�'q�h3 ���H��U� aA�N��5�	�'4T�����m�z��@H�B�bA!	�'��IRH�"��ѧ�.��(�'��8놬V1~^ �'�)���	�'�Rذ�툕e��-z�eR&*Qa�'c�x����g�`�����`�X���'��q��N-3�L<YsA-\i�q�'�A���]"q;\iq��DY�N�)�'��y�*/Vi�);�	��D'̙H	�'~n���N�; i
Ĭ=�$���� 4M��snX1:���:]OhXR�"O�� GI]=&�Z�%N;�d "O���"��PA@�(�%��6��YK�'(G��	
x)�r��t0���'���*�Ô�2b� "#�4hHI	�'90ઓm��I���C#�ۉv�9X�'���aBB�b��<��K-:ɮZ�'��QhD�Vh����R�Z�"R<Q�'��� �+�9�ʸ�"腘&�DL
�'��pA�̦6 �\3�$ޅ Ґ�I	�'�0d�a#08y>�CqO�:kZ
�'�Zar-�"d@���fD;-P���'���#����ٷ���\c	�'>8xVj@9GIP=i6e���p��'�4�2ȶw���P��Ը*�'$���C��E�!�g��+x��Y��'����B& �h��ǅ"��'�&�F�4#쌱@�B�H��S	�'>�|`dL3h0}{V�@ D�����'I��c�h�2B���0��"Bڌ�Q�'�� h�&)\N�Pc�ؕ+*D��'4Lq �`Ɔ"&6�X�B6r�Ƽ��'���*sN�2U��v�\7�Yj�'�=;�gjO��*�L�!�4 �'ۂ�4�ғg������P^<;�'2d}ÕZ$G�2�k�S�-�@��'��1��\�:Eh� ��$5�8��'u�m���
S����!܃km$Hr	�'�(E���B�(����![�`��	�'��QeaJO�d4���6	�(H
�'���3`��V<���P
�' ����!��,��R�څ?z���	�'Jh��ҍP�xԀ��
�LZ�%p�'ޱ�Р�
Q��'�Z�mBP�[	�'�zͻdg'$iX��P�8���2�'7��P��3B�=�398=�p�'�X���/U�^Q�3!%7*��	�'�m�CKиy�6�H��^!|<x�'�p�k�⑧_��m���6ph��A
�'�v@���>��㦅Vb�2��	�'��T���5$؂�qsm�Vt�q��'�B ��]b/ˍxx2Y��'c�d�Ĥ��|��g���Fg��h�'�H)�ÎH���� ��+A����'T�f�ǯlN�Hx��:F��B�'�҄�`&X�w!�  %JL68Y�5�
�'�v�0��¤���I6.F��@	�'���2w/C"I�֑Irm��,x��z�'R����;f�>���d�1*�:=��'���C�/�L�+����R�8K�'s����]z	J(�W"O
!�4K�'^��G�t������4���"
�'�qs��@Y�6	B�Jո-�9a�'8����H&$��ɉ刚(t��8�'l`����R(-� �7
���
�'1�u��D͊Iwx�֛֡X;�\�
�'᠄�G�9�إ8VCӛ (fh��'�H����]��$�E�ٰu��<��'�4����7\B��%*Q�m%�b�'s��P��A�H�U`_�i�v�R�'7Zᒰ��E�z( �T�IV��0�'��	0���mi4���'�N�,���'yrm�!h�,~�RT�	L�j��'+��!@�Txt��Г)M=rR�i��� *i��� �y^�x��F�>CP�G"O`j��_zNT�kEf� &��"O�ps ����������7P�ސ�d"On]#�)�
H#5C1�G8f�j"O�)	䓙�\p���S�,S"O湰�h�<����VH�i"O��a�&�V��p�'Yug�A��"O���`�a�>ٙ���Mojؒp"ObtQ!��Q��,*�D$b}��q�"OZ����ДJ��*$�C�8e�$�w"OVA3��ϹP�*٣!��.c�	3b"ONXۦd٦x$�V!=q���"O4zQ�Țu&H�2�N+,��I�1"O��Β�_�>u��.��E� ]+R"O��i��2@���h6k=4d�	z"O�L�%/XE�X5{��mM��`�"O�U�3W�=Ԍ�#u-(���"O��J�ޓ�f��a���C)n��C"O�}Q2�UpN�ᛢa��T�,T1B"O@�j�*�f$�� �ʥy	-�3"O���	Z ^� e��'q�$�"OZ"��M��%��B�?��I*"O0��Ў�0�D� �C��[���
�"OY��{K�H�`mۨ�<�K0"O|mcĲ$!��(�	�$Gl�H�"O�س%�N�tTH�0H�!�Vq@"O���LT�w�$yR��j�5HQ"OΩ�ˎ�^@@r�(��Z���x�"Obx��/EH.xQ���H�N8�"O��U�@�آ3ĆB�[s���S"O ���3��A�Ř��Hz�"O��#��0X�ډ(�B��~�s�"ORp�$*�-�Bq�T!� E����"O��C�B7"Ϥ(�6�Ϯ(A�"O.)�2�H�^������Ґ�\`�"O p���2/J�a��흦a�>M�"O�<�s�3}�i�SNǈr���9�"O��`�l�
<�Q�!R�>���&"O���f-�*�4a�\,ej����"O��Ȓ�[$g������ţOɌ��"O^��r��]}r퀆 F�����"O��
f�J��"�P#oj��=1�"O���!%��t)�<�4�Q94{���p"O�����ܑX���ktIL�Kp"Ob�Q �[<d�����]=C2�`�%"O L��еp� ����7�X��w"O荘�%�W�\<����0B�:R"O¤pS��5n3�#c�|)�"O�@6FԻ`wZU(gce.� ��"OV�H�N�X��Y�BΐƮ�!'"O�|�S �&
�}Qs��Rd"O�$�6�)��#�o�S�� U"O$3&f���%������K"OĔ��L�J����c��@����"O4��	Fm8$�Vƒ�j�c"O���T�Ifi��D�,1��L��"OH�
`�-J:Y�ᜐv�����"O��"qg�z������xľ͹�"O$*%�	u$X��σ�|����g"O������Vo��`�#K91�t��"O��J��S���a�� (��Q��"O|] W��6Y�<!pТ>tz�Q��"O*4:��3r���"��ד?X�(��"O&\#�C�-�"q"��eI����"O� ���6�eҐm��]+P�8@"O@��%�ՀK�����I����g"O��`��#���RvƘ u0p;b"O���7�� �-j $�A�e�"O����N9Cx�B���3f��k�"O�iw��")0���g�3>$i�1"OL���G	p`K����R��Y�"O`�H�d�)�5fE$Z6�R0"O�i��̈́�c.F�3#ͻ)6̰�"O� 1�no��u�D�¶M�ty"O��s�	   ��   �  �  �  �  d*  V5  �@  �K  �V  �b  �m  �y  ��  ?�  ��  ɝ  +�  Q�  ��  �  e�  ��  ��  G�  ��  4�  ��  ��  %�  ��   c	 �    �# �* U4 �= �C CL �U  ] Cc �i �n  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^�+���������Q��_�P��I;Tf�����a��3�i�L�C�I:V�Ł�
Ӥ<��
�f9��C䉼R��Ӷ���a�f%y�ϓx�:C䉢G�"P�͍f`��{QK�E�bC�	� ڦIAVe��y�$ �`N?hŀB�	`j4��f��W���d��"C��?0��C��|̩#�]�z,����>9�k['	U�H���#�~X�V��C�<��
R�2��*6a�#" �]�q�z�<���%T���2��>�&պ�Uu�<��Z�},L�TTT���Ze��e�<���[7 �:ӧ^��D�Ej�{�<��	�4&�Faz��. L:W��px���'U6��j�4{HIi�J�=<���!�'@�<5"ށe�L@�B&?K�y��'�AC� ]�h R�d�2v|3�'�R���l�2#�{��L"5��`[�}��i�ay2��L����kh��պ����y�C�@Y��c�o2bX<�ْ�Z��į<�K>���U?��X&o��@rJ#@�g%�1P�'W��4�� �$��򌓈2��Bu�=}��'�6䲓k��_�,���펫��t�	ۓ���w�\a��G�r(]�~x�
�b D��*�m͟&���d�-p���cѤ>}��Op��S�O�.�@�,��(D�(�Ɗ4p{�Z�'q�&�ĕ۪��fh��e�����C?)Ց��F��'��-C5��9ND��h@�	�0���3�'K����KW�("4#���Qb�	��|�h*|O��C�3e,N}�ڕ���>щ��~��'�`�PuE�nb.� � 1B �
�'�~�re�0̖y�P�	0��)A�}R�)�Y�s�2�s���O�Q��a	�|n!��<J��AS�ϴ6�2��aP��1O|��dA�9�#�'�65�nd�q��v�ayr�	��&5��=nv!��&\[���y��'�A�E"4x����UA�|d�(��'��EIO�Bc��$GU,{ ��'k�8�*�I֚���j��{���y��'�,Q�߰n/������Rщ�'�*q����� �C��h�eO��� �=Bo�]��nJ�$	.���'˛7O�+�h�d���Q���ݾ+0���ȓ,N-��B�����FhdZD�>�U��$x�����[f��Q�+R��pǦj�<)�ʂ�a�(q���¥c�D�bH˟�͓�ا����`Ԋx�L	{�,���\�bL%D�����+ApbC�;`�����<	�S�? ����-ϷQ�<=Q cۚtu���O�u��D��^kr�[p�W� v~�q�K G�<���@�B��H�fD�?T@x��� Y����>��T8B8�b��4��(�t"�Q�<��/��L1��*��7X�*����<���S���l��J���髴AT�Q�B�IS���4E�82"�[��E7^���0�S�O�ʜ3&��^]A�T�W��@3"On��I��L���򭞠,�jPc�"OԐ��b�>ZҁC`�N�>�X���"O�A��P�޲�$f��Ѩ�y"O T`�*O6/LLI˰E�M���w"O���Pk�*ˈ�Jq��X�)Є"O��8�,�/f�P�Z�.
�:H��1"O(�D"��2},)T`΀,���"O|-A$YO��9�v��R���9�"O� X2eb�����,�I�4"O0|sȐ�H�tZ��L5x�"OFÔ���($J��1J�Vb4��1"O6��DfC�Z��Ƙ_G:�Yu"O���eP3*T��p2EX
n0*Đ�"O~�%�#�Y���G`��"O~�@�h��x�sc�0b(��"O0���l�) "�u�۴-X��"O�x+�O!�̨���TT����"O�%3�	�1�V�q�-ӼVb��"O2��"���!T�F:wG�,�"O.pB��/E��c�m�@0��"O���d�7�^ #',	�w*�L8@"Or|{Ӊ؍6Q���<}"��#"Oz�X�:^KQ2fkD���˟��yr�F�c���F��q���@�R.�y��')��(2��'l;JX����:�y���S.8h�ČM��x`����(��,HG�׆%���X�`� a�Q�ȓ{��2�h��a�!�Q5E�Ta��TJ&���.W�8��!�9����I�D�˳+�|�4����Bо�ȓa��(:�C��(�+ǳ!�܄���|6�ڰ]����`�
"���ȓW�� ���*P�	��*&����J՛���U�Rt�K��f��\�ȓUn�p@���Q�4�C�	��*�� ��K��ѡ��ml���7��gN%�ȓZ�*���!���YF��La�s��i�(P�t��+M)�l�ȓ[V�Tav
N.l�idZ
!� ̅ȓz��%�ttQ���WB����ȓn�
��Ո)cW�;s,]�/�̇ȓT&��cK99JyK���1Y��ʓsՈ���m��y`�U8�j�8&RB�	��f�y�@K�{��c���*J�bB�	�i&0p��Х�=^���(��yB"M�v݀�� �\=�,���"�y"�T&�9"&E�Us~Ȋ3�^��yB��>/�-y%n�?G@�@{"լ�yR�K0�r ���@%��bf�"�y��J +�n Pg�5/���J$e� �y��'::��! �ܜ"����s+��y�◜f�x@óⒾM.����I��yIC�d���I�X6�; %�:�yR�)6|�!v�Ӷ%�L|�흉�y��Q�WH�q���K����y"e�:�ؔ#�o��`J�b/���y
� ��K�cд� ���&W�4��"O�P��_>(ލbV!�0sy����"OP��ƃD5	�# ��wb��q"O�����:�Yj�.ăzO ���"O@)���>bɖLz/ԫYN�sE�'��'���'���'��'�"<xŀQ�6:.�1�dJ4S���1s�'jr�'���'���',��'Z��'d~D�ǄI�H6:����T�C�h����'s��'�r�'[b�' ��'��'��|����Y���ڥ����~����'a"�'�b�'���'���'r�'¾}B@��m�thg�r�Jf�'�b�'F��'j��'R�'���'��E��/��z%9E&D�THX�'���'�2�'�2�'�'L��'�T a��S[;��S�%R-5d�����'er�'a�'�R�':��'nr�'k��)�f	�s�Q�F�|p�����'B�'��'���')b�'V��'/�q�ݳ9�Y���z�2`��'9��'���'1��'5��'�R�'�DA�逯 � ��a��>ċ���?����?���?��?����?����?)'gٕ,�5�`�*EF5�S��?����?���?����?��?���?���.zvZp�g�SIh���)�?Y��?���?Y��?m|�`���O���܍}�Ăbi��	]�pĭ����D�O����O����O~���O�lZß��	�1J�u����nʡ �	�>>��+O��$�<�|�'5�6m]$Y6D�/J-:�����zfV͙�����ߴ�����'�Z�И�*��l�X��F��g?�<��'��E�0gA�v���Χu�4�~B��%[��HA0�<l�@�"�d�S̓�?)-On�}ʒIJ� ���&�"e�,0Y�D�����_���'X��oz��1��	/T�Y 0�OlU�m	'�U͟����<ѮO1���P�/oӊ��x�f��R��)����F�?`J��I�<�"�'`��G{�OF2�NA,Ё�@�Z6*�Q$@:�y�R��$��!�4z7p��<)�dRH���˖�E_ˎXI��1��'���?����y"V����a��%��Vh�'A/���`�5?����a���Q�'������?9�I� ^����*T�+��A�Ԫ���Ħ<��S��y��S�9`�7>�x����"�y�DxӒD�՗��x�4�����L���}�D(AA�ҩR�K��y"�'���'F�T�оi����|�u�OW|@�ϐ�s��7�R�,:$!�Jd�	hy�O�"�'���'����=�ځ(a)*Q��+e�!Y�	��M�����?���?�L~Γb2���O6�����.ݏo��X�R��zߴ)�&-#��)Q-e��KRNK���;��Ԋ �f9�&-�=8��ٿ9F�hƨnҾ�]��?�@��4
,OR�a!�J.��CB�i������OJ���O�� ~1�5�N�<ن�i�BDy��O��P%/�u`D�A�0-��Q��'�6��O�ʓ�?�W� 0ܴR��V�'��U��O�Sx~ib�g˒$fĜ�Q�˛�4O�h���'6b�;Ba�4���D�H��ݿ냋����ܻ�@�>o�!i��<!	���4������4hhR Ñ84�����?���N,�����˦q&��G@X��i���F�K�И���ē6��FGz��iņ3� 7�;?!1Κ�o�R�0�@F-w���H��ۃdd ������&��'��O���F]��i�D�7������I+�M#��@�?q��?�/���9�g�!-@�xp�Џ¦�B����O�m�?�M�f�xʟf��Q-�#l��p��
�eC��w��ʁ�sӎ]����PO?�H>Y׎ʹG@�@���&K�v1�2(�u<��iz}��<pn$<�A���J�m���S*X��'(7#�I���������.s��IG	�3R,�k�"E��M�u�i����a�i�������AQן~�=�pX��,ه� |�r�Ҋ6�����$*|Oi)��Я8{�����#z���̛ݦ��tN����џ$���y'�	�qY�\��iȊ�
FŽo"�6-[ݦ�H<�|�)�M��'�i���B�d�Lc�.�*�l�a�'O*l:���u?�O>�+O�˓_����Ӂfʁ#�����U�ቊ�Mc�cN8�?Y��?y(M2`�r�ȶ.O~Y�Ђ�&��'j�/���bӼ8%�t���#`[�G��a�a�Cd,?������ߴE�O7����?��.�Oy���ؠv����b�<�Y�Jm�ĹŅ�#5�f������?�i��Hy��'��|ӆ��݇J���!� #W\DbL<�I!�Mt�i��7mU��7<?��n y&��<�Y�C	@�&�ȥ��(v��4&�Ԕ'�b�'R�'���'̺���q��4S�A2j_��0BS�0+۴z)ZU����?9����<�w!�k\���+-�d3R��z��ğ�o���S�^;�,�n��Hp���	�xIa���0��� .��J��O���I>a*O��hT��P4nг���?�X����'��7�� �����T��l�t圉7H DAN��<�d�Ц��?)�U�@��4yx��!{ӆ!��ۺI��h��c�����(��~�6`����?iK�ӟ^ʓ��{�? �l�W�F��ҥYQ"��@�X��=Oj���O���O��$�O��?�$c*%!���X���X��L���@zشkϧ�?y��i��'���t�F5��.ޒ8a�|��*�$�����|�'K�
�Mۘ'��L� ��
L��br�O)K]���6,d"e����,&��6�+�D_zy��' ��'�Ү�(I���Y���#5.��$٣C�b�'�	�M����<��?�(��I���o�噁�G�/�$���� �Od�D�OV�O��G�\Zef =|V��N���<y$�79��xm�P~�O��l����!� M��F)/�A���(��I���?����?��Ş��B��Qsph��L�b,�����DyS��f������A}��'�jH�rcK�`�^�s '� K�8!��'<��3؛旟�ز$�1W�q�A���fR}ʓ�e_��01O�ʓ�?����?!���?q����	�3qv��h���A�E��2�mڶg��	�	џ��	S�s�Б���3'�U�=ռ�I�$Ց�F��$&J9��z�Z-%�b>	�sm�Ϧ5̓/�*Uj�̞d�4�A������ϓd̔H�&��O0��I>�.O�i�OB��:G��"%��	�=0��O�D�O���<��i����'��'��dx�R�N�4-A$t�m0�|��'���?����tӴ!$�`�e��[ⴭ��O���p���|�d�	�Y(�0�-�Ҧ5�(O��	Z0�~��'�(p�S"[�j��u�,N�q�9ȧ�'lr�'���'��>��ɇ(��a�U�H�`�"z�Y�I��MC�AP��?�FW��|���yWO� -�a��H���q�P�T�y�@|�­o5�M�Lج�MK�'�r��NU��k�t�@�$g,��ӤC�D}�L>�+O>�$�O��d�O@���O$�A�1"gV� H� ��A�ĥ<鳰i*B�"��')��'#�O*2���R|Vn!1c��S� �<=��b�6�h� $�b>!X!腨c�\�T�/ڰ��EcC&@J\nڪ��-sr�'V�'��	/
��
�F�<[��&����؟�������i>1�'�6-·w�$K 9F�����m�Ȫb�X����e�?Q�Z�����H�	2	f"����x��H�b9���'��U�'��u��|r�;h,|k�)�F�L�Q��E�?�<���?i���?����?i����Ox��:4A�j��by��)y�'b�'{6�6��I��M�K>) �ҧ���9�GЁJ��ecҥ�2�䓚?a��|*�� �M{�Oț�I�$- !��z�8#����\�nHr�'��'1�i>�	ݟ��ɐgc�͉SE��Z��5[bϯo�8M��	�7G�*��'��7��"�f���O��D���ND�)X��R ��m��<���O*���O��'�"�'vɧ���'$x�"�ԈT�B3���?5E 0��42�:���i��	�?����O��O=z �M]�F���-n�����J�����O����O��<�6�i��`"fM�t�x����v #ŕ&`�	�Mˏb�>���iT$�y����c�ˏ�l���u��z�֭k��dyb|Ӕ�l]��^*�T�~�80�����!4���<�(O����O����O���O<˧L٫%e��;��=c��B?+ݖ@IҲi��qU�'���'��y��x��n�V��0ɓ�2��52���'~@F\��Ӧ�IN>���?=�
t�Ul�<����M����ጨr���'��<�D��R��ߡ����4�(���>S��q�<f�ڽ�$�.���D�O����O^�fO�&&*C���'�R�	)2FFd�����C�](�*��f�OB%�'�D6K��QpO<i&�μvB�W`K�P6�2���y~���6���c�G����O�������R�Q�T=�A�Ӈ�'�����$�j��'b��'V�ݟ��Bǡ20�P���8��}�� ܟXK�4s��y:���?�S�i��O�Ύ�qÜ�� ld�Q���!��������4n՛���#?J����d�6
W	F�I�ni�PA��+��		1�l�K�m*�$�<����?����?��?�Q��7�.)X�K�H��][!���ܦ�)���˟���ٟ�%?�"!\u��i	�#� R6�M��!�O�m��M㳙x�����#y�f@
�G r����'$L U�X,j��i�2˓#a����ⱟ@'���'~*�`�J�#��Q�'ױƅ��$O��'���'H�OI剆�MbG�?�w�+H
1�i�&��@KU%�<���i��O8E�'��7-զ�3�4,�����LTR�0�	��'�4i���F�M+�O�L2��H�������wHԺ�M&�,@FlE�4��'R�'���'3"�'��2! �*�2m���ˉzd� 7;O����O>Hm�$q�d�uۛ��|"b��;��ڴE���yãńi)�'�����R�Rd�����G�6 (�R&��q�]��x2�Q�OޒO���|���?���j�b�	�gj�QSdCZ6A: j���?�+O�YlZ�����?Q,�>ha1*�+}"���e�Zv$�v��|��Od���O��O�S":��#+ӥ����aY0f�\)��n'Z��lH~�O�j�����Z��}�e��N��3"��^�B���?9��?��$B��O_剸�u�*�<�Z�Eʒ)�8�!V��#P�DXݴ��'f� *�6��4��K񪀶/�n�R�K�"�6�
Ӧ����	͓�?���E
[���}y
� �	9po��\"���f�Con�H?O|��?���?���?	���iϚ:l��[!�ȇFF��3���
~ZmZ%j�f�I����_��83��w��e:���u�6�H�H��`�]+Sy�|nZ*��ŞdKD�ߴ�yr�ƴw�`�2���z�r�p�M��y�+>�i�������OL�R�xh�1
�	Rv�0��,Z4�$�O����O0˓O`��h��;F��'�Rf���4왂l� �.�p`�C�n�O�'{��'��'F*m*pa�* B� �QF��gV�a1�O� �qʛv�*����i���?����O���c��z(wHK"9��i����Ov���O����O�}b�W��b ��o��8hHM4�T�+��vIًn�	��Mӊ�w	t3�Άr��,ɷ�h�d�h�'x�'�¨�M�搟��A�����e��y�$��7d��{0�S�脀�pc>�$�<ͧ�?y���?	��?�a�/A��-��n6R� 9#1#�0��$\�Q1c�y�h����&?�IF�>u�"�q��T����q#����O����Or�O1�X�7}.��CÓÄ�ˀ��y0�6�2?	���zK���e��|yB.��\Sf̐-#��I��E����I�����ޟ�SIy�oz��B�1O,����I�{~�1�X�q��y�?O��m�m�#m����x�Iǟ���FE*h�"}1��I�2�i���ۄ �4�oZ^~�Bn,�E�t�w�H�T(���Ā�@�H�b�i�'���'/2�'�bZ�b>�@B@نI�V���ĭ��X�Qx�t�	韜��4��'�L7-<���+L=L�S"^-½�f��S�Z�O����O���Y�>7�8?)��_�TD� 3���Vp�!�n�� .cT����$�(���t�'%��'���fGP0?A@	���O��5���'ebV��
�4hO0Hϓ�?)�����fB���/�$�D��"�[A�ɱ����O.�D5��?IR �Nq�.x�1�L�MH�! �	A$����AƇŦ9��d͇X?M>a2/ 9I�y]��)�+%L� L����?����?��Ş��D���]��jT�\b�t �`ڕ"TTŃv��.Y�D���ǟH��4��'\�ꓝ?�[�6a
��a�ɬ`Pj����?)��,(6�B�4���L�,j\z���@ԍ8�1w@B4�1��ܦ�y�S�h�	ퟬ��˟�����O0���e&V�I�@��K!k���+c���A� 	�Op���Or����٦�݁X�葱6�Ӌ*粘��fF�V��	ɟ�$�b>M����禑Γ	���Z��$_p�+
�=���E�4@�Ǿ��%�Ė��t�'ǈ���#O	+��1`�E�
=p�I�G�'xr�'rR���ڴ��4����?���{��!��	W+B~^�ۆ
�0�p��b�>���?�N>!���))%~��d@�7<q´1��P~�� op6y#Ӿi�1��h��'2�(N ��u��k����I7�y���))�� �a߽]��r!�>a�b.n��d�+�O&��Zɦ��?ͻ�ƄS��9�Tru!��P:1�5��vg�ZYlZ�-s�(nZB~���"K�d��Sl�$S
׻]�����W�d�TpO>�,Oޣ?A��7��@a��#���鴧A~�Gy�N�z�'�O����OR�?�@d��W�\�r�'×x�6��_������ߴx����O������J�7� s�2�|a �Ao-�v(�<a���o��	t�Ivy �"�ya��I���8����YS��'9��'�O����M�����<�v��`�����H٘u�w�M�<1��i{�O��'Q"�'��M�,i�� �*!:'̘�����]JҽiL�	D2�ۂ���H��9R�$<�C!�%lf�8�c����I�G(��V�	A�,w ��q�T����	7�M3�\�d@sӺ�O~,;��
�=R�`́{x�ѳF��r��:�M�R���t�U�v���XVGՋ��\�P �"�����_0��� ��O
�Ol��?Y��?���(A"Gŗ;�Ebt ���M����?�(O��nZ7�"��Ɵ��N�4oj���H0��!B��!б�D����_}��'S��|ʟ��5�^#km��b���-Bh�:�どj�~��1�o���|�租�'�|Z�蝉z��m��Á\_�Ի��&�$;�4. l�PWk]?B��)`ď]NP<�! ��?1��E����}�g`�"�&#iR�Cɨ��<�o��{ю7M�즅��&IҦ��'�d�P1b�i�-O��9��J�4萩ӓ@�߄�P%?O�ʓ�?����?Q���?9����iױs2Hz���^Ҫŋ�O�3ڭoZ�Xx�������Io�s��!���[��Ԕm'�9� (*��x�"�ɾEB�i�O�OQ���G�i��?����S�M������ ��D�)d a��dК�O��|2��C�ph��շ4�x�H ��64<eC��?1��?*O\�m��4b�IП�	�/z��󂁂(甡q���I���?ѷQ�����%�4���R�R �[AmY�{ !#��'?��B�2ZV����4�O��D��?�W�C҆U��L���L�"�t�<���Y�܅ʡo۾(�$�QMY��?�3�iY�5�W�'>�n����]�yX�= �/��7Z1XB`F�X@�����m��M�"JV��M��O(�6�� ��� 
x rk��;ʅ�&G� �Љw�)��<i��Dɏ[`$��
�tK�,��K7)���)�M#����?A���?���ԇ]4���m��$�"��!�9s��?2�fr�b&�b>5�d��%>,^�E-�8&�X�Cp
ĮJ�=lڱ��D�: BQ��'��'��=+���ՈŽ_Xnd8�$�t���	ߟ�������i>ɔ'P6m�|��D�S��"�f�( L��2֮�I�����I�?�s[�\�I˟���:C	�Tb��;{�x�:����{� a�#B���'�T�B�O���\�5]�}���Q'9���RO���y��'
��'���'	����-.�h�[d ':�@R�](+��d�O��撚�1?i@�i�'�f��0	Q�t0��R� X�B��ӝ|��'�O���cU�i��I�.�2a�P���@C�kC�Z��K�jN� �$:���<ͧ�?9���?�@C?[��x�É=��x�ɕ��?�����$���Wyb�'�ӆP߬y����&B<�g�as��J��	�l��u�)��$��z}�k�iD�j5�ͱ��L9	K��OH�n�R���Di�џ�HG�|b�A�n�J���j�^�kS�Ӄg��'���'��O,�i�w���	��MS����H܈�@̯P>�-c4��1�b���?ᑳi�"V��*��D�O|}��E�$P�������HQ��;2��O��$�%�6-w�x��*Iƺi끟~�����L�?�,��v�Џ.�J,�����O����O��$�O��d�|"�O��W%�ap�@Ҕdհ���H9כv� �l��'����'��6=�Jqц��au�)�2 2z����צ9�ٴ`���O2��jӽi9�Ĕ�9����t�H U�
����T�'��$�׼ ��J�O���|���9:F��B��4V����%�</B(�����?9���?�+O&`mڮqO���ݟD�	�A�X� ����j��$�1��p�~��?��_�L
�4gԛ�'񤕡V�|d�tM�[D k�HX7���pe���P�X�)O~�!����	2J�"��rH�:[TlL��,�% �X�	ԟ���ϟ �	y�O��B�&OVL�!�dP*El��T�'B@qӺ��W%�On��ܦ�?ͻ���[�)Q�>_^!ɕ&מG��Γ����k�t�m��B���m�G~�͚=��������V�[g��%L�e�K>�-O���O��D�O��$�OL�X��[8B�M�;bR��95K�<�׶i������'u2�'���y��E	p:�	��>_����_?J�n�w���y���'�b>�Xp�V�b����c�#-|��ruj�=$a�+��7?Y�jðwI���/����C&����C�.v�@��Dd[�a��$�O����O��4���1����_��ybÁ`ː��n��N��y22�V	�y�j���C�O��d�Oz��fB�)D���n�s P�1��o��A}�(�G9�'���2��3�������4䪵ӵk��<1��?���?A��?i����7�,R#'.+�� ��µ��d�O�mi���>y�6�|2ߟ9�̙�����<����R(�'����$Ԡ{��������aN�P�l�2rNN��[�)�"�D� u�O��Ot��|����?y���h�0��m�@X)Dˆ�&�6����?Y.O6(o�+}6���0��R����3���v�.��� ��$]}��'iR�|ʟ"ՙ��;Ѹ}9�ʊ����FR�z����wӌ��|z�⯟\%���F��X`�K�aȚ5�*7��ڟ��	�4�	�b>��'s�6mV
FIv p D(<���A9w;��S���8�޴��' ���?!��;1~J���%Y�G���B5Ɯ�?I�{��i0�4��D��a=h}y��TIO3N-B�h�g9J�+�N&�y�R� �	̟��	ٟl��ӟ`�OS��c�oٔ8㎈��ڥ@k^�sR �$�7O�D�O�����ͦ�"���׊�>k��+uj��2�rh�Iӟ�'�b>m��I�E�)����K+���2��ӱ�vΓ>t�S����$�ԕ���'��Ru��W;�|"6eUѾ��'T2�'p�\� ڴy�����?���c����FF�]�8��m�u�Q�R�>��iӸ6�w�%⤙A&�K��Ш*�B�'*�@�\��e*�T"!�|u*�O
!9��{�<��D?NHʰ	��-<�E+��?q���?Q���h�����<$J��C"Q:b�d0�c�����¦u �b�Zy"E}����];q��ڄ(f��ǎ$i� �I�L�	����G"_⦱�'��	��iZl�E�&B5��3��F�)������4�T���OH���O8���*R�Cs��m!0K�FX1x���������y��'hR���'�и�Â	S+�T3B<v=,�1V͢>Y���?�I>�|"Qi/]�D3�e�'5�tyVWO)Bu�ܴ���Yo}r�8�'��'�����3Z?b��XA@#7~�����'2��'�r���V��bٴSvU��>����_uL(�"I[�|���r�F��Z}��'YB�'�T�!��^Tݬ���$��	�A���oP~�ț��V���]ܧ��+��ڟ��Q5��59�^0�CCC�<q��?y���?���?����̍;E\�Gݩ\�T1�udAm�2�'|��p��PY���<�#�i��'��kagʷQ��9�o
M)����|��'��O?`�q�iH�	�Z� dE��6*�sJQ���)4%$�?��"!���<ͧ�?���?y��Iv�|��F��!q�p4�,�?������ϦY2���0����$�O���xCW\Jܡ��<$�0��O���'���'9ɧ�I��4����ӿl�֜��Ϟ%�) �*߶+R��F���<m=���Z�5{��H&���S$�Ace�ƃ&�.9�	ݟ8���T�)�Sry�d��UM	�'e���3n	�\
�]�S�8yԒ�D�O��n�x��#��Iߟ�@ӣ�$~�ܒ��5>�!���ӟl�ɲ,���o�D~�I��(����M�I���h�b��E�3������7��<a���?����?����?�+���3t��n	>�x� Ęu����C�����ǟ��Iߟ��C��y�4`72��#*�� ��Xc�`P r�'�ɧ�O���0�iH��JJ��ÇEצ�K�k�h��ԏ
0.xx��A��O"��|���҄���0(��Q��v�=���?���?9.O�1m�8od���?)�D��"\�|#�$�<";`e����'�<듒?!����
�ܩ���}��`�h�B��,�'��E����)�6��]+�~B�'����Qg�>Pר�@�H�8=�"	Q��'(��'�r�'��>���T%�Y!'&C�:D�C Hp��	��M��-��U�I�?ͻJ\�ą8ac&d�3�A�`d"�	����ܟ�B��
���'s��h�L�?����ԏ�9[D�� �<�:�KH>!-O�I�O4�$�OD���O�嘕��%e�X�c�-P;C���<�'�i�fQ��P� �Ik����p̃x%�"&Eǖ/��@��.���O��d'���_d�%��芅0+(��c(�)V��}{�.M�~d�	S�����'��X%��'Fd�U/I�YL @��Ŗ89<�v�'���'=����4]��شo(]+�J��05f���P$4S;hΓQ{�6���X}2�'�b�'O��#�K^�X8�%�?[2B��4K\	s֛����Am7�Q>1���gN�#��ڠP2(���B)�	����I�T�I��	t�'F�Ɣ�d�9"�� 	�(sf.�y��?���(���� 3����'t6�*�J@O��G��*Q�E��G�Z<��O8��O�	��7??��Փ%^�S4Ô0d��U�����5k��b���$'������'<��'L�q�n
�@�#&�\:\0S�'�b]�(�ٴ@䪼̓�?Y���I�"E*$�G���$��`��XY�I6��d�O��#��?��@�Xt�ar"D0B��{�����O��%��tėw?N>9��V+H��Y�$��n2�B�@�?i��?A���?�|�(O�mکh6|�'�M�
ܲ�;'���A��{DDgy��Ӡ��;�O���l��N �D؍(�fp/�����ORԹ�oӔ�*[�91�䟶�Ol�}���-��d�L<z|D�:�'�����0��ϟ,��ҟ\��K��(>��zB��/M�J��V)��	׈6͆8mN,���O2�D0�9O6�oz�yR���U�n�G,�>�bd��o��?A�4b�ɧ�'E�`Xٴ�y��+<n�9@�:�۱��/�y��F�#&1���
�'�i>�	,%�VQ�RHA����b� T�h��	��<���P�'��6�[(IA�$�O���
�,8p��X	e����� S���L٬O�0l��MK�x�.�"m9A��^�"����K�����=D��4k��ϗPy1��0+��Zy��D�0Rbp$S�Gѿ}�!˥+R hL�$�O<�$�O
�d �'�?Y�j0�dPR�IݣQΐj�)���?�S�iB��r�P����4���y�b��)���kH73�Fh�c��y��'��'����ĵi��	���d)��O���b��؈A�U:�L�NC�p�G�n�^y�O0B�'i��'��'��y���K�Ei�:�	�,4y��,��k�
 *��,$?!�ɑE$
��f�-tڢ���I��DǶ$��O(�D�O��O1�X%�Ht�<���)u�	{���RP�D)Gg�i~��*z����I�S�'�則(i�s��p�`��3�� �&5�	��H��۟��i>I�'8�6��U�:�	�q<R�	�)Qe���2�Q�|�dUܦ)�?)�V��I�� �	���pA��?P��´�VI�� �`�Ц�'D$A�s��?��}j��j��U���]�f�1s��J�"a�g�ԅ�	7ڦ��G��6�^���ǖaCj`�I�	��M��M��n�j�O8�x���*|���i�&���O�ɨ�Ms0���ďC�9��V��d�я��X����������m��:�Zp���OO���?Y��?��c_����IC�hKs��4*�(����?+O�o.�I��؟��	W��D�g��лE��6,�(��%�%��DW}"�'	�|ʟN}7┌2�1��)���yW��'g#�Ǩ~����|zWL�� '��PԀ�rv����^8	���1�Qß��������b>�'xL7�H�OV�y˖� ?M�h���0#w��jve�O�$���?��]��I-�12S���I��-�ub��(x�4�	�<�Cɦ�'��!@��?����`2�8Z��a஁3l.��qu6OJ��?���?���?�����ɖ&F�����)3�����B�+4@��n��#��\�'��������w��3�┴,㪁{��͹`kߴD�f+��)�V:7m|�� �##��9bS�ɺW��r�	��1O���3�٬�?�!�>���<�'�?�vm� �֘iBBDlM�+L��?����?i����dL��8`������⟸хO�\xz�;���[�`��3"�x��h�I)�M�`�i�lO�9B"霈.��}`���a��I�P� aE�:-Z��*�S��������K@�<-����$F��n�����������t�	П�F���'g*!�E���h d��:Z.("��'&7��?�Hʓ4��&�4��0�u"��7����� [[Jhs�5O�Pl�<�M��i�p)�q�i���� 
���f�O�N��ŨA�[L��1e������˃؟ȕ'S�i>���ʟ�	���	r'd|��O��]U���2�GN.4,�'.7M_><��O��d(�9O� � .t���Y���	�t����H}r�'02�|����j�~�	�eV�6⼱(�d�6|�\���i)�I����z�O����<�-O6�3��9���F/�]�XP ��O����O��$�O�	�<	��i��D���'|RA�GbΈ?-�3��L\��x���'!�6-%�ɋ����On���OhL�u &Q�zp����-GH���ʹ~!�6'?)e�֪|�|���׬̢��0wO����V&��Γ��?�pV2P���#��L�����"��?��?q��i��˟��l�s�2S��P�qO�+v�3����$;M<)u�i�X6=�D�k �a�$�g���Fg
�7Qd�[b��2<�x�$"R�gu���@�ry2�'Br�'�R�ћ	^�P�ǿ]LV��W!L�@i��'��ɐ�M��*��?I���?�(�� �FY ����a���tpA��8�)O��DpӖA$��'K~�����%� �;C�I4���G�/{��[޴/�i>	�#�O̒O�A2���.BW�0�/�;q�( jFi�O2�$�O@�d�O1��ʓY����Y�%�$�ۗ蒃�����A�P"�'��al���DثOX�o�|��`��I
U�nxh����7����4�����(��f���h��	�U���<��*"у�2�( ��P�<�*Or���O����O����O�˧ot��� ބ+P��8���.�mJ��i�T��0�'�B�'��O�2�c������ Eo��Ev��2���doډ�M��x���?�v7O�Hإˈ�TR�݉f���x�2�8O���#Ŝ��~R�|2^���	՟(TȪD�t�Y�U1-e��Zeʍ���ʟ��	}yR�t�, Ж*�O����O��2�`iN�")'\��+ `.�	:��dJǦ��4u�'i��	�n� D�F�;��Z7� ��O�q* qD6m]H�S�@���Oh�	�	V  ��IWj�);�=� ��O����O~��O�}�;b�|A`�}���s�� �8k�-���i�s��'� 6�+�i޽��Ȱ x��DF9n�8�������Iঙ�޴`�.�[�4��d\7�M��O|�X*f��'-�FU��ֆV�0��T�|�V������@��ПT�Iǟ����	b\P����INY�!�Sy�|�>��c��O����O8����(O�ư(��Ή��С�IӣWJ|��'�J6��ݦyrL<�|���ϥp�����Tm�� [aLݶ�L#�-B~��m%(�I3�''��4} ~D�UnոgU����g�������������i>�'U�7�K�7Ģ���9miHi�Ӆ�)Yzh�i�+��Ĕ���?A�Y���شA����|��D��"F!�T�8�Ɋ]X���E?n7m%?A���#3к��$��߭�"�J&H�41����7����q� �Iٟ�����	؟���i�
xq�؀
���p��+�&�?���?�b�i9:5��S���ݴ��r�`�
��� Foa)Dfaj�� ךxR�l�Ġmz>Y�O�¦��'�X1H
�n]*�R"h����հ`���K�p�	(%��'N�)�s���U	+�"`:��U8���t�4���vdӀD���'�2V>���B�o���0ĝ4s�e��L>?��]�d�۴b���;�?Aҷ��,��a�nV0i�s�X%}�^�!֦B��+O��O��~��|�$F�@�L�ЫF�v�桋���3�x��c�X�:`�R(BIt�)@M��T|Y8��H�"��Ozym�`��YF�	��M{�i�!Z3X�YV�̪����3���g��vKfӚ	��Ns��Y2���F`�?��'��A"�J�,[��BeN��-����'���y����hZ�2����E�-�<�`�	�Mku���?���?����r��N�' -������6�E=m�Ll�M���x���+GA��V8O��aA�E��U��G�)r�ъ�5OR��`��~"�|�\�����`���G Qq���5��ܡ!�����	ݟ���UyrBgӘ1�tL�<���B��+�m�8K���rrI��P�ص	��>)�iV�7M�e�ɱK�ȅ�Efݺ9^	
�%E�?��wsz����y��|B��OȽ2��*�)C��"�B"��|�9B���?���?���h��n�C"�`7爬
�8Z��@x���Y¦}�3C!?)��i��O��$j���q�g�]�xQ�������O6��O��3h~Ӿ�=^�����?�y3�X�.r<iQ�ɕ5�x���]��Ty�O7"�'e��'A��"=,5��/&��Q�������M�U�P�?i���?yI~�+b����G8�� GlШBXJ-�bQ�`�	П4&�b>�f):� 䰈2â.54ِ��Ҋ��}�d��-k�I�/�� �'Q�d$���'uv�Ӏ��p઱H���?9�V���'/"�'~�����P���޴&��l��-�^�B�fՈ+��Z���NX��v�&���[}��'��'�R�Ӑi�,�"�A6o��"z�T�M(����!� ��T�)��r�m_�d(Q����(C�9C43O���O<�$�O����Ol�?5ؑn�p<DMy�D �U���vf�Cy��'�7�O����O�\m�t�I�|g��Ӏ� ��Qa�L2���%���I��擳 �1lA~&�5^@�A�]9c�N����Ŋ9Q������3��|�S��������ߟ 1�D��3_�,(�S)S1����G؟L�IIyboӐdɰ �OB�$�O��'F��T�։{)�E�E� _�}�'�b��?a���S����1��9AƧOu8B��Ci��U��dT��O�Q��?�t�.��
 ��ec���b�04-�5���$�O���O ��< �iUJHBb�![�q��8�LL�ӉH�$5剛�M;��>��j
��9�D�d�.!!"k��4b썡���?�D���M��O�9Z��6ʸO��	��o�.�
�:��/
�Y�'���ϟ$�	����� ��w�T�[�K�4�G*�#��q��#c�7-Q�-�L��O:�d&�9O>�mz���!��'{�=`GHrOnp���M��i�O1�0eBf�r��ɚFr�����;g�2� v-1::z�\ �ċ��_����$	��U��D��R��-e��)[�И��-SJ|��!("��Eխ�Tອ�u!�2aJ1C�	U�j�٠�)�7gc��r&6�x�IV��`�j��$̕r6��&��<s,9�Lӊwھ0�gf��g���AF�e�$�(mJ�xi&��F�]>u<a�v͐�x����V�1�^L����9��dHӥ�	�2i#�lǡ#ݒ�0mG�)�hQ�+(���[���N�	P��/�	�i�&/|��z�% :�$��l�)7>��I�m���$ �V�^IÀD�?bP+"�:�6�O��DC�^��уÄ�Ɣ�g@	�!�LnZ۟P&���',�y��}"���O.�H)��\�5R��t���M[��?(O|���g��Ο����O���IAȀ0,
��P�4@p�u�N<�)O&ѐT�~�N��IE@(��\���q�d��M�'���T n�-�O""�O���m>�yJ�n�9�ni�p._�rԸ�oZyr���O��X	��̨7��,Q��'l��Ժi����u�p���O2���&�p�	&uۀmy�@�$B��#ƅ��p޴*�Dx����Oм��� B���A��>��Q���WƦ�������|'T��H<���?��'���z�-ۃ 6T�M���d��}b�8��'�"�'/b�P�9	AlXSk�sՋ,:6�O���pjc��?L>��:܂X��d��X�^��4�$Q�D��j>��ן��IƟ�'��)j�A���>����?Z��Y1��7V��O��d�O��$�<�*Of`��@ߒN5tH�c鞼�pt,G�Lg1O0���O��d�<��d��h��ɐ)Ѥ,��F�e����"װ{��Iǟ(�	~�	Gy��$�����*�jd�p�Wm+�k�"��{��I͟��	��ؗ'�,�##%�)���x:�_�b!�G����n�|'���'��蠋}"�M%}��  ��jE�h#��$�M���?�(O2�"�O~������S-}����I%YFl�����j� �N<	/O�h��~B�JМ-��,�e J�* \ç�����'�F]Xэz��M�O2�O��,�R��7΂�aCH��G��W0�-oJyBcN��O�����qo�=�P��;e�����i7&�xӃm�\�d�O~����%���ɧx$Y�#B�oj�Q*Ɯ�Bxzt9�4z�TtEx��I�OF����K;%��W�Vx{L��f��}�����4)LQ��ǟ(�OGB�OZ)i�m[�b4��2_�@�d)�aHJm̓ 
�Q���t�'#��'����;��3��	k�e2�k��扑Yw��D�O�t�O��|�C�5� P�.�7�0�D)� /�Oڜ���� ������I�t�ɿb�6d�7gA;��U�ǈ�q��p��c�RyQ����V��ޟ���B00i�]�u�pa#q3S��nڹY�@�?����?i���?�� �"��䬈�sqPqS�,q��t�U� �MS���?������?�.O����i���3�_5gQ��0A��+�0�O��D�O���<��N�i%�S��3����1�2ѡ���؜�1��ۇ�M�����?��x�H
�{2���cU�d�UÁP�E��,T��MK���?�+O�@G@q�4�'��O"�Q����Z���	��-݂݊��"��O����6a����'6����a-M]�lIF�*@�^\l�zyrj�0R7�O��D�O��i�j}Zct)��n	�~1T���Tp�ش�?���]#vHY�b��� ^@�B0��8oK��x��9K �FDǮX� 7��O����O���`}�T�4�P̂\J|)[Tȱ�ɋ��x�4Sr ���䓎�O� �%E�F���Ȏ\.H��L�+�"�?Y��?��& ���{y�'#�dY�Gk���o@)efy��.��f(���|"a��P�P�d�O����SЙ���M����7�U�A>�=lZ��������<)�����6!�9n�N���b	.gM������[}"BbY����֟���ey�ؕx�Xzf��l���1�aR"x 0�M�>�/O��D>���O��DG_�? ��P���-��&S�z�	�So�T̓�?	��?I(OzH2��|����3@7�Q!��|���B���%�'Hґ|��'I�d��-j�˙=&���������0�Е�ڥQ����?9���?�-O$�����f���'���#��2(b�YQ��<0�0|��!hӀ�$(�d�O��d��"��dY���k)B��ޚ>:�U�`�r��D�O�������_?���Ο������0��������#^
b���L<���?����?�N>	�O��@�P/�t��5;���D!��۴���1!Ϥ(nZ۟T�I���������*1�s&%J�IK��A;�����izR�'Ith��'��'�q���1�S5 b|��i!����g�i���k`�����O��$�� �'C�	�)��eB��A
Ff�y�(H�%����ܴ�QX���i�O!{�K��I�L�;��1�>QԏR����ȟ���5�q��ON��?��'C�4���˒$�D����F�xI�}B��'B�'�B�'[�HB�c�Y���E�FǤ�eF���h6��O��+��ET�i>Y�	K�i�Y۲L�v��hCB[[����&g�>�c���?�/O����OV��<��f�gE$i�~+zQ�w�P+��:a�x��'�B�|�_��S@F_$l\4[�gK��\� �z����yyb�'M��'��	l�> ��O@�*r셮$}�m:��.}�	�Op�d�Ov�Or˓S�H��AE�����ݣ�.8�7J
�'��� �X�0�	��IyyRk��'@��0S1�N�2J�M�!���kC-�����i�	Xy�F�H6R�~Ӄ 19���	��(n�L��� ]ݦ��	֟x�'Qj����8���OR���T��&-6*�<U�Sj�?��8�ՕxBW��h�!���%?��'b:�[u#S���e�@�ZmGyR��(�*6�@P��'���"?��M*>�~���AR�HH&�Lզ��'�8�*�'N������)�F���H���a˞4���M; I��?A���?����b(O��F%��j�H��8>D���߼yAZ-aشyG����(Xw�S�O�Z<ZC��@2��Z�).-��JS+tӈ��O����Zhh�S�D�>�a�y����o�Ԫ����Tf�1O�}3WC�d�'�?Q�'`-귡�<xÔ���T�M�۴�?��ؒ��$�_���DQ�*�R�y��M7V\��@NF
G�J��'pV�R-ڸ���O����OfʓH��swʑ�6s4�xC��u(�s��9��'�"�'�'��ItIܰ	�$��%����p)�Ft��1�d�O ��?��%��tH�-��#��%U�6��Q��4�MK��?��r�'�R�8,�۴qL�S��W�l�i���U
v��'�D�	zyr�'��}K�_>E�ɍw���0��+a����$X���%�޴��'H��'G
%���-�ē {҉bqe,t.NM� 훖#S(QoZ���'��K�=��S�L�	�?�X�(5)���/��M�(Oj��Or勖��Y�1O�
������>>��J���2����?�`���?���?���2*O���*� i! �Zﶖ?�8�۴�?�X��,�x�S�H�f�����@a�YK�/Zj�4�mZ���{�4�?���?��������_d�B�Y���Qa��6��$�����O(ʓ���<���,�Њ���+"?����L��Z<�58��i@R�'�҄�./pO��OX�����	��ʄ(䩂 ��XB6��O�N�`u�R?�ß��۟\2`�˯h�F��R�̜Z*E�p���M���(�Z��$�x�O��|�+Z�#�pqx�!Ӻ6�b�q!�ܡx�0�6 �%1�����O���O<�7x*� ��Ɓ�r"�)aox`�r��&��'���'O�'���3Ԃ�;E
�z���3�KK78Wz��0EV��T�'���'�B]��S0�ׇ������$L��n�d�&�JP�%�M�(O���<���?��c)d��I��a怌8��`ƋC>��Q�$�	����IDy�e�$~만?i�`�!��\�.H�G��pj�v�m�ȟ��'���'"�I��y��'��L4g�(l��%�1dP<3у��ou���'Q�\�8{ �	��)�ON���U��R�6�c���(fB�`D�_}b�'/�'���OZʓ���Z�e,J�����P���L�M�/O��ّj�Ȧ��	������?-�O�.�G�4��(�\� c�CV� ����'����yR�|��I]d�n�a��%v_0,c�;���M�(5�v7m�O����O"��n}"V��C@�|863�進-�.���]��M�����<.O��$$�ş�gL��52|�/$��L�
<�	*�4�?i��?���9=��Iyy��'i��K�-����1- �X��`�OϏ#�&�'3��'�иq���	�O����O�h���`1"<8��?s
�i�EæY�I�:S�]��OH��?!,OJ���4 �㖃q8Թy��G�GH\��iC-�<�yrX��I����ayA	b8���重V��]S���,t�+F�>A.O���<I��?a��M�=��	�*9�9#�M�hʀ�p��ZI~b�'��'�BU��Ee���t��ki4Ո'�}�d�u�?�M#)O��D�<)��?��~�R��cƣ]><�*�@�/��k�঑��֟��I��ȗ'J�E��N�~����W�D���§T	|�>�z�@VѦE�I_y��'��'�`q�'�S�? 8���EH�.T�	����DmR��5�i1B�'@�I�l���󪟐��O���At����D.S�Q�X%7F@�`��'���'���ɼ՘�y2ӟn�j�ƀ/���1t<Pv�xR�iL�ɥF��e��4�?!���?���P�iݥBn�5l$��0���BS$�c@i���$�O� �:O���<��l�9M�6YY���1>�c!����M�n��D��'�2�'��g�>!/O�i��aj��h��aF�X�a�H��
�y����Vy����O��Ps߅i�prD� N�QdVȦ���؟���1�,�O�ʓ�?��'=�E:�D��\`��V�e�4`�4�?9���?9����<�O��'��������O�.�i��ݠH>$7m�O,�)��Zu}RS���IqyB�5)�`�00'iN c.ڭ�S�^��M#��jF��̓�?����?��?+O����=v+v)���L�d��Y�@�:.���'l���'m��'
��'U���Z7�-Z��}�!#�v�L���'��'��'�rP��0�݌����%MZ��7lYq���т�H��M�,OH�Ĭ<����?)��`���L�x�z��ۮM��+�eO�e�E�i�B�'�R�'��I���񑭟z��������(X��#�1iv�iz�Q��	����QZv�B�D ȷ(�IH�+OV�K�̄�^�7��O��ĩ<�`i	�sI��џ,���?}P2�#��'�y������d�O2�$�O��?����΋z�TH�"Ğ�H�l����ӄ�Ms)O���r�A�u��ɟL���?ѓ�O��%7��A����`yN)�3J��A����'iR�[�yb�'m�p�'z>5Qa)��"WjAs�$!5鼹n���.�+�4�?I���?��'��Ihyr�	i��xA G�^�`4��r�z6��!2�<����O��Nu�rY1GA�S�@�`'��i.7��O8���OT���!e}BQ�,��`?Y�C�M���I0����QC �_ۦ�%� :�ok��?Y��?��gʰi+��X$�P�tm�TQ`Ĵ��&�'��I���>)(OD�D�<!���2��:=i�l:B�Lb�\P�	����I=5�D�I۟$�	ӟ��Iԟ��'��Z��Ҽ��j�g4iy4!	a(���D�O�ʓ�?1���?��:2w�}A�X�E��V՝AB���?����?)���?i)O���a��|*��Q����{5��r �idFVԦ�'�2P��I��\�	�8F|���1s#�>J� �Ǆ	\/��nZޟ��Iҟ��	uy�j� �'�?��Z���1��
X�/�8؞�l����'���'����:�yX>��%�\���1ZG��?τi	���ȟ���̔'2�"W��~����?���N�Ve��
T:R�5F�:n���Y�����,���IGP��j��'��)�+���G�s/\Qh�˖;�vU�ث��� �M����?���ڷ[�֝3x��0�ݖ ����T�ESn6��O��F7����M��'q���014�.� ǃ0;���1�i7�(�։}Ӟ���O����ʼ�'v則�d���<�v��hL�tn�ٴ8�\��?�)O��?���-L@���ID8q�����N��Msܴ�?I���?�a�	���Ixy��'8�d�6�����&58i�ᇏ����'�Ɂs���)J��?1�6�,�a�^b��l���3v�b}jS�i9��<m@ꓲ��O���?��G��u@6��N �4�$Ѳ5����'�v�c�'������	ڟ(�'��� vH�V���ǀ�>���U���`�����O�ʓ�?����?�'�A-�fa�u��+�l��lF�2�Plϓ����OB���O|���v�O#���L� �0)(���VV�V#��M#,Oj�d�<)���?��� 0���'ʊа��A`��@ b��ISᩯO��D�Ot�$�<����k�Sܟ԰��>A��MsU"��|�$��Kݚ�M�����O��D�O���9O���O2�M�K#���V׀5����iO֦����'j�%���)�O�D�m��	�07p-#�eѽV��Q�&!�m}��'���'�Xy�}�����\LL�D�N��qɴ���I�/�Mc+O�d��K��E�	ٟ@���?���O�n�1s��G�IY������e�v�'���
��yҐ|�iS6�i0탹`W<|��UG�v�I�-��7��O�d�O��)�t}"P�x���A&#���y�lƣT�QS�����M3"���<iL>ь���'�� 9�e7^�4�7A�,]4�u��x�,���O.���2V.'�H�I˟�r��ʶ](�vY�&J�.Ug:-�>�u.S^��?���?�+69!T�U�q��t�b.Gi���n�ݟ��'�P,�ē�?y�����F�{�(̳d��T� 0���d}b����yBU����⟼�IUy�W�ljH�z�ɸ\H�@��@���&�4�D�O&�d0�d�O$�D�MB���)S.ֶ��ɋ��X�@4O0˓�?����'#�@P"�3���@�ɚ�O�P�7iA�vU�%J�\�h����'�l���|�!�z?!U�6;$��ׁ���8d!TjVl}r�'���'�剂S�80�L|r�-�[�2d���,�4��Q*(��f�'c�'Qr�'�dc��'��|X{��CY�0�b�ɍ	���m�ğt�	]y҃�,�������2s�F�3�@�B0Θ�E z�����@�����I�f�܌��i�S��B]���z� ͮ���5������'���Fx���O��OL��%�L(��
����`�!;�X�l�ɟx���"���Ij��p�g�? ��0$%�5o�*����&+e(0�G�ipv}��yӞ���O����,9�>	$ř�E�α!P��#�Ԩ90ƈ:]���T��yb�|��I�OH=���D"o)`)KÀ�"pldZa�զ}�I����� ,�J<9���?��'���@�Go��x���<]����4��Y��ӕ����'�"�'6��gF���p�i�
U�]^̍��c�����0L���>a������gގ_O�1x�M�8F�ԂbA^}�.�f��'���'��W����J=6�$`��L�0��\`��з^�F1x�}��'�'��':d�X��x9�����%\�8�1%��y�S�����X�'��������^1+��L�)E��(���$f���'���'U�'���`���ʄ@g���7�_8	������D��@[�6�iQ�����&]B�~B��(�H�p�����b�B1b��M���䓝򤅤4%b(#��x�d�/Jx4c��O�P���-�M;����D�O�##�?��	�0�Φ}P��[�p�� ��V��,���xR^��3��J!�c��eNL��q�G6���#&� *��o�Iyr�Д�V7m�OX���O��j}Zw6�X����
E ]�F�/R.���޴�?Q�b��ϓ\��s�P�}��O�z��.�-z���R�E즥!+�=�MS���?y���rS��'@�� b���o��- P�H8<����gu�D��;O��$�<���T�'w��$�رP�b��m��
2��!G����'���'6��0d�>�,O�������%ʌg��i0c[�8��ɰ	o�F��<9�D��<�OB�'���>L*�� ~�"S�C�IF���'��\�C@�>�,O~��<����D�Öb����7_[j��1�̦E�I%���	ϟ�Iɟ��I۟��'4B�*T�� �*8h��S7@��jB]�����O�ʓ�?	���?�0�L�_)��P�rL\��T�L�x`����Ot�D�O��*�`��C:��0���gO�M����.\����5�i���䟬�'���'�ҭ!�y��O�<��8�G�pa��q͘�U�<7M�O���O �d�g��ួpc�'�bk�c:`���T�RQZ`���cP6�O�O�$�<q%��I'z�U#��~�N��)"R�iC�'���1.4�H2��2���O��IK9ye�,:�{���b����	l�T�x�>�,���
�K�e�������;zt�m��d��Qd�<�	Ο�����?�1B�0�-�9gg�P�Ӧ�4nRr(lZß �'2X�h����`�^:��:Ǐ��L��lH����Ms����?���?!�����?�(���n��6���.<�\�C��GI}BF���O1���ڕ_���H6"��8�Ⰱ�3%�^�nZ埠��ǟPi�&ӕ���|���?�bH�xzx����s��@y��W��O���'���O����O��� F*GZ}��k@�u�"u����@zE�'�@�'�?	H>���R���àj��L ��D]�'f����O����O|�d�<Q�"��	Ԍ�t'���bT��q�L.���?�����?��0� i+*ѐs�1�
FERV��I���?)���?�)O�t�3Hfj�)�?3�4�E+ �T�!k�>!���?�M>)��?�pO�w}�I>���r���(u*�4A��'�2�'5P�@	�eP���':|Lt��
S�`��h�2�]�P,�ҹit"�|��'u���*��',&	��g�7OB��)�G8����4�?���$�:�Tq$>��I�?I��LË��r*&@/�J�$� �ē�?9��Dx����6&��2!�!��!!M�e�s͗�RHE��d���ǆV(��Oa(�O�̩(p/���K�@��"%*O�\�5��f�^Aq�A�/*�@��3���Yl���vk-��B�֍0G���D[�u���1#C�%>�0mh����E�0%XCH�q<z��C��d6�xq�]�?E\�{%�)7 aۀ���E��FC�]d*m�<Sx\���Z�#+nY�S���,-ifm;*��g��DX�����Ҷ�'L��'�2ft���	ן� 49[谵9�j�6E��1�q#�=J���DQP�Y,�����(O20�D@�?�p��'D�%L��E!���L� ��+ʇJb:�Å�t6��D�'����6*��l��E�3@� }�d�:�'Fje����?a���<�t,R��YH��B�:��e���O_�<	��7F��,��fn<x���4O���'��7���lZ�� 9A�Y�?��+�e�Y�\���П�����P�7�ݟL���|�G�\�O-h��I�'��c%@K	C:d��FD��K:XX����<i���)H%z�i�N5c���	��S�^b���N�x��:�����<Ѱ�N���I\v`�B�!F=S	8L���o��D{2�ɴ3�|MS� ̖�.[��^�?�B�	�[�j�2&��#G�٢DdG�M?�牔��ĵ<a��_
(�����O��T��lR�`s°[v����� �(O�2�'���Q{b�0�%�^�D  �L�O�S�h n���A�OΒ��%���P���<��M8_n.��&�@U�N|���ʺ)���f�T8\6���S�':�0����?q���#^���q;��aOP�S�@��y��'�N�����e��Ju���0m|������� ��פY�
јH�`JC�rB���0O���Ήt}�'��u�L)�������7C"��%�^�ER�R�=B�H<��d�f̮�iW��7"�`h�S����'��2�͘�o�~�s�gC CQ��3.49�R���)˷q�3�#�O?���~꨸��M<.5;�mO1;K���n�O4��4?%?E&� j!�Fv�*$2�N�.#�: �2D� ���l�D҄��B�[6i54���V��<���'nhd�$hx1*"�����	 f�8=B�T����Iϟ@��%�u��'�B/�_v:�a�/��BbtQ�+Y+o�<����܄+Հ�!�P���hOV��UDE?�3����
�f4�ЬX%^,�ty��+D�ԁ���
�?���ɖ(^��X��	��@�ie.ю��	�OM����O�=I(Ojdcs�F�";tP��oė(Z8=rg"OJ2$�$3�6��'I><�x9H^���i�<�����p��h�
V;��9�ѨD�8�`!���B�'�2�'.�ɘOr�'��e�f�%�(dAl�X�ft�s�P�4Y^����ߩ�p>�'�KV�h�zva��l�;�.Q�r�0��o��E���gW0��Y�ቬ|#l�$�O �iP*�R�2��E勿_4��[Iئ-��gy��'P�O�	;$��BG�7tV x��1W$��>�ųj�|��)�#:��,�2뒼_0�d���bܴ��D�1Aʄm�쟠�	v���1C8Q��.$Qp88�	�ap�P��'��'��yU�'I1O响2<ԉ�&�/�"}��%Y�C���<&�T�O=��	!CM�ӓfʽ]w �@���T9��S�X��b D��M[퓞J��B�I�����C�ڻ^��1�&`�P����d�J�IPgܤ3���94|mɐ��![�~��!39��4�?����IO�a�����Oz���o湐E5QU�d�Ua����ORb��g�'Y���`�0
Z���@H/`hE �E;m�"~�ɗ�:-���ܕz��Up�&k��|�1����<E���/��B�?G_`uK�����ȓX@PRN(J�.�Xi�#e�lhDxR)�S���'h,�����!A;b�qsm�����'�v���!7�r�'LR�'?`�]����;^�4RgQ�d��qc���G�������DK�OP��W�[1QX�PZP"�#	�D��L��}��ON.�M�ehϸ"%��`�K �~��,�?�	�S,� �
8����~����ȓw��Hp�I�i2��@��V/G�����)§h�,m[G�i�T����L�(&xؒ`�S��]�'���'�B��a���'i�)�	e���'�
 ĂV>1��ȇ��!���[�]c^|�'�a����b����դ��!�d�(
�Q&�X�I!PgO>�d8��	87FI���9D��h�	�>O\L	�Y�ډK�7D�<��;5~�Qz������w�D��}���r(6-�O���|:�������31~N������,�7����?y���?��i�6N�BQ�y*�Ȑ��$]֌�R��b�������x���=��
�韲��84D_�(��<��M@�l�	u�����a� �P�&* ԩ� oR����?E��'���"K�0r?j���9��(�s��'��)ئ�u��ܺ`,��e|�y�'�zQp��|Ӛ���O�˧V�\`��?)�3B$�ҀmOM=��4͇'����S��6�?ٌy*���j�.�.K0��啾LsJ!�D�.��xGx���'�2,�c�	̐�zT��2RĔ��ó8r"���O�4y-�4<�P�)26 ��"O09���8�@����>/0(p�%�ɺ�HO��&f�qxRJ�
p���.��T����ҟԓ�i̗m"��I����I���Xw��w'n=	��ؾ>ɨ�eB�3�$�K�'�.YB�f�*$������<�Rl;���y���)�Kk��$Ӳ_i4��BB�`�̆�ɴU���2�9	����H({� D��. � ]��ş���t�'[���Sd�WG2a�l�(�*�ږ�=?a���<n��ՃC���e��B	܁��ٴu�Ɯ|ʟf�N.T��׽is�\pA�2R0t5K2�3��T���'6��'3�m�8kr��'	�iޓ
�>9��A��3��Sc�W��EÌ�0��P��e���'5"M�7Ɗ�RHE� ��d����D+ؤS�̘�kR-:��8��' �̐��?�B� ����@բ*�2��d��?����s��xg`D�H-�1�P�ZQPK�k*D�D('c�0+L�F�)A��St��ЭO��Q�ڠ遺i��'��3� ��S��*p�0D�T�#� `�`�M�n�N�D�O���:���4�|Br'��(^9т�	2�r��^�'��]`���TS�`H�r��iQh��'`KpQ���G�OL�}r�lE�<�h���"Ӎ9��h#���W�<aG̎n�p,�!�G&uNK�Q��RL<��jSu��h�c�2���qfC�<!B*R�1=���'v�S>I��oß���şP���Q�qdd ���
6i�H�b��1h����I@�S����[�Uc࠙TEp�QFLA{,Ȧo=�S��?��x��5��e�}��h�̗~w @��֘���"�W&?o��&��z7<�s�$Ʀ�y�MLh����yq���GO��O Fzʟ��AĊ��\FF�@`ʗ�m1����OR��=r�Eb��O����Oj�����{�Ӽ�D!ՏO�~��+&�����]A?a�BNx�T���S>	���;�Bv��h$g��T��
0�O���T.�(U?� c��$tR�Kr�OH���'��{ҏ�t�=�0#߀T��kG�2�y"EQ�y�Fl3��T�n8��[��"=E�DC�)����6@� 4�����}�$c�)���'=b�'�����'��5�L��g�'�B�+�f���+T �yg�2�p>1�`�Hy�A*^(Tx
$-J� v���0�p>�5��T�I�7���i�"R���]u,B�6y%�E�c@�$}�*��#�+B�I.8�u�@��!	� UKǦ�	JT版��'4�q5�}�
�d�O>�'j_`�� ̈́*b
1�ܾUÞa��"�	�?����?���=^Ҕ�S�|��b $�����ǟ�*�h��T{�`s�Y�H�Q��ȧ�ɂo��ei�G�b[:���?IA�]"^� �`��B,�J��.ʓ5��I��l�Iğ�O���Q�5*s8ij ���x��\C��'{�O?�	9~�J�����d��ATK;X������_�I4�z�!��B��#� 	8B�D�ɠ�2���4�?���)� ג��OB���#@)VYS�M�A`N�:���r� {W��O�b��g�'G��q ϑ�A���gb[4�sD� 1��"~��.+�ε�W@q�ղ򈔆E���"�\ڟ �<E��*H�*3(3�<��W��x��a��r5Qqj��*H��ࠋ]�R���Fx��*�S�T��8A��ؔ��*.�L�+�KC ,b�'��8
!	�����'!2�'�N���]�T�q#�@��14~�4�O�J�8�{V�iW� �� ��f٨�zF{�E�$V6|UoԥH;�&�I7��o>�4=�+κp.P�aޟў�pR��9p�Ԣ�k~�zlb楟�+���O`�D�Oh���Oe��H6־9�p�*">��
�'��I���1M����bIҸ~�ܻ�''�S��[�L��̎��M[�j�@Z� ��ȚkTj$+���?�?���?1��Z&����?�O�����?9���)h�:�*S:�5ΏC8�tiδ<���جq�@!*��H?H �D��w8�< ��OF�d�&��`�T���Rf��4e:�(�'�0�	q+D �����+&���	�'M�"D��_�l �L=����'�Jc�|ɕ(ͮ�M{���?y)�@�!�ы$a����MB�f�8����.]�d�O��$N~t���A�$,d4�捃��'S$6=�'.�.[���'���u�v�EyBk�jPv5�T)Z>5^ȫT���Z"GX�ܓ�Y�u��yJK��(O�@;��'<��'�BZ>�W�O��`�gE>w ��0�+���|�?E��'+б�p�ǋg��3Q�Ͷj7�)
���'j����-����-�eqx�ˊy��'��y"�L����R���Q�4��E$���y¡�4h�AC�Ϡ ��p������y���i�� �*K��@Ȣ���yB�T<y�捪���%&�)
g�_+�yr.��Pty��&KZ\�BÌ��yBoV�K�`Z$��u����w S�yb U��h4�ED��n>�E"�"D��yr@EIp^h����!7[��H���+�y�%�Wr0dI�D�Ѓ��y�D�2����,�O�ժ���,�y�m��d�3�Z�N�H,3�&4�y2NP�=�*���KZ�[p����y
� ��+r�6�*؛e�ߔa��d��"OpYa��E�'��n,0)r�"O��CDb�����z�&��n�HH�"O����$f��8#%��G��tW"O��i��fɫ j�/+�bf����ybaP� H���׆!"XN�Av�Ƿ�yr.�-�P'�X%Ő�!�B7�yRO/T�.e�G��
 �6H�5T��yr ��x|8ĨT�̛rl�t�e�E��y��T2� �:�j�-r�ha	���y�� �_ �\�+;hRL8w ���y ��X�;�xʴ�I	j�x0��'���qb �G7�q��_�R���'��h�>I��9:��U(e���
�'���1�ϩC��m�(Y�0)A�'�8]����\�����R�Ze �'�*����30���J 6&e�'��q�A�f:�t���V�*�vI�'r��1֯P2��qc E�(p���'Üdd�Y5p�!�N���*�
�'ն�{a+ŦA� r���� l�	�'~AP�םQ<�=JbÃ%FU��'��|�W�\����j&E�t�i�':R�h�YT�4��)��mԘ�9�'ƨ`U�Jf���)�. Џ��U��>]`�M>G�C�_�8���� D�PdK�y�:X�C��*XB��T��p�S�O3���%�&_bl��' ݢyx�1
�'�f(y�B � \�p
wɆw�^	�I�ȡ��O؞,)��D����rhੂ�%�O�@;1�e�P@���M <{<ؘ�J�
�,��"O0iyd��Z�c`jE�~10b���C���D� _uDN� g��4�-'��yrM�9�p����.�v��eh��~#�z��O�>�� ⓭B���F?]H��G�9D���� ՗<���{��� l�U{t�$�$��E�a{� ��&(���ύz�4��R2�yB�	0�i����$�x�beN�y��ߣ	��b1���"Rq�a���yr$�7C����O�NC�	A#W.�ym�R���Pe�]=FD �u铄�y���fs�2���9CDP�u���y�/R	+VT�d�N�6��(���I&�yr��\�
�Cܶ(Q4��@ƀ�yRfD�frm�0���Y#���yRC��~*����
����B�T5�y��ٚ/ȠJ��
b�ʵS�$׺�yJE/d�����Y|QKG#���yr)�QQ,Q���M>v�Ц���yb��N�]���G�t��\��iU�y2�O=Jp"��T'a���ic��y���*mp����')��e�h��y��&�$�b ����T�DE���y�&��]�t���՜��|��@N��yϕ�K������؀���� �y�_/R��=�G^��NX�¬I3�y2M�!niPm0�fԄ��,���L���=��ʀOA�4��n��(���(�j�3�E	T�d)��y�<+Ag!�\��(��X�.��?��+և<�D9��Iݔ)����$j�*]tl)�"+�}�Q�l٢)?ڧux�m@��:Z�|����<u�,��4�&�D��'�(� ( �Id�iI���	�\���'	mb�}��O>�`7`� Պ��b�50�Ȑ���Of�JЭI�.�hpC��{x���c�ʿ*��`���PGm�<a�'x�O�a���Px��@�Q���� ���E��p���b�9~��G@9�OH�c�w2ʘj��جR�Xː�C6�<�'���fz��ɑHq(E�Cѡ=�ڹh&�ɞ6sX�I4���w��\��C��~���&��8�Р���ḑx7�O����~5P�jG�K>�V�b�%�'K_}�N�qXi��RƯ
mhp��+⟴��찟ф�^�N=�<0 �4e�eSré�T���@Bܓ~��(� Hҕc�E��i@PGDFz4AZ�*�=� �� �4\���a�O�u/ �5�m��@�CCT/��O��͏6ԊqV
ų5�Z�r�xb��#떴:�ҡq�J�bFZ��I�c��%�×m��c���f�x���2�N}��%V
&X�~RdD�~n~�(B��Bz�d��F%���Ǩb��|b ��tHv�Rh\����+ċ�7&�z H�l��y'Z�!p<�cI�
3��é��0?�TI��B,!@�X!)�Fi�R��5wPZ݉Gn�F\5��l��%�\r�ݍX��b��IiFh�V��7�Z܋Cf����׊��Ų	�e��H0��'�4�J�S0�7%��Pa���!IF��ק��-��M"�qԇK�w�FH "R�Q�)9�(�,'�8�{�e�4Br��>)���2P��X*����MD�<�`/75�����~PD�(��?H~2Q��H
\i���A\�BL���T� ����3aިC����ȫ-5�A(�#(�OD(p�\�)3$i���HY<�)�G�"W�T�6K���<��B�Fp�)s�D�I�)*�iӢX�� ~�x���	b������LT�%O=�O:��'��9Y�2lr��I�%&Ҩ#�녊h�� �%�c0���L
U���Q9O�E�dV�"�L�SC��+UQ>�C��O�� �"�v��lS���"�d����7�Bd�P�_�i�B�aP��lvr]$Տx���C�:x01�����5��D@�{T������Y�Я8Q�dJp��7+�h�B��K�
�q���j�X�҉*@C�$* �7~��eHt��kh�@��[�F���E�`�W���}��PA�	��8n,��T��9������SE(a��O�DX1��Y�"n�2Q�6���@F�7W0��i��V�r��:d��,r��V���+ĩS#^������@X�t�xԹ���H/��;��	=c��	���'?�	�Oj�x�C�Wv�Cӌ�Q?!��H�9슴����&&Ř	ȵ�O�'�N8i��L�r^`U���A9�U�E╱b@���p �(~������E6��J� !��K X�m�TlS����D}����)vڄ��ރ`��92sA��y�L�%��JB�w���Ɂ���i�څ��Σ <�80�OP!��@)?�]��l�IKbere�Y�
������8��G�`@���
�*!�p���X&_>E��T;�w����B%Sb]h������9��MH���ƥFm�,�F���yjņ�=�hO�p��H�Kx�Щ��֧>Z�ca�O L���@:�|<Ӓ�ؕf�~����'���2�뉶D�5��܍m�&q�H#64.��`Y���X�GH��?aG�	K����S�۬U���zXC�'�^Ěd�C$q�Qr���H9�}"	B�;m,�y�O⭡�A�dB�S��)&
U�<̬�C����59᠎2!"�~�)�:DyX�fJ�$^�);p��;R���I�g?��Fɡ3����I��?i��wOF���a�	�l�#��ʏz���+�'�~�sR&��m��������MK�/?�ky�H����u��Y�D��2ޟ��d?)"� �qʹ����(�Xe�l�'��4Ѧ�X�`i��k�)2�I"�*�4Y������E;@�P��H�zw�&�?U��j`� j�(bU�^��OD1[�E�:N3�91�0��Ӏ^�p��ř)MX�8z#��&4"��ɦl-}J?���V�H����E���y&�<D���LC
8�n	!	n�\���)jA4����0��Q�t�T*wMBO?i��V����03��-gD�93��Wb؟�H����*��!�Gď��>A2�*6�PȢ��:����e�c�ʡ`G�:� D}�b��&2c/Ϯ_���*������O��2�8�v�@�F1M�Ԕs5�i��t�ԅ����xsՏĄ,��,�rB^����RN��J ��e���ϑtR�'��-����?<4����X	gUp$�M>�O�.i)�h٣X^-A3��<C�Բ
�'���`f�HJҔa�
P�H ���T��*&V��� E)��~���B@���1��A!w�Q<����$���(�Y �'��@#s���d,�����y�0�A�gŔv��I�,�$��U��d��+	+~�*%��H.�I;�l���i��Iu�y��ɚ<!��?��k��As&�����f��
�FQ[�ب�/
4J����L�J�����xҡB��į*��%��I�0��R�@.T�^��V`�<p�*�=�T�VL���;��Wb��0Lҟ֝&`���2�X��a��3!"B�	�\hѲ�ӫ'����ǋ�*%R��ĕ6m�:�xVCY�8<�P&��L����ţn�� �A�ɲ�&e2�d�VstC�I"GU
�J��'a� �b��9�n$pP�P��^p2�
&��-���6�B��	�F�����;���u� �0?���ZINZ2TѢ�����7TD�4H<1`�$A%�;?�Iy�e���4���or�cd�G��=q��!o��Յ1]T�z��v`9��.�6AX���#B"i뒁Ҵ`���>���0D�� Ԡ�pa�1�]qfE*f��GE8�?���5gFP�`2���<�Ԁ��a�3��'e���ݢ����zs�]q�j�J�`��T��!�����$�P@S<3�~A�(��M���� �1Od��g̓!*\�t��(2i%��l�1V��h��I�GA4[I�qqǋQH80x�D�����%4}rA�$U�� ,|z�*u�L�/ (\8��%xv㞼��ا�g�"(tjH�H�Rw:+AH@�H7D��nܓ����
�cN�
vG�#�O��ю�Y�(��Uy;��"t�Iw�xIu�%D�x8Nպ+i�X2R���=�`�
��b�Љ�%�W���;bQd��`�J2"(���"D�0q�Ö���	!�ZAϴ!K�!��xD@.u[h�"�;˚4�1��z6m
�Pl�Ob�G���`S�P7��3��
�R�c�����&6Zܬ;@�d���l�B��?J`��%�^)X��p��
�%� p��:�(bd�.���Od*��ɀٸ�����,ϓKS��w��KhE(0�p!"�O6D����LE�L�X
�6�h�"*6�I
S��DO�c"qO��ʝO�Nt"���
<���`�� ``���'/*1H�ID.+1>�2K�%(�� �딙`���%���'*b#}n�:X��|��d8T�hX��.A�������Q�@��y"
(�� rL�
�XCs�F9�yB���پ�P1MV>��	�y"�����	څy�"쉑J�24���e���!��т�>�b��|�8�Se�l�qO܉�2B��0<��HB>p.Ta�(�f�0��#"�AH<��3�����L��N�Se����qO� �m�
^���GB�\=��X�"OZ�k��D�O��6�$<��f"ON���m���T�*$�yp"Ot�#�.:=i�Dl/_�0�"O����"H�u�@��H���Z�"O�-�d��7�BK ��x��LY�"OTA�q�A�:+�<�&_�,8�u��"O�I
���7� 	� F۽A5dK�"O�����=�2a o�55�["Od��Q F���2�̒4B'���t"OT=hd�_�]^�M��Y��:H�@"O\�SqF(m���E��4��	�"OtLs��ԑV��놏8=��A�"O��b5#^0yd��[�d�{xLi�"O�iI���mh"���A�r���c"O��x
�?.�b��7�L�o��#"O�:���>P'����@�&T,ӵ"ONu��H$ �U�/p(؉�"OJ��cF��s�"�.e�Jpi�"O}�dHU>FP�E��\�|��"O�A8�/Q�0�$�]<�'"O�	��h� W:��#^N��!"Or)�OޣynV�:��h�Pqٔ"O"�T�8I���J������ �"O�3Bh�u�\Ae���$��={0"O(�R %��z2����AE��c�"O�]"u�Rm��,9!d�)���p"O��%��+{���r[,M��Ip�"O8��'�!n4�A��ۨy��e�!"O���ϴSW<[q#n�N�q�"OH�{3� ldA�d���}��S�"OK�U	p�1�)�T����M2�y����lp@j�C�v��b�ɸ�yB.�$'�m#Vn^;R����"��yb�ԑ!4F�3��E:� �YA�����FC�e��  �p��ծ��H��=_4�(�4RKF��7�X+C�(��S�? ��K#\�֤��4N��I��4"O P"�!���C�nɄ4)�]�d"Of�Qǥw,޴��M��'A�MjW"O���p���7���S��*#(�i�`"O����-�� \8�&l���J�"O�	��E!�R�ҥĆ(�@��q"O�a�5h��M�0�η5�Z��"O���Bu� �b�D%�8s��{�<Q'b� WH;�A��O2�a�P�b�<q���'I���f϶b�q���c�<�g��=/v�� �K4So�yJQa�<q�M��+.�h�� Q0eV��#	XZ�<��ށɺ(�F�?j�1���_�<鲅�4K�ء1�D��r"nA80�\]�<�N
1��qZ�FE�4?�����V�<q�ś�G�"d!��S�f_��C���V�<a1�����D��c�H�+��TU�<�V ק4b���7R�0i�R��\�<!#���8"05� �J�~������B�<��j�|c�e��4��)����A�<Ɇ�[$U��*�c�)�@��؇ȓf'����jW V#@�P��7���ȓRv��CVc.�h���6Wrȇ�V�P�ku�K�	G�p!S�R�E�d�ȓ~��1Xq!�q5��y��'�T�ȓq�<�b#�$q�l���@�x��y�ȓ*~d��(�N��iѓ�P"Q씇ȓP�N�s�Cx��b%���w�����̴��+@�G�}r�m$D�n��ȓn�ěv��HC��Ip ˇ��t�ȓ0������iaj�	���`!�'ў"}j���<vl�w� :*���&�w�<���ٷv���i�cQ�o
�i���w�<�d�N#.�tܚ$	���`i��r�<�D�X�h|���<F���#�H�'^axb�\�J�\��E x��
R��y�c_L���h1a�%� ���ʃ�y2�v{�|["&�?0a�	��ybd�2r��sn�����c���y2l�r�m���T#:����L���y"FU��DM�"��?;�Kķs �͆����6@�`G^�i�H�0|��C�I.w�xp�˳	*���Rl�$�RC�	�cw���4 D�Ta��
�q^tB�I�Mm蹱�#E��SF�E�n C��\���aJH�zf ��mD�J8�B�,�bK��[�T�5eĦ��B�Ɉ$W�� ��?Uo�a嬁84�hB�M��0��ܚ Oޜ:D�B�	)mԤș2���H��q%�^�B��>NA8�j��(8���3ǔ���B�	,i�<��ʉ�2h��8F�Ѯcf�B�	�:�,ӄ�<�����i̴a�C�	C!��q'HԄ\�$����2�rC��>J��Psc�4\�R{f���FC�I}|8Y1�H��2i��R�kBC䉭R9ȡr"�Q�{ ۟k�F��hO>1���"z�vDHbd�! H�94�&D�8��G�${�tITM�)*���"c/D��q@�W�p�*�/ߥ|ʄ��  *D��P�
�7]��tq4��9DTP��$D�+!��%(K&
�?5��,;c�5D�8�"�S�2����c�W<2�J��.��p��(+�?s�R)���߈4�TY:�-D�� �آЃ\���p�y���"O���RE��{+��!`8d�����'0qOx��T�[5*���a�n�O� s"O\�!�ˈ�K��6��?~�4�ʴ"O ܡ�o��_���#T���BՀ�Ȣ"O��6$E4G��(���S��#"O����38�q�CH�ȡ�b"O`����ɰ�L�s�L�8��] �"O��@3 �0l$���y�ٱ3"O�)��ؾX2��)@�U1dL8:C"O��R��/��@����yJ�p� "O����Z|"�������X�W"O���卟�7{�U!0�� j|����"O,�m����X�N[�@��E S"O��Pե�Ju�6�B
B�H4��"O���;=�\ytk��c���C�"O��@n��r���qa�e���1"O�HC��&����[�$�b!8V"OL��4�! s*�bN�R��q�e"Ox=:U�_�q8���cK.2v�s�"O��3Vm
��>��sS�c�1i�"O2��K9q��)9OC����+�"O�0ڀdQ2hp���D�m�,��"O� ��lљ>@aD׎k�0���O��dU�7�j�qH�%N�c��/�!�dYU�����Κ�?��X�&��)�!��
��x���B�V<�{ aA��!�d��W>�Y"2�ܘY�X��͌�_�!��F�BYr�˷懩1���q�P>4=��)�,��IK��
�-`��;C۲(�RL�ʓBּ��[��P�� Uy>U��r<PU�oη\Ixp�OT�/��y�ȓ&<��k�� o�^���Ҕv�4��ȓ#��!�.�`B�l�U��,-��J�Ԕz�GP?}߂��⌜Ezd܅ȓ ��#"��MvJ���>k4��h��Z�d��ۈAK0�#�%Dp�<�P�N|@�j�B:��`���l�<�qOW&�֘��ω�kp2�Z���p�<1F��C> k��D�7�桪fA�i�<I�%��⬐!�������`�<���V$h#�S�Q�`Q�)O_�<�Ah�:ᘥ��A�F��Q aNv�<�$h�&��C`��'��Ҳ�n�<q�Q;PI4�!D|��v$�`�<9v���*�ctc�3�2�`��[x�<��9<��r�� ^����vĕr�<Ɂ�*pK�MÍ!m��"DU�<A�U,4����Fd=Z�k��SQ�<Q��L�r�Եz�1f�*�cV��O�	j��8䌈#o�`�*eBQ5(� ѻ�	"D�0�ӱ	�2h2� ���=D��0Ej��x���%ہy�� �K/,O�7->���2�hP����X�q��/n��C�Ɉt��@�o\.�vX�E��=�=	�'~h= ��
]� @.�?b�m��Rx�37��IO�L�glC�8SDe���������O�A���}��P�ɺo���"OP�%j��lHW�����"OX��W�I>oBM(�K8/f|�2"O���'�NM�$p��ϥ����"O
�jB�J��f���閮�,��$:�S�S�q��(Ô
Ś"�}��ǙrD>B�I�/�Z]����o� �	 �?&Wr�O�=�}� v�!�/?��H6!�U����W"O�Yòb�!in(Vχ�hF"�R"O�馡��o�1�U[�0���'���c�V4���*��I�rnT�#���#"O4�!ׄıiAP�h��T4wjRd���'\d#=�� �N� ���g�%��e�_�<qD�˫I=�P"���,���^[}"�)ҧ�z���F���5�]�5h��,�D&�ON�c���=��l���!���"O��U�X�D� �;M��d�"O��4$ǭ"b]3C��:�²"O(��HB�!��r�c�z��K�"OV���ʘ4/ne`��La>�Z�"ONı�c,X�P���g�J����"O�#' �
���HS'P�2�`��Q"O:�a�B5j�D�j0%H� ��ݳ@"Ol�q�e͹?}��0oU5��4�b�i:ў"~nZ�Kth\@e' �oꨱ��hB04H�C�	&b<��P��%���P7`�4��B�ɘR��-�1ڦ����  Dg�B��];V��'�I�1It��c�,B�I6tRU�o�.8���w�� )�C�	�_� �� I�15L�t f��{��C�.*��c�("<�L*�k[1XU�C�	�QA�Y����
T��C��C�AI�C�I�?����ub�n��`�B�x�~B�6Y�F4�f��.��A���E'x~B�I]�~�:7��}���է�ƲB�I2vtt��� Zpj���8B�I�/��Q�cF�&6� �
6shC�I>U����Dȑ6a�uc6(�&C�IF�4�F�K��"E��&A�
C䉶4���NZ�qx�E�e��U�C��
_���`hB�!��ԊE�^'<E�B�I�0N:}� �	*fh��,ǿ��B�I�8�� �� X30��"`��;b�C�ɥY��� ,EVD���I8X�C�	�I���j��>m@2E����(@��C�ɛw�ؤ�f	}�"�+J<m�C�	�^����JA?\D��k�e��:�fC��0Ր��EC��U�0ʛ�Z�ZC�Ɏ9}T���Y4+�*�A�1"O�iL^��R�����,�0��"O�p���`o\P�&��]u��3"O̭��c\P̌ YDƑ�^i�"O�q���1.��#����}#"O�ْƩ6��B�䊋�^:�"O^@C�)�=)��Q�N�gϊ\�"O���"+�;���[# ļ51�"O��$D�%$�l;���
��P"O�;�O\M��F�Q(�T3�"OH	z���+�lGD�B��!򤝖,�\��H���O%m��ȓ0�� ���A��Ր��͟q^��c�t���\�b=Ad�.	@���A�E; � ��f��iҗ�N��ȓ/͒d;T
ОAF	��}*T�ȓ]��D���H�C�CV8n�X��ȓq)H���J��4���cͿG��$��Hڨ0���	�����FZ�И�ȓ$�bF�Q$:�勁��[��q�ȓ7E(���'l�� {a�2&˺�����TXт�P84�E�ЮP�:��ȓ0���hgC<^�-#wa��%��e��S�? r�y�)J�$��E!!�	��* "O�9`d)7?=v@�&��Y���y�"O5�"ˉuK&�'lh|���"OP�W�>_�mxC��Re��;�"OV����VI@څ�Uk\�O��Bf"O�`�SFޝg�|���+l3D���"O���������P[��S�b���g"O�H��&Q2F�{r���9�"On]� �ξGpSH�]br9a"O����&^V�1K�aIwU���"O �Xg�B �.�s!��J@(5��"OK��z��5H� ӦiبP ���ya�;nh�Ȇ�ɯ~|��@��#�y2)	Wk0D�3E�s�j�w����y"ȝ!�\�3 Tnh<���+�yRʑ�b�z�g� 9B��E��-�y�LS.�pA��䉌�d\cU+.�y��n:d�f텀C�|�q� ��y�,��=�sB79��08Ԇ�<�y�/f9�,��ӄ6s��H�Ey�<�e�H�4뒤�qn
�|Z�8�@(�{�<q"Lb0�x��I?r���:��]u�<c���E� ��c�>ǂ,Zc��x�<����"sV�a��ݤF��5�GBx�<Q䏓�$��)�i�"/�h�0��w�<�4�3s(	�I�F�x�!H�p�<!�RVEna�i��|��U�NS�<��֚N�����4Ȉ9R�y�<ag .\�QS�_�=v���"@�<)fOJ&f{j��� �)�A�A�<q%	G��ʵ�7��PT�M�% �B�<I� �8ǲt��g�H#�Mp��FU�<� NR<9��voFP��� �a�h�<i�bm30��E�hIS���5
�C�	*bh�0ˇ ��x��U�Ýj�B�	�b��� �K�(ٔy�,�7_:C�+:�*\�)F�`-`�9R�{(�C��i����5@rXu ��ں8�C�I�J�� $��R�bGA΢�C�I2I ��NV�d��	��B�,9��C�	a���D��1-X�MP��>'��C䉱b-F�� ϖ�-��5ȇ��k�C䉸o���k�H�4�UH�%S4SB�C�	&�P��_�aC���WE��m�C�ɾhjf�K�@ނ	Xި��#��*.�C�I�k�J4i֬��ր�f�u�C�I	1��ZU�	5c���Z���'_��C�	 t��\�d��[(��Ŏ���C�	6r`�-	A��64|�ٳӯ��4�C�	?H���S�(6m��R�J�8�B�Im�U
����xqbc��+5v�B䉿d̛u�Z/K�@�x@�A��B�	�C�����A6��X��ȗy�rB䉌(��\Sb�;H���"ǖ�.��B�	�
�X����ƍl1H��@D�Fz�B�/Jڮ��Phe\^�E�Ĝd*B�	:?
.��HN9@02P�
��	,B��(L���A��g0	w��l��C�	�r5�Q��l�@���	S}B��=`�$X�5���f�(A��Z�	 B䉡c��)��0\6�$2UkZI��C�	:f"M�4@��V5�Q��NЮC�ɪM�DS��`*�T�;6�C�	�4�ba��DطG�*x�`�Qh�C�)� pkuD��8I�ykf Z�A�����"O~,�s�Z.��!�F�h�"O�a�/�Lu��+��F�KTf��D"OL��3bG\������	B,��V"O�Yh��=5�Y1�I�<�M�r"ON�󀀱Q����lL3.�V"O�!�ը���s˗%EW0�A0"ODa�� �@HȁjeL�z��9�"O�m�&,U;� ����${����"Oz��mػ#{*�r,ݐ����`"O(�ya�ωb�B 1fK�$`���"W"O�0bզƚE�:E�UE��)�H-��"Oz�V�_�S��es�yú�Q�"O�` ��kb��6�L!_�>- G"OF�t�5?z�� �b����B"O�Hk��R�����@��{�"OlYz#�̱�D�"��>�T!�"O�]�@Hڝ5���` �x�"X��"O�QR A�cl�5�I0B(�=8�"O:8�4���Ut	r�ˁN
��P "Olͺ6�'��e��g�t��V"OF5��!ۺO�������&;�"U�"OB�wiβS˨�q���|u($"ONl�SE� f�	��JÖ	�fir�"O`뇌F�s!\y%�	 k�����"O(ĳ�F�-�	�eGC*�\bP"OF	zG	��vːl�f����@	�"O*�Y]0�ʥ;Bk�f�x�"O���P��+��9ӯ�}p��R"O��qM�1,*(�gĜ[p�Q��"O�E�D��*�8A�&�'Bq��ѕ"O2�F���_�H ఏ�#8o��QW"O��`�ѣoq��#�.^/6�r9�E"O����K�Xd����FFR47"OL��E��5m��В�n��(�R�"F"O���4?:bu��m=�z��`"O �k b��" ��UmS�v��"O�36�
�>y8'�

�R��"O���F�/P�� B�!I���ˁ"OT�Pr���nj��cg�ܗB��4;�"Ot�NQ�(`Dhi�+� C�,�G"O$�b�
��_��PQb,J�H��a(5"O��+�$ծ|>��SLJ

����"O`*��u؄+	^�q��bW"O����U�E�l�K�<�@��T"OȀ�mΗ���,7m�:�"Oh��UM\���!!��8�ހ��"O2�*H��UO
��2@�2w&�""O���`e�;��a���� ~�����"O�E�3儀i�l�"���:F]�,2�"O��;�dC��q�F��3eYz��"O~a�牚�sJ�axK�;'"O*�+�폼)/p9P�`�&/��)�"O�u�r�;�����	A�G��rs"OZ��c���E���0�٠{��:�"O�h8C$T*X\xA�Ry��2�"O��p�@R�16�pك{����"ODX��OQ���b��gJ �YS"O���UbU�0(�k7h��>�A�S��F�O^�i�N�13�R�S��^7��c�'����a��雒�-(d`K�"O���O��րХ/��u
�`b�"O� ��
�<:��(�CH�^	��"O����#Tq>�)�� �0�T�w"O� $�"DEȍ"���`d�Ϲ;�$�b�"O�P�� ��]�>���#�98 ���6�IL�O�j�Z�h��J_�Ѐ�I�y�"��'yr}����Ե0%�ru�m��'st)����>#2x�b�	4ĸ�0�'�`�sM��-V*H(��%��\#�'c�-:�n���싢˗�t ���
�'.��0Oܦ(�� `R�P��`�	�'���tLѹA�|���%̐��m�ϓ�O1Z�M:T|D��1bݝB/��k�"O�BD�T͙�&_�*��Q�"O��g	�79�d�X�FաI�r�[�"O>����,��1X�fT���aBA"O̝A��5R��Kw���Q�"OP����Ud�.l�C�\�_�x���"O��g[*v�� 8�<J�6�@"O�)���
�.{B�
�H&g¼Xp�"O, ��A"XY�C�n�p�q�"Oz��B.|}���S�7�N��"O�p�B�37C��r#㝾�8��"O9BvM�89@�q���A�ĕ��"O����搇$��6a��~9�$I3D������?"0��#�T���6D�T"�����xys���� D3ړ�0|*�� �j�Y O�.-Nyˢ)@_�<d灠a�>��ъ�*��C���d�<����:��k�,@&a�|X�rÈa�<I �͇aD }�畤)��i���\�<Y�V6	�<0�HC�;^P5�5M�O�<�t���O��y���"���
5� L�<�$	[�>U�3���J|J�!r�<17$�� f\ �2�[(�̅�u�Go�`���O]x�#�Y$O�AX�O
�A���
�'�8yR$l6T�b|�ᯀ�0Y��	�'_rDcW�ݪ+?L��(Rڐ�	�'G�z4cц-�$�p�
K\61 	�'5\�cC_�w������Cʬ|I�'�|�gx#y��Ё���J�ў���S��
�Y�B��PP)���0�@G{J?��mLxVz�D��4;W��" D���çGe�ze����s���E4D��aVI��j1 ��	f�޹Q$/D���Ŗozx)bo�����0D�@� K�i�X��CٵH���� -D��S��ذXw<��s�R"6{�U�5D��㡍F�A��&�07}<Q��4|Oc��iBC�#)w���w���z,��b5D���b!¦	�
	�q/M5q�P�Q.D������9`4���y��=�K*D�� �h45_ȰZ�)=m�tSe&D�Tj��	V5"�Ha��!X`t� -#D�dA���3(��M���ʗlV����!D��� ��.5 ����!& �G�#D��4.X�]��!M8Eh��4D��2�鐿&"r����M�h��1D��#e�X�	����ݍ1*�ѹ��.D�k�������˧+� }��}��+'D�� An�Y̸�:@�D�^�xYb��%D���W�_&�ra	��D�p$�03.#D�@���S	V@�	*��C���qZǆ?D����oKB쑲@A�L�Y@�7D��2ă m�I�矅Q�v��� 6D����'̬#��"�.R�-Ƭ���>D���r$\
��-���f�)�!f;D�� 2QB�55�D4!�C	�R2"O���0�W�{5���7f.R�XU�"Op�"G=:��P�ǥ�H� ���"O��FF��u�q��ڙu�<���'!�ˈV@�R��G %����,�8�!��I<+Ö��Ƃ��c��	c��gw!�.}�aÒm
�u�D�
t!���J�`$r��D:Eo mI"��_!�̝���RUcOhU��q��	��!��ż?F@K��uT��A��R�q�!�7L���`�I@� ��t�B��>L�!��?���B���:�P�b!��'Z!F�pvnęU�cCkâU!�$�Au� ��o]�A=�jA�ܣ);!�$[wJ4��EH�U7���3+� vT!�dX�z�B�����.V�\a��@V�|k!��B�(N�D[r��wm6Uq�M)%V!��,i���wD�
��X
V)̎zF!򄝣k6@T鏀[�$���Ř��B�I>i5b	�Ҁ�'��	cd
W^B�ɐLh�B �^y'����#�%C-�C�	.;]~�0dG�ǀ�BR�F<^h�C䉇u@@eŹ]-N9�B�_���C�%Y� ���>1�g�2zpC��eג,����^�`F��yRC䉱����F"	d�B�5m)�B�I��LX���[,nB %*���}@�C��xU��իGXU91�	�D��C��%HZ�0�ě�To�Qh�"
��B�	3)Bh-�ˑ�".�l�"���EՄB�d.��[⦅ zJ5;f.U�(B��/�
�[�C wHi
V��Q�V���??��J%:��1��d�f���EA�<Yգ��Z���ZWl��8Pb�{�<Y��C���2�mǸ��)Y�/D��Q��Ň%�����(�z��5�2D��x4��bjhpQH�?Ct�t�1D�h��'�'SE��� (V*><�p�2D��!�d�&Na:�aA�;:�
,!�/��(�Sܧ%�z�@���6��Y8%� _�b5��.?��)�/-�蓇�<E>����T�"�f�!s�,X��![�\@��	� ʓ�OO �1�k�=�j܄ȓ&S���&ظf9>�%,9M^����G��p����%C�q��o�*���S��M+r��?q����hqqv�V?0P a9��5?<1sW"O@�r#M�s�h���®4V$�"O~��Z"K��@$�U'PX�S"O\<��KP-E~ � �d`���"O�%� '�PGh,��)p�ۂ"O&�����j�2g�5ROd����IڟPD���%Q��1 Ɨ�C��Hb����=Q�yrÆ+	�!u��@`�8���yb�_�?S�8W���J�|tk1��y2�ɷ$���৑5B=T�h�yҥ�	F>��C,�9�x�#_*�y�牨h�P��4�5>9^������hOj��_r<2 ��
<dt, 3��M !��47�ة����S�TY�*I6�!�D��Q3DI��g��%��-���B�!�!��n���Af$�9�j�8է>
�!�d[�g��*GÃ^��������!�˱0eRU��-Qvu�p�%��(y!��_I>����' �P%j�Eלlv!�� ⥒4ݦ5�X+����r#�I"O���h�>��K��Ŏ�2!�"O���#��6���l����8�"O� �W'YY�4uӅl���b�"OV����6bнz��\�Rn���U"ON��W��a!��/��EY*�a�"OJ���j�2U��A�^� N��k&Ozy�)	�x��]��F0v�Yà$D�p �@7!A�<[U��{RP$Y�!D����*31ȜCA�7q�p訓�!D�,:S!Fj�H2�%�;+W��+4`!D�lr��l�"	���g�b����>D�D�v�!|�: ѳF��6s2��`f'D�8�2DG�2)r���<(�AE, ��?���ɔ�K���FG�Zž�#��H�T�!�d<9h8��d'�v��}�U�x�!�d֕ݠ����7$�J����5c�!��?H��t�F��q�� "agʿ
��)�C��lP���C���k'C�d ��'䬐�!(M�b�4��U;z�nia�'��1gϚ%@8����%B��eA�'����S�z DhwD�@��<�
�'7�1��l��{/�)CR!�
br�U��'��ib��?�L@�!J�Bw �@��hOx�=a���xy����I	ވ驃 V����O`���S��'7̹+�"B���3�	ʓRX��	�'�գ�H��*lZd�uK� ����'2�� %x4�Q�5�! ��@��'�BT�u���]y"U�I�
�����"����)U.2 �\��%���^���"Oֹ��H0��9�$ս�x�¢Q�PF{��Ƀ6^��`Y���:F:��o� ��Ty��'�Z���!��g�8=S☤2%��'8�`��I���ŐV��;.�a��'��z��Ӧw��-��!:Qp�M��'��8� #�07�\�З�H�J7:9��R�)�D%U�$SV\�r�0|�x��/E��y�OX�!S���Ɖ>>�2��6A���'���'Z?MS���!�>����It�&�$D���H܋,��L���!���-$D��R��g2����'�-�*\���!D���vfH*҅hDJ��:*25s��+D���`��&8'��Qȝ0N}jPc�O\�=E�T���<b=�2��?(�����W�!��ƳS@�<:�� &� u(�"/
�!�d�}7��ѐ	Q ��t����ў܅�I��̃DM>aH�
�4.��B�I,�P��� FTix�U�G$�B�I��#ŉ�)�JA":$�C䉆5:t����1y\��d���Y��=�Ó=0u9cL�Q�>��d)ШL �)��m�
�J!���%@$Ar��U����ȓ.�̕h���e�VѠ�*˝$y�=�ȓl04����J�E_�a`�EΛj�ņȓ{������-�ͺl@�v)�ȓR��PQr�ڊ0l�X��(v����pP����-]���B���7^Q��,������RR�j��ԁn/<Єȓ\&)A�O!��s�R�q��l�ȓS����.�4q�� 4�����f J�턓L:��h� amPi�ȓ7�^Y3�g�p��d�	0���ȓO@\,8�&�4�J�� aN����	v̓X���;C�.^���"�D�i,�̄�S�? �	S���s�T�qi_6h��e�"O���4D�?Z�8�q&�o���s"O*q*1D 6�$q�8}_PE�"O8�1�/];S��m���Y%�W"O*`㡍�5���צ#�����"O\y�lZ����$�`���g"O*8QVϕ�u��q���(v�0�d"OZ�D�.�HX����cmj�"�"O�ѻ���+v�=�M�DR��)�"OPu���h�X��薢86�h�"ORR0��-+Rd�zv��_@`�"OJ�R)�"�B�H`-8�ͣu"O��`�	�3*yl��S�[=�ܸi��\F��jN�v)�̲Ǌ�<��!&
1	�'�� 1��%W��4j��6���	�'�t����ȴԂ���L��O��h�# ���ȁ�D�h �ȓN(��z֧ �Y6��HS$^P�E�ȓ\V�!i"�1\AQY!�L���i&X�Js�޿<`��P�Ff|��F{R�'�?�zU��wIa���Ęhް��l7D�X ��Q�XxL�g�A�e� p+D�x�Sb�8B�9�FA�K(D�d
�Ɍ�8Ra�"B�}�e2D���G�K�AҠf�0jh�|���1D�0�Àtä��l��F�qb�9D��hq ��.���̕�p%Δ�+3D�X��W+w۲��b վh8,y�*3D�\�dP�{�*���!�6�S��1D���Fی?0� 0�ВH�$��D�/D�`�U��(:��[1/O��P��.D����<5�� K̭#�*	��.D�, �&J:,n���7o�)�<�!p +D�D�BI�=����Hۇ�塢�=D����^X5�I`�X���dcdc<D�`2gb��<�$t�U�H� ���
6�8D�`�4�X�_^N$cPʇ�x������6D���l��Z���P�ڕ0ac3D����÷+�,�	��
A�(��2D� ��%Ix� ���\�r��Yr�+D��ā5|�,չХ�fQ|�"�-D�\	BΑ|������-Zap�.D� pb�ݓB:
-��FhX�DH(������Aa	�5x�R�j�i�=L��S�"OjUh�O��A����JCT|f��P"O6���I�D�BH�щ\�ik6t��"O���WbU2mh֕؇O�?H_���c"O��{��7mF�҄��m�u��"O�1ҢϜ(��4j�e��E/����'���2��@�B����Ȏ�&���'��	�
	]��A���9#0���'�"�#��^�5� ��,U:s,���'C�ؑ�V�_�<��&��k[�T�	�'6
C&j.II���K�4c����'m6,�� L^��Ŗ[�6x��'��T���no܄����Y�����'�0)�S��O0f�1E�� �ʓW\�Q�����(��?�,��ޔ!a3ƇyL��D���������H��Q=A�%�Խ�ܘ�ȓL��ԫ��9O�@�Ŋ�t�����Pw6}I�]�unt�#�N�g�r!�ȓ��b�B�K�P$�����FP� ��T�l5�+��R��JK�-�H<��S�? ����E�4#TZ�i��f���5"O0�:r	�U
m��GJ�t��(3�"O�A�Ǯ��l(��kf��\�q��"OP� �B	[�ޭ�@�R5;�]�"Ot�/!7��iAdT<Fɢ�"O*��5��FJ�8&d��&JL�"OV����:WК�8J r4��+�"O~���'_h�6�-r���*�y�̃@�p�Ǣ̴��{�f�y&�"���aR,�?�Y��,���yb�q~.�a�@ 7
�IȐ�A�yR&�v,�ـs�8��	�#ֵ�yr�αn��
!��7�l��� �y�[9_�ޱk k�0�rq���	�yBK-�<��rn0bd�摓�y"��'c��qI�Bz���)�Y��y���88���0x�D0#�@�y"���l�lĳ�"�1�F�A��y��9�bFaM	���Kk��y��Lfp����oreh2a��y�e�U�$(էL	�mKR/��y�G<�M[�a�� ��c�C3�y2B�V�,��+PsFz)���yr(��#e�[` O�f!x�#�*^�yb��}���3aJ�6Z�va�So���y�M��+B���	�(^n@���ƈ�y�E�%\����v'\t�Y�S�yB���Y�<� ��x����e�;�y�NFf���)�fעnbj�pe�˻�y
ʹ6�*Q
FH��z�~����6�y��,)�BDаu����m���y�L�)'�	k0��=l?�ȁ���y��=(.�!E쓳2��9�C[��y"@G�K������b������W�y�c��\09K½TD�\�#%Q�y�M�N�������6�YrS�<�y��1�t��#�f��t�.��y2HŶ����]�V�ɀנ�5�y��,%9������$=�<�(vM���y�(����@%:6��b�I��y�D�z��R�:�HB�%J��y2E� ��@P$�,b���$��.�y�JP�#���Ō۝Z��M�JV�y���hknD����d~ys7Hț�y����z�
)��V'aTh:'�	�y"��O>h�!mǭјhVAM�yR�N�1F�!�3��ݳ�'���ybC��ɱ1�$�ܐ�o�8�y��o|lD��c�;(��1{%e��y�&΢�Lu%�2�`pU�G"�yr��PK�p��	�eQ��S��y2��)&z�p/�i4�w��y"�;H� Pѧ$�Qb�]bƢ�yr�� #��X2�Ar���e☆�y��*��JF;?�3mb!��3C��;���|T��u���uK!�d( ��ID� zp)���H�J8!���.5����\�P����%U0!�DƦtA,�{�M�T���V���K�<is��KJ�{!kz<�B��C�<�W���j��C�lA;1�,�� �[�<i��K�W�ұ��N'����T�ZZ�<��O�P[^2�����ܥK���S�<�1�^BMh]��NE "��Xkk�P�<� �Z��$m3� �|�B=��"O�����1K�]Y�e��C���(�"Od9�V�](i�8ѱ�b�/}�X�@"O���!@���@�2a'T�wfu��"O��i.Y�,mZbe�
j��@��"O�u���p0�LSQ�ٓ.���"O5B��AX.�g��K�}2r"O��w+��4�2�z���y��Ls1"Ohh�����T�<¢/=7�H�a�"O�ZƠ>=��й�-V�k�r��T"Od��a�j8^�K�KކY��}��"OLt� ��l4의�t�0�8B"O��h��X��(��䏾�*��p"Oإ���bPb���jD�`�Lʁ"O(�!4A,~8Z�C�J��j��`Õ"O�z#��?��)R�'��\�@t��"Ot]*F�?m{4£���4��2u"O>tz���1~	��r]�:���I�"O�|�g ��l�R���W~�{�"OHX�څ�|��mV��W"O�1���B�*�/�	Pa��c��'�ў"~z���Y� [�W;jh:p۲�ؑ�y�E�ЯĔc�8�
�%U�yh��
����a��1�����y��[�=���P��W�n`Aae��yrg��zݘ�zp#-PHb��p�R ��?���H�,x�2f%��7�)"d#	�'�XE!�eX1�4�1�%*���'�P���.'^ ��7�d�̨�'���$�Z&fd����#m�x��'�����@�h�(��[~��'��=����/&��)�i@��B�'�­�$IϽX��i3��T!4	V���'�Ը�歎0W� �N�'vL���'70@R&�xԐ��xUJ�'�s���}�-r�)��{��uB�'�� �J
@R�x�s�+tJ�P
�'p��B����-��z��'}�]��E�(p�|Q��te��c�'("y���rh��됇A�c�D�)�'��)���"�@���dc���J��x����e�,i��lʆQ��k��y/�07sv�C���!2��#�?�y�(.3�-!)	�'�B�b�]/�yb��x�>Ypeфwq�	�O�yR��dˌ�Xb��h?�y�щ�>�y"��{~���f.�� ������������m��g݈j� �'*a~��{(v�Pf��r��ً�͒��y��ĐVnҐ�7�I�r��gױ�y� L<�1�F�o�v��`i]�y"X�)�F�:������K� ��ym���4TP(���qcNi�	�'Y��!�D
�����@�g�u��'AB��Nζ�zlIufژXȖ\��'�!�$�7q��Lbf��B��څ�[� �!�d΃B_�M+�ft�7��-�!�� [F�a�B.�,�)j��3,!�C�PL��d�/�����	+!��8�2��Wk��gMH����O!��B�v�t&	:���@��89H��2O�S���>���(yeTm��"O�T��l�p�i���hxp�_�tD{��铴D�L�ё/C-T����r�ޝ=�џ�I{�π $,�� �?�r@�"��e(yv"O|�y�&�:XְA�F^�k;0���"O�A�F��7��1ˑ�{#�T)�"O�K���1h^lE�c�3�P��"O�a ��x�x�Z�+%+<	J�"O���"���)�@�OΒF��yb��(�\��5�A�i8��@Ǯ��y��P�ޭ�D
߈v��Ƅ"�y��~�� !,��u�)+!����y"l�UiJ�JblA�pڤQ��y��<)�\HcG��n	D��F�*�y���T0D���Hi�L .!�y� A�Y�����8����D��yr��+���$�>b�2ѨVCY�y" �b�e#�_�S�P�bqK)�yb$C�k�, Kc�M�.2�#����y�`�5l�f���c��hq�gû�y�lY�V�N��6! 1go�}c!��y""Qb�T1� ��X���{��@��y"��:�B�h���E��y���9?����
z,�a��jW+��=I�yB��GV���mR�jӺ�+�����y� �@hQ�Dj��`���ȶ/��y2��[�b�℣��X>��6
�y�KB�cv�؛X�v�xŭ��y"CR�o�����Qm��J"��3�y2g.[/�����HV�0�ѥ���y"��+H\\�a)G
��Br�1��=��y�$M:��͐d�$&"��gP8�y�eK4(t�Тo�.k0����W��yb�̲%���;6�t�\u��B���y�؟y�r��� ��=%�%9�+���yR㞍D\���d
�f�|�2T��5��'�ў�OE8<
�H��Nv���U��,A���	�'z((H��T(
O���u�۶h���s	�'f��� �9�ܤU [�_R؄�t�N�K���-}�:X��n4
	"m��ZҖ]b�\9o�@�Q����!���ȓ3Ֆ�#��3���ҵ�'p�H���p�����ۇ�^r�Z��5b+�n@���8��Ո��S��3�*���nʞ܀��|"�)�10H�8r�$L�^������
e:D�O��=�}J	�qi@����6�n!��a�<���6��hdF>Yf�E���r�<)��4C�j 0��$bq�9XH�<Qr�H�d̨آBI�x��[s�@G�<Y���6�Y�A� �mv��lAx�4Dx�����Փ�)�J���*;�y�Y!�0��lM	jٞ�C��)�hO��𩙀4�	�3��p����)i�!�d]�{�P�0D��L���E�D'{�!��C느�1F<S�	����g!��2f=2�`�>"���mU3L�!�D�9�^�Ó�_	j �Y8J�)5�!�$���L��d��B�ʡ��od'�'a|R�T�?�����l /����g%���<Q��d�UT�����Z@�P��W0!��ҶRX�@	"�V�e^L�k��J6<�!�d	l��K��7EV��#���!�d�>.�3�'׿v�����Iş�?E�%I s�q�o֖H�h���Ly��'E�O#|rr�V�ri�Lk�D�a�x�9��QQ�'�?-K7�V�8�@Y�s�[�H� rs2D�Ti��4J�nA�p�1V�Ji�c/=D�� �<��q�졂�5'r�z"On0�D	nh�b&�"{.A"O�eS��L 	�(_�xhI���|��)�ӊv��)�d^2+z�Z��1�ʓ�hOQ>�(�m�J��*���l���B��Ob�=ш�	J�p�ѡ�͇�{P��bW���!�� ��ʕ�
2?f����ŕy�!��
Z{PL�e� R����D�ǋ#�!�dS`u��x�1-�4p��ȝ$c!�d@<�D�h��X�)��:��Ϧc^b�)�'u8�C��Jh�p��B�.���'��"��B�kUL!��i[c8<�
�'̶p���P)'�ڠP��T!���'K �1�Ŕ8[�	�� ƁH53�'M�I�۱h)�XuEҜ`]�q(�'��K5�S"#V�@K6[�����'�xu�� X�
�E[@�j����D8O�A�D�]�y�h�3�B&|�,̀$"Ol�2$��?"�0��rk�n�@�;�"O�Q�C�?#�Ȼ�`ș!�T���"O�:��X�F�D��r��/qE8�{ "O�YFƃt�h�Z3#].s�5V"Oʐ�c'�7!;^A��`ށC�X�c"O`��Q�&Ȃ
����&��+��'����}׶����q��1y�C�ɸv�,	�,6NL�v�R����þv` ��T�9� `�wHթ%7!�$ʭ[�Ʃ��댤<�֍0�F��'5!�$�>%̰Y�e��&|��  ���/,!�d9c��0�4F��aÉW�M�!�D�(,�8%AU��s���z����{���B��d��b�<	�H6���s���)�Y0��^����'ϙ�9=D�Q�'-���b	��Q���P�J�C�ɢ�'g&�St�PV�8-�ЎQ�j2���'�4q���{Gh��G��dK$���'4�� j[�,nlmDB��U|�-#�'��4�W*�0Ქ`�EH��E*�'t��9q�OF��3���I�����;O��Z��CR�4A�M
^Jr"O�H�̜�F��,��8�w`�
Q�!�^攑����?��`cE��?v�!���v{��qբ�	 ���Z�`�!�	�^���F�d�V���M_�f��}��'�d�8K>�1��m̑��-�ROU�=h!�]h���wK�'[�u�m�ў<��	��Q���6��eq Iv��B�IM��@�Bق	������bB� ��ph���(?�~��o�`�>B䉚cZ@m���x�dE�	%D�NC�	}5$YGn�j��#3��ON���g����AA�-�ƕ�����i��f?D�tR`���kF���Ѓ/��h�>D�H�r��}�V�c¦�)/�t�p�;D�� g�UM]�m�� �O�t��R�+D��;p�� �lI��K����rJ+D��bS�X>fv�i36,�!N�]zr�'D�()ĊI!Y�ٻB�Z*$�M��'<O�"<��gY*�N"�o��#�����J�<���ծ6|t\��fѸ45h�RB ]�<�sJ�U��-���7e�* �Er�<1�Mgx��i�ŵ[�)�K�k�<ɴ�K�j+����	.yvd�A�`�<A��Ykb���Õ/k��Z�BX�<� $
��G�_Bl�ѡ��7�Fh{�"O�=(�Bz����3@�B|�106"O�Y:��I�1��;��Ez�t"OB���-�k��M�,�I�"OQۡO^ ��`ss�@8,�"��B"O�i{��̊	b�%��n@��ޤ��"O�YƊU�w
N	�P,�ܵ�E"O�ACFLܑW���3�*��h*،��'m"�'��I?������C!Hk���w�<���ȓ}�=S7�_'~ �ElɆ,{�ȓB�y�7ǳ9F��@�?aX����|zB�e��<���G�Ȑ �~��ȓ8���:qˀ@|�E�ԍύ#���ȓT��QSv�_;�EB��[�H�.A�ȓ	y�����!�"t��:$���]�����V�7��D�7g�Ԍ�ȓ^���á��ȉ�!�3^"�(�ȓe0(h��A� �ҩ� �ڮ1� ��ȓ�VA-̜MѰ8.�<�s��k�<��E7qV��H�o��@-�e�G�k�<iJ�Ka��`��X&
80��c�<q�C��p��D�<��[�ɐb�<�4�Ԑ8P�e�5��6-���a�<��/s����'�0!�Ry* )K_�<aK���hzP�8!Ė@:�b�s�<a�O�=�h(���$J��h]q�<�B!#(i57n�D�Y�!	j�<��j�5 ���ǫ�(5~��P�p�<�3�����#a����0�l�<9�N۳w�n�2c�dv�R��K�<!!2lЉTn��K������CP�<q�%é}���3��z�ȁJv�N�<�V(߹Y�" A��Rx0!��I�<!7	G�k������V��(X�@~�<�4�X)�9	G>ϲ��rGIp�<y"됸�W�4(�$4h��p�<i��M+Ƅ��FL-iTXA�m�<����%s(� �� j�*`�sn�P�<���
tּ�����:��٨���v�<i��^ |�]��MÕ(���[҂J�<iQK;w!�i����%�t�F�H�<4�F/ာ�Lε$�B�E�<�3Cի2E&$�0��;k�@!�A�@�<�D͟	�髰��f,��3K�~�<ᇉ�TU�T���Y���#�Ld�<�O� ��`z���4�,���M�k�<���Pp����IHv�]���f�<`(T )���f���� �A�H�<AQ��	"T#�&Oplh �D�<�QH֦\x>$x '@�b����!�B�<q�OԤh�i�ŋ(R|�k'�|�<i��V��mȣ5S��� �y�<��EtH�k"E���@��eGs�<af��+�6Er&댉���q�&z�<!��o�6��2��>G�(���}�<�c�Pe $�F �:sL�0$�|�<��b�����Ra&
�r2�I�fv�<���j\�XJ� V.k_fـ�,Fn�<t*C�)�`{��-KS�EZ b;T�삵e�AN�< ��U���%L#D�����E M�l +��.">�p�l#D��S�ՉE��	�1�?v�TEӢ7D�X[t� ��0YUo�	�zX�(D��r�n��NuXx�wDF�-xʓ-$D�� ���aB"!�b��1��	o��a�e"O�联`J�`Aژ����n���k�"Ol����4���X��Ӌ@~��Ja"OJd!֡� t� ��D8nh��U"O��	�D��Bޜ� F�H�V��V"O�R(E�ij�c�o�s�H�Pb"O��seo������
N� �"OR��a�\��y�e�݂"�h�bs"O�h�˯f�t�Ε*-9��"O�K@G/:��Ս�!F��"O0��9zoX��2�
J����"O� ������� )H1iW"O^0�N:�)� Թ!	��Sc"O&X���7v��q�L�d��Q"O-����|�����1+:�zt"O���[, P\�A,C=P��8�"O�y l�'[ <��+B$ �`	��"O�-�B@Ϋqi�	3@�T(_.,ڷ"O�}�D�v��0���2\�"O:�X���:R讽�i��A�vr�"O$��P���7�L��(͍ �:���"O�M� �ߢ,��(��f�_�@�"O��ЊZ���[�&4�v}�A"O�R� �m��J3�_�n���S"O�1�g�mՎ�IE�/��pt"O�v����g7p<ҥJF ]�~�ȓgK4��!)�2y�H�c�L!Jd���ȓ)��5�O�;�R���l�X��6��e�šf�"͓�gJs�⹅�����kF�qjݰ��^#M�}�ȓ$~��w+�O(�h�)�W�(��^��9��9i�a�v���$��E�����$Z�`�aYw�����b�
�J���-!:YH�!��Qu ��D�\��O9%���A�d�؄ȓq����CG�w� )���.��ȓ
B���C$muv��p��	f�D�ȓ��9`J\��i���1�DI��PH ��.RdmA1GR.G T5��q%¨Qem�8p����#�1���%�V�
��W�%G�#���[��l��}��ˠCZ�&R�2�莓�,�ȓ'��TA�$��OmZE#4J���<��|��� �^\x�r�j��E ��ȓAWF�QDضh��ȊEf۟�$��ȓ$�`b�e�C���甚Id����<���H��K/6�0�G*ܼ8\x�ȓW�v9V'ǘR���`W������ȓF�t���}�@@�3@�ņȓ>K�H��L�pt��1N�Odp��ȓ�.�XFb����`����Z��+�" x����L�Q�w�<J�1�ȓ޴���N�j`rQb�;9�����f
T�nˢ�
�ҁ�5�h��%�	۠O\��f��A.�.$��ȓ`� ���Q=�����ԧS�� ��g��8a���*I�L�B+YT��Q��^Yh@S ����ô!�
s����>=AT��`.�$8�!&WR��ȓB��� ���4Iw:�kV@�*x�̄�	�xa���^�+�㈱Y�)��4��)���+?.lP�d$�O�,D�ȓ r�	��$w}�!�Q�u��u��(�Ұ�%S*6Y�Ayb�?@����S�? ���Ț&r��0�@�_�Lr&"Oh�B��J��τ�|u���"O�\��fC�\pZ�AsMV4Jt����"O,i���P� fX�0��նLnrM{Q"O~\�/ؔ�� �*Q� ^��#�"O���B�I�4�8"$�,hY )��"O��*B��c�T�D��IK���4"O:��C
��J���)@�\1R�B�"O�m��b�����@��f���"O� �Gh� +&��)w�O^B$X"O�;b/�&�lء���9H�,у�"O�Li��('��9Җm��/���"O���Q�՘T��kQ-��v�&"OƘ��H�x����R[K:�1�"O�-;D�2�
�j��_0Lg���"O�$�f�V6K>�p&'�BNh�)"O$D��N�ip�HA�W	f�� "O�y���~D�S�U���!��"O��D�+4X@�"�9� ��"O��%f�H�PdbW���y"j��"OT ;�N߼g��t@ꘊ\���"O l�h�X���@�d�� ��"O�pѶ Y0��臯�c.8��"On�������`G��9�`M8�"O~���"����G',�¥2�"O8��(�! ��}�Ɓ�cᆠ��"O�����t���y�V�8�F��g"Oyzc]�d4�p�����t%�f"O"��'��#'��p�LĠ,��1A"O�i�/H�@B+F���2"O�E偏:x����R�	�~��p�"O$p��J�-3� �B�͊��-�6"O ���n�+�Y�u�'O漴��"O�MÃJ�02��a�GM<�X�3u"OzX��W���Kܴ!,+��_�<�!�|�����E��D\��q�<1+	�M65�H�7m��p�T�s�<A�Gӿ{�Е�VG�v�X��gA^p�<I�*	I'��8�mӑy��Ҍo�<�p���w�z���`]
ښ{wOi�<��L�v/*��"��h��0�Rj�<TI�X`�s�=�����i�<)���TV�
���"8H�ȵ�Ig�<�!�W(e����l�\�&�HSĎf�<a�/T�Z�PA��G�aa�h�*Vd�<)5��E��- #���PED @Ī�a�<1����-��1��s�@��#�]��X�>1�C"b�lŲa㘗A����T�<��b�<OЈm���F�&�.����QHܓ�hO�O�bP�	-dNF�pt�M�#<�p��A.4�܊���(rGJP*�M.8�&%G�nӨ�=�'0��O�С�`�3 ���F��V��}#�"O*y�� Ǔ:�����"[�bxH9�BW�DlZo���O_�QCjR�vS�a�� ���	ۓ߸��$ґF즑:B��=2���f��S�<9��Ex�Y�3�:��i�F�'D�?�X�Z�[�jH�� �R|�`�N"D�\*w��d�v|����ZU��Ȣ-?D�x#&���*�Avn�..�Y�@:D�lq���K
- ���U��7�e���O��Hkk�;��!1@�6k�$Mq�'`����4n@:ի��&-L���d-<O�SF�Ӫ��J���!D<��@"ON��`@��ntqӪW3U*��"O� �0�)Sάݸ�ŋ'�5�"O��('�эk�	�'/%�3b"O�qІ�N�}����SA˗]l4j#"O򱲁D�?�ZБ'#�$]MlX���'t�b㊜')�E/EN���I�C�<�����1�py����\��E�ì�?T�O6�=�}R"(R�r���!~αAm]U�IN�P��ɟ�-F��IB@��`���R��3�Xl��Q�4bp"�CB�vB�I!s�0qr���y���k����>����ie}r��غ�<	�1���<	�JY"p:rԓ@>G��8u�e?�
�(����c탁PPS�h��v�܅ȓQ�h��]	k��2HK4%���H��l�umB�F&��:��4T����/XBQf�>Оp�BN7z�p}��7�pl��I�#ko����1{�@Ʉȓn�L�rю@ E���f� ,i�2e�ȓX���ܼw`��9�BS-]���'�͓�M��'�� ��ф4�PeYaA>|xG~��� ��o��
�1|*�j��$8�:��U�O-���<�O��zх%�xx˛�;�`��r�-�I���p�SG��	6�΂t4��tֆN��t˪<)�MS�]���#��Т�Y�`�Q���<�۴��훶��3��'|db�%U�U��|
�kX�w�J� 
�[��P
:
^���ֹw e�a��S!�xAF����e\9�e�rOQ�����8u� �S�J_�5���튣3~B��5��h�Lݢo��x	�I�e�B�I�\���Ђ�54n|��oƨ#?�B�ɲ=���'(� yMJrc=O�Ft��%C:�D�B�F ���i�a�	]�����?����4:�X��(H�zNT`�I���M�?�����Iq���`����V�"٘L1U%�[��b�"O8Pbf�ִzr佐GK�����V"O(${Sg�	:�*)�ƹ��'w���=	ߴG�\h9��v"԰�ץ��n/Ԅ{�O�8�gZ�5��#���34����>q��X t�O���i]�T�f�#�ON*�tX�"Ox�W�Q"!��0�d�� ��T�|rΔ� �ў�Oa![N� ��$��a�&]�p�	�'��5��(̯HKXe��.������$D�<h7o �:��LZ��&Q͞T���8��>��>9�'��3$�P8S�/��
1D� ��l��|� 5'�
@�݈#a4}r=O�c���~���Hq֐�m_9*ٙF'i�<� �L�iE� �VcPv�5�tJ�n�	P��Gyb�x��=��U[b ̩ ΄2�	^��y�jO=5�ԑ2�%/hH ��ȜҘ'>ўb>9����(z5��v�I8ĉ�c8ғ�hO�>I������08�9K��|�H#=�;��,Q��%�������3#w8H��[�>I���I�9��1M�ڠ��J����A�{���C�@�3ܰ��B�VȢ$dUЅ��5i8��}�<1�J�.���k�7�)���|��hO�O�����Bݏ:�@i��D�vY�)��'��b7gK/+�� '�-^�����'�b���n�eq8x��T�l(�'z�4o�e&j��E��>},�'qZ���&G#~����1���p.��
�'�������\�YA��@E5`
�'��y[���AJ(� �=5��i
�'���ʒ�J�8gԸ��nL W�Y��� ���q���Vzl���A#F��""O�52�@�>sz���ˍ4?�h8�U�>A�'�O�(����2����!	A���`��*O�(���g�` �3�J�B���Ӊ}�i*ay�hB�d�,A��Q40�:U��n���p?��Oд�K�$�z�c�<���;"O"eǎ#&��v���M�������OT7ͷ<��O�Ӎq6��Ea͞f�p`� \̲B�vK�([L$�KE�.6�%���Klܓ�hO�O�pb5%��T��͑a�R�?�%��'Xɐ��d����IA�/���M)�Ĥ�TG{*�<�b�)
D�&���ȏ:X8!0�'�Q�,J�G�k!ޑ�F�B���A�$D� �0�?�*�DA��mz�:�l"D�ġ׋��MW��U�"JLl��g?D�Ƞ0�֔2�&��2W�0�`�<D��`f�B0xM|���H�C?V���94�hy��j�Փ�KR�#0�L"3bOB��Iq?��{��)�?SKB�e�%/<�Ӷg�)��yBa�q�R��Y"��@~(<@�� �BqFx§<,ON!��"��GU�榖�20Д�A�O��I��h��Q
v��9HZ�	�טF]���j�M؞L�F��$K�ģ��ݐ�0���%}�]�%������GT�4�Cv#��ȋB�Ùl'!�dOV�t��.6���"�\86Q���I���)c"�� p�L�K1�ǈK
*B䉩K�$�i�E�R�rd ���U����'�~BN[�]���z6h��Yd�B.�p=��}r��N�P�֯�$k�y���^��y��w;d�t�� |� FDǦ�yɄ6!� 5@��A6��q��y2D��D���ܐx�B�qVk��y� �{���/Y�p����y"�9}�(���R�i��4���.�y�T>x��1�A,�a��C%b'�(O@p���ԟ&�r�f�+�
G^�w�!�1"O���S�m��LC��Z�$S%"O�����!P�� �N�3o��u7�'�@UDx�8 �!K����v%���C%�y��O�Q�n�c����r�*@�C���IN���O�L)#��4�ا�]�y���'�~Q�ƀ\�l;�	G�0��&����'�R���	�t&\��+^�q���?x>�B�ɣw�i�&ƠAطf�n�|B�ɓ$8�9�Ci�6NjU`3"�)^d���,��'���Ȇ�G5ڰ5y�kE,'��	�'~U��i��Xiƕ(e�B�$2
`�'S����ȩ�����E������'n��e��"s2���i7D�Y�'�r�
`
�	�xq�R�ʝr�Z�y�'	p��І�:��$�fCO���I�'�pd"�*�uJ�;C�Ԧ
i(��'�`x���;@j5)��Q����'��`�r	�c��uCe�̶C$�%��'bL�kU�f��X�d���l�|���'�,	B�§|��sD@!]�h���'�إ�,�	cW�m����$N��]	�'{.���<=�0Rc�Nr��'����gg��G\LB4���n<��')��9%��3�����ܹ ��4��'z�Y��	Ϲ5���\%Fu����'Ɯ��ԧ �x ��M��pJ-X�'��A�!¿Ov�������o_����'T�# 
E��D���K;nn����� ���𦑰|�T˶@�Y�Zm�g"O&5�`��.6��a ��Y��y�S"O"{dƉ�wv�X�����h��"O�mSe30Zy@.�T.`��"O�mx4ɒ�R��Zp�Ѭy>E�"O�����X�8�}YBMס|�%1"O�D+�〯\�bE:-�:.$�f"Oh��hM�y,�"�͍2��Ӑ"OX� ��3��`��$�`��"O��2�� d��h�*�����P"O��I�o
Z��!�pc���"OJ	��_�F�̕[׀��3�!"O��6W��� 
J.��p�"O T���ÜB9 yӃ��{�tI�"O�s���n.NY�G�>W���*�"O��Z"��)G٫��}���w=O4��$Q>=n�ݢ��ݹv،�"��ɧ.V�a��.@�Ҡ��/�
A�C�ɼZz~Lsv�,���TЉ,o�C��pd1�F%~�i�5�N�@;�C䉐/�e�V&1Gxr�F�N֤B�ɑS����3�2$<�y	�!E :~pB䉕e�"X�K)�v����1l�tB�I�U����D#}��� QZ�B��?tZ�ls�d2�� ��7q��B䉤g�6��X��p�mL�]�`B�ɏt?���������A��C�<X��!͗3����#�H�:��C䉂P�pP�f�+�|����Z-�ZC��6"�e;�o����2��V�/d!�J>4堶��%tf�C��1&i!򄙔�����)L��뇦�"I5!��ڳM��M�L�n+*p	+���!��T���9V�B�vfѸ��,�!�DA�SHD��T�ڂw��3�P!�!��Cxx��t㝄��d!�?�!򤃑!֮5��L��rm�Q����!�D� ���9f�
d��gA�%`!�$��}�n͓�&=w����w��B�!�d߄ �ơJ��Źc¥��BF�[���0@k�~�OBɚ@K�pB�\k���|��
�'e6E��C�R�0���n�4x�@�I��B�<➠F��'�U*@*�Q���A�P�)����'����+]Z5x��.-�X z����M/a}r�2FLl� �<R���di7��=�Q�8L���/���c++��h c�_�A��!LŪ!aH�Mz@��2�[g;h�?i��E"��
ٱ-��Ԛ0"�-0���ڕgS_�<�;d���X�ݧ#X2���2���s���+�g?٤�֊� p�f�J��~qJ���y�<���Yf ��%�U���y�O�ҟ� ��Ɠ\a}RK�<��}�6��%.�����%V��0>Ve\���´r�t�	 �qҢZ�L.��	�'Q$E��Po �C�Jl5N�h	�'�tQ���И}�,��Q#�#Yx�ܛ	�' |1�f��5Ej	!'ڞ*�r�����#j��#}b���"�F�#PB��Y�Z����HY�<�w̋�rb�b�LQ1(}jŚ2��<9wƁ�e��"~*���h�a��1+��m���[�<��H���~�#4C�C� ze`I~r��(����ɣ]Cna`����*t@Q�Q�T��N��$�f(�:r�Q>UD�1��
8��1V���|(!�D�?�<Ab�M��-�`��a��.e�d�G��KOQ>9��,�Brb�2��3{�, ��!D���pJ�8T��MU�:p#�}�0�3��03�qO?� X �ԁ��Gr\�%@64�hA��"O
|0��3,ơJp	��;�x����>Q�`�ڰ=A����b��%=�-+�J^|�<�Ё�(��H�&n� �P�K{�<ѷm�2������D3�B(pq�Lv�<A��]�wF$$�כ��u���e�<�!%	�4H�"%�/N��L\�<�t��01*l�s�Δq�����Z�<tǉ$vn<��B
�MQ>�C��N�<y�C�4t�X[fFԉj�-h�\�<�$F��O�<=9��J�N~�Ax"��C�<��@FA���˗E��K��} ��U�<����Z8¤
9D*h�V�I�D(l�'�:���e�����-��Q
ד~���sS�E�v�����O�9f/�=a���tR.l�J�s��9��Z@��[||�HFF�=��Y���"�I�<��M�� ­J���G�	eg�D�K|��e��]sK��9ؼp��E�h�B�ɧ#��Pq�&�=��	"�$K�`B��tkh4�íݡ0+XL�č ��H����  �T3sC�pt��l@�C�ɓd�`�4��6��<��"�	�$qKƍ�J)HE3��K";-t����bޢ>�w��!Ǯ|�УMb�i���mx�t �AѠKn��	'a�~opI &��9���@e��;��d�ٰC~���Q�*�)��.J$rǰm�/&�d
�qͨQkr�`�rd�� ���PGL;
�i��t
��kF�A�V��b��H�<Y��NQ���vB�>^����E*Ʉc��tp��ɾk,�ųE��]��tP��t�ר!�.��fPu�`	߁G�l��J�<J���dC'��y�f�\:X0J��1�Q�l��}Z�.\�l
ҕӕ��O)�6�_&��QF{R'\'���Ȟ���h�3/۟��'w�m��r?�5h8��X��oZ!y���e@
1;��;�(�{��"�-
�8��IA9R��}��)'�{P��	~�z�/�	Z`9�2"�z?���!X��+H���H�-��<F 1ü��׺z�=x�����i�
�Q}���2|��O�>�r�%)U�N1�𮅤��1�E+$Z��*�n���Bx�A��[��z҅��V�@)�Ў�?��rM�O\AǏ�.&k�!Sr�Եrw(��`�>Q�(�!�	�%PiS��<����b�hH5c�T,a����%�<)&N�Q9�	���H hd"ꁒ`�b�h!�� c����Q�����AY�d�IXw�� 3�<���f�~g�`	�5��;>�(' �.��aΝ�|1$�fd[&x<耨�Z�$*%��("��bU�7�O�h��F�+N�"Ѻ�cW6z���ٔ�OZe*�IW��~b�R����9���H�$�̻;���H��Y�j�ң�B>��A����$�7�)sb9�Yl�`�-���A�C^�Wh��~bdV*e��R�мG��|���INv��'C���I�=��� ��
\M�6r��' �����\]?ɓ(��Q��֝�W\����m\����q�I�î�O����#w�b-!�N�?�$��)2�D(R�K�R�D��	�t6��!0�A<0.�H�dOԂ1��9�
��!�%J�{����-ɻ���Ӌ,W>�+�P������1���>!y��w�^����(1J_S���)�KK(2�5�0���x��i��G`���2S�i��Ȥ�?OF���0�%�p��}���:�y�FV'{njF��'`/�Ya&��p?Qq&�\��-I��
�
�Sj�2S�D�{��F����I�0�� #��r���ܠ�p�8������)�to:��̋J�<a�Wd%�?�\�y��3�'L�������I(p��kѢ)qέ�h/?)«��DW�sI~�=�$��3�����[��G}� �q�O�XS��Z�q�R�@άr�؋e�Ѿ
"�ˡ�0?	!fݮ0l�!���PV�
eh8������%@Xy���t��p�;P�B	@�*%�Cf(D�PCg�)V��c�ż>�}IL;}�g��|q�)��v>	�p@�zSh�D��(ዑ�;D��B��;N�UNC
3bYbTM�#1�'d ��H�O�g�1Z��eǙG{|8Dm�4O�XB�	*�dJ�%�w�(�9A�-pd腨�`J�BP-R��'�����\O��A��$Ap��sQ0��^�Q��7upˇ�B�G�mC��� [�9�ȓJ�>�:��*V�����@T�5�(�O���AA)ym4Yç�J�PP�O�Q�ʅ
u��K�6��u0�`�S@���Z|r��N(Q��Mp'�/���(S��Y�~&�@7�ЖK[��IpH���0ѡ!4�JSnN�>8 j�!�7 ��Px!�ϼ5�������� �� l
�k\�+ �H|x
��ޘĠ��Y��L���S���g�!&`]�$'EyǢ]�HP<��_��95��"!nI���F�T��9���\5$���d8au <����9I��x���jNzeP�-ʮ4;�O�y�⋍�4}�8����>h
��]��m�֟BHy�_&@�p�c	U�Υ� "O>���W�B�k��?C�4xe,�B\Q�H�:#��Ă���S�(�9��Ġ���ug_�fGڹ��+,1��Ƭ�q�<��U�xX��*l�ł�%8�B� ��F�QNv�qf��Ud��o�	�l�<��'Ŝ7]<��A�A%}�2Y⑮{���J 	^�J�l���yv�r�+O#�4œ�&M�6;�/�.B��0�=�p>���"�\Ԉ�O��~G����F�nܓ"��]S�V>4�� Q�B�U��+�̝����͌X�Z��\K�q�e, �!�dV$�Z�ےAն^M��K5ˏ�fru!2�8/Pa��Ě<U��sf%�^�˂U�_O���s��΅�N��mP��T&)!���"H!��*W<�pӫ��;Ő� R�B�j<�R�# 0� mA I�D�O � s��9�1�r�a�Kظ)�X+���
� �[P�'��5�rL C��ϓTm�4(3�òM����)V��{��	ß(���[�=Ǽ\��x���D��mV���Q*<M�1�Z�f��Ov��F	Y1$�c>7�R1e8XL��#�3cH�izb��O-�`�H�c6c䘧�0?1O�h	
�s�L `�̈��;r�PĐ�0O��/@�Mk7���
<Dg	�F������y�����tI�
ݛ[�T�̉��y��Ѧr��m!�! m\����X7-)m:wH_j(�pfDT�u���B/ðy�v�+᫖5YtP1pƏy��Є��v��Ԁ��x�j������=�b��M��7�VMa�@+ʨ	��`Q�'Htl��H�T,��kr��{'� ÓG���2�^�PrB�Q�!0&�B�� ��T���%^4�A��@Cxz!N�e��X�@BG�x�4�sg����),?y�N6:LI�Q�
D��`�O�%}�P�1Uv�T�Z�&�y" l�wT��1�%ڽ�yR�"q<��p���4||����J7�d!�c
�E�F\�G�G�Zg�p ��aXc�t��rq�\��/�7e�hta��%j�x���st�t�E�}b $؂-���GEդY�h�wFb��U���<𬠊#�|�B�2e4O�r,��.<J�!��+�I2U#Зt��Sٞiq�l\�L�Z��UG�$y_��	>w��5�22	#�ݛB�A*��M����`��&���������S�O9(���"ފl��P�(^>��(�����(-��l ���B�Z�Y F� �D�@A�|�	�>	bǀ�!���|�<1V�!�n��#�Uܒ8�0*X�<�J�?�n�s�)}����)XRP�b�؞W��%P��EXL1PS�Ŵ*Є�q��W%��� ��b �`�L�J~\T�'� b�՛"����'��B�H
��'����F+J4>=�XZ�0'��@	�rF`�Pu�C�|�׋�>#�Ȑ�u��p� ��<)cbV"J�b?mӓ��?
�:=������T3p�0">����y�]B`G*�5i���(&'�7\����1JdB�I�o��1�%(�½�ei�*r牛.xh�m�Z��S�O�(�y��)�<����n� !�'O�a�7�J�b,�B%G�.,a�m#�O,LP%�O[R�4��Qq[B�A�b?| 2���OJ�P��	�'@<�J��Z)@��""'�F�)#�kƳA�6�*�
O�+c��cjxD��Z`�(r�vc\�!�¬�q�T�A�eI�x���Iw�F�[�"O����:iR�т��wdj}�;OJ��F�ܬ+�*�qO�"~�AƉ%y��͹����0��f�<a����Kp漒�N�)=�^qD�j��4Q&�*¨<,OdY`4�5(*j�(��_�f#�lH��'h���(�!��y�񋟪�P���8 ���t<hPoV26�D�s�U�T���~��
b��(�����E�FՆ�4�V����	� c��2z��ȓf�j�	J�r��$��Z]j<��j?J�Ɯ<u��2cj�&l�|��X9y��O�C��P���R6�ȓO

�B9/w��5� rxņȓVL��*�l��cR�y�G?����ȓl�l����&'������F��\��S�? ��z��&ᾰ@t����T�0"O���-��B����3C�$#تi�"O�hj���o�ݲ`P$nB ��"O,�r
��k�(�9 �bCp�(�"O*� F�*��]�rC� DI�XR�"O��8+%#q���'A�%L68���"O�A �,I{��}����Y#l8at"O�e`��O�G��|j�͘%��QS"O&���e#�D,�@��4��a)d"O���FM6�QB�+$�Iې"O�4{�n4
T�d�1O�'+\1�F"Ov�ˁ�ߦ]����sn�O�\p"O�T���?omN�����R�zr"O4�)B%�G���R�l�#L����"ONU��-��H5n���ƪ-\��"O�}��Iԓ
4j��ɕ���6v!�D�;f��{�b��l�
l�$ʀ*!�/#�̌2b؋P�<���ai!�$½�65�b/֑`�����C3&!��}�J5�5b,&Bȑ����-�!�Q����a0�U wf �@�H#�!�׆YU^�eD�x^�1fa!��ju¤(�˃9''�d�/�85!�d	&{d��Q�Q8;��KT+�6!�ۧs��r1�� �� C�#x$!��Z�M}�ԯ�8QU��wm[�9!�ې%�T����v�D��'��!�S�1��iyD��y߮���D�i�!�dV�_�"�34J�%(��<B��D�*H!�D��zXpIG�$9�$u(�B/3!�D�a0���bO��6&��x�!�)J#!�$�`��s&"X������R!�w�x�i�D�5��pU	>!�dNH��,��Ӕ��PҒB�5.!��.W��R���"؂(��a�/F�!�D�(�>��t���P
�%�!��N#S�F�9���*D�L�[!xS!�Y*Z�Z,yC >$D�`Q0.I!�$�Y��6�N+hf��J�<^!�D�~X�J .ܿ;B��E&HK!��ĭU4����Ⓩ>>
��%��<�!��-��Кc�3|�u�*T�d�!�اv�|t;Rώ� A�+f�Q��!��!fN�ҏC�&f��8NS�~�!�D�+�\%�R�q8�LR�,�>jӴC�	��PA�@/K+-l�'i�H��B�	�f���ʥ�{t�`��ܵv��B�ɡ<{��cWK��*K�+@!�8E�B�I�A�%�HI
��7R"B�3�f�r��m���/W�$�B䉳7�@�KB�?�a�$�d�B�ɠd�N�Жd���Nm3���-�:B�Ii�aR-t�R�!a+�"��C��)Vw�}z[�Q,��A��C��C�ɠ4������z�a��Wx�B�	�u�=(Q���6lq�cc�#\-�B�I��z�]�=_"Az�)1Ib�B��`MH%ѡ�'/�����7�tB�	A}��5�ƨ#� ��M m�BB�	r��L�q��>O��
b�޴E#^B��&.S�Y%�G@XȰe�ҿg|C�	�.��H�H��WY��Pdm�g��C�ɻ P�%���=G�fԀ��)]�bC�	/�t��#�ҝdɛ6ȍ<�.C�)� 6�	g)�f�,�Zp*W/���;D"O�����N�PYx��6ݓ0��r�"Of%@��3"�.��U�تl||+"O�\�5"�
-W��bP��/^���"O@�a���W���Jd(UR��C"O�1Q���n�\��gC�r�f�"OlЂE��Z��h�U��	�daCV"O�ؠ�ӫ]��B�Oc���"O�5�e芛G� �*Tg����j"O ����N��%�'��Q��"O�a�����t�]�U&��$�d"O�mD�#!A�����X�|�B�q"OҜ�Ĭޘ ����So��8�\:�"O<��l�KӚ�*��Ϣw��њW"O�B�i[�hl����˞)*?�iQ�"O\ݣ@$ܭI�9Q��~�A�"O����H7c��͂p�מ+aq��"O��Q,�v�Hا$��k�:I"�'�!��ڢOD��I�����/=G,X�׃�#8�C�I7��X����
�9
!�	�Q_Vc�<aAI;SZ\Q#.-�^5f���-�L�M�fBN�!	@���bS���ό&Z��Aƀ���F�0[��`��O$$M6�3}��*G\�Ј�lS�OtH�����x�hp�-�U��
pj�̪tHyY��p��X X��0�*|O,�FhF�)oVy���i|(`��'m\e�uk�op0H�G��O���'��Q��i�	���>�Q7"O���D�ӣ~jF�jU	��y���C��|r�I�|���#S��K!:�}�&V�Y���1��ԨH0"�Y%l�i�<V���5��gT�G�tEYC���g9 1�0�"��d��I.�?�'��i�$#��=r\��O���2�'�08��ǭ.6<�t�1@,�9§���h�C�8C2����_.92��4RLآ��ʱxe�OpU)6�-�~"��5QB��SkK3{`�d�)��dcq�ׅwi�4)�hD+-�!�$G�[ ��� Q�H��Jf��Ppz �U�̝�~�NP�2����3�@l�T?���wy�1G�\W4`�����r��'�$L96��?{G&စ�V+����b�1OT	�oBaմ��Ē���'��ZU��r����v̔��L��ד��=c��*a�牛$k��"d�` R��Ŭ��Y��-G\�P�b\�.��7iJ�|)��L�S*�	2���qO ��gȇ k��]C�'/D���HM~�*-5���o��	��`ݎ�yb��4��ZV��)F	�e8f�@.[��=(Ӂˬ�~r�0nf��=ͧ�b�]�D@
Q�!VW�0��I12٬B�	IAF@��m�dH�І��[���%��/H@"BB�koL ��dNl|H���OA�D�N|؃�(.��z������ G
K�<y����Wz�7N�_��@hU��W8PP9��ƻu�0��%ɈD�����
�cD�Q!"�?J�r�� ��$� %q �!EU���9�49�O�Tk��;*�c��ތ\��|�1"O�h
VeC�Y�f٪`��."Y��Q$��'bP>��-O�l)'�QM��|Z3�����cT�d�A�%d�I&`�Y$"O(�g\�L˒��3D	9;8����B  |�$�� �T��?�	7nS�e��g?Y��î��Qr��b��t���y�<�ԇJC��J�ݺ7��u��;O��O�}���z�g�ɾ*$���CޣO�9��E�'��C�	Jt�P4j�0a:\� ��:��p�׉F����'^��S��Ą,�2tuw?5�Ǔ���pE�pv��,��JR��ꥯ��l��܅ȓEex��˪|��!�"�ڨi4ħO��{�œ�W�$|�ç0�x0��R�g6<����˱I|�чȓ,3��(��3o�n@R��.&�͛B��M�d�"VTT���L>�`��y�x��R��"	Vj<�!��x(<!1�ο��ma�e�
4���Q�/k���kZ�U^��$]=.�z�Cŉ��UZz��eč*S��x���&�BA��
Q~��?�7A�?|2^R�j�!��:�D���ӑZ$<��N�9��#�B``nI|qx��� �PR�D�(x�2�¦�˗"O���釧^#��(�/�O)�(���H��O+�<����x�.�zhXk���u������؋��xr ʶ"�����eU�?�ZAP�
�>"�d;2+	O؟tҳ��kx��H���-�g≷;�����H�3�ɪ�"5������y�Gϻ0���z�� +�(uB��<xP��'��#��I+dE#�����<g��yCn��l9�P�V��<��>�u+�����ْ�̻HRH�E��Y�S.$}�ux�
�V�|�p	-��B�I��,��.��P7J�H4��$���HH�9Ꜥs��A��b��.�'��D�?/����:`� �8���� �'�ڤ�7H(u�4�R�E]�~�R�"��M�}� ��S�FU���Ʉ/W��"?Y��S�Sئ]3!��e�x�S�e����w!X/�ֈ���-K#^���M	�[�>$�c���"��e@ ��9ٞ���I2[v��D�{HT��5��^ ��2��H,8������#���{��,��k�p�ɷ-Խ8�aA���!�d�8=����s�IK�)c�kB�,#���Sʈ�?��8����7�&�Bb�8<����c��J�-�s���
)]r"�*7`��,���
��& !�D�d�N!K����U�`F"�!a6��1��n�!H��X��O^	@����1���z�GQi�6u �D H��l��'�!as��)&^B�ϓ'�(��c@29mi�VFéhu\�K"�� ���P7jb8��&'�x���$A�^�db�`�,��!ۄ�
?)߱O4)��xc>7M��jԲ``DZGfu�!� %Q��+����6R���V�0?�C!���8fY� /6� �_�>6��1O���"��M�g�V�.���L�Px��'�y��K�?ϊ̪WL�
@2���<�y�A�v-UbG�ۣ��(��E���{�b�'p��°�˱I�\ˏ�4٧B)����䜚G�^84R�ɧ�&�����b�V�~��!Gk���ѩ��.n���)O�p��(q/М"D��A�N�'&���'��Eީ�I�<@|���0�l�P��L�
�!���d��Q�-�%{3!�=0���A钲������r����H9Q�v3Sq�@yTJ+?1r�>`��P����YY�W�!���S6j�W��N�(f�8�
p?�<HuK�8�y��Q̊�pAA�i9��B��64�@�숌���Cήs�BU����/q�FQ��\0���@��<R:\�c�4�(����]5�ܚ7��~�.��1��q&���X�~^�7�r�Dp��bN$�2���+����aҶw���R�UH�ቐ���[��VH����l�+O�H�A�d�?F�8!��I'%9,�ɐ����b���<F���mˣ���.�m���5/��S�O��$�U� +Y6U���H)gu�����2ZJ��E3�f��h ���6Kk�6ȵm�.A��>�w��n�}�|�=aAM��q�0�a��M�5-��37bm��
��S�u?��HÒ>E���E4)D\S%�KUVL�1c�0δ �4T����	1J>��+и&���N*���p�@�I"i�?P�J�
��W"Β�ē9Zİah�b�R����J�R,��ɥJ.��b�N�剱P�@�����6$�4P��#�kS3#�qO�����ϖ�k�^)B�)�<e ��a�	Q����m�G�q�T\[���>o�(5�#�3!��DxG"O��ɂA�c�L�Jh��6_BaR1O�u �M���yK�"~ꑡ��������"c�!��YG�<����= EV�h�ɋ	_\6,�3(�t~�S��\P��|8�D�M3t�X�Ѩ �_���9�O��b#�ók�\��u���kd��/_��S+�$�Pxra�	Wb�q4��	r	j#�ē��O*� a
�0'�j�2���JQ�>I�d�K3toX��dV.�y"�X+u��aC_�\� ���N��yB��1�I�E�@@���*�`!���6+Z}�p(�.*H4C�	:m~�
��5(���$!�3y,�'Q���Bf/ay����a�'C�v3�I{�덹ư?9�h�058���7�R�CTL֕4�@T*W�#4�88&
ٳ_��h��<�4G/D���5�O0������C��P��*D������~��a��EK�|j�����)D� hu�Hz�\�1ǟ���1#qH%D�H�!	'V|�TE[�d�D�g D�� ��Q����9�A/L�;�"Oȹ�T@V�ei�P� )�-�2\ �"O\�8�+E�f��WΛ�aKEP"O�`H�g֓*)��L]3�.���"O�Az�i�%�8x��K��k����"O�T
�׺>`n�r*D"� ���"O��9�,�>t˖�2��Qsl@9v"OtslR4���P	0@`�]��"O�1����+�h�"1'�4�r���"OĽ�B��:)��@c��.x}L�	�"O�\���&H\����֕ZS��ib"OhUH0n?o�pM�5E6ld� "O �@�+�!%��(�k7'E֩�V"O"�A��
<UBHcJO��Q7"O�E��-�z�.���I;4"\%9�"O��E��.U�8�)҉ؑZ<Z�`1"O��hIZ�za�לj
�qp�"O m��厾5�, èJ?Q��p�"O�S�)Z�4V�5CT�J7�@��V"Ob1R��.Ş��p��V��Be"O>U˲��	E��]:���AǨ��b"O�Z�Βi[�=��C�Iˆ�:�"O�Dh��A� ���V��P�S"OB�&��'=o���E�h��9Ov@�f_?_D((0�@�~�\,���	�h����>w�� %R�)s.B�		$��^ԲP��$�HA�B�ɪb~j��$�#v��MM�w*�B䉪-M�dh��\�	�x���$v�C�	6+h�a��4k�P"�/+5�C�ɉHO�!*�l�=�r�q"�,}��C�,'s����H_F�Qc�R�t�rC�ɾ`��2��B�z��w퓬��~���>%��)����!�̦Tct�!"JZ5��*]���hJ%f׽#�%������L���;�B|Aք+��)!g�$+�<�+	��dLĸ�)ؒrpa�$+�r��%�T�K�%���3�gA2C�%"�"M��PB˙�Cz ;çO�����$v�,�0Vɐ���Ԩȑ}qnIjwc���!�Q[>M!�hȨB���f9���$��"����1\�am$<�3��QM ��?qH~�hN�|:d�q�^�9dj�ZQÛ ��0������S�.�2���ӱa�Mµ��,�i[�哽q���4I�Ԕ��գm*�x�'�Z>���nC�����.����J0*��d�&DO�Z��Bi�����	��E2 �r���|x��*W�K�i�R4#R���$9_�(@˟�6-/�S�#��X�D�}8&��'a_X�1r�
EIv�ؗCB~�Q�  ��U��c�2j���рһ$V^� �x9�	��!��BF��ʉ���q�<�%×0��գ��(`��	/`ལW	G�Q����)�h}���	\�J�F��!��Q��y")R-mD�aT�->@r�����=��y�&
}�� 4#�\�H��֘�y2M�5N
�) R�N)"��d��
�y�ꂽqg�]���X2)�p@����;�y��U�\l��TC#�.E��d��yb�MC��BJI�h�.�;��%�yrLF�H�Ā81`�5��D#�	�y�d�k�T��E�'�Ȩ5�C��y���.���K��dq,�)cF@�ȓ|S� ���<*6%�r���]��a`���8�$�(��	uDĆ�O�(����%F�LE��'6_�^Ȅȓ�J!��"#}Q��BC�i��1�ȓS���W�8�F���O�Q��U��V�$!�7P� �P ���>La���b����(-��sda�6�u��<����� �,�P�덖{�BL�ȓ5P��:"^�И5�ƣ�!�����.{n�l�@"�;T�˵C�����S�? ʍ��e�3w����7��Kt� �"O +�bX�aS�T��mݿmOd�E"O��÷&C��h!`mT�~�&��"O��1��I�0eb����V�k�"O)	''�<=�Lj��@4}Riڄ"O�d�"�:R`B�����q 5�U"O�X���K���GX��2�"OCo�(�V$	�Dւ7V�T2�"O�e��+K$*P�A)�dJf"O<D��j�j(j��8I����"O ����++�8�qQAK�z�i�"Op���S4�� �(Q�v͒U"O�)����ʦ�3%��d݃w"O�)ڶK 9�a@P�N�J��6"O�]Ju΂��x���@��7��TX�"O��`��] a��� ��{��<�w"O�@�&�~�"!�t��|�����"ON�Q �g��˷��k'V(�"O8�i1��3�t�-^�z�D<�w"O�A��ʛ;M��d��1���D"OD����7��(�'��)4UB���"O4��K�;#ț�M��o��9:4a;D���%[�<i�mU0�c;D���
{���A�w�
1QsC9D�����ՙ.  �[�'߻%Y����7D��G�ܙ�@��3���t���#��2D�����\�ka�IQ'i�*ef����/D�I!l�K�(�1����=0~10� D�`0q�˩"�xUT��:_�N�S�?D��+���$m�s!�J1Ne0U!TN=D�h�d�۞(������/F�B�� �8D��)qNA/0ה�%�B�9Rը(D��
G� T91�n�0b�Ea$�(D�DR�FG�y*��r��]EbAJ��1D�dH��˽v6M�Gi�&4�2��.D�\��-D-B��5[��M�Z�MQw(0D�`��B�qۊ��c��f�Ҝ���/D���Um��	K ���P~��v�:D���HJ�f+�u��e¶
]�A�&9D�T�Q��*{ǐ\0$����a�1-6D����1_���S�����=ˁj3D��ʧC��n�98C�uz~uE2D�hR�%K��]a�
PF9�P&,D�T˧�² �p����:$ur�*+D��)t�d�ʱ�"��-�8�ǀ+D��q���Ҁ�K�Gԍ0�0�V�*D�,:�b�M��tq'#��$��q �n*D�Աj�t-���W��6^�!���'D�,En�2��`
lۢE+��%D��x��V�E�0I�mڕ[ے]h�+#D��
朳0J`�� UIb)�#D������(�K�.m Ԋ�!���:*�Թ��\'`�qq.Q�J(!�d	,x�T��@�MoPZ!k�;�!�����SQEJ-f>M���=~�!����`�$�3p�p!Q����!�Z��y2-S?S�R��� kX!�N�t�Q(֥�p��Ks�^d!��	�����'Ͷ<x���4�!��/m��bQ��#���WJ�!��UFl�{�D�/w�0c`�ZT!��޻VCݓ��I>�2=J���z!��%��M�q#�U�~p��Z�P�!���i�d ��fR6r;&PH�5�!�� f�FK�\m@Ѫb��7?�)�6"O*���-:dlU�F �C�$�Q"Op��sE�<��!+��H�E.= q"O0���Sc�	�AG�5x�I2�"O���т�(8:H�4��%G��<!&"O<(Д���X8����A�=>�)�"O�%�W�ܭ|�Xy 0K�?mج}��"O�a[��	p�]�W(�6a�&��"Oh����o��I�`爲e���
�'�4)�a`�%	z`�q�hP�'y��K@(ɋ	�J܊�',�8rPh=r���p�-4hl��'�����@�Y]���GD�9	���'�=���
?��"0&���A+�'n�!c'F�y���C���\�	�'n<�$�B#EgNXj�"O�~`�9	�'���p�9Q���1�R�u�|܈�')Ū���?b��=�pɊ�$耕�
�'�Jdct�J�C✘r�E\?$Rh8
�'b��' ��v��g�K,2e��`�'�y��EK�8�⨱� �>$pB�Y�'�"�� �:|�%�3����:5��'wd5�1���*�d�0�<͓
�'P*M�s�FE\�MK��/wZ�  �'k0	�u��$E��S�b�!n�.qz�'��Y�s�L��]ir끣����
�'�zp��/^y��U����5��N��yb,ɕer*�8p���7�ŋpaQ��yr`��XŐ5�Q#<@Ѧ���ybIɠ?�ʕ�r+����A[�ko�<��!ć,Xn�;5!���gL�J�<CG�<��*H����h��A�<�p�ɇv}�؋����8�WDe�<�2쇛Ip\zE拒��G�c�<�tj��d���*V��%c����k�]�<q5O�-̖"��<����Z�<ٲ��Wє�{p㍓FZ4�2.�q�<��N�����B!Ì]p�T��s�<qf	�'o/��0��L}`����u�<!���>	~M0DȎ�H�H$;�Dk�<ѓ�G���o�4c0��qf�<v�H�V9+ N�3U�-	t��j�<�s�R�j�`$�� �qRhZ�kDi�<Q"�S�Qе�B�SI�*���b�<��-P�`��C�N�[��i�y�<��OA':��L8񯂡xcBe�t�Nn�<�k�*u"��j��z�фnLk�<A�J�4���jf��9
l	Hv�e�<�q �.K� !��F=1�\��0�^b�<�s�m�D|�@P�S���*�_�<��R<t���i׉�6���'G�]�<Q�IG�H���/Y8�]���c�<)��YsD6d�4�\�*X"�
�Y�<9�"�	]��l�aA��7�:MJ��ZR�<�$�2�tT��)t��9Ь�P�<	fR�14T83t����Y���Bh�<!��ϡ5JX �O�0�8WI
c�<�q�X\�Q���L7J�!S�`z�<�6���3�\Aj�-�y�<a���&\�r@�W��P�"��$r�<!d�9~|��Ř< �e��dg�<��e�00��Z��^���E�g�<�b�q�BP*��O
A��4����a�<�$��!Ca�\�Ƅ;��q���E�<� ���cO�q\)8B�ʺw�|��"O֕�W!�XU�����<h{@�(U"OB�v
�/=���GJnfHm�A"O�����S�D(I򨛾?|�X�"O�Y"�,�P�⇂"LK���"O���-�M~�={�'K}�|�"O�,q�eΆB�����?� a�"O��hK�"9�,�j�opDT��38��ϰ �
�a�H>>����ȓ-��8{�@ P���H
�C��0��p�PtJ��X�M���[��
��ȓd(<�����!	�U�W�1}/ⵆ��8HzC�1�r�sOX�VA�x�ȓjʎ]�6�Χ��˴��+YvM�ȓc(F����"�����j_(n"P���zF`�٘"QN�:�b��Klm��ooF$se�m���U���b�ȓXtԩ��B�|���1R'�'O�D�ȓf��I+��#!�x8� �W�p��bV�<x��J4N�d�ɚr��`��a�E���F?�f�@V��s~|�ȓy����E��d�H���d�0�	�ȓS�ؼ���@�+�r���ݡga���ȓsf�7�M��M��(3u(��'բ���"�]�6P9�M�)�T�b�'���@,L]�![ �T0L?�,y
�'5��c�gT�~1���ԯ�r�l�	�'�H��$�(�:,��AR�n�*�S�'�J���Y��X����([
�'v\�I�R*|!qJ! �#��5p	�'�X}�vk�!4��u$�g��	�'�	!�T�cTf��Ŋ4!?��Y�'�J*�IʗJ��ɂ%����J��'�nxC�C�ht4<y0厶#�`�2�'�x�����w�JE�G,J��x�
�'�B���ҿP0��դ[�<'L��	�'�a� ��#^4���Q�֕4%ܭ��'��m�/V�D��ѡO�0|�9�'�`�)re5Oa�$�RK�(r#�'�`�C` YR�B�r��8�Ƅ{	�'s�-�.� I��3у�.d��{�'1`�e�Ǐ/k`��@ɔ�(Y���'����ҁ�X:ՠ�!'�~�k�'���FDʖ�Q���.f�k�'�Nxs�N*&��1� �?!;��'�0{�'=^V�5p�ꇮDb���'V،ـMթ2�����R=+Y��	�'���"Q���zXT�{���=.��0�	�'x&(�s�ڟ_8l9��ϰy�����'�*r$"�u����)�8��'����n	�i�p ��(&�]�'�Y�gjL $��%� '����'�b���^���1'քP\�h�'����  ���   �  Y  �  �  �)  M5  �@  �K  �V  8b  �m  
w  �~  �  H�  ��  �  '�  k�  ��  +�  ӻ  L�  ��  ��  9�  |�  ��  �  C�  ��  ��  ) � + l �  �) k1 �8  ? ?E +J  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���CO|EK�T�!�UjA�Q��Y�	'D�X����(�ت�H�H����g!|O�b�c�e]T���`�lY��!
��y"�ݔd�R®ɜQq�d���ɡ�y£-gnm8Vʙ	P,���U�W.�y��^�Vlh�'���U�F0U ȼ�y��-���h�bU�vI�����y�Q�lI�Vi	{*��Ӯ�8�y�,>%I#�gU�����A?�y�uDQ)��F�J_
b���<�y�'N�9��� D�ni(�+w$��yB��22��,���H(0x��s�]��y�� 	�1B�\u���Ò�yr�6(�4���\@�*a�W:߰?a�'�j�'ѱle&�S)A%
��Y�O�Ԅ�	�`��9Q�K�i���Q4!-7fB��  \6�i��@�L��,��Y�b��B�	�/)|G��:Wа��f	��B��.Bf=���ȂS�(H�g�/�B�	�Q��1j%��2Z��+"f��i��B�I?,�T�: 	Ҋ?/p܂�ON�"mrB��)�đ�N�6�ZAO�_e�C�I�k6���o��{���J}zC��'CGQ�F����T�V$ț�B�I� �X1�&i�FJ�����A(.�4� !���~J�D��]�!z� ��&|rwjN�<Aa��-6��%r�)�[�n��C�G���0=	�,]�ћa`��e~��.@�<qЀ �:�Q��W8�H�9t�B�	��a��g�O�Nز$���B�I#����`�O���H�f��pC�^0��6��? ^������.�ZC�|(n�kB�
=O�B���l�L{8C䉖;��A�6�]>� �uB�(�L�=�.�f�$��,N�tЃ��[0@W��ȓ02(0��h� ��g�I�IF���+]�T�Ge*`
$X���ҀL�޽���^İa�_�S�q���0\����� �1���I>��� "űq�D�=!��)��̤r���9�֖��Q�vJI�Q�!�Ƭ@�͑t�>�ʔ����Vў���)� ���p���ҷ�C�<:<2a"O��xC햭w���@��;��tr "O $��*E�gD|���-
<���)�"O�@��/ư!�"��6�߰A}�11c"O���ǋ�.�n�������{�"O�u��ΎA��@c��&q��H�"O�\���]�J����;=�  c�"O�!!_1	�yB�ŭp�bcV"O�͐��؋�ܪ�i��>R�h�"O����6f�]2��- ���"�"O�e�V �T+��C�֗�Z��"Oe(� [�I�.��5��D�>	�"O�}2��J`�؉%(��$ߞ0
P"O�!bT�Wi��ӳ���1 Mk�"O�S�M�T�RY*�[~���q�"O0]�
5%4�৮���\�2"OPi�J!lUBgN�9���г"O�P�'Wi�<՚��U�(l�P"OPhy������P��`���e"O�c�쌋S��c���~}���b"O�Y�a��W�!�CE�=	&Q��"O��Ki�1UX=ڃ�Q	| A�"O<�*��	g�vm�FC�m��u�7"O�p�4���-U�v��v�xs"O�D0�#V'��=H�cOV؈Bt"OV�ȴ�Y�k�Y�V�<]�0�U"O: ���^8 ���8'g�5V�c"O�)2U�u��`#�f�;&��U"O� �^�pYRl*��,{ʍ�U"OX+�bޡ�V��6�^�zw��j%"O��QCf���ka�0v"O��1�V�䃤�ߚ>���z$"O�I��v#Bx�j�<v䠖"O���6"��^����օ1�N���"O,�:�V��^�����a����"O��A�d/#W�� ����':�Ȇ"O����L0pZr����$��8�!"O�sE��0�01�ׁI�,X:���"Ot�Ib�>�X�a�@�\U���7"O� ;�H��Gp ��%��}�~;"OҼQ��&!o�(����/d �p0"O�A��L˕:������G�
�	�'�Z|ZMNˌ�AҤ{����	�'sZ�˱LOK).|�`�v	z���'�8ٳ��
��x�eʱnئ0r�'Ap�D�K<Y^����ŝa�`���'Z�}0өٮ�`(�E��-�	p
�'yt��T`_�>^*��DC@�N@	�'��tГ/Ҵ�,�C$ˆ!U����'P,��BIC�$"C��N��m�'�"4���/^���Ȃj}T�5��'�]����.°�K2��2u,�z�'��1�d���f�a�c��#U �c�'�e�s�+&�J�����f�`�'�
	�p�T�qb������2b��|b�'I|��a�У\�hA+!�&/�Z��' �hJ���i�!��,R�z[�'�fb�.3)HL@�ǂ�V]����'f����*����+ŐW�$���'˂�� �՗\f��
W$E�nF%1�'�TЗJ���Xq faP�M�(���'͆����pID�[�F��I���Q�'�v��[+4��yPE�@o,xK�'��0�kL�T.�(�M�`��u��� ����ӧj�P̉��1Y����V"O�`�����lN0�z�ϟ�Z�m�"O<:AY<Sn8����A�ua�"O�$c�VF����lكX'TX
�"O@dT�b�JT1��@	����'$�'��'��'���'��'*�d�V�L�Tn�p�]�V<[�'�2�'���'���'xR�'���'�^8�3�92�l�2��3D��͘��'?��'���'���'wR�'���'1�p�F̄1j� ��/(����u�'~"�'���'���'9r�'���'pp��A%��t裲�C�U�8�u�'+��'�b�'���'���'_��'%J��!���l��	Y���;���Z3�'�R�'3��'D��'���'���'�U�#�z7�Bt��؇�']��'(��'o�'�b�'�r�'	2�
�BA ��Q�+S��Ay��'�'�R�'�r�'mb�'�b�'L��`U�)-T���c�חlAЕ�U�'���'�B�'��'��'K��'�j�� ��~V����-���W�'O��'���'��'@��''��'A��8ң�9?��sg
�FH	��'��'�"�'r�'��'��'мjao�3i̜���T�-���R�'���'��'r��'��'��'県�`J�K�80���C�|��90�'���'���'t��'<b�cӐ�D�O6� ���B$����ׂ;"9���Iy�'
�)�3?���i�)	#�J2r��Hƈ@G*��2F��
����æ��?��<��sڄ:'��W��Ǐ�$SE�t2��?���Ŧ�M��O��S���K?��銾�hJ�ʔ�yH� T$3������'��>���qݮ���\T.UYbc1�M���u̓��O��6=���͍[4��j���cD�?i��yr^�b>�	Ѧ��h���X1@�(bY���C	A&/�&�̓�y��Od���4���� ykx4�2�B�h��M3C�Z�]��<N>Y�iT���y���#Z`J�C��R_��C�HL,\�O���' B�'J�d�>I7n���E2V	_"Q��y�Si�Z~��'�ba)C����O�`e��!��b�|�����n����(b�Y�,��{yr�������D�<�����V���Q�P�j%�$�����??շi��O�\.T��U"rϛ|�+�=#�$�Op�d�O~"��y�Z���T��R
���$���i1߹B�<xz�$T����4��D�O���O����r�m�@��.-״A���`I�ʓD��&�T�H�2�'�r���'ݸ5����&T�6��%��*1Έ���>)��?�I>�|�RF��I�j|�W�B�{�Zq�)ܹH`|,�~��'? �: I͟԰��|RP�D�փ�6h�c!G��8M���c��ß�����D�	���SPyr�k�X0��B�O@8��eJ�_�M�p	]?6���f/�O	nb�,��	⟰�Iʟ�jQbB�Y�����������P*\=��n�W~âp�X�D���w,��B�4$*�Y��bM|Bt�'���'��'r�'�}�D��߂l�񭝆A� ���O����O��l�B��'� 6m;�䄢Q� LZ�$�-s��ۍ�^�O����O�Η��7-=?1��Ҵs2����<7��A(���vLmk7C�O��{K>A/O���O��D�O���'ð]c�%(���S�,�a&�O���<�r�i�>4���'��'j���:9H�՘=1<HC�	 ���Yp�	���B�)r�ن>L`pk��J����6O0m���Ē���d"�ȟ,0@�|�+-�С�SH��ʈA|�2�'�"�'���D_�0��4CN�G �&zo4�[��π���$�.�?��+��ĐF}"�'�ιpSn�
A�	��&Ê�nQ(��'�"I� @�f���]
U��S���	�h?��:��!_�!c��9���oyB�'���'�b�'`�\>J�:=��~��a��d�L��aشN����?����䧉?�7��y�̊�(��b�z)�`�C��8jb�'Tɧ�O�r�!�iX�dԋ5��HYE Ң9E|	�B�	oZ�D��x %��*d
�O��?��e����r��2$q�x@�nĉ!�P͈���?���?�+O��nڃDU>��Iޟ���=e,���� WN��C��0�*��?�pQ���	���'��2��߉ld�X�#�</D�m�bH0?���C}�[۴՘O�0���?��$"9&5��I�>YDa��F��?i��?����?�����O�ql^�
�
yHU͐�Z'2\i���O��oZ�=��	�	ƟtAܴ���yׂ^<G��l�v*Z*f�����J�yr�''�.y�<ql�i~����{�0��=G��Ĳ�o˴2�����	�tF�X�c�|�Y���I����I�	���*�Y�����H���EV�Ky��w�bAx�l�OP���Ox����|�NMx�!'6/��[�kL�@f���'��'gɧ�O���2��C'�Mj&H�8v�	u�Ѕ0x>L9�O��*B!�?�rF0�d�<�
�m�*�d�]z ,҃h��?���?y���?ͧ��$�զ�q�`����ƙ�w62L �k�@T�D����"�4��'Q���?�)O�y!VO��u�N��_n����Je�ܴ����6\�q	�'{R������ ��(t��U�P�bj����['1O���O����O��D�O�?�!�/P"gd.ԉ���� �t+�^y��'6^<v��	�OJ�lD�Ʉo����j��N-�skߦ;�E$�,�����*��<l�c~"�8�dL�cI�Onl!��CYbA!�j�E?9I>Y-OL���O����O:��F�S�]��)1���ָt��O��$�<Q��iז5*�\�l��u���+z���5��~�!PFb�/��d@k}B�']�|ʟ�TQ��.@*��! �[�=HC�NMB�V�3�i>��!�' f $��1e�Y�^���!�) A藠�ҟ������i�l:��IyrDq�F࢒�:$4��;T���Bd0V`��X�͛V��q}��'��,xrŅSxvt��.W�(Y4h��'��"�ߛ����Bq�X���~R�I(e�r$q Ş�m�
���,��<I.O��D�O��D�On�$�O �'UV�i��	J���c%j�-���iL\�Y�d��B�'���w��L��Vm�I� �݇C
d���'N�|��$�B4R=�7O� ��$�'��t;� �Kܗ�y�Nhv����f��'w�I�\�ɣq��4P �A{14h���UyHr��Iҟ��ן �'L6m�%5��$�OR���Y;d�(�O�08)�$+�-À�t��Od�D�O��Ovu8�n,��<��a�KA�������yP�"3��oZ���'En���H$,vK�e��v�h�EI�џ|�	�l�I͟`D��'�di��&�/�4k�\h�'x7�M+=��˓ ���4鶴��Hŷu�NY8�GT)u+��=O����OT�D��_��7�4?YU�ۊ/6
�i�#r�i�4���Ԥa�D�/�H>I-O���O���O����O���0G�ԉscC[$7�D�r�<��iL�(��'X��'���y"fΰun�Jw���D`�w�M��꓃?����Şn�M"w
2[��aVI[�'"�BТ�:o���'M�����w�|�Q��!���&�h��ƔMh����ٟ���� �	ǟ�Uy��v�� �g��O��ꅂ��D��S�H&��)�<OPlZH�l�������� �5��
�q���v�(�Ǖ4�@El�i~R�
W�`Y�So�'ƿ�W��<V�����A4�,ġ�<i���?��?i���?Y��4Aj�b�Ю�a.����+%��'��e�p�h��?�0�4��1�p�#Fŀ�q2�t���+|�XK>���?ͧ4}���4��D�6��af�,<��I���58c���~��|r_�������쟜����qj��,9��i`�C���	`y$dӲ���*�O���O��'wg$��%��#P��c�X�Tj4�'p ��?q����S�D
QtXC��+���cl4}� ��:�旟�S:��D<��D�z�1�HVq|,3�S%�����O����O��	�<�бi�r��^8ܑN��x�=�_�9�� 럄�	��M��BǾ>q��zt0��i�b�P
<�"(����?A�뉋�M��OԄ#�ۺ��J?њ$A�`��i+��$su���Gu� �'��'�r�'�B�'d�S�W�ҥ/��#q/� V8�ܴ|�B�I�ª�?q��J�'�?1��?ͻK	XawEl�v�b�㐂A!�x����?�N>ͧ�?��%VL�ش�yB�I�[���S��-J���hF?�y�@ۻ<�8�������D�O����x�>��\�}��HӤ��>vvn�D�O���O��rC�&+F4b�'��� ��mJė,;�HM�` �%9��O�I�'*��_$:�D·K�u]�Y �h��4ܺ�{��"լ�&?�k��'Ь���^�
͊�m��w��=�b��	����؟l�IF�O>���p%*`ɝ(�~�Q��"N�R�r�|����O6��妱�?ͻ0xI7�W�f�H�/C<B��HΓ�?����?q���1�M��O���oQ.���"�.�7&@o���"g�SO�R�O���|����?���?y�h
We�:�rA抆�<0K(Oto�1P�v��	ß���B�ß<$Ϊ#�\4Cg�P�Y6D�"�!֧����OB�$5��Ɂ#=x}I�߫4���%'L�
�"�ߗa�h˓1M�D����O�!�O>�(O���g�\2{�
a�1��,{�P�PcG�O����O��D�O�I�<)�iz�ĸ#�'��i�Ef�$l����d�F9�#D�'�P7�-���OЌ�'���'���Z���@
�L(�H���IY����d���?Z�e�e-�?&?���:c� U��?5���B��<�r��ȟ��Iԟ��	���	E�':���M�"��!���n�6l����?I�(�F����'��7M*�d��$>9z�bD4C:��ҙ#�"�O����O󉗥i#`7M-?�`-�d��L��oԂ[��<0��&o�����	wy��'c�'��D�L��a�ŏ��&퐶G��B�'��I�Ms�&�?���?��'�r�ON̰�Bo�+ �\��ʐ�<��H���՟8�?�'�?�b���>�H�b���@���F	?6-�	�C�V)8k*O�����?�� �d��3���j�@�fZi#훫�����OH���O���	�<i��i���¥��y�� )��Y~��A.,Xr�'6M.���O��'0�I 3h�cW�B�q�Q҇AȘ,_�'�r0���i��i��bƂ�?y�U�� ��r�b��� ���hq�>O���?i���?���?������ȗ*��J��	9Y��u��HD�\���mZ�^��)�������R�S��������*Dt��x��� �N�V-@��?A����Ş
j���4�y�-�2^�;� X&Xdy 	G�y�Ũ3�y�	��'�	����	0� ��60�5�GAڨ.>��������ڟ �'�b7�B+�����O���̺g �
�c�SF,��k�(���LH�O �d"�I/-�XM��M�jJf�jp�R�6Ɔ�j��� �E�zm���O~b���O����@��A`������%G-& ����?����?����h��d�3Db���%��>S�*9���V����������S�\�Ɇ�M���w�p<�$Li�� Ci�k�ڡ�'��Q�td��!�'�� ���]�?)��,@Bbؕ'R�@F���/vX�'F�I֟��	ן�������	!�<̹�Ọ� usF��m��'�26�Y
�(ʓ�?qL~
�8����éh� ���-# D���6S�D�	̟ $�b>�	u%�6&��)�/z݀!Jd��w��Db�	+?I�H7��d��䓵�K�Ve	AE,O t�5�DN���ON�$�O*�4�˓m�VD5��ݍw���z��W.~�"A��� �y��nӔ�|�O����O<���W�6�Q)DQ���:<f�j�x�����tg��P�>9�ݸk�&�ӧbݕH�xQ���͂nbt�������⟼�I��<�IR��W��I2BާR��⥆K�E<�Y��?A�CF������$�'d7M1�DT�#/R���]e/�T0�B+&�@�O���O�M�a�6� ?��/��3��#1��K�� bΌ@AoW7<r�$D�	wy�'���'�2뛗|�����XT
*]��f�(Y���'��I��M�� >�?q��?i+�*)�S�5q$���I�,L�ZTsԙ���OZ���O8�O�S�N����g瑝_۪�Vh�1��l�5\ �l��4���B�'�'&aW����нZ3k��Qb��AG�'"��'�R���O��	�M�G�� o8�*�@��)��+���r&�.O��l�Y��)���Lj�͐�K�z�Zf&_�8:��3�ğx�I	%�$�n�z~�������L��S1,t��BA���R�B�((j��<A��?1��?a���?Q(���f�� I�J�RD͟"m{Ĺ�EG��5���ɟ��I��$%?��������<��L���B��\u�dbp�D�O>�O1��	k��kӖ�I�,.�Qs�.��]�p1�c�٨�|�I57�ұ�U�OD�OZ��|��,,Ʃ�SG�9�T��a�2�%(���?���?�)O�dm�8}�H]�I̟$���_��+���`]"�c�G�.m��'�������$�OD��<�ĝ�*I�E�6)E;/r�%�1�\0!��	�v�PaCA�ڦ�2M~
�����	�����1�޹�bT59������	��Ia�O��a\܂���<tH��D�H2q®m�F�H�΢<Q�i��O�N��)��T�#��d̔���Z*$���OH���O���l�B�2�~a���?Y1!(܂Dh>� d9+��@в��G��yy��'RR�'���'G���*B�Z�	�q���z �i���+�M#�L��?����?�L~�d�ҵ��V�aAn
�C��M�`Y�4��П&�b>�"�K�B[V�y$��g�~-2�O �@�)E�Jy�Ȝ>���Ac�'�
��83 _�n�
Wm�F`Ā�I��������i>��'��7-�.c:�$�Z^6�s ΍U�	����c��H����?��_����ɟ��ɳ#a�*JU1��p��	&`hL��f ���'�P��H�?��}b�;[! �����-���I�*�4Γ�?���?���?�����ObP��ad��g��xS各��٫c�'G��'oV7�?7t��OL�o�X�	(D�ZE>9�7�(����� �S�	�X�i>]����1�u��H�~�P�P�!��aѺ`�g�\������'�%���'nR�'��'������K	���C)���\�s�'1Q��2۴;������?�����[�;@�R��R5g�z����[������O��5��?a��>�b� �%�'m>��V&\��XfJ� Q���|j�L�O�@KK>��ҁN�)'їN�Zp��-���?����?q��?�|�-O Hn��K��$���1B�y�V�6����D#Ksy��t��㟬y�O|��J�5}�x�Ӯŋ �Ԭa�� !YM����O� ��g� �Ӻ�.G�2���<ի� V��=����7\L��`�<q-O���Or���O��D�O�ʧQΰE �!�::(t����j5(�$�i���S�'���'��O�B�g��ī������9B<�@�DA>q(J��>�)��t��tmZ�<�V$��kD�vj�dJN�� d��<���Fm�,�D����$�O��D�!I�X��nG���j�8���D�O@���O��F���-K�~�"�'����>�<�Ӈ�
	}%*�a�,Irn�O2�'���''�'�T�Z�@��-�2��p��	N\�	�Oe�C�Z�C4,6d�1��$�O����� 0��qv`@�
;����O
�d�O"���Oڢ}��=�2���`��}��	f_�ŉ�	1���81��'�<6"�i�5�bg��,3�Y"Sk��"i���c�j�������	dXbPl�n~���rs�T�g�? xt��M�g��� �f��;�'���<�'�?����?����?�6'� LXr��R�B<L�B9sڀ��I��M÷.�3�?����?�J~���3j����A���Ԫ���N�<y0V�t�I͟|&�b>ź�m]�[�x��P!DL�զ��B{�H�ŀ�uybDԍB����*��'��I�w��4���Ƥn��C4-�#A�0�I��8���H�i>�'�H7M���"��.���	y�ʵ���
]���V5�����O}R�'���'�|�wL_�/$�1 G��4}HόF��f�����%E����+���{���a�`��+I�	Hb1O��$�Od�$�O��D�O2�?9��ΎA}�(dH���k"��ҟ�����{ٴ	-R��'�?Y��i��'�x�bم�1��*.�a�@�|��'��O����i/�Ɂ|a^��  �E$��Pe��n�� �`�)a	��.�D�<���?9���?�d�-E�AǎvN��ac-=�?����D����
 ����	����O���c���>���Ƈ$?8�A�O�P�'�2�'4ɧ�Iʈ=�E�ǯ¿}�B����2g'����׈w���ל��S-���h�	�	����!Ým�"`��sn��IƟ��I؟��)�SPyb�g���0��W�|���?p�9x��O�x�t˓&�����}��'�derh�F9`�T]�:e'P��dG_�M�'�����!��?1�%[��"�f�Ja.�iы��:���x���'���'�r�'k��'u�S*�=D�iGn9iU�ŀe#�|�ٴW�x����?q���䧢?��yg��q_�k��׊KϾ�kM	R&��'�ɧ�OX����i��׽	lٰҢ��H���C���-�t���x?v�O���?���+�K��;Bd0t*ō=T�p����?���?�*O�ul��8v0(��֟��	!"�8 +�7��Q�$ ƾyi2�?Y�_�8�	l��>�&��m�l��Q��ȟ!����'�E�6	̟"fCT���I�ޟC��'Z|}��h�/tjsōO,�4�@��'�r�'�R�'�>u�I���h�7E���� Ӣ��;4���;�MsR�ۑ�?��z<���4��ڔ��>���I�_�x�6O��D�O`��ۇt274?�!��u��S�f�8��՞gj����!/!��&���'�R�'_b�'��'~V�$�Е
^`�SCFo>тU���ܴv>�}���?y����<��>q�t1��Fטlm˳�w3�Iퟴ��^�)�SB�$9sAk�*��9BC�cJ�Y��
+����'�A`F��ş��֞|"P�Y��;�� C����M��Z՟t������	���~y2l`Ӱբf��O.����X�´���e�<Z<���3��O2�oZt��d���������H;�"��XC!FJ�S�d ��$���l�P~�LHN݌���h�'�3��P���b���#���<)��?���?���?Q�����v�X)���P�?*:��0��	UB��'��!v���)�*�<��i�'
�Tx�A�E�0��e�$�|��'{�O�j r�i/��8;��q����j�j���k
��ࡡ\�7��4�d�<�'�?����?	������C3�ܔ~�]�׷�?�����Q��=`�/�ޟ �����O��90M�����ˤlH�h�N��OPt�'B��?e�j,r��Z��1�hق�`6��qa$����R��$���`KU�|���B�:H��,�@���$e³&M��'�b�'t��T[����4b��1(�C�ۘ�i�eŜOhD��U�X�?��+W�V��W}��'���A%S5I��c<���F�'\���>V���tɴO%q�V C�j�F�zuCF&�_�3>OD��?���?��?	����)�"�"5h%�0+���Ė�Lɾ!oZ6�ƕ�	�����{���������#k��^��E�J�`H�a�]��?A����Ş=��!�4�ybLѠw�LB��L I%��0f���y��4D������d�O���Jv��ebΟJv�-�6o׼A�����O����OL˓ ���#	�;��	���c��\P���N	I��iS� �x�a�	���IH�	#uj�����91ȪPZ����>�rb0U�@D=>;z��|.�J�䖭�?�る�2��ǡA�_�.��Do]��?���?1���?!����O|!�ă�'?�<�!堒3oء��@�OF�n��K�X�I����4���y�O�7M��9a���ʝ�����y��'f��'_��hP�i��ɿr�&Qi��O�4-�d���_z1`�̀��(	���R�IUy�OZ��'H2�'V2��u�>�5!�)h�n� ��Q���I��M#��T��?���?�H~Γx<��A�D?hy���NN�Vg�	qS�������&�b>�QSM%5+2��M f�@����=6��SFly"���sc����
��'`剰X����L:kĎ��|�x�����`����4�i>=�'�B7-ѽ9����?l�hH�D�@y���T�o��$]֦�?�!U� ��ɟH�	�?����*�;7>(�R �<�*��ڦ��'�@2����?��f����wL`����[��wm�vp��K�'���'�R�'WB�'��f��AŖ6I��Z`�K"3�����<���0��f����t�'7--���x�,1�Q�јl�6.��FN�O�$�O�)�R06??q��e�? �H'V�#���)gL^�H�iu��~�|�V��S��Iϟ�)w�	@<�\
@W.�n��3��П<�Imy¤jӮ�{�d�Ol���O��'C8.E1�E
��XQr��CVH�'�^��?1���S���g$.�q���2G��΍�N��y�Bir��i�P���xg�Q�	�l&�:��K�b��)�D�,Mh0����D�	ן$�)�Xyb�~�.Q��"��c��ꗀ	�r{���I�u+�H#���J}��'Ov��F��k~�m��
�9ͤ����'n�O�_s�������욚t_���<9�J�R��2�1E����uE��<�,O�$�OD�$�O����O6˧b�R�!�o 1w0mP�@Qm������i%4Q)��r��'���O��'`47=�ĥ�c��qzl!ĥVL���%@�O
����	�ʐl��<Y'(�L(>p��?TD��"'X�<Ʉ"E����T����$�Ol�䂗q�"��G��|�N�zwb�����OZ�D�O��=���L^r���'�֟L^P�Qgs�����=}�O���'|R�'��'5l8���Ԫ?�֙K�K�	@#���O*��LΜ,���[v�/�	L�?	v��Ojp�c'��JJ�,PfK�
9h� ��O|���O����O4�}��*�X���C�XG�<�V�N�(�t���UЛ� �'��'��7-5�i�m�&�� ���u	�Q6���g�X�	���ɸ"2ԨlZE~�o��mxB���r	���οRI��0eF��_L`�E�|RV���Ɵ@�IܟT�I��
����Ѓ�R�h�lu��hy��j��}3q+�OL�$�OR��H��_؝ A��O���r���,6�"��'<��'Fɧ�O����K�S�����7Z�Hj�jH%Ū�s�[�`Y���� �B�Q}��oyRd�&΢�b� �.\oT���3S|��'b�'��O��	�M���)�?��,92Y�픭GH�H4�K��?q��i��O���'2�'5d��F�p�N�R��頏-�Qb�i���>v<�P�۟В����y�f��2m��t&ְ�6 �	O �D�O��d�Oh���OL�d=�ӝ�v��T)���J&,T-���I����ɥ�M��F������̦u&��b�A�R�.3犨��钰D�B�O
���O�V?�z7�9?91Ĕ�2��IPAcX�${P��!5-~p���Ob��I>�+O�)�O����O�#��ܪ,W�	q��p�R��s��O��D�<��if2��V�'���'��S:,��xQ^�=���q��u�I埐�On�$�O.�O�ӂ��91�J�$���� (8q����UnZ��4��X�'��'�,��-�Z*(M0�M�ryXY3%�'��'����O�剧�M��˙=V�*x��@�
��x���&4Y��{-O�QnZf����	��C#X�LE���5��5'�`g��ԟ4�ɲ1�V�o�z~�(Sl�t�SK���$f��+��wu:�	�
�f��$�<����?y��?����?Y(�@�q�+6�ť�5"1(��dk��J�6-̻w�����Ot�d%�9O� lzޑ[fe������Y�d�"Q�PCٟ<�I|�)�Ӯ.��n��<I��պ؈	�7I�2T�*-��+[�<���� s�>���"����4�����{�u�Ǩ�2M^�� �YV���O��D�O4�{�f�&���'�Mξ@�|�QK�,L�!H�'�!"��OVi�'�R�'��'�m��cשw}�C�X�}�d���OZ��<!���@C��<�?C#�O��C�I�f��q�׵
y>M���O��D�OV���O�}�~���F��FtuRuh����S����ٴ*Dpr-OX-3��O��ۖM�J��3E���Y�Oŭ���O���O�%)��t���Ӻ���G-��T�)B�̻�(f�0A�k�o��O����O�*ጥsO��ԑ�SC�����4,'�����?Y����OR��x����W.����LL<}�4��!Ⱥ>q��?�L>�|zv��h�.6fK�w�j@1��B���i/��a��
 @���$��'%|��	4q�p�ӛ6�z	����.�7 !2�žP"�azk; �=S�%M�y��{�f㟼��Ob���OB�Y#��]$f��W��|�0ĭ/���3wnsӖ��
��v%��J~J�;Is�p5G�]�Z2��W�L|���?��[��h���#��́	��B��?i���?aQ�iyt<�͟��lZJ�	?2R,RD��Ȅa��ȮT�l�'������擭E
dnZS~�O����Gy�xpc+,�e�⓬}���������/�	}� @!lK���MRk['S�#<Y�it�@U�x��g�ԁN-Ab�bw(ǣl���B�����L}��'�2�|ʟN]�F��?�����R��4�Ǭ�E�z�D��}����|BU��O�3M>aԎ��`; �4Z[4��I�D<��i1��J�
րl�Hl�G1~
��۔�9$���'��6�!�I��$�O2i��BW�i�S��9��-Q�'�O*�d��F�6M5?��c���oyZA���6 ��z�Q�"X
�y_���I�j���OL�J7�	p�/��B��ߴkPČi.O���(�Ӣ�M�;1�`u���(B��R��?Ҫ���?�H>�|�%�K��M{��� �d��	תl�j���.��l4�E9Ot��I�8�?�f:�$�<�.O|	��ۮv�b�b�L��;�����'�.7-�+ZϬʓ�?��h��=ی�"��,H���K�FƷ��'����?!���`��he�!<f�h
@a�4 ^��'z�T�$E@j�@�R���T�ǟ�R�'u"�ᡦ�B�z|��a��R�'F6��#M�.p����!`���Y��'�7���K��F�4�L4P�����I��ݫ�C��yB�'\B�'��x�i��iݵ��A�?�Ȕ�1P�u)�Z�D����KU� �'��I@�'Xrt�E%�|�X�p�TF�d� �O��mڥT�Y�'Y�����N����T�j;�e �ɏ�m#�T�'g��'|ɧ�O�t`p񍙗QAD-�ELD�Mx��dY�]�QQ�P��9�IO�d~�EP�VynY8"�
�)C`P�I�p��&�̹�0>�E�i���1S�'U8k��ׄ]6�@�d�*i3bp�'�j7�&������O����O$�{�ȟ0:
����c�Թ�C���6m"?A�
�C��������ɿ�ժ�6���I�
 i��P��<i��fE.`$D)CKVE1�A���-B��?Q��:0���)���
Ц�%�����}��Y��Vΐ�ᐡ�[�ԟ�i>1��������'lv}A�#'-m�I�� 2s��4:I��'+p`������(�I�76��N_�TU�g*QW�"<��ia<�$�'���'��d��	���%( �2��#��U@�	�H��Q�)���=a�8�=y�z ��jř.���9��E��M�[���m(�d>��R�c��O3!ԼB�ËHQ!�dTᦱQ�.�<�	8���)[�  �	#w0\�'��6m!�I�����O��$� .H�%�slh@	���Of��əI�
6�&?�;H�-��'m��I���(�t���U�\fv����7|O��1dFL�E�����
ؕR*.�a3�Lצi�m�۟���\�:2��y�o�7,��4m�>>�� eR�:}r�'�ɧ�OVy�p�i\�d�!F�l��G QK^b fo�0V���:X:���'r�'���\y
�/uf&	��H'��]AbkW4�0<��iBN�y��'���'���G�ԚCF���/�MЅ� ��x}B�'Zҟ|��C�Jb�`�#�#@�"��'�]����G>g���Ju�\�$?e���O����)_�6���
d����(X3�j���O��D�O��d6�'�?!uo�4N����L?��E ��0�?aŸi�Z8*�W����4���y��
4g�D�Tn�/	c���yB�'�r�'�|� �i���	As�d���Oڜ��h�!2� ��@[|-QQ!�n��Ey�O���'R�'���[�#i����GN�yXr��%j��H%���MC�͂��?���?�K~Γ��H�%Mh�VYs&+�'BQ���[����۟0&�b>����1h𝒴�Q�'��:��'se�41!&:?�u�H���M4����ϱj�)���S�1�Tazp�f˸�d�O���O��4���\��Fie|B��g��<���c��4q���+�j�X�O*�ēW}��'\r�':\���!V#3�*�c�č�� ��v�
�K�����(@��7�t�Lg���ߙ�򇑹B����1�5��uSu/w���	�,�	�������� ̠yj����AN)S��sQ�v)����L����M�V��?���'�MCH>�B�l����1/�$jd��;b�����?9��|�c'���M��O�v�;1��YX���% w�MF�� $��M��yB��3 PX�r�+Q֡�V�q���0Z5ᄫQ��횑΂�A��8b���(*�q�qD� f��{7�>\��ia��"3�b�0i� @Ɵbi�3 Dp}2�ƻ^�ҡh0!�3`�	��fܯArl��5�݋c�[3w|��eF�R��͈��S4p��ӆ�&CZ<�tm8o� �j�N���߱{�1RM=c�n�@w�2_4&��j&[�̠��l�	b��S�ԧo�^�D�@�9�����F�%l5�Q�ކ�,MS�Sʆ,yÅ�"M��b�;�M����?����21@�+ḛ�& F�Gp =�r����'���'�����D�?��+?��)�@̈/�j��q�`�`�*x��i;B�'���Ok����� ̖\sfŖ�:})V`ަ���ҟ������%���}
fm��P����� �P���%¦���۟�M���?A�����_���'t@(�	�Z�QTkB�!\\��j�z���3�IO�'�?�FL����/�V�AՀ�1 -���'D��'Њi9�ȥ>	*O��d��0@Vz�6�y�kƔ*�<��e�@�Oƕ�W�J��������{�L�'���3���g�H�Jq�i��dU�\Jh����O�ʓ�?��>��@�!�	z]XL{v��&�
��'kީ��|��'8�'���$��\��Ųu�m�FȌEP�q�Jɇ��ĳ<���䓥?���.��U���-����K$z{$A�p*��?�+O��d�O���<a0�T�}��C<lY��11
�+�x��q&��l���]���G��ɟ�I�>��`�)H�� �^�d�h#�	Ǖox�'�"�'�[�0����)�O��R���%�W ��e�O�9�Ir��ߟ<���O����u��փ\p ��� D�|�� ���#����'��_��c3�A�����O����2�� �M�%H?��� B����1�xr�'3`�c�b�|2ҟf܀�äa X�0@S-c�8�@��i��	�e�h�!�4�?���?!�'S��i�E`3@�;"��@`_N�����v��d�O6�-wM�O��>]�a���La���/ �%����iӼЂ����!����`���?u��OʓS|
���h��C����%��,?��A`�iO�T���'b�'��p���#n��()��V�PF�9�qi	&�n�՟�����̀�a����<����~B�Ls��у�*�	���C�HA���'d��|�'S��'L̕��T;a������\�O��` &�o������C����'��	ϟ�%�֘��Q`�  �=���˘s��I��N>����?������3�¬�@(Z��z0�-��I�)Z�ҟ���b��RyZw� P�`�ʀT�>5�QQ���4�?q)O��D�O���<AH�u���ٸw4M�5#� +=.�0��[
}��	�X�Ii�Imy�O�⎖q:`�����Z�;�B�kw&��?A���?�+O(�{ƣ�K�Ӝ�\{ �1k�YB��9o��P�޴�?9K>�.O�	�O��O����Ҥ�)뜔!)X�n�����4�?q���d�> ̾p%>����?ט��x,s��v����C�Q��Of��?����<��X+�m0v�Nz�y�F��h�osyR� ��x�X�Ou��OȈ�� Y⒩\�r��E/Z��loZ`y��'��e;�)-��i��Q��� ��0
Gd҇T��h�4~�pyJ��?)��?!�'��?Qӂ�Hzv윞�F���E�����"|� �</"V񰦮��s'D頡��5E~��'���'����X����ɤ9"H��'�1'u���+�1��a���\�'�?��'��'�0K6�����%/����4�?����"��d�L����8��27�]�<���@�	Z��$����>?	��?�����d_�i�����TB}&�sdHÒB\8� b��|�	Ɵp�Iy�IFyZw��Zv�
�8�VD�'c�NX�ٴ�?iK>������O@���B�?��T�<� ��E��T8)�a�����O:�t�	Gy�f^�MS��Îp��y���!$�1 �l�s��Ο�'"g� =�S؟`�1���u�8��)�9��q��H��Mۏ�'��	�zB�Orl*F�N:b`P��EW��鶸i�bX��I+�4�O@2�'��\c6�� �ֳ/�͉��d����L<����߹vI��]�GE���Q�ؔR؊�b�E�*�f7��<	w�E;|	�fm�~"�������|�g�A�@� ��Ƥ!���~�N��?���@��O���M��"�}�48���R�W�@ER"�Ц�ѭX��M���?I����P���')�X��C�b�F��%(�<R0ֈ���g�,c�9O�O~�?��I	�L#v�C>4��A@Ϗ�]�05y�4�?���?� R�ZL�I~y2�'���0_�%rD��mH�գ��M���|"aN	�yʟ��d�O��׿o�9з؆P�N�X6��m�XmZ���sHѷ����<�����OklY�y��R d�C���T��"eݛ��'vN�1�'���'�R�'�Y����O�X��0��A�6N�	;��%b&����O���?�-O��d�O����f��:sDC6c9��ō�7V]�}F6O0���OZ�$�O��$�<!�K�\�I�V9D�!�َX� �E
�m\�FZ�@�	kyR�'"�'i���'�r�R��II�t�		v�,])�'v�����O��$�O�ʓ
�0���T?��i�ň��	�TP(��E)�Ę���iӰ�D�<!���?��,����ܴ9�L�8Ć���<�m��s�5l�����	\y�ʚ�qN\ꧽ?�����ƋI�>1���
ZV`;�՞1�����P��韸jS�l�@��y֟@0X`�ް%F�d�����fOJ��i
剦d���`ڴ�?��?Q�'`O�i�Q�3i�$(@T�*S'@_މ)�.h�$�$�OD�k<O��O�����i�7
Y��|�`�#�vѾm@7M�OH�d�O��i�h}�R�Pwg	~�&�10�R�<�{���!�MC�^�<�,O���$������J2r#���
C�B��@u�C��M[��?a�Hʢ}�Q���'���Ov<�e��[��@�b�I%F��e�s�i�b�' 2L��yʟ����O��ė9J�h�4���Q������"h�l�џ��Tȕ����<)�����Ok̟�a��Q�<������9��I�(�p�ߟ���ɟ���֟��'�L�!���M�*4����[��	�2��듕�D�O���?����?ɷ���$���牃�l��9Yѫ$� ��?����?����?�/Of��\�|��� ���IJ5`e@�#K��1�'32[�4�	�����0x����3�ʀ��؛�
y��#�vxڴ�?����?q�����בg�l�O�Zc�|� #V�~� ���0M�!!�4�?�/O��$�O�$ѭeB�$�O��I�R���Ϧn�J���aF� 7��Ox��<I!�v*��l�I�?QH1��y� ��w��%X%�C�A#���O.���OΜ���T�'��)�;�
�@��G�xH�]��_����*�?�MC���?���2S�֝�s9�1�:sM\ᡅ�s�:7�O�����h�$Zg��'Nq�F�i��[&.R}� _+,x�aKոi�4��ĎcӨ��OP���(|�'X�I�� ��C䕂s������3��lH��i}���'�Q�����D���Dc�*u�0�B+X��H��?��?���܁G��zy�'���p;�E��'V�����M��f�'���29"��)���?Q�p;�2��?x�H���5sjv�jw�iU��)�p���$�O���?���؄Q�g؀8|�1�4�ԗ"���'W����'��՟��	v�]"��!ã$Z�͹�m�=�N��p���<1���$�O:���O@�����7b��1��g�I`��˵��s|��O����O�$�|Γ{'xi��0��8�(�9~��L�P��,�D��ði��	ޟ(�'���'y��V	�y�J�v�b|��Σ0��qBB�ޠ��?����?�.O@TH�|�t�'�b �5���Z{�����W����m�D��<y���?�s!b}ϓ��O�u��-��I�:l[Aa�*h��l������Ay�K�u��'�?���ʷ$��e:j!�aėk�:٫Dȁ�l,�Iϟ\�	�, �io�Ԕ'��ݟ�mjv���]��K:nJ��������Z�mZ���	ϟ�S����5	�>{hL4I�Dtzd��i!r�'� ٰ�'����y��č+�$3�/�ݪ�FV/�M�F#�=���'���'i�$ȼ>�-OXAt�A'0���$TE���bI�̦��v�c����Ty��	�O������m�L�z�bG���a�&��ƦA�I���I�!��T¨OL��?1�'�8,�UK'(^�H0��.v ex�4��1���S���'9��'Jd�i'B�6'[��C�̂rw`UX�y�F�d]h	hT�'��⟜�'�Zcf�a�;4�,т��
�JLr�
�O(��:O6���O����O$�D�<a� �1�H(�o��X�i4�ܤ[-����^�8�'��X�<�	�\��V�Xh:�$�!jHxf��{�n-��`��	���I���	`y���9[#D�^6�]�e-4yھ��6�B/�,6ͧ<������O��D�O4P��5On`�3�Ͽ2�����:�X�@E}��'vR�'��I�i= ê�B��ϿmB�0���LVA��F؜
��o�ɟx�'���''RnU)�y�\�anҾRVl@ ��ڝ5Z��s �/�M���?�+O��:&i�i���'�b�O�J!6C-!� �)�)�D��D#��>���?���w��ϓ��9O&�S?$6p��+ܚ|G�$���N3�
7��<qu��-/t���'-��'�d�>�;<>��ٟ�8Yf��Zn��4�	�Lu\�ʟp�'�q��H��J�"@]G��,"���i/h]aQihӤ��O����� %�t���X^�1��H�u��BՃP:���۴�� �����S�Ou�
D4%��v�ԢO\z�� ӻ	�7��O��O�pr'!_{�IןP�	z?�[�`?��cN�%�`�9�B�Φi'��������'�?����?���c)ve�E�J2R�@P�G��	�v�'�\Aƅ#�	�4%��	 �zT��S�&=`% �.�"I��J������$�O���O��z8��A��k���p�I�EQ�m�N�bW�O*��:�D�O(���(��H:p�^?q�,���Bדm��ّd��O�˓�?���?�/OD)��n@�|����%A�f-��`�/J�\k���\����%��������(SٟT��"�S;D�ó�[1,%+Ղ���$�Ot��O��~}�%sW��d�T;[��"@�I#��PR�ؾ:p6M�O�O>�d�O���2O@�'2尵G]�&��5$���MY�4�?Y���
-���&>�I�?���KEw��|yr"��N���	�`�!�ē�?���~gD��������1Dd�h�pg�)ej�K���7�M3.O2�A���aB��<�$��^��'La�UC�?F($!�@t����ش�?��%X��������O�]�3A3�����ތn�5�ߴ4�LW�i�"�'L�O�b�@�#��#vw
�"���F�^�M���$�?	M>q����'�؅BF��~蘡�$��l�zղ6�fӠ�$�O��D7p�V�$����ğ��T����#ب�ҔS��ʕ��i�'�)��.%���OL���O�[ ΁�g,F�䪑� ���%o�Φ)�ɔ�^�	I<y��?!K>��: �-ٵJ	�r�܃��Hv�a�'� �|�'Y��'�剹3{4��d�R������,�h���@���'�B�|R�'���6'����2�_a&��+�.iv����'���I���'����w>�
�`�w&ik��V�Q��ʦ�>i��?�H>a���?	��<I0�P�h(��0-�Q��)���׿3��I͟��	����'�~}˱$3�	�	¤hy�fʃK�� �'��2:^�m�D�'�Iʟ`�Of\`���H���f�|�D��t�i��X���I�3g,8�I�l������'D�����}*�ӂ�Γ��I<�����:[��ݩEZ�I#�KR6�T�iD�g�7m�<A1m�<��'�~���
T��x�W��'��}�3K�qgZ�C�/y�H���O���P�	l�'y;�$z���n���z�Y�&��ش�v����?).O>�	�<�O~�1�PE��%��N*a)�H;A+�>aBS���O�r�P�%�\�3�+��W����V!��
md7�O~�d�O��iF�Rl��?)�'r����󞴫"�@,Htq�ۓ�?9���?�G�E�������8?�d���M�*[�6�'�,�z��'����d&��8� $b��W �XJg�P7wݞ���Iԟ��	🼗'�bxywnQ�X�f�2vn-U��L��C�wO$���O�O&���ODK�)ԃrw�]8E+�OS����K��1O����O�d�<Y�A�.]�i+ʆ hsGW%M"FiH�B4*��	ڟ���V�Iڟ��	�	3(�D�|��cn�  �����~^�t�'���'!b�'��Ē�hB�'S�I�2Ԋ��H%�E�0bZ,��F�'F�'YRP����=��c�*�����2�Ĵ1&�ē.z�6�'�P�x��ħ�y�'k�20�4g��X�1av��*'d���i��OB�(���?7�۫y�e��h���=��`)T!�&�'~Rn��'���'��I�?�����֘�� �ga@%4^T�ZG�ʵz6m�O.ʓe�P(DxJ|�W��9[�%��'s��������yp",USa}� ��i�$ȩ,תJ䶬�Ɗ��y���'i൰���-W6�k"@.cH�)2�]%��҅�F�0.�0���-}2��#��#K4F4��C$w`�rgoCS~�ɚR�ݵs�@�۔�Ԥ'�$����'I�����[�&���jFGV�i���ڻo�0 �P.3�N��do23����OPF� *ٻB��Ђ�_ A��'"�'���ԟl���|�@ą�6���/XaV6ŐWdئ!6\�-˶R��aucӗJEn�S����[-�����
_|~,ڶ���u~�d���T�(H�8��K9]k��� �=��O�IA�G��g�h�mڰ1a�H '�U�L\R�'�ў��?�t�>zfx��6-c�����d�<y����XGLA3 )q ��J���i̓���uy" ԫd���?Qw##O�\�8�%O*W|X�Bs�J��?q��'�����?��O��D1�H]�h�ː¦����fIh��ѻ�����E��1O i��	�(k��H"�L?�Eo]�1���	���yI@���a8�@b��O����<�ķM�hi1��޷c*@cQ�a̓��=�"�)��Qt��[�$d)EϗX<ձi 8�;�G��k T�뢋��t���'c�	-l�.�өO����|B�/�=�?I�o�Z/� ���9�h�c�D��?��� ~���H[6A t����]H*��˧T�)g(9@�@� k
�k�h�O � �[`��Q`ĬO9 ��#}��J�2d,�L��
��b�i���0��'(�>e��5�N�u�$0X��ҏZ��C�)D��C,h��'�����$Ga�'D��	�7V�\�p��i�l1{WD�>Q���?��nU(nr��?q��?ͻ@�pq!�Fe�JuR&䁪9�*]x�� ���!5�'�x�pn�����c;��(�:ݾ�[Ո��$� �AՅM/�٠�'݆���U�g�	r��0A�O�2j���CM8MԠ���O~򍇚�?ͧ�hOF�97L�1)��R] x'"Oz`[�B��7���)��b�L�u��L8���?��'��ʀ��|s��Ӵ�V4j"�p� ��4J��G�'�2�'��x���I��H�I�bf$���<{��I ��$j
�%�g��+Ϫ�i3�O
좁B^.�,�!g�Ɂv�� N�A����9/��p� R�\Taxb,�4l;t�6J��p9�x��(t�NШ��?с�i-�^� �	M��"p�Jp�E
�+�	(U^��Γ�xb�����,"2J�/Uތ�R.����*˛6�|�2˓k#H����i���'��k�h�HS4^�l�r-�џ���+w}4�	埜�'�b4A�+m��ţ�X�MEE��J����=l�X�a�I[8��S�/%ֶ(��m��l���")��L^(hµ��d��Sl ��D�2y���'L�	h;H�1 0r�Z)�d�܃fb�$���#8���S���L���$Z�d�(C�	��M÷�V�e~��b4�C��y��n��<1���08@��:�l���e��'N��C�ɫˎ��%�φ;�|a �	r֜C�I�>ܞP2VmȌ(7��Y���d�tC�I�RV��Ac\/�L���P/x�NC�	�H�|�zԫ[�V�@C�	�)q���g�@�)�n�s� _vC�I3�*@��,�>*D�K����NC�I�[�@��TK܇7T%��I�:@C�	�b|�����_fy���X�C�	'?�~5�ЍH:If8�s���.^�B�I�;��*�N��Gkvx��E0|W�B�I��±j"�կo�b��UI^.:��B�	6wA�T�V!G�N�śP�$��B��%AL!g�K��2|��o+:��C�	>!���`7��N9�dc��4��C�)� <�q�h��-�H@�c�56�<M�"Ob�@�,P��J���6�\�p"O���"�&����`��Z|PHW"O�����L�p���j;�蔈�"O>ظ�cÀ\�����@�q0"OT)��M5ht�2�A�_1$5��"O4�3ՌT$)�� �S���K��s�"O������O#&=��ǽ��U�s"O���%�
_&:�X�@��2�ҳ"O� 4Ɩ�԰�A�V�;ˈ��"O��ҋX�,N��kҁ?�0�i%"O��Y e�t_6Q��JJ$�<�86"O⸁S�A�JYx��gLO�$�e"Op��G'�9k0	�d�Er�{S"O��Ц�{���R%�%D> A D"O"q�'k�#	��Y�s��aӞ�{"OPiC@�N�[�n��0�,v�t��r"O�d8�F�$i,ȼ� �?d����"O��p7�RP���bJ�!i�RÁ"O���� �P��#G���b��"O��"	:�tR��T�]� T��"O��f�A1^O��`�ŕ!�ڱs""OV�sj�"�����Mz�Pj�"O��@
�E�Ph��S
P/��I$D�8�Fk�!R��	�i�o��q�g�&D��1Qj�3"()#��3HS�X��&%D�L��ļK�HX+B��$D{�l��'8Z=8�MI�?b��,Z��d��'j�}��%(8鋅
�5�
�"�'ژyÏO�o�̀u�U����'�t�`5��M��������F���' ��(�흪un8be� ��'�ڡ����j�D�':�`��.b��L��	i��dE�m&��BF�4�"��b�݉-��~�b
�ś�a5x�D*Є0�t��E)��?QփF3L����g "�y�(\| �-Rz��C��D�1���	s�����B�����(Z]��bbX�&�!���t)���@)�>9[����@�.D��NI��	%�H0y��S%C6��x���# ۮ�bA�[�JB��t���#��K��|3��\45J���?�?�O�5�~Ғ~�?�6��Njd�c޼�8�W�҄�p?�!���@xdÇ;`v� W�D�jE�"L�Ol�CvaF�ܰ>!!�]b�1eJ�,RBA���^��T�'��Pl)*���9����!�b�p�'��+aD�����H�Ez���
�'�(��D�)fz�1�<	6��������'R�>��BKYa��Sm������nB��u %	��O�C���Q,͟7�T�QUB� ,��9��(q�"�:Y|,�"HV�k|D$���|-�&@F�+�D%�]`���2�[H� #G!�T^6���]�N�[a��4#uHxc�䝑L��U&����l�c`ĩ���	����Hj���3eh�6o� $y��"O�ݪd��mOn ��#ڊd���l΍
=���⟬jD��)Kq��'�{��U�� �O�f�rXs	�'zy�Gru:-��|�${E��[���#S�Âx�(��C	?lOnqB��ȼN�;%F̼�=!��ɮcs93��8qsr�X����n���؁( �W�4Q6<�d�����O<uPq��h�O�P�9�.�di*��2
��H�0E��O�UHmu�`�Я
q?��ȦW& a��S+@����,��L�>��T
�4Ef��T4)��3��z"_�tq؜CAk��1�����Pyʤ����D��#���fW9]�hp#F�t�r��cf�d�\P��O�;��^+][����ʁ*��]
�E���бm�Ja�F|�_�Oi0��'\<D� -%+�h�B�Z0~bjD�@�Rk��P�
�&hd��#�V�O\<E��>	�O�W	�'f��!� P�2Ql���K4��'
�]Ɇ�T�O�<0� ����i[3P�Bո2#Zed\ �fڮ/&B�)]�s���|�	�4�.͋�T9Y�������i&l?���X#k�@H(أ��'K�������n�1E,t[�-�$}`�۳�p�>�y��@��YA��}na��'��Z���5$�`���<��㞰�燛36�h�)�ā-��|���O�#C��N@�d׷oQH��ዂR��o�?}���;���E��'01n��T!F�Ъ<���X:�,x ��-�b��I�r��t9`[�x2.!	�ʀ�U�
LK�(1�ȍ'@#B����;�Ш´`�#�\x6&Iʁ�Q%�$��h�J��CΠ[�G�RA^v�p�����?I)��8$d8�I�uh�{.�T x���GJ�3�4��R�i̓sZ4��V��Wa�`J��){�ds�fP�x�a6�G�T��5��L4e㞬�O����g��~���d�1W\�`��Wi�Ɓ!7?n��b!��w�n��j-6�\��u-�)�qO(��'N35�"�rh��<��6�'s�S(� F���Ǜ9�)�2+Wq2�	v`�_9<��2E��
�
Qp$�!�&u��_Q�j��d� %�| fcB7p������^*@��'3�5+SÙ'f�. ;�I�|ffL�0E�R�xa���s�E�gb�$)��4)Wˉ&)�O��8�/L�r��0��H�F��S 7d����S�hp8��"I�m4�1H��Wf@6�'��$H��.D�6�+�(��LU J7|r��	���>q����n\�cS�y�	דc�|����$!�pɳ�/�X�R���P�N�J�Asޮ�ON�H�I,3^���q"� Y�A��D��(l�i�B�Jp����&g]�O�x��I7�"����+U�0�)őx�KK�!i��t�X�e�:ء�G�8<�E�N�� ���X�a��x��F��V�����H�U�h��G�7x�DYe��{��UXч���ax"�E��l�0ODc4�T	d$E�14!�I�J&\��8ED�ă���:��٥�Ic#��Kk|�̻@��y��\��|C�D�	�~(�����.�R@�t �H ���0}��x��G3
1VM>y��WJ�Vj�$rlL�
���iܓY8U�pK-Bi�A3��$R��%�I�	��bL<I4��j�n(�A ](�~܂@��W?��E��J���I�h�4-�p�*���YŧD0(�%�"D#\Ovћ6���`��=Y�k?u�z|��4Ohy"�αQ3V�Q#��7y�vЙ2��$r"Hը6! � zڄ���Qi��ф�Im���`��Z�����=/��MN+{�F���E�F$�e�V���CK^;WF �3��@�B ��hK�T	S�܆&�L�#'퉎=�0���4�5B>�� E�'= +@��1 L>)D��&u�0)J�+I*,q���Pܓ#P8|(@�'j�Z��io��ϓ9�Dx��4�]39Ǡq����'�;p��u�H�e�܈(�08v��C�^!Xc'�T��t!�cT	4�d� 2�[�V� t�$�n�p�(���.R�v��fC��T .��ɨ:<�u���9[�&Us�G 2g&d͆�:H�q8e��L��-��ۙta��̓68�Ȁ'�K���K./z��p�)ʧ��g+	c�8T+�j������(pqCA&9\@��h
=����"W����y��t�B���Un�a���f2$30�ą�w8���G.`!�W8/ �r��K���ܸy��:�	� N��e�� �|2���� f�#r�u��?�(ONݑ���f����]�U@ƥW����6��hC�\{2����dߤ�!�$�<#=�ؖ���!$N��Ã
����qV�
�-��Fꄏ��Q�%"��H�7�
2>���&l�5<ưiQO� �y���=k��\�F`�i������� (ݱ���.��Y�2f_�����O���<A�HA�}�@����Ҏ9�Y��B�V8����*Eې$PT�Y@�L�i�,�P.|�I�%b���0�D�6M¡	�.%���*�$��<@t���ڰDyb��*����"�=dh�=Bp��U��S3S�H�"R���G��9��C�2	�zB�2�l��햝���� ݜ�Z6рix�f�'-e�1J3/њVJD�\ccĐ0nF�)�8��eޞ>�����'���bǭP��4�cW�)9�Uِ#J6\Jʓ1���Rm3�3�	�$$0	�p�2,J�|�pJ���!�=i�l@&N�QGD�`Q��c�!򤋽Urbux2��)�d����$E�!�Ȑ*NPe���P/�]Q"�)Q�!�$ރe[j��҆�9���
TJ!�D�?n90!�[}��%8@�VT��=��I7�э5�ɢ�^�a���ȓBhD�9p�_+�tL� �Ȳ}�����m�T��b��2|�Ir3H[�,��ȓ<Th����Ĝ�"kE�P�40��AC�@5�H�L���%��a��e��>ΩH�Q�t8�(Ч+��?L4؆�S�? z���J����[p�¹ 8>1��"ONxҲ�N�μ�P.�*1\��T"Oh|����_�d��5��?5 <��U"O��1��:e�RU�T�٢=>��!"O@<Q��:Uup,c'�C!(�����"O�d	hY�})&���N�����"Ouɶ�b��0A4^2-��d�"O�]�gԩaM��*��G7Hm�"Oꔘ�.[��=C�#�'S�luA�"OZ��L�?L%�)��%J}�<�'"O����L��=��a"� "[l&"OE��P�0�B�� ��ta�r""O�aX�L�;8�Δ����VWd��"O��heK �6q���<@U�h8T"O$���E]��%�Zi��]���\�y��DT�<Кs ��I�y�c��yr+����ذ'F�I=P���'�y���\�D8Q�X�R9�.޵�yb�R
^�pR`"֑F��� ���yr���H��jp�Ԉ>��]k�y��Z�'�����N�l���۷��5�yb�Y�1�p�a�ͨh�qJ��<�y��A	y�!�%S._$�1�g.�y"N,@���Q�[�f,�+��͢�yBH�9���)[\m� �b		�y��C�UǦ�ZT�V�_����1o���y"*�L|����"[ښ9(��Ɨ�y�$��E&�Q�M�X�:�k@$��y"��><�(
� EP�:�#@���ybH�_�����
P�5XW���y�,�dIb�ϔ��-
��yRJ؝@T�A��Bvѐ���y2lX�"�@��I��f��!���yR��e $����,L��<��*���y"�S�H����Q�8A�ȝ����y��S�,�u"�̆d�,��q`��yB%��K�8��D�Gd\50!J[2�y2���'��{��b��S��p��'Z���"-�PӃ(� �q��'~*q�䅆2D)p�l�,:|)�'���&�%��H�ˌ�_r��'s:�('��Iy�-B7��X����'�`zE��,e��#e��?��Ek�'|4ĪF G�*����82` ��'�`z�#�.^�u�_k<�
�'�I1(C	/��PG��jYx��
�'�X�KF!ڨjs%���K�
� �'-��qe�V*y�(H�c��%
�'brD��@�TD�@�a�b�Q�	�'��\)�
 E~��h0��|?vS�'��h�E�u^��kǊܷ'�8���'h���g#�b��A�'���b���'�L�K"�[�_���cb�� 9�4�
�'pRi�ξQ@���,AO��r
�'v\�ӧݒ>�t� ���62�D�
�'�0"�D�I�"#�O��c����
�'ɰ��ʃ���ذt�\*ad����''l�ȧ얇�
m
�I*�M�ʓHx��銿bX�p����\J��ȓb��mz�fM�AZ� Htg>i���ȓ36�r2��/&�H���N4@I�ȓ\[�h�u�9/���%hL���e��n��a� D�JQ|EႨӽ��Ćȓz+\��uB0L��1��=_:0���S�? ~�:d�"Z;�D	����5��"O,�IM$\0ƵAc�D���õ"O�Ԋ��X1�H:���3'����"O5�3*�p����t��9n�t=xA"O(*�@DL�6KTh�7I����"O0	-ܘ+�n�ѦF�'�,e�Q"O��C��?�(��`�8kh�9I"O�$aRXb�����o��rU"O*��ة5@�<����"s�4�V"O� !�D�l�����ͣadP�!�"O�H��ύA�]�D�5%7���Q"O���aR�0�0)@mոm%��c"O�M�7�Y	W����T�~,��"O\袇��.Wp&tIċ��a���b�"O���fA�pҼI�v�ծV���Z�"O�D�J��N�0�ʕ�J�8�xrb"O�H0�Q"-l��򭎳-�ܡ��"O�D���֟8|آ@�WK��ܐ"O�ݘf��"Z���o�� �u	'"O�`2%k�^x��%���T��"O��)ӊ�S�'pz ��"OD�(u�h�1+�^�(Z�7"O@��r�
8�������N�9��"O��	��ʴPoV�ӄ-A>+��"O�t��G�|@�$c�E �)
�"O�R� �Zܜ\��c,~��T"O���(�?c���_ ���!q"O:,DɃ8x:�z�k٭�p)��"O�k ���3�"��'�Ǒ{���1"O�� `OC�Tu �o�~�hb�"O�HS���\j�J��W�w��A"O����GٹZ��4��%�`�ja"O��*Z$�b,����G�f���"O��b��ǜ� �<O�x=��"O��������;�D�����e"O*�7��*$�@��nE�'�sb"O����O9G�:9s��1��k�"O*$00��1Th\��l6:E^eȇ"O|@5 y LQ0�I�A �Q��"O�@���oi&��P�T�F���"O�I�v��"f�����N���S�O���ȉl	�!R�f��`/f	����&�!�Ē�"#��*�'N?��1��F!�DX�[���`���	��W��?h>!�>w��P"��A�Fh}{6ꊶ6>!�d�@ ���g�ι_��� �
,o=!�DD�|�L��p�>��e��g�[.!�$β7�!�@���\c`u��2�1O��=�|��&G��c�	.G��d�$�]�<�C@�od�4�1"�{�jQzƠs�<���,��X�&��'3����Er�<i��Ε_ ��ig̝��B5
�b�g�<!%	��\n0�h�D��Y�fe�<���!k~�1R6��zF���c.e�<i���d�� B&]�H���:�n�V�<a!��#!�2����;D������T�<a5��I%z��5(ӳJy��1��l�<�4o]�$�r�b�wMf!bS�Fi�<فDq)��aF��0�d��@�<i0 ��FL�+e��0n��(�'@R�<a�*�-x�j`�p�+9������\t�<�e�P�S�`���ADP��%�p�<�'��>����, db:� 6��o�<9���$�R-��Pm�����"�m�<� �܉��͍a��}x�_�F��]4"O�u����/S5�D�$S�x��"O�1
`M�ga���@�)l�H)c�"O��P�Z��x�r �9w�hx�"O,�H�OQ�P!����F�A+��y��7lxL,8���V>�i���ڠ���U���OF
t�m��B���ȅ&I>yl
��'j	 �j� PHqT�
`��Q��'Cz�L�22:�BAA�-�����'��bˁ��,�#�o�4��5�
�'����"�T�4L[��; d��'���c�%�\��ؙ�Y�,�ȚL<i�'�ў�'!A�]�gJ,�<ȡV�\�SlY�ȓ L�Y:������3	z��ȓ;~��E��S�iaKCA��Ї�0!�"�Ý?���衧�I%F ��h�x���(ܡ]P^� q�\;Xr�Ň�q �Ȑ��@�R!B���}Q��ȓlE0�k�R|�9�mѳL�IDxb�'��Hi���3@��-��N���i�'6�����P����J;�Z|*�'	��P��F�v����3_߸q	�'���e���QEBC2g�H��	�'O�|A�F��B�VM����&���k�'3�l�uf�+L�Ҙ9t�P�R��9��'O�Zea(o�L�scV<K��|��'���X�ɇ�| $����=Y�Z�'�xJ KӒ07�J�B�V��\��'�B%�����+�懊S ��'},E��gS&�\a�A#�X�-
�'���!l��VxYq�[�{� 
�'��=R�b�������q�ȹQ
�'�r��(�06Ds��øm�
�'K������C�
��#[ވir�'��P��(�
>��!��I��\�
�'��@�e|���q��$;f@tx
�'NT})S�8Z��W��𶬄�; Ĭ���$4rtA��S�dmf��ȓZ/�)z�Ԫ+
���� �|<�ȓE�a�C��0~~l�bDQ�L����CB|X1�M��
�L`�ڋ.���ȓ����l��<hC&

_����f`��5�H6+���b,�c�
��ȓb�f))ѱ�aW':Yi҅qqD�f�<�����6��rD�1=	�ѢϚc�<u���H�z9S�&1Q�.�p#��`�<Y`F�O��`)�G[�'!��%U�<A4 �f����̒+sN�l�F� S�<)�L��1�D�+Y��Q�5I�M�<���.eNN�
FEռO���)hF�<���n��ES�E!uSd�IҢ�~�<�����T�@]�2�@SX�,�Q�<Y���RƘīݝG�M���x�<��&,;��i��K!Te$���}�<�j]�A<��� �p�7��C�<A��|+n��⓲C���"�Z�<����kPRô��+b�4d����m�<qQ%�*]�s#��k�ӱ��d�<�h��9���Is�8!bJ	��y�<9R��g{Lɘ�K�4#��|�mQ]�<�W��oRR�z�fγ�>R�Mr�<Q�P	ZfjH�3*md���c�r�<��C#���EDޫ&�E���v�<�F�L��\넯�-�>�)�`VG�<� ��J��-�F�1�� AkR�h&"OTh;�4�y���8��5�"O��K�Fǭf|2�Hb��&��h��"O�z0ʩY	�ِ���6~�B%��"O�h��%Ŧ�J�#J�fx	3"O���h@ ��t��
�O�2�"O�I�%j͜N<�aÑE2ba+6"Oh`��������pXV��$"O��d��\�FRИx�L-�"O�4R`
��DE3Q!H�&��SW"OH��ۺ+��(�F�n�����"O�q�PiJ�0v���@�ǩ�2�34"O�s'��/O�ez"�#d���z�"OZ��ƻ\,���W��V���ȶ"O�!����n�������a-h�q%"O4�s��29�"h���.(���V"O��+�A_�0����r�P&`)ĬP�"O6Q��-�k� ��PAU����%"O>T!G��<x���ϝ?[�P��"O6��"8j��C.��LM�\��"OH0�0�Ř��,�nv��R"OV,�t�ωw�)����R�*�@"O�]3VBZ<h����P��0��"OD@{5�EV̱�hY_���"O���fH��;Q$�@c%��W�h``"O������ie��8 b}�:Y�B"OTzrā�^W������>Mc $"O�=�b�։S�\�2o�bH��P�"OXY�"��EH�"D�4v<�"O2������^8��!�T2�p"O��Q/�6p
�i4�K9#p\��"O��4��zG��kD�d�8U"O��{_���4��D���@4ď��yr@K)�\�c̄S��!D�D�<!$���E
��:�h
#�\T���Tv�<����:�����]Khx�A�g�<i��U���C��,؃��c�<A"�� pht��۩����g�Ib�<�c�� [���
���%>�0T�@[�<!R�a�Υ~�b�zA)�Z��I�ȓ2�͑Sd��Ű��B#�<����*		�b�P�hA��h�*F�����n�I%�G��^���M�b����i0�����Y�i L�Emo��� ����!e�L~��c0��Z�͇���ъׂ�1Jm:mۅJGh,��<�.�ç�Z,q(�(��C�+�>��ȓ$�Cƪ]?|�p�� jyP��ȓ��X�ˌ��@|�1甤H$�=�ȓ_� R���wCP4��钥�i�<9%�O
\�A`cX:S_��q
�^�<�V��1?!q�k]�;���R�<i�dƱ�
�����Y�Ȓ@(�P�<�a�^�T����XV^��X��_A�<�윪.- A�t�ș���P���@�<�&L�c�¡�a(�5�����^}�<�b͈HA��b�� x���M�<YF��G�F��A�޴"�0�d�e�<�'+��i����MQ�����b�<���̉K�"��S8.��ynz�<i�� yWT��&�R27<���_�<��Ȟ$Xn��&ݣ�.qa@^�<��Bu[�yBT��Mn���r�<qi�|O��1C"qrX8��NE�<� ,����\$��(=Hbb��"On�k㨎�1`B��D4"qڅR "O���c 
�n��i�'Yb\�X%"O�`��Q������/E/\j"O�@{���#cQ��"��S�}��ik"O����*�"��������M�T�Z""O���@�ZH�ͪ`�nJ~5ȃ"ODL���� ��iX���RZ���"O�,��*J�<�d�iӧ�+@�y�&"O�@�FKM8z��M!X�+,
��"O�haŤ�wV��(t�)l� "O��y�MHF� c �7�"�H"O00���4���c􅂅0��G"Ot�c�.S/H�]J�$_�Y��)��"O�U�kG�L�t��\���	6"O(<�&�<'c�c`� �E���1v"O\$j�E3|UT�s��$j�	3�"O�14%�.R[��Pv�9@g�Ŋ�"OR�2��E6!���'��#��%�"O�� �Q��4K5� Aj� Є"On�����:������2
��	C"OTU�a�ؔ^�`m�@i�=2|z�qe"O:�xp,p��ͪ@ϡhg���u"O!Cc�2Q�T�C�GG�bx���A"O
X(%C>�.���F#��e"O,)��ߴIm��hׅF(�4x�"O$�`��S��~�(��H�D��p� "O6)�ciN��>9p�I��^v�$"O�4���ߍO4|h�IQ l����"OP�)w+_8��H���P
���'"On0��숚
�PlSFaRE�|:�"O8��6��!{%�� ��^�d���e"Ox��⣛��}+�OT�9���["O��D�
���T1�yͬe@C"OV9rFc�hPJ(�	U�z�4p�"O�DS6�/9�FY��Ew��	�"Or���h� ���QE�M(�+�"O	��eǕ3��Y"��z�>��u"OZ�P�&����qE����@q6"O`P�G[0Ye.����-	�� �"O�I�Cl��iiCI�?J�
"O�=����Cu
��'�
2�D�[�"Ox� �$Y�>nV��AΤ9[̬9�"O��Xs�يc
�ҎKA� zS"O ��E��g�zY#E��#!��� �"O��ҷ��!2��j�C˓ �r���"O������+w�*�	����m萹�Q"Oj̐��Ă[ ���.N���J�"O��R㫛�-��y)𩟛��m��"O������x�Tu��i��L��U"O|Q0�@^5l�rLQ�&�l�,Q�"O��9'�<E �)1f�s���Z�"O�5���*M�X�NO�W���ʃ"O8�z&���n�D��
'b^�QV"O�t��!�y��� 9|��0"O$�#uo�;(V@��ǉ*���"OT�Z�aݵRN���ک4�N�"Oz�g�ġe�0����Q�E���p�"Of�q!���^&�!��Gդ���"O�9�K�6-��| �/���Х"O�I��Q�L�b �ud� ��V"O��H��Ж d�J刃�B��Y��"O����A��4���ӡլ3�"�P�"O��#P�P4d�RuI@Ý|İ�s%"O� �h�h��p�-�o��l�x��"O���4�� bR��I|1���"Ody�'a��Q�h1S�(�	|���"OH�r�J�<;4��a�&�2Y����w"O�B�I�[�ʑ��%����C#"O��J�?e�"U�5$P(/�б�A"O���E��N�+���-&DՓ�"O8�Ê��_�Q���9,l��"O*$A��W�Yz�H�� �tJibU"O�x:��lF�z�΢�f�0�"O<E��( ��v8K��^7&�NHX`"O�!� �T�j���E�ܰez��JT"O��(Č_7H6�H�R��}\,�U"O<!)��S>���� �zDnժ�"O.cU� F����a(��(E"O�1SG��`J��1@�1<�����"O��J��
���ȚE"O`$ځ��LhQ	F�>|�e"O�1a���(@�.��цR?J� �!"O��֎)��S��>��E��"Ox�� 55c���1+G(��1"O6�ٵL�"��Iru(7B���'"Ov V(�
����H�'sm��bd"O��� a�f��q��#aj��A"O��R�hI�,�7��jH����"OTh� ��[XJ���&��}�LY	�"Of4*�ßKu"��$D��!�ڱ"O~�
%+_��y����>�J4�u"O���/U%K�P$h�a�
DӘh3a"O�@Pp�G�F�<\P�a�1#%���b"O����؟p�~	� K$����"O.T���_�3��9�#oW2oДYE"O��Dj�gG�Y���'#axM�"Oԍ M�^�1Pw��-np�|K�"O��q�+�[c�mc$L؎	>iD"O��*Ε�߮\
pMϠD.^�"O�xJ��W4b��!�Q#t,t��"O*PC�NG7EO�$0�*��v,"O�e��B�$#��p�JZe�<)�"O��0@-6�0�S��cE����"Oʙz�y3Z��b,�/+䦝�d"O�8�pC���`	�kI�m@��e"O�(�w�69$k�?R|d�"O����/ ����)͏�@(��"OV���M�p�E.�{��b"O���hT0�j�Ö��(E֮QC�"O&���ץi�D����I�J����"O��j#^(*�0S��l����u"O\؂��\$2>��"äR�?]�9"O���ȊnW�P0S��4�:���"O�1%��75IPF����q�<���3&
����,9���W,X�<��£*A��x�ɗ'~��d��`�W�<�O��rBVHb3�ߟe��T6�i�<��'<�Θ�"�X�41�©�g�<�s�0[�"��wE�R�|�����d�<y�D�z��9"���&kt-��+�`�<��:JĈ�q �����#c\�'�?���D&w�tۥ̠#����!�>D���@&Mx뢱��^{{�`j�=D��:6��{4萃!_�L����'�<D���W	IFH�� ��ȋ ܄e��'D��w�׼r�6� ®�0p(�3�$D��aìZ,Ľ� ��o/�$p�.D�� |�RႥ<��ա�停}o�\�5"O4��_�SnN �dE��yV ��C"O|��'�i�` ��jB%m:xa*W�'4�ɮ����Ǐ	�i4Ր&���w��C�I!h�*�z�IH�N�2iy��A�\O�C�I�o���¨���*��@�B�o�pC�I)O�� � �8^l�D��@���B�ɘa�(�s�V�2�\h≞� ��C�I�&R����\�[~�� p��"�C�I1� �C�i�+X�����Y��B��>��@����0���o��9(B��44�H���9<6��W��5"V"O����Nì,D:![P�æk���"O��1gI�+H �����r�A'"O�x�O��~���!e(�:D�����"O4�pd��{T��2�f=�~��d"O�h�aI���sU�������"O���5,ӏ@ɖ�p��Rb���"O�p�f M���8�j�  ���u"O蔹⇃�#u��O]5TK���"O0C�n�1Xxj��w P!H;L�(�"Oi1�D܊=U���w�X,Q,���IF�OҌ�Q$��?BF4�m�% `"	�'�(ە���¸�c!�hܻ�'�����*ʘ#��� s�(|�`I1�'% �`#S�q��<y�`֔xb����'V����],1:����X:T�y	�'�d�3"k�0Hox�� L��(��P�'A!���?5U��i��u ��b��d=�'Db��*W�pu�����3T꼰�����1���9_+�a8rAY*~�U��p����9:���ч����q�	V�����(�eFS }��8��C�[N>	��9D�DcgH�~a�E� �EN!Rf�8D��i,\��)֦xܠ����4D�l���]� ��U�6��yZ��1D���U7E2��p+\>H\9�Cf5�6�O������\C ��{��!�c"O���b�'�<Ȫ� "c� �:W"OF�􂄸Y��2U&�u��@�"O�!Ə�C���b;���iR�'c1O9��6�&Ac�"��VqX"O���s�Ȏu'Ĉh�c%Zd������D�O�TM�2��	��I�F݃*�r��	�'.jlA�I7j����#�J	�'�jكRK�m<������*�JP�'��T a�[�[��Qo��Qk�'�J��u�N�E�}��o>7�L+�'~%+�
�x��ɒk�A����'e�3W	-j�b�+r%��|�����'�,JA����;э�,z)�p��'�X`Qӈ�?m7����qi��
���y�s� Y���C
�����y����Ip1'L�J��KN��y2�+.
� �$k}�@@B$��>y���y©\3�|��1�n�F��6@���y����ݣr��4b$��Y��;�y2�J3uQ�cV@F�h�(\Z�G��?ɍ���/?��K &����H[/2�ډ��#�N�<���\����5��/�^�	tiIΟ�%�\�����IR���Wm��r���f�޻F
C�I�B"zl�Ģ}@�|��	�X2�B�	�wAsd
�$m����Ř�*%�����OB�$c���B�R�l_�y�p�Y��`��6+-D�� @�0���Q��:�CS�ju��"O���l�I؄�s�
ƫ���"Orl	`)̂L�*p{��[&�b�w"O����C�#V�%����
;����"O��aH� ��ň�0'VDx@"OX�B�9�J�x(��cZ�bS��'�	zy�5O|X��aZ��ܙjQ..=��"OT�!'ꈦ$��� g/V��vO:գ��]�:i� �L8� 0a�l�O|�`D��'i6q!@L�1��<�"ʓ�u(0�����?q�B�I�L�����"L��S��/0� B�I�\5��l�8F���9�-�
.��C䉽|���:!�Kc��0��#Mϴ˓��O"�D�On�	�Q�������PnԡI1�^�@�vC�I�&�jE��|��a���:�OУ=��y�cL>>���ʌk�Bq�NS/�yb�C;3�`�yGA�.^����L���y�N�&"TQ��䕇iZe�C���yb����a7�v9�4���.�y�S�H+�h G,�%@��j�$� �yR P�KL$P02�����D���y���4RX\A�� �T�Ð�	���4�O�B�鎅/���8"�ӈr�"��#"O�E2a �5'�&݂�M� @��['�'.ў"~2 ��?��!�fSQ�̐�)ƫ�y,�>}��x@�X%P&��h%i:��=y�y��+]����VK�!>olL����y�W��\ ���4q��{F�֢�yr@�72,0P�4-���2fP�y��I�4�\1�;2���S�D7�y"�]�@<3����!1��<�y�<=��L�!8�(])�J2�y�I��r0Q��C=&c&�+�C��y"���;"\Pcc��h�0F.�y2I��`!z��N;ž�P�ԁ�yI�!uNd�Z⁜���;��ɝ��O�#~�BhG��X�����lj��ۘFU�$:��?)�𤃁o#�t�DI�9��8��*j!򄙽\Z)⤨Z)+xE�w��o!�K�adtD%�٪}&&D����6I!��O�M�2d���I�9��Dk��ȃma�'�ўb>a2��2A�l�v	B�e �H[�X�<W#	�Qp��pP����<S� o�<W-w9 �!��э3��=x���b�<�b
��CZ�1��=�Ntqn�ܟh$����1W��e�0V�F �$O�egtB��+O�Lف��F5(�b��:g��=�	çHV��i�,�Ra����mh\�'�	F����`��;��� ^ Ta�M>D��B� L��dC&!-�>I�Fd<|O�b���U���q�|'��-$8�r$j8D���H��K�x$�g���/YD�`#D��BNJ�^Ց���.���B�"D��:���J1�l�S��3d�-���#D��!䇿h�н5��i��� =��0|�!�:d�h�{@,��y�i�l�<٤a�"o��<��5:b�p3��TA�<��T~S�(��N�8Ȉ��P@�<I���#G~�W����p�y�<�V�B�M��Cd�u<�nޏ�y͏�`Hd�rK�.~AZ6Ĝ3��<����-aI,��0`ʭ@h��a ,�g�џ E{��ُ �;�.�9h�EB�(\/5�!�ę�~昹+���z����ǔp��I�,�?E�� >%���=�\8��2��D��|b�)�-�d3�cPvL�5r�闰O4C�	��q���	�x�`����vgnB�*#pdS�
%J(2�YÄ��M�>��;��90��r�%���y%�ѯedC�	�q~rU��a]�S���EaJ�.C��>Am����׽˴4ȥM�'	�*C�'8�9��5���bA��.E�2B�I(f�E�̐�M������&:<��=�ÓxӼ�Ґ%�a�@hW[
Y/���r֩q&�͔Y��#נR�ȓ!��*�xt�=x�n�("q�e�'g��f�)�Ou��L��:"�,S��ئ[��X�D"Or��O�+Q�}*�D�,�E�"O�gk� k�t%R��]���z�y��'�M� �K�T��GMl��a�'�0�Y����_KbHR�hŶuP\K�'t)�@ʴ]�4a��a�@�`4��'���X	�Z���6S�P8,����������s"�D;	M.��
�E�Uǁ8{"�[�
�9u9��ȓ!�\(@W��En�J��̎O�F��������u������R�4���6��D	�̀P�(q�3�
2�����̮i��:D��-�1ʟ�3���ȓO7�Փ1�L�@��q��4H����E2�Y1�C�&#�}���O�����!H@�؀X�V���aB�����<I���=n~P2&#�h�C⏗N�<���]�;���CQ�X6F}���J�<a��X#%�$,ip� #7"�|[�mGI�<a�̍r ���!
�G�AC�WN�������$�(Ru�A#�0��Ts�H�:Bj��ȓMfe�ϵ?��x3�e�6K��`��QM��1���uFPY���
X����Iq�`r�4r���8u<�i2��S��8�ȓ"����g�?&6f`��Ϗ6�$�ȓ+�,�:FL�j�Z`�V �B���sO��7d؛��X!�i�r&��ȓs �xKT
Ě/ژG+=F���	c�xy��L�$��#�X���ȉ��!j�.9D�\ɥ ߞ?�4Qj��!:�n�{�/)D����m��j�(�C���t�x%�)D�XDƿY��
7B<rN�0��)D��2f�ĥ�qI_eb`���(D��{v
�hR����[#�� 0d:|O\�$�O@��@Ш5S�/�E��}+���C䉨?^x��D��du��M�a�vC�	wZybg��J�R	�0J�\E�C�	�	V�x�W#äa{�`�n�>��C�	���qS!W�O$��x��M.�C�ɗw�DQ�H/����E@�IڰC�ɏ ��)z@���8q��*��C䉵dw���@*�E���bD��;0O����1mbY�U�4�d|��W�HP&��.� �
a卧=�� [�n��x��ȓ`v�qʔ�ПD���ߑ,Xm��"Ob4���U�-�$��A�Q�dh$�80"O$�aQMW.<�|4z��[&T�06"OƬKf)#7.$����1<#R���"O��[���5�~��b��.ܬ��OLѐS/��#�A�A��%�<4�V`1D�p�.�]h�� ��¿6}
,Ȑ/D�4�!���F\eA��D� ��g$7D�� 6�*7I�;ϖ�ǋF�.p�Y�"O�`�f����:4-*j�B�"O�Y��R,5V$L	���.G��$B0"ON�����_�����dǉg����1�S��@�j��K�ǡGE�U	R���!�d�=i@���M�E;�e��^�4�!�dX'C�tQ�њ-v(3�(M-!�$��y:��9��f1���U.F�Q"!�$�#'��I3�E�v+6II���@7!�Ğb��hr�٢a��k�\K1!��&A��͈t$�%UQD��:�џ�F�ĭ�/p�(�ե͂x�P��֒�y�.\�,�Y�q#*e��NW��y�Ü�(�*,�1AUo�����O՟�y�*ū:�6�P�Ռg��QP��]��y�9#��f鍐r��M2��6S/!�d�*�ڶA;[�l���Q�P/!���0�������&q�h�"�噻((��)�n�4i��BߩT�̉��4�*	�'��t8��?Ul �{�K�4"�k�'��SjA#N��E!�iL"�.�X�'����cKO2����3�E��'���a��U�z��RB�2^�1@�'�^�g*��?��`KO�/1V:���'!�e�P�Є~�^E���;+�HA��'�$l)`�Ƙm�H�c�F�@��'���	�mB'?Pp�3�L/0��P�'��D+� 0G�40�M��|���'�~`0�>���S�h�-��<�'(�I�D�K3V\\�Y���xj24�
�'���� J "��d�J#x�J�����h�<P��)�+�N�\�suo�i�<��$N?'@q"���4���"O��c��\�#}�M�!�O&.<ȣ"ORTa�B�0#�u��0� �V"O�B��ƚYX��R�nŏ{�Rɉ�"OҰ2��p�|���L*k���j�"Ot$����c'�}H���3�2�0"O�)c���W�L3K���P"Oj ���0M�\�æa�<Q�"O���
92�jQГԜ+�z��E"O�Ɉ���
K}~�qďR�e�.��F"OVS���])d�YEn e���*�"O��@u��Cڄ��G� �v��1"OP�a������t�f¢\��"OL�E�:��hc��=���"O���C̑=�T���ܹO��\�"OHy�'�P�le�ir��ȞE���`"O6	X�,��1 Af@+zz��#�"Obу���I�����	
Svp�"O����H�p��A�s�Q�WȒ�"Ot�bJ^�,�d�[��R ��X�s"O>IR��B�ȃ���7�h��b�'����"�kõ/bJ�i��j��B䉝��U�a@�a��hi'�W
��C䉄KaJ\��i[0DE�����
#&�C䉁M�%�cE�6���+C*��NB�I�|�����]�h0�4$Ԧ`�C��<k�zŨ��5VQ�&ж:��C�	 �*��冩-��ı����	�B�	>HNT��!j���ҕ��8�B�	�$�� �N1q��8�0b�(Q��B䉸�Ь��@�8Ǝ4 �"��B�I��U��˕#�|<�%��5�B�)� ѹ��(dpЀ7)Y��3 "OH�����pt�1�H�J���"O�x��K *�=���@8&�T���|��'�pd�6��_�z����=b����'pHW�U�Ԩ�#�B:F솰��'*�!3`�X%MTLH��-<M�`��'���`�9�i"��Η-t�a2�'�ly����*����/�Y� �!
�'�HIxd됫%�T��#�Q��8H	�'�t��"ρ�56.<�5* 'Y�D���'���T��TĠj5%� ��1�'<�9�F���?����	�/��`Q�'LB�����F,Bi#r��2O2�)�'�HX�Q�Zd(8C�	ՊN�|	A�'�����0cL���S�Ȧ4r�'r���5@U�_��B��Gb�X�'�͚��F�7�\�Hp�߭L4JQ����?O�����a�z��A)\�!{�l�T"Oa�ԩ�xP��x�E�<Hi�3d"O~q��iW0��-�ŀ�egf�B%"O�Y`'G֟K�Lt��O�c��0"O&��E�ʞFv�P�Ta�(g9Z��@"O�LzÁ(8 88VA "s� �"O �8�`��<�V�Ǻ��
k����O�=��'7�PÆ��o�h������H�.�0H>y�'m~����� �� S�u���ȓ]xf��c�x&�)d��'
��ȓB����G�k�f��Y*J\�X�ȓ;L��C�)=��Z7A(&����c���C�	]A�Ց� ؤ�^���z$m�Q@,J`�=�!��\T��SL�eh�+]�Y9�	6j���b͆�E�Ⱥ�/Wӂ� d�Opj�ȓ2.�p�g���M�0@��S�8���`ߢp�E�0�`�{��E7�"�ȓz7��ɣI
"xS )���U0p�N5�ȓD��T�DG�jK�5rP�_+Qn�`�� ��᩵��(1I�����.�݅ȓ}v@�T�K�`���ɐ�Ǽ5�ȓ�B��㣎��q�kF�����ȓYH��

�X�� @�����ȓ~cVIp�H�a��(�1|����=@��Q��T4%,5��a��nՆd���|iI�W��h�!��MԄB�I9�t�H�&µ-�4`�@Y8�B�I�O�&1��]�5l�(����E��B䉺�R�b��Or�;�l��
4�B�ɮQ�|��+Q�v:�� f�N|B䉪iZ0��q(ͶiJ�!*��c�B䉫�81���'[n�`b��>)rB�	�A;�����E�I�V���B�Z�tB�I�HQ��Z��X����w��-y�B�I6�3���c��) ���"VF�B�I.jz=&DI�r�!A�Ř�,pB�	�
�\���ȓb(�!�2`�79JB䉙s�H�v�G�Cʊ-�V+v�8B�I4Q�P�GX��}R1Z�<}NC䉞�Č`o	\T]Z!S�m�BC�I
8�Դ���N�F}1G��?f��C�ɪr�T����!>�S�j9i���d)�
 ��%�F=����w,��Q�Du�ȓ��8qD� �P���֔P�֩�ȓN[8�����Cz�Ѫ��E,����49NDb��>��'�Hv6��S�? B�1tmZ��"`���4FJ��"O �{aӡIX�葮ǧT�6e""OJ4B�(�̽#d��[���"O�l��K�)'~�8L�d�Tx8"O<�w�Y#9��4��̢5�ִ)�"O(�؄a��$�$�����"O����+c���i) 5"���"OLd�e�>���8բäQ&q�4"OR5��!*��QLE/?���"O���#���[�P-�˝�y@���"O�9�@��9�,�����#'�=�"O�Q��:h�d (�*Y,ò���"O �!f㋂
0��5�Z�a��4�r"O$`R�4d��y#��:�(��"O�s���88r�XJ�@Ʊ9�d���"O��P��@+ ��ؙC���6l)`�"O���Ʌ�/�V��XN�t"Ojp�LR鼘8UN��fr���Oh��6���Qb�ڟ8����n!D���Tb�$w3���w�َo��� �1D��6G�6s_�Z�ח�`e�gK1D��pwk�5Y��	��$G�T=� 3D��p"�6!D�#�=l}�|`�&D��z�n`����b.eҨ�L$D���2�܅0�|U���%-�� �<D���G��-�P�w��y���;D�,�v� �`�d��sA�9[�8D��*�(B�gTi�&�N� ���puE6D�<
�k����Rڎ,�����.D��9�*ùQ���2BW PL��ڕ
.D�8�0fO�uM|����<k��:�&D��jd�	X7�X�� �:֌7D�D�s*G�g��8R /�N�H%-4D�L��L��:}�E�q�01;d�3D� !4 U;�A6���h����7�.D�h{���0jr�c�^�+d@���N8D�@4�XU� $��D.�$���7D��R&c�'Nl1Wb��gf
���� D���A�"r�Aa�
���b�?D��[��(j���I]�k���w�;D���BĄ<b\�A�G(pċQ%$D� ����7~"��tlJj\\!��!D��B�΀�w�����l_�\0HG� D�h	4ퟹe�b(���9r��8E#>D��2��E�P�"�F��:3��ջe�&D�lZ�AζaR�I���*�LA�w##D�����<V~@(r�tQ���T�"D�Dy`�X�4��Q	ûy���O"D�@����Pv�-A,�T�4ۢn?D�<aRZ6]l�3�Dv9��C�=D���� �(|��yW���>*d��K<D����̕����.���[��:@"Ojd���9t���x�0%�1"O^m9g��,��G�S�Y�r��"Oƍ��@�o�V@yċ�.7��"O���$	"V�H�d����9�!"OL�cԋP��6HK��[�3p����"O���؄~�<��#�/mJ��1"O��j6c�/+Z�(%L]5Ei�"O��V�!�Y��� k.��"O++;�n�Yg�K,�(���!�O�<Q�.�'Q��.pd��Q��K�<Q7�U�$�%��u$K�`�`�<rŏ�6+N3����/�$�rc�CQ�<� �}G&mY�
�d�..�X�;�"O�kcd��'1����[%_�J���"OF�s5�]�w����JN��NMI�"O��K��^��ex��!n|��7"O��A@F�S�N�;P�ë���7"O���WfU r&b�餤_�����?!�$
3���cZ�U��1��%W� !�$�f��4��Fh���re�&!���>0�ĂY%}��	�Q%LV!�,CT�17��l|�ӵ�APA!��<`D��r �ŔR�� J�=!�$H�>��I��H:=NxIC!�d��_ 08�b�m\� )� ��W-!�d�rZia3+Z kL�|'�>{"!�$B3@��Ԅ�^2v����@% !�����q�Hx-��
"�%f!�2_iH"W-�#i'J��0��;!�!�D�&*�u�a��:�Mr� �?!�$�X&��b�F����@@��
�'�\iCd�2GL�U)U%d�84r�'�P�a�X�z�(����cg�%��'��:1H�"}��J���/V�!��'�6��S�γ|'Vmu�=`�f�[�'����p˨,�܂��ݼ[sPh��'�6�aO�S���(DAѭMn0���'��ek��μs���83#�\b*��'e��6�ѽ�(�a3)�	[	<ER�'|�� ��]����b�]���m��'r3�C��Jp|��"�\8z$��'���%�0>L���Ӑ5�FH��'����LΆ6�^�H���<!P}Y�'������5���ɵc �c3��S�'��P  %��i�$��t,8Zq����'V�)��-L*��=��(S��셲�'8��jG�Z�22�BC�3�0e��'�����J�'jR9��`G$};� `�'Z�e2���4q|��w@�:{UT$[�'�T�WI�AcȠ�/C�D�0�
�'���fiāѮݰ�'X'<IB%��'�&x��J�y�8("���=~��<S�'�p�Ef����YV�Y�'��(D�@�?H��@��L0F
��'�`٤mËt?|�mZ?/��j�'�*�ku�"7��]k�AG,�p�Z�'��Ȑ�&Y�Y��d*%��"�n���'�h�k(��XA,�Aq�:%Z��'i��[�JE9r^>���)(vt��	�'۞9!SbE�@���8W���D9��'�6 ( ���8`��ږ��.����'�,��`�K+&�����̄[�'��yq�S�c��!����v�xA!�'�$@�D#*��-�Emχ!�Y"�'`i������z�+	��P��'��� � O,#���[DL8k��@�'?��(�k��Q����ۼ��%C	�'��D�aڊFkR�	����J�'ö͠���?��s�.\�d�̹
�'A@M�s
J`Y�4hU�i��'�0QO�,q��q�G��|���'�,�Pe�ЇTLp���*��#
�'����2e�(y���S�#�::
�'od5�"��q�<]sv�!�z���'G$|{ҡL1��������	��'ނ0���ߕ��} E.�_��8X��� Xm��aK����B�͐9��U�a"O�;b�5�L��f�J�+��1"Oj����W�.1�&��-ZT)�"O��H�b��]$:��C�\�OXQ�"O�eQg��F�qU��/nE��#"O��P�� ��X���&b �q�"O Mj�e��Q��3��/W�٫�"O���Q��<s�`��Ng�ճp"O$D�!*����3��>#[�̐b"O�bPf+H<��kB+S�,X �"O"�W�u�����@�A���6"OLu����$j�LG��0*q�2"O(�����)2��Gһ>�8�"O~�Ѥ��H�Nq �o��w� �"O��D�bɓ5⌽E��M��ᖇ�ybǟS��W!?e���1�y�j	$�f@8��X�	ɂi!p,]1�y2	�\X��K���t[��0�y"�>q>�y�f�O 5æ���yR��V�jIƍ
���P!
6�y�� �3��t��C�	�4(�0��"�yrAX5$�|Z�(�9r�<]A��ޙ�yR�ҵQ�p�i���qӀ)+T(Z��y�3Ղ`��ąb�����cP�y"�*d���oɗ]�.�C��9�y�+�r�������<V�ms2eՍ�y�&E�b��೗^�L�ʍ��6�y��:Z��$@���>'R�Z���y�G��x���+b[PQ�Gj^��yb玠V�2K �6S��\h�N��y̉�v��D���]G���r��V2�y�/1_�թ�f@4o�T)�� <�yr$�0Q�N����]�8�1�L�yR�V�^�"͊@��X@���j��y�C��)?<�+���5r�qC���y�+`V%{��yr��:����yro�(@���ʄ?x�����7�y��[6!>�×eUiwZt���"�yB�ǘVJx����"sØ��*���ybcp�)��͓�3X��fQ%�y&��W�h-�f�̜9���j�IT��y����	�\�s�&@�8k��zc@�yr'�L�K�ě�@�J]��f���y2�V�)��ʊ,�\�����y⤚5x��J�:ˌ�����yR�M�-uсg�ɝt���P����y��W?Knn�A����lF�ْ�-�y�N׬>8�%�ռR,�d9&NN��y"���D�X�4I�U�pQ����yB
�"���B3fW�Д!&Û�ybǉ�?��`)բ�=x�x!�h��yҥAv1���?�`)4д�y�'�#)�������R�(P�U]���e%<II�,]�	[t�'f[�O1�T��_��8 �'�#8*x����H"��q�������X�hM��@�HӼl,��e�B	�!���d~0{ҍ$f�]�ȓ7p��s�	!��pk�Du�XQD"O|EY�N��zNr��
��܏	!�D�"C�!�"��R:��r�C�:!�X�
՘T��	H!s��i����J�!�dJ@�(�q萨v�B4�צ��c�!��	�/2�`K�Dq
�I"&]Ar!�T�!_ld��o�}2��2$A,QT!�� ����� ��s�ҍ0Z6S5"OV��Gdޞ3�j0��Kɗ$4�tʇ"O�!�S�$D*�lR�@P�kh*�"O.���<:�� �DD���X�"O^t��ŝ<^��3��F��Xf"O�Da��`I�ȴ��5J	�I��"O��X�HʪT�ls$��7>�b�3"O�9 S!���R0d
3�l�"O"U���~�4$���@�
�YT"O���©G�b݈	��:�4=*"O�QwNͯΤ�hj��1��E�'"O\u����{ >̚Ab����(�"OPI�cV,#�>���*>�h""Ox��flڇJ��b���KM�eA"O�tA���n��Y�F�DL�ڦ"O��H��M���'\*��R�"Ob%�T�L8D���+p��@�"O�x�e�%3]�X!i�?xV���"O��"
W�26��j���$��Hf"O:Hk�BO�	��S��Z%!��"O�u2��.�$�C�ׂT'���"O���M�|(����9mb���"OR��5��~��Z���tP���"O��I�DO/��CA�3J�<`8U"O��*F �5�BY��E+Z5"O���?M��t��<H�q�`"O������{3F\@��Z�+ X�c�"O�qr��Q"�e�4LL�X� "O��#B�B�B���$�\��"O�S�	Z�p�)�4>��R�"O��4 ��w�K!E�F�;t"O^}�Ge��<$���eH�H���`q"O6l�Ř�����E���R�0X#A"O2�����S8D"���D!T#�"OD�0���5� �T��D��"OV���>}c����G�PN��w"O,a�"��>*����<
��T��"O �����4�VDx�kS���2P"O~]H& �x��I)�� 
]=T�R"Opx��#ʥhw�bՋ39�H�"O�вPl��%���	�H��F�̕��"OBd��	Y#5xti.��>-�1�"OE�g#=�xu�a0L'��2�"O� ����"�S�n��6��5"O&aj��:���y@��/S��2�"O,�3n��qJ �@L�a���b "Ohy�E�4G�(�AŦF�t5)6"O����@:#)r�	��A�}�V�"O���2��4jZ��%̓�8�@u�"O:)pAI�fl!�#W.��7/�!���U�:�9���4P�)��@O�!�dFv�Jq��i�9w����BNU!�Ӂ��A��[*��baZ=!�q�ve�D^:�����4#�!�Ȅd���Dv�\��k�,�!�ߓ�D����!n��T����e!�
�<���K'�;Ķ�
��@�!�d��|�ơH��[9G�,��6E�S�!�d)uj� qeځ?����#�j�!��	rH�3�R�F�� ��Ș�!�d�T��-�Do�]��c�k�<
�!�Dϙu��H2%^�����J��!��ë��hZ���
�^���h�Y!���r�`9:T �-V��
�J��/�!�� (<��ؘ ]�D��.ضK��]��"O�|��6�H�#]-�^iل"O�Yg����f< @Ȍ(��d"O��#�2~^�Q�H@;����"O�z�a�<P���֞*-��w"Odx[��І*�h�1F��E)�А�"O"���C?Z�B�┾ �`"O=�	�k�J�g��\��:�"OTd��T!Į�E�<yx([�"O�(ʴ])K	4���B�|���"O�Q���X+�,@K��9���"O��*�%�f�!��4Z���&"O�}�G�E�Q}LE��H�scz�;�"O��Qၻ�dh�w(U,G\��Z�"O���c��a˒��$���A��z�"O��{(W�cS Ef@-H.4uB@"OB��1�e?�%{ ��ww�0�"OJ9��$]9$�����ۼN�de9�"O�T&�-[ZTd:v瑱u��LQ�*O68��b#kDh*D+��Tg��	�'���UC�;�^�2"/��E�b	�'¼i�-�3Ġ��π�jZ�5��'�V�b׈�<B0i	'�iE|]A�'�}�5e��]qڑ�-H�-��H3�'PzA��O	0|v��E�
��T8�'��`�f���z2���Są���i��'��U�'��dH�(�wF=�
�'�f�Z�4S)s��~� l��'d8z�� z�La�bJ�"�Бz�'#@pp��"z�&a��!{���
�'���s懖�N-|� ψ-bF���'�X�]��V�xgA8c:���
�'��Ԑ��մ(�J�0�
EM��
�'�j��0C?�z��X==��q��'���cv�D�B��Sc���5YL�2�'����V�Y�w��ibF�3,�u��'�j$���?
3|�
��ߏ#ެm�
�'A�T��Aȝp���Y���(	�'�^|k��;f� ���� ���':�����@I(`9��*��
�'�*�� ���O:�Y�� ��q%��
�'MmaUfN�T���U%	-�T�	�'��Z3�
#(����|ڜ�	�'�����7i���������'9��!�NK�e��4��&Ư|rX��'B�K7	�(z����u!�-�h*�'�����	�H�a���-A�\��'$�h�ݦK�<�a�n���'(����f�2�D�zYH�����y��̫D�R@)4"�-9�@4�U@���y�,��%<&�����=8s|L#o�=�yB+��`�p=�AD�+����t(ܳ�y��η+��k�휉0|�4jG��yČ�7�����'����c�G��yBeh��r�e�\���0#	��y��ǔ7F���AS.Z��#��_��y2%P�?� (�eGY�uYrOI��yB�
-V�ԁ�g�0?FT�iT��y�B�G؜�avL�
OR�\��-�H�<)��-8Z��bD͉LJ%2W��L�<	  B&ˮ�h�Q�m����`!F�<�d�='��a�Y�h�䐩ŌF�<I�g�	`�`� ��M�h�"��E�<�ņAL�xA�ލVGX!���z�<� ]���,)'��&�ț}�����"O�!ö�K(h��sK'X���"OFe��͉e���2��j����S"O��b�(/�AZ�铳7� �*A"OⅪ�W,�d�1#	�	T�F`��"Opj�n&E��|)0.�k�\]
�"O�ȂkټO�>��qk_^���{�"O�ᩱ�Ą3��uː*�o�=�!"O�H�U�K"A>� �虣�L���"O��P�2���
��U�:e#� Nx�<A�I��
�q�'�͏!ti���v�<��.�"z%bdӰ%���@��u�<�@IM���RD�^�=���7��r�<����2hH��� �Q����LS�<!��Rr$�*�ǋ<�azDo	P�<�,J ��1he%U�fJ��!h�R�<�sLOWh�9� !K�3~x�!�I]g�<������^��@a�48� 3sg`�<��M��/�0�J�� s�N��q)�_�<A��~�v,��i���e:S��_�<	�%Z0V�{�Ϲf��a��[�<�WA	*��i�V�H5��Yӧ�<Y !%;�`y����^Hk-LA�<I5,��k� ���
'z1�b|�<q2�M1&��4�ڹOLP�Y��Dt�<yCL]��41�����?�zq�7�RV�<��]Z�D�3�N0�ኁ�V�<�D�\&{�uI��	
!��j���S�<#ża�Je�b�*6�X��PX�<1 H�lЁ�*���e[Q�<�d I�N�藺Y`&*�M�AZB�ɧ4]V 6,��/����|B�	�/=j�H��R"%Z� ���R*�B��d�T��%A�� Ѥ�:8M~B�#3}��!wC	,z�ʰ��Â�V@PB��?x��e�b	X�$ ��#J��$�lB�I�-$�1��I��aZ��B��8L\. �ǍP2���p��,:C�I�@|Y��ڮA�`�sG�M�NC�	�-B��k��M�7�d\�D�8ehJC�{����,7mFkB�W�0C�ɫ=J :@�� ~�h&9X�C�I+KY�dӴ�56ur�����0��⟀E{J?9�ô?�� �������H�O+D������Mq��8� �V��zE��_�'M�>�	0gi���N$I�0����@#�C�	P�N͓�2��)д(ڡX�f�I(ð?	�X/HsH�q��6Rd��@��^�<Q��C"�D`�	�.1}���l[�<�Ӌ�&b[:L11iϟ^���c��@�<��n�-9]N�ط�W�KWJP"2��|X���O�4hU�:~Ex�0���,��,b�=O��=E����*�t���Q�M?�������y��/N��h$.A�	��@�-]��'Mў�Oت��K�Z��	����`®DZ	�'�L'"�6b��Lhq*�
El�4����-O`8�1[&Xv($`1�х]�J���F^����"� �u�PQCãG�5ij��ʪ�y����\��4ENa�$	
wρ��'�ў���<��FS4��r�4$ X�c+Kj�'�1O8���jRi̢'��\ ��79�Z4qD"OF9�C.Hw3�!� �ӹ�j1�Q"O��s��TP4�f	��,��D/|O��WZ�w���v)̜FO���O 0m:� �Mq�OB"4 黐�P�o;�9��"O�����S�4	geE�7A��0��O���#;��EH$�=N1`�E⍸&�ax��)�5���b<bh���#�ɐM���ȓy\p�7��`�;f�[����';�"=E��o��3}f�8���o�f<��f��yb/��c ���*�t�5�⅜4�'�a{��Q�+ a�̅ o̩*���,�y�`�G4����,q{�:����'ў�'&@R� p ���d�ʵKP Ƌ�y�l������EC�
��P��(O �IP�'(p��R�Z���q6�O����R"OV��ԁ� �h��~Ѵ���T�F{��I	.A=�s��	 �yC�+K!E!�dWL_ā��hʾ���(BɁ�v�'qaxB��@��g��@q���22"�5{� |O���?)S	ug�h(�O�d�� �W�'2ў�'?��͚B��6��e�V_�:�t]�>��[��ҏ�	,_��Tbcb�|�U{Pl��4;�'�ў�>YB3*��j=�q��ę�j�BI��i&ʓ��<ya�ύP��%`��sJ�H�aT�<�T�7�O|=K�o
0�~�����6x6�!�"O�Z��r�X���Ή ,wލ�c"O��C��C>0l]:�OZ�Y�`U1���Y���IC8).`�S�O�����{!�$Ӌ.��e�%���f9&�!�dH��H���MO��I�g�K��f����b?�a���IT��*��{�вEE6e��z(�%�:�p{ (ѰEH��ȓ{ۦ�3��K�d;&��-m� �������O��}�,�à�D�A��%��p ���N7f���G�5�1�^$�f��<��'���T?9AgȄ�O�4���P's	��'�hO�a��=��X4E�>(�� ��j��hO�>�9ң�
�p|�!.�QaȄ�*?D��bP�N[x@ȴ��" �*G�;?��i��{ڤ8x�R6�60�0�2�߇q���hO���Wv��]�ވ8(śF����C3]F�D|2�%>(�ͳ�%�&�Ι���A�Z{&c���'�?�d�����c���Q	��Rŋ/D�ԙ���3w��a3�o�u��-{"L�ϐxR2{;8���0>�Ʌ/����O��1?�b?�"�D��4jPk�7Ql�7J'D�8I��ܿn����/ �V8�9$#d��'1O?90����W���`��0}�v�!D��IvG
O�E�UlD�iL����!D��csB�4(np�G�E�L�ʬ���<���?���@\��v�^�v�ʶ�έD�ў��ɸBN~mh��:!׾��-n|"=IO���� �YL�5�+�g�䛇��ȟԄ��k
"��5|+轁�V-��%lZ��8}���i�|�pc���#4�����'Y2�mHF����	
�z���jJ�(��[����'8 �X�Ԯn��6$mFT��
���DD�S�&ň3��#-�����N�"?qOZ��$�0K 
�B�6�Ғ-Ύ!�31�(Hp���T�*� VK�>a8�J?yۓ0��x�^�M��9qL�&T� �@�"�����'1�<�j��@���1NҫAC�ɼTh=�`�)yr�u���8<�C�7#a�l�6B8<j��Rѥ���B�ɺ|	v�D��Wb9h�03��t����P� ^ر��]��L�w,�59!�$�)b�F����S:D�D�C�[�i=!�� ԑT$�{7�u`$��IqT��	y�����R�1���3so���fH�#�!�N�.a7YN���t�8<���'*1O?��?@g���CC��qC2`�s�/M*!�?YY�e��\6���F�ִI�ָi���F}bD�^�A#@1v@�z!C��0?�*O|���n��,�8�9P�((r&��4"O�Q���=�^@:� خ;i�&"O�ˑ'
�0�&a('�r�!��"O~!1�ՌE���j2��"O�$�P�B�(H�����h���d"OƅK�iN��a�!鄢�N�;�"O�쫱��6�(��A"G �-;V"O@u{ud
&@|4" ���Z6��b"OLP�������U� 4[�p� "O��S���7`B�ATm��iD�QC"O����H�4BRb�P��/�>uA�"O�d{s,Q�A���2i�-UT���"O`�G 48݈��p��(C�&H �"O��z���"qPQC�Y�I���;3"O�u��Q\v��aC�V�^�%��"O8����"1Q�ڨYC�9 �"O��d�.R ����I��#!"O~%2'&޿Fl�����ʔiV�(�#"O�dұj�^�.��\5Yt��S"O�ՃU�F�6x������ZB��W"ORQ�O
vH�K���,Q,RQ�"O��;S�4���Iׂ�l ���"O����Ȉ/�|4���_�,�:x��"O>�ґ�ߌ&�X�4.�
x�L�	�'X4d��
�Xh�]�ƜxT����'E�c� ͡%Yʡ�5d�����	�'�ܽ�uV64�b�r�տ SLT �'�=;e)�M��qEIЯdЙ��'ʩJ�F+�����1"N�2�'��$���6�0Y�
��.�B�'l�L�"LE0&��k�� }��\��'���ٵf����f+��{o�H�',���	[�8��,�F�>{{�]	�'��ڂL�)���U��<�ؠ	�'��
��C>��C�E^��� 	�'~�%Z��BՊ ��v�@�<)�-G�1fF��ǲr8���lAy�<QE�/z�v��&ᐮ'*`�2 �s�<��l�`�N�u��"p�H"Ad�f�<Y��ŧ}�d���CӠ�,��N�e�<��*�tLT��f�K�	7�);�f�<��I��� I�4*���,�E�x�<�'�̟aJȕc&B��nlӄ�_q�<aC�~� P�*��g�(4H�a�<��g�2qN\���O�
,\ؚ�W�<���99 ��`�I	st:D��+Q�<�Ñ#a��HiD�y.�\2��TT�<q�ĥm�@xe�vI� �]M�<���¶zx�"��8j]�T�I�<��(���bHփ!j.��BC�<u��`��90��N�	/L��!j�Z�<���@6[e��R5��6
D8�P�^�<�cGX'(E�d��C�4M�\��uE`�<W%P�"B@����@-d��uu�T]�<���Y�T�\��B��C���(KV�<��,Yl��QP��&�>����T�<��b�"Rd��sd���w~�����N�<��-�-+�q�/��%>�-���GG�<� ���+Q�0Kб��
9|�Z�s"O0m��@Y� ⬄;d@ʟl1|���"O4�H��I�T�����N�`�;�"OF,��G.��PB�픕����'"O�����"�`mʃ�b�FA*�"O��s�h�1G�ȝs����ԁ!7"O��Q��8X@,��ǅ�p�b�A$"Oh�a&'U�f_X`PvFWJ�M�@"Or��M�/�I�q�%QrL �c"O&�� �T�`4�T����"OJ���S�Gx�*ab��p��1(�"Of)���2+م�ׄ<t���"O��:Q��������Sy��Z`�d�Tv��"�j*ڀ�)�jY��1O���MY��$1'GG�`ev|�&"O�<!1�܄X*е0��
Vi`tJ
�'� m�2*k��<93f�;5�����'��Er�
7qX`M7�K�/^�T�
�'�Z�z�A�m�^D� ��S
��X	�'tFt�ЎK�bn��37"�1��
�'w��r ��[8�a[� ��P�'���A�֟��0Cn���PmY�'�N�00i�:p�f*#&�.*�!��'�*x!�J��"x�X�0~Ա
�'W���BC9��3An[5
3�!�	�'h
�" �A��D�H6���,�z�'�@�4�	)]@,XV����^��'�hq�eBW�$h	[5*�?u��`	�'X�=��#s�$*Y�tDB@���y��]
j}ti�0��aZb	���y���"S?������7M����f^:�y�*�T���sDs��:�K���y�̠%\}���6&zJ<i��y"��j��r�
�$�qG��y��G�/�X���B")~~��p&��y�h�����{c��#R��
��y��'���]�28^��FȒ�\���'�>���4Z�~�j3Eކn�8P���Uå�h@%I!h�*>�U� ?D�P�/�=p�H	�R(�m�F�@#;D��"���61Qhtr��O��1��<D�x�/��KQ;���cr�:Bd!���UK,��I��4ؠ�@��/Zq!�$��sYH����?d�%:�!K�x!�$ �rU�w�$P���ߌ��| �'���a��^�@�^����ɥ��QH�'���E�9y|<}ڐQt ����'ᒙ���р-���$N�[��m@�'�m;�	��A�u�çG�Ih����'�8T��#�%4�(�pF�Er��'�a��i��`٠�AK��b
�'�PA� i״�-z�-ϟD�Z	�'���҅��p��sꌮ9��T��'>�"��D� �DA*2�2�Tl�
�'���C7��5�*e�B�͆?[ʰ��'�P݋��7TϞ"n�@��	�'g^�ҳ����٦�?G�>�ٴXx�5��;�Ot:�	� n�ЊuL� k�����'�f�dhZ<f�I;G������xxg"�$?��C�("S��Um?.v�eLڎN��c� �5�M�Ν2"�ӫ6���`܏e���5�L)�C�I�ZG����38�Q u�߹R��-��D� Z��r�ZUG��O�L����<Ø�q$��!&���@Q"O0a9��[�2��WJD(�$�DES ;R �%ɓ��p>�D-"�r�3��$aZQa3
M���� G�3���1��O� ����U�\$�@�Rc�[P��
4"O�iP�úY5 �i��x�����N�{��-�D Θ����:Ņ�~�Xi��
U��m�C_��G{���T�bΜ��Lo�>�T@��5�Z���&̨��	6%m�#|�'xY��$R7E� ��f۴.�`<�N>���''J�EMP�� [4�τ&,��f�DS�
�� Nq��T#��e��T��-P��ѓ�F	�V	��I�>m���j}�,�sUؼ���8�C�O׎��O�]E�E�!4�袆�Y P8 ���'��T��,*�	^?����%@�2/_%o�ެBP��<q�)ʧN}J�ba#v'�[�(�->�=A4�y�s�7�'CB<��Nӛ9�|���[�'��0&���ߓ�$�@�˒�X�00Ӏ�7.9�����F�*���O�u��,�����	9]������Q����7`�Y��B≨~���bHA�D����Rj��Z�hes& �>+��bTLω-��\��	�.r���Ћ"��홖c�a힘�K�vM��{l���և�$��K��}،s0�Û	z(��u�!s��X��'�2�H��C�4˔@I�o����&��6�*}ta�3M�l��jk�>�@��R�A�b?5*SdLd�j�a�ѕ?Q`%���6LOv��
+�PR�'�=�2��8X�@,�'J7 ����X1+�N�S��Fq�$Ò�ܸ��[B���V���H�������.Vu�<�-�+BU�e�;�'[@��y��]�֭�eF>Mh�az#ؒ4���1 hXr�����&63�%Y��i�$��ڴ��V>M�t��^ƒ��C��|�̙����H��E�>!u���|�K�WVr`�Vϙ�W�y��i��W�X��po׽J�x��☯I:�yS�-��tٻ��g�.K?�qsM~�<y4cC9}��(�r��8~]����ڳF68��')�+q@��W�����¹x���"�$r^c�M)��N�vLX��m�:SC�@'�q���B'�ߔ��?�b�s����R��8���2x�| sqg�p��xq�D�0z_��W�Ʊsp�7*KER��3{�h(#�Gt��Ddu��3uU�6�<�8`��0���Be�)�I0���ŧ>Q�Q>�+5��9��J6��z��跩��^LR��c@+b�`���
z�2E��D>��D�
@� �O�6ʧq����ݗ<LB<ң�Hc�!!g�lB��'�´s�O܆����bKbdc�i9#�(}�1�J���E+�bʳD�l\���������?Y$+F�>�B�� ���{�+;M�،���U�;��x��V�;�@��,��=X���
P�1ti�3+��L�ؔ˃�5�T��)r��X���W�U�z ���~�����6nu:���l���pcIڿ[���<}k� �-�}M�e(��)w�������D^�#����g��B��y���I%dI��ɛw���.00��e��G`���'�Dݱ���TB, *�k�cSD`#����y=�m!�C�W�f�"v�71-�u����֟ j�F�aP@d�Oa�`����	6��`D I�څǥ��<9�fSh�)!�I����$�W;:�Ah�Ֆg��]�H�f�v��`��~��'VB�$���y2�M;lpq�C�6�M�Wn�7��m,�A�O	lE̤I�mΠ��Om�i�Bלk�& H �ϝ<� �k�Y#pɩ�/���a}"����wN�z_��C������a�	�}���I�Mn(��O
�P�ˁ�v�0a.;B����"O��ې�ìzlP�"F\��5�͏��8���f)s`a|k3�\R��(:<�M����,��=���$M���[�`�˱� e9����&��	�ȓw/"����׳�X�K`Q�g>؆�d9�	�(5=|��'�z㮀�ȓĠu�7�*N�
U$�!7�̆ȓC4��eJ���DR�'�1�ȓ �,�B8K�P��a��<x��a��j5�qҀ(I>��ehȲ�8��ȓ<<��R��ym�4��T�b���hr���f�C\�����f���O�sQi��$�t5p	�'ugҐ��.�=l��@����{�`��'}8YSW�??b��8��1n�H9X����ĔH�������?*�t	R��%���L�8>��ҭ�<-��*�LS69@�D�Bb�2w��,
���A�:y�S�dy�hH/a�%�=�O$����1�ܴ�c�Փ]�0-�����,�h "S&�SGzEҬ����!<��)��ѣ���a��ˑߔ�1�/��s�D"h�5A�����X��#�<�7��P:tHV��?�L�' �h����|��MR�#:�!�C�Un�>�Z�j�Ɵ(�Cؓ:�P����'�ѳ3fV�m�D�T�:A�r��J��8fb��$8Z�)z܏V��Ot��#�W��7M(i$d ���h����sG��e�R��)l(t��F	ǫ8=��CM�bT�m
[��T�#������o�ܰ�����'T�e"�i�� &q��'C����p�49[r�t��,t�E��oBw��t��^?)��m�h�&i���ZZĐQ�VH��-�6�S>��I-���#�-�&~�OXLx�ʏ)���b��3=q*��T�p�vK����ؑ �S�s��b!��	4�Ӏ�\l
p� 
t���aI�~�Z���'m9r�׺��=AW��2||�uH�/wҮ|�toR�v�t(#+O�U��R�M�A�ɟ�����}���z�B���"]´�d�ЏQ��m�%>��c��6KbB�RTHZh���k�@X'8�Pä�)E��	æő����2�@!�'�a�SO6J`�]�wlX�*8-��lP�G�^��T"Ov�"ΐ|�\�Cv��M�
�������>��IS#�)�C�_j��nWz��cM�y��h�C̸@!$��I<M`����&�!���{Kao�!:@��Cm��A��Ĉ�y���	���0��Xό�H��uRL��<Y���pXX��ao/�(�,�;���F�zipB�49J��ȓY(��&� D58��@[d�`,Lj��'���������8L֘�� o��]u �	R�"D���6��f����瞫$mx	7�A�nA��IVA_���>aШ�2�j����ǻL3uj�KD~؞�h�)F�OL�Ig�b9�H�1�~t*���:%�C�I37���k�^@ZD��`���hC�39d��蔃ɹ8�x� [�C��B䉡j�|�!H��Ahv�r���J8VB�I�۪�I )d}	���m�.B�)xz���t��-nࠠK˾<�
B�I%��a+�iUS�LK��(IH�C�*2<0�A��MQ��A���`f�B�	bi@AB�S�*T�9�n�61+�B䉪�nh�'�xR9Z�Q/3��B�'0�TU UF1�� �� ��a^C䉘O�0+bgӛ`9���g�RC�I��y23K��s$Ґ���"C�20��
Ec�|��$hu��<��B�	:�T��`/$!O� !��'{�B�I#Oy��6���(SF���B!��C䉔8�ظzFa�&b�NY#j�n��C��-v�����3J�,�c"QxXC�	�c�0A2��S7Uz�E�ǰ�`B䉟{�����W�,��'��m;�B䉉R?�8У'��8]�(fn��m$�B�	6��)��	�`���cҪ��B�	�"����0"&.ʾ��vg�DW�B�-~�����a��#��H`Q	��7�,B�I5h�v��w�!%��#�-l�B�	b&�y�%k��-��H�� 3E��C�ɖTTx<�sL��8�p�	A kB�C�I:R����{L���r��7�C��"}��=8��R�k������<sܦC�ɩ~�z|�&��4=L�gy�C��-�^���%ۂ"s����U�X@C�	�R�IJ"�W�@*�rr,F;q?�C䉵fELQGo�T;��r��%�C�I�j� 4F]�	��z�H�9lifC�	yx!A�o��Iٰ���PC䉕n����g��	���f�'Wk.C�	�n��h2�h̫��A�&�	%5zB䉋+>0aK�N�2��@�
G��B�Ɋ^#���د;���r���:C��5yV�=��@�=R���[ �;$B��-�١0��>]f0� ���Y�B�I0
��	V�`�b	�W��C�	�N|���A�g|��ua�{
�C�I,j�"�UC"R��򵩝�[Z:C�$N���k��e0�4�SCU�8p�B�	��Tt*�+>s���֍�xjB䉘=���!������*o%LB�)� �E�++! �)��ĺV>��Jq"OT����[�v��ɊPKɦfN�PK�"Ozቢ��1G��s+E�	�dh�`"O�Tp�@я /��JQ�OS]���"O��ڇ$�#k�v�@�&N_��"O�e@-ݳ'*����ԕJ;���"O�mBb�.�؈���X�G.�EAV"O�xJq/Y:O��8�n2wԱk'"O�A���$n�p:��,H��V"O`uX�o����hA�;���"O4��� 2�A�%ʜ0�\ղ'"O��@�� #��@J��O�T�zC"O�xjb�7\����@ �0P��"O^@y�E���u��@�ol�(9�"O�$ 1m�:e�"�`pN�D����"OԄ���p�=�SB��D0"O���#ҘA`�-R����^���"O��"�l�>�aoLḤz�"O�d�vg�[��M��
��Ȃq"O"���-&A:v�;SL� x��u"O�$�S��$� aC�K�L�$L
`"O6A��Y:N�9�E��V�����"O2)�,�k��b���\�a0"O*5�R!� ����f(բT'�q�"OԈ�A)���)#�	� ��U"Ov�а�\
t��T�υp�1C"O����RT}0�*���'Wm�u�"O�"��|��agi��(#:\c#"O���I�n��q��j�:*��p"O�����8r��� �.�	ehX�"O�%�ؕC���e'��+�J�"O�]@��ѴB�l��m��5�X��7"O�5�F@Cl��yT���d�"OJ a�X9�� ���h�u�W"O~q��R)jB�$��ԕ+�U�d"O 6��Q2�Q�Ƅ,�f�:�"O��kcFJ�|�Z��'��al굻�"O��q�Gǻ{���ū�(`l�@�"OddNM�&����pjߎ5�X���"O�D2vL�u0�A�����0f��j�"O�Ặ�_�vE�٪0g�IA̤�&"O�m��o�	�@��1� *O����E"O��9�iz�1�&�؞/j���"O����m�
I��S4��2m� �5"ON�B�O)0w�%jvn��"���3"OR|�f�Oaz�DM�M�(�"O8uK�@��-�а !Kݕ9����%"O�Bb�!kـ2 �K���t�d"O̐��ǹyhR�k��*1z<��"O �cU#!I:a�%��)Q��s"Ox4Ӄ�I���3%-hd�|3�"O���A�$n� �A$�H�mjDj�"O|(3A��1%W.�R#�њA�X��R"O����g������v�B�"O����~$����

���zc"O�`1f��V6 �Y R�XW"OP�e�N�g6m��Ϋi�9� "O�T0�b�d�������|	�"O�yt��#;찇���S�Fɋw"O�HUd�b�ԊՃ@}B�[g�i�.H��Lx� :�iC%_��P2�A8&����*\O��P��Έ>2��Zp����KC'�D�C�V�(}`Q��,�2*��*>.��`�C�o���<�@	�	l����#�J\|a.�� 8ک��ۄ/,⠆�S�?  -���o�LA�c�֤tX�Y�IS zq|H�N����(2�g~r%����{��.NHbuh���yr��,dȘ!��Lǽͺe�%�65��F�~ԇ�I4z�2��w�ʂ���H��V%8��ė�fK�u:�'��~��T#g@U ��ǌ��`�=�yBfV�p|��"�-�h�PCץȘ'�b�ː�֦Mcl=F�Tْ.>�mR`�T�&����3D������H�� �w�II��&"Z�Ę>��LD���$�*���cیX?�ȗE�7!�D�%d�z}!2jҘe�e8&D��6UjfL�!�,�Q�p�����$�+1a2�[s#�m� ��	�M���`��u}RjL�f#&)��/Áxy��[G�˰�y�Ų]�B�A�]�{��H������'�����k�OE���~���Q�[Ҫt�
�'IL�����RT�:�#)\=�]{�'7�p�n���T��.S�,Dh	�'ۦ]�T�H�D���үס��I�'H@�)M�$N������.�
�'����,A�xa�|�%��J	�'� �c�Ғ[+,,�U�ݦ���j�OҐ?�qOd=E��O��&�8&%�d�� ���"OX�B@�z�ؒ�D4E�]�d�%`�w��mX�h	�唘%t�	�E�ts����� LO����;:�����'Ovh�e,�Jϸ�x4�1إ Tf�<)��ݬ2��+DaH�5Ȗ�2Ԋ\̓4̚�bt��A�ڣ~j�fQ��fi�f�)4����aa�\��1Sjh!���B�8O�"ꁅ4�n5#�I#&�@�z FL�T��x��6}��L����ɧ5�x�p�F��� �A*RJ��lrc(�&q�$HP��D'��D�8¤I&��#)┹��:S𩸃�['b��(�428��`G*�~�Zcq��(W���S�W�ѳe�� |�x�R`Z�gs""<������%�7����	DM� H�-���'<5<�S5�B��$��Cua�����_�t,Y��R;W���6t2t�rr* >����Z�2b������_�"tc��.wN�zf�L����hĖ �t`g �+da���� Kz�RpY��JsH���M��Bp# �ȖU0���'&G3B1�dڰ�Ķ�dQM�4�䡣|�QlT=43�1��$�>AD�~jH�5�Ю���F�	A�� �W ԟ�ѩ[fh�$?��٧�ў�N1�D 
.�LLZV�}���jԐsO �زNŧc.��O��'	s�	(�A��=��EA�f��0�Cᦒ�<㣍]a|����Sl��x+O2��Ǩ��_F�0�R���L��A��|� �O((U��"t�	cV4�6Ƀ�Q1T��Sm��K�v�dQB 5:C�	 i���8W	5Zز	
�f>>״���ȏ�u9�H���[!SiJ���K�h����ɴXڱ�hL@��='�>@���/t��D�V�'�6X�rNP-p��L�'0@���(ՠ23�e�n�59��TG�8�V	�pi��)D'Rx�g�Y�9����WT��S7a�l�� %��Cg��o��4��S8jEZ;@���JI�腄Q�P�|�b핰U���DQIX����0Ƥ4B��K'�rMr7(�Y�'�Hbw�$�g~r�	|���Q�
�eZ�h�ڝ�y��@"zs�Q�*�/dh�qEP��,�G���0?��� �
���U�hi�Bp�<aQFA�q2�����[<ܐa\d�<�2 �A��P�3H*)zi��g�<1��w��E��)Tl���0��Y�<��IA��Ԩ�Ջь+��9�Hh�<�Ǣ�4��{�G"3p\�"7�2D��! oE�:Q)���D�&�p-D�ؒ0�ӈ�4u@W,C�%i�,��6D�XY��	) U���+�%G�l�7�0D�@c��dt�iq��'�
��c�.}�D�)L\�]>	��CS<�ق7L�/xY�j�o*D����쇠5_���P�ݓv��X�@���`y��].g�h�*���yRB8[����V�J�hU�ۄꀞ��?�t⑹X+��G#���<��6�Q�ONqb��0x3�0Ӈ�<A�ɑ9����'�4�R��ˊG�0�э�L��8Fˑ+!
����52�:��O.𩛃+Ҁx�4�(Ͻ�`a�B�;;�(�ǐ|��9Oj@�/"K�0h���I>��M:1[���Х�� ����-���%TO�1h�_>� ThZe��~T�FO�rN�X���'�lԑ���<e����	� ��M� 띒
O���Fř�%ٴ�h�(�%�~��7.��	�&�@ⓘmV��k�
��M�W��Ք��PGC9V�TQ�"N�y����'⋗;�a�RC�!�����f�n��ΐ�,;�8��OT$��k�&6 ?A�,��?{����
~ ��7-]�ocڸѹP����K}�e�Z�3�Nd����u���� Z�� ��	�
p�*竘�P�� �����,3(�@��A���'R� ��^�"�#:��%a-OV�;D��K4�P�'�����M����A~�[�O�I�p���w�N|����E~j)�����oE������L�4K��"s*R� rtA�"$Ƥ(��@j���<�u�J��Xi-��J�&>8u��r��
�O��8f��H��Ǟ�҄�1� �@���L�;�O�<a� Y��ڋ�ȑ�QkD�s��	ʦ�`���]&��')�� ���Uc!)��X� f
�H�0˶"O0l��/���RQv�)wnd[uei���@�����5jQ��K��O�d��/Ӊ-`@�YN�J�Ʊ��I�2'�bgǖ�L��d�|�N4:�S���ء�޴d��Q�/�<@� �8���e̜�UB'��5a���<Qg/�0k��3@�3�'{z��lú���1�Z�����O0����6����5{2��[���B]��'�`���hq�+�
K�@3!.
$bLD�1��)D���� Xcj�^b�ek���y4�'��>���\�:��頧C�8q;1�GC�v؞,.�#g�剬H��A�R/�s����'��S��C��,�5��.J�/���'���oL�C䉾
L��l�.<b�����o�C�	
0��5)��G&�w';#)�B�ɪc&M�T�ܳ ����	;j�B��;N�[7g^$6�ᐎ@+�dC�%r�1���aU��ط���h��B�>�tI�M�2�ֽcVF��5ӌB�I,v�@d�B@�Z�Ja!�.�)��B�I!+�0��4J�>�6q��)G�B�	�
�ʕ����B�켰��"%�B䉫"����Ϟ�9�҈ٵjҧMz"C䉦'�ĊR �����o
6�<C�	�t���i �ƌi�h)�N�n�(B�I�J�iS��E��h�*�Q�B�I�2����s"U;3�������!��C��`^�C%�� Q���Q�K�0�PC䉡;���� ��e��=�Eƞ$j�C�	�[�"a|	���39BC��j��;'-b<r(2G�PVC�	�|���	c,ʸB<���0�C�ɿS�lţ�Eٮd��=HaI?�B䉕U��( �Ȳc@\�{�'_�{��B�I�b
(�t�$K*�id��PD�C䉥<
���S3;�H�@�N�"n:nB�I��X���'�8hR4 Ā��.9@B�iլ`$���l�
yaCP��=	�'�D� *�I�%kA#B��N�z�'�h��2e��I��aP)h2y�'(��p%���v� E�w��f��(�'b6���!�B�T��7j�\���'
�izC(�%��H׮�l"heY	�'�h4p���L�zU#�л
����'zz ���L�R����)��'�`<��;]n1�+·m�a
�'�d�&D�E4ސ�6dV�k�	�'>��z��!H���3�^d$}��'�>)r(�v|>�b# сY^��
�'��x��������掸�����"O�ɛ�猡/�4�C6G���5�D"Ol�[#�_�~�	��r�^��3"O�4��' �e��1 �Y�O2��{D"OȜ�n[)K>mP�@Z�����y
� �hr��4�ެ[P�@�i�A�"OL̫V!�-:A�tN�!>$4k"O4iSb��V���"TL"'����%"O���æ(@��a���6z����W"Ota��
0`(z��P�X��4�%"Or��1o-Y r�  %}F ��f"O�ĹUcI�u�XDY�!`Y"�"OFt��d�[zT�ٝ/���&"O�D;Qg��PUIa��
lDa�"O>D�V��+�Q#O�w�B��P"Od���k-s�xɈ��K7~�\���"O�A+A*�$hG�U�bK��Rc��pW"Or��4G�>bTI�u	X	r8���"ODL��-Y�6���.�7L&��"O\�c�xGLAcԍK&E\��6"O^QPÞ�
U��	AMU�P�"O�����G�j0��� c��E�G"O�Ԉ�h�:C" b"�H��AI�"O�$��d�-�U��OF&�zSq"O��iC�V]�|2��r���Q"O��3LE�8RҬ@�K�V��2�D�*L�H���-ι6�*}($j��"�1OhM ᯑ:}��qS�ê_q eB�"O\�	*O�X�$1�Ŋq�<"O��`��e��8����f�A��"OZ�{0d��O�X�h��R�vI"O��$.�;rx9#t�U�6�V"O����F��0H�	�c��(�E�I�x�,G��' j�q�+�}��&2R{ �|y,Yi�'���,{���ccޫ�,�'�� m`ԧO8P�o� @������O�aу͇wS�*S(�ˤ8��	 2��5�'a​������~���Z�Z��1X�ኡs��SΗ?n���+��yX�Kyb��I�6
�LM	Э��H|飃.̢Ӗh��'.A2�k_�t`��'d�:<��Ңd5�'8Fܼ�I�")��`3y`��q�[>j�`X�P������(������!&	��u���Z����b��۟�|�ԟ�2�G y>�]`�Kƒ��i�Q��sy���C��&�f(�1mߖ�a�Ԡ� ��]	��U��Ri�Tǀ̠��Y�����M3��
ⱟ*���+փ��/{��
)��W��0��fN<b<����Oι�4����0|R��,p�Ip��P�)I�����ٝ��B� yƪ3gva�4L�6Q�"9��� ��aɃ������A9\�˂'�g�)�'5'F0�d�������cܗ����#�"ah����=�6��6#����*V�R	�l��(�u�<12�M�@c:��l�&��3q��n�<�$�Ml{�=
�7�9`��^_�<I0)@/q�(�$=w����O�\�<��j�	���>!��Bb�[�<1e��\1��;��X���p�$k�<��ʪМ�I��:#�2�kR{�<�獃
sjƴ��d���B�Du�<�#Q�!khъw��&��@s"�\�<��N��Z�R�Jpm�	"��h��Y�<�։X�|�F2�iQ�a`S�<)���-�jYC�CɈE�t!���O�<�rcR8=�"��AaS-,�X�(���t�<!��O)�&]�#E�&gJ80ag�p�<�(D�?� �0ؽ.?aR� VW�<Y�%j�V��/T/ۨ�1#RP�<q#♉Xt\���*gm��KT�u�<a7%L?{`�H�n�' �P䋒�R|�<!A���`��Av����h����A�<yk�	�d�:ҫ?$��:�aZS�<�1��tk4�@��;4�� �b��F�<i�h��C���xfɖ:�R�Y�D�<��/T
ƢE+`��DT�,���k�<1b�Մ�z�ǋ#�H�P�	f�<� �!��ˆ=Z6DX �'U�K�"O�`�ѣ��t�x�����,T��2"O���M���V ���Q;#"OfE�v��M�� ��ȑ,���Z"O�7��nX$��E܉�
Q�"O�ԈWIˊh������f�Y*O�D��-<.��1���Z<���'�`��@�tPH�cW:V����' ����O�i�����,V
h
�'��!���C�"�+�k�0z&��R
�'�R�$�O#����"g )I��k�'l�EB�-I��=�D�5wށR	�'x|�Q�>vޕ8T�݅e��		�'M���ԝ;<�X!�(�V���S�'"�,�ԇ��6�A��B�c����
�'/x�c�4~V�=��(�.hR�0
�'�J {w�A�7��5 w�.o" ��'R��r�M
�E�6Á-�����'E>4��#*+���i慓"Oo�4��'+N8i�F-�"A�E�M/B�5 �'��Q�)C���0Y�?�xI�
�'?T�A��,��d/�I0��*
�'u�}C��ظD64��Dƪ�z�J	�'}�IblDKJ�C4`Ԛ;r�q�':�(��N-p��C"`���`��'JzA�����D�x���Q�S�	K�'i2�g`1S(p3s�����
�'!N�y���m��ْI�T����'�����6wa��'��	TÖ� �'�,zmÀ�*�W,�!Q�p)�'���PU�D%�f̓��Tk�X@P�'�b�����)�Б�C�c+�0��'s��{�MM�U��K2`��W�����'��}j��!OJ�pS$!�g��;�'%�9B@��?q����)D�O7�xb
�'�������Mfm��j�D����'������8 ���p�D�q��	�'���Qel�40�@pzᥜ��6D�	�'!���AbD�0��Dçʞ� <��
�'WlI�&W�*"4�Y4m:qt��'�@��2�Tn�ơ9J�&qޠ]�'���#q*��5�$�fY_SjY�'��EP -�0��=s��ͱU����'¬�0�Z�OJ�Y`o$���'}���,^�bi�F��PH��Q�'��p���	)�`�2� ¬q��A��'�����6 ��R�O�W�z�'<|��$�N��]w$�{����'S�Q�L�L�|�AMʄk�� p�'��%�!A�}�B�����9\i$͓
�'S ��w�R-Y1�A1�*�=@��k�'ظ�;&��{e�4)V`v�* C
�'�dM�$�޾NB�$&�;����
�'���n�i���H	�6`�	�'�P���O������RIt��	�'[�|�$oE�"�
 �c׶v]t�9	�'�A����<(3ĉQ��U�XP��!�'g
 �Tn�F�z���?y�5�'(%q�k�i�n���C����'������_�F7H�����#cN>i�
�'��(asHҙd/�Ȋ1��W�☪	�'ی�Ѕ� �͚3��B���p
�'Md��D���ȩ�	\%3
dL�
�'�~���Ϋ�:C����05�
��� �����iΰ�HG��9�d� 1"OL5z'��Lk�`˓����.��"O"IC4n�$��>y����'�x�0$�|��䘕�БG"��'��H�i�n�^��ʍ�D����'��i25��h�:�Cݣ6Irp2�'͞0[TKŦ1�n�c���#(�'�l�BE튖?���i���6�D;�'����-)!P�±F<z��ʓ���	���[�r!p4h B��؇ȓG��$k�LA� ��Pj5d�u�ȓ1��s�g��O�V�;�R]�m��rKd���o�e����G�� }ZX��p0�`�"@��N��)��`��u�R)�vg�!#��:T�d��ȓA����j��u���G$��I�ȓS���Ԣ�&6�CŨœ`�����Y��h��!"x�+�~f>���jx��7���a�F^�!��a��i�P�١W�$87쁽l�<@�ȓc����L��5����8pL�Y��n���aM�62y�=bwG�6sXFH�ȓA.M3H+Q��Q�'�(���ȓL&��B���m�t	b!r�n̆ȓQ�d����,V��QR!#A����7P�3!�D�B�`��)^����:rX���.
�;�ґ��#��7��ȓp pؘQD _zP�ۨj�����b�4y��:�PD��$�l���E��؀��%��q��B �5�B��}��p��F�/ExNa���#[�R���PYX�`�c��l���ԭ�Y_x���&A@ͪ�(��u�["�3��m�����ۓ�r[��S�M�R�&���a��u���F�\��1�DJ)i�NŇ�z8\�R�lB�!PpܛE��%'dM�ȓ}j �iߑF6B�k���9W�Ԇ�"�X���ʦ*��5�D�B�&�(d��i�Xj���8<�����15Q�i��S�Y��Ă�@����7nN�l�ȓs��٨e'}P�� � Z�����@h��;B��d�,� b��p�,U�ȓ���qAn�xE�)��h(^��a�ȓ/��૕�ItL@	���n�����*�$�kM�WTh]!FMSJ<$�����u��O�*FxPwZ
îч�7H5�5雫���A�A[�ve��<0�)[Ŏ�^���@O� ~���TwBEk��Q�{y�ฤȜ<�����1pe�;<R��`#�T�����J6�33	���q7c	�s�Є����� �(S�H�u����7�JQ�ȓG�D��:X��)� ����l�@m��B��R-�f	��t����ȓJf&��O��v�R]
v睬����ʓ�H�{7	>N�l��4V����C��8Z2���n2�	ۤ%�-$2!�DƑ,����E/x$��e��os!�D�@��h�AR,'(,Ր�n��-Z!��ŊCDD�	um:Ljb�B�͗c@!�dوS��eCwL(Wt\l�RC�(g�!�I�h���(��;_,��$-,!�P�
"͸C�ϑ4OL1��� ��!��=E���%�*I��f%@6!�� 
Q�hV!�X�CH�gHV��"On��r�E����~D��J�"OJXCbL�I��0Z��ҁ-�p9�"O@��Ѷf9F]� 
�7\b���"O��A�۬8��P�kH�C]j�I�"Ov탆�ܷ}xx�B�J�?c�"��"OF�Q�՜�d9�II�"����C"O�hXހݨ�ᗕ'�ѺU"O.0�a���D��E�AL�X 37"O x8U���I+�T���L��j�"O:U��k]�]NP}�b�ݿ$���7"OR�� "J�j����@���eif"O��u���Q���#��_>!��`p2"O��pdJ�	&�FI� ۷f�R(��"O��$�
&7��q[��-'�l�"O;�FǡM6Pt�1]K�L)�"OҌ��jZ�{v%!A�	jU��+T���1��cXVI9p C9FʺP��&D��hr)��9A�}�B-��w������&D�|!��ʦR�P���@!O���A�$D�,{"�?!0�x�f���L��H"D�@��셝G�4�q�=Z�2AsQM?D���$ �J�v8cdJ�^��YaW�(D���@H:���0Pp����0D�а���x'(8k���4�!D� �C� 4Z�AI�N;�<��"D���Aa�	U�4�K�*7e�V=2�*,D�8ජX��j-�M�9�BI��h$D�Rs�B5gt�=��þq���3'(D��JD�6�8��N���H9�n'D�L)�C��%x������BEnt`�0D��a!��+D�\�tM�5��x9Q�"D�|���Q>	<Hi��P�+e��y�i	�I��x�u��"L�9ۆ���y"i�,�0(`c�=�`�A��y��ɈE��h�g�	,kN��:��H�yH_���5z��10�kč���y�B����tϞ"5(z��46�B�Ʌ@���b`o�7$+�}
d�L��XC�./y�!�P�U��x�AX�g�vC�	<F.��F.-x�	���C�B�
C�	<�tȡ�E˥y�Q��V���B�$uޭ���9YVu����1v$�C��+����s�,*�$�PA�Ԍ4V�C�?x����bOw(��Z���r�ZC�	1�.1�W�6#�`s&/9�.C�>�b�� P�fC�h�f	G�69�B�ɭ!�	��/�18��Ż2,!1vB�I�}���ɀ,U�������,�C�I0��+ ��*KS걀c���Iz�C䉪q8Z    ��     ^  �  �  �)  5  e@  �K  �V  �a  =m  �x  O�  `�  ��  -�  ��   �  C�  ��  ��  �  X�  ��  I�  ��  �  b�  ��  Y � B � � �! �( 6/ �8 `B J QS d\ `d \k �q �w z  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hģ�%�it"L�B�x�'�6,�pvb�q�ΚO~��Ey��|Z�(��-B$k�-Z:y乲6�	d�<y�+S�
���w�þw�����k�W�<�WO�,�R�"2*ܥu5�@XI�<�2̖8��"�m\�)p�ESG�<YƦ��S�T���m�<`8$��'o�<�q
44���rT�.U�X��k�<�T@),VzH���F0��	�1o
h�'a�DĚ�GJ��aj�(K�f��tO��y�A �GЊ�/����(?N`�J���x��}����b(9����;TI@챗�Jn�<9��6?�]�s�ߟx�r���B�<���4V��ع�V&%���*�v�<�T�D�p��sn��U���`�Jn?��'�a|�n�1Y���#hF�M1�i����$а<Ɉ�DJ�ax��E;z��U �o��!�$��x���He��4v�&���0�!���
b�Y&���V{�.".!�Ă�o� 87Eӥ�bI:GMf,!��@��͢�@�*=�X�2b�/!�䆫`ɶ�(�BF+M�D9�eh�#x!�D�3vLZ��?4��pÐ�B/:+!�C�L��0(���0�s�%] 0>!�$�I��HF� ^ؠ2�"�
r6!�$�v��Q�DTv�Ic�?�!�$�� �b�
�M�%ݒ}0�-�#�!�$�(���ŕ'q4��­�#�!����2�s��T�x]J����`�!��жU��¨�d"x4:���2)!�d�8�N��3��\8���ŞW$!��?&B|��:y��ңkɱ$!�3��̒Õ�w�x�+��P!!�_;3�:m�'o۹a.0(ՠPQ !�� �a���,g�R�(FP�P����`"Of���L0/m�`�1��M���"ObmR�$�r�D5��X�
0@uR�"ON�J! �Fi3�0�z��v"O�@7'��bC�L:� ms
�""O,�톋M���(7�];yfth2"O�s7&O;
��\���H�J9��"O�X�uB�[L�x'
�ߚ`��"O �!�y�(�@kM��ܨ7"O���R�����Vi��X��L
F"OJ`�$NAHz��g�׃��!�E"O�{P��,uEУ���|a"O�8�
�kOԅ�o��^�Z�"O
�BTK�8 >� �Ο�X�|ez"O���ЬA60/��k�m�*OU�"O��zr��D��/8Y���5"OJ�I�dϙ�|a)��\	A\��@"O�)2dk�os`��*"�kv"O��{�*�5O��qi��-z��"O����B�T �B���Dh�@��"O��J0�X��r �dfY�"OhMxC"O�i��  ��@��N� 8�prs"O�,��F\�B`']Y1:��"O��(ҫ�}o�i��FP�2h�"O��t�׿W��%�!����
`p�"O~;f,�|~���K��b9�""O��* �Y���9k��F�6�, �A"O�qZU��)Ty�Gb�	3u.-�"O��S�F+�!עC`ry9"O��x�IK�d?xEㆁ�>x
�"O�0f �H�����(J̐�:�"O�hiU�'#͌�R�N���"T��"O&8���� ��K&MU�vI|�"O���E<�6uJ�	FR��w"O�<Cr�;U7�Ĩ�+ �2���"O�q��H�9��A���u�y�"Op�" (�[f�����`=�"OZA��b�b���h��ڪf缽�"O~�;���A������2�T"O�Ёd��<��EyQ խg�R�A�"O���2���,0ZTCG/��@4��ؠ"O �*'���;K
�)���{�&�
&"OnU2���f$�u�ϰ��  �"O*��Շ����$�
+Xpjx:�"O��xUi	&FY����q��pP�"O�풁 �����(S�Y�.�y�"OH��G+�%V\pc�i�E�Z��&"O�0A�/:�V �#�86g���"OX�b�X�`���'�Q�f�@���"O��2dC��m��I%�1q֨I��"Ol�s#�S30���q�I:��-�W"OnQYГ2hpS��"n��q�"O�,`A��$rd!kX$K~ 4"O�T��fI�D��1I%��e��� "O�d��)WM���SbTP ��"Ox�ҤL#wʘ��̣AQXݻ�"O�x���X5K�&���h�f��$"O�l2�L/t����%4��qq"O����ʌ@K(�35� ��D��"O��P��h'�Q��㎺i��h�D"OR����4N����<^�� K�"O�Ƞ�X�tS��$e��W�0X�"O��
��dI`�Z愔%~I��1�"OLa����RL���C@Qڐ���y
� ��0f� �"ii�b� ��=�"Oi+wn��)���A �ó���"O��)��чPk�Å�M�^� �"O�C掑]�Ȁ0��~Ttb"O���7Bz���I� ��zr�8c�'���'w��'��'���'p��'�ry���G��&
EƗO]��W�'SR�'��'b�'�"�'W��']���o�N��1�͆�`���B�'��'�R�'s2�'���'j��'Ȧ�2��h�Qaw���O^��C�'�R�'�r�'t��'��'��'��܊��0<Nn�9�&{�ؔ���'2�'���'i2�'8r�'�B�'����:����w-R'2���CU�'���'���'R"�'���'���'٢Ikv"�+L$Pc�,ݝ�Z\���'�'�"�'{��'���'Mb�'�`d�j���9�CB�|U�ڴ�'i��'%�'v��'���'_��'g�1��جtZb�XE�A$V�>|0p�'�r�'/��'���'�"�'���'м�s�T*-8�a�vdP���+�'�R�'\��'�2�'��'0�'$���U�#z!)�c@�24=c�'cR�'r�'Ab�'.��'8��'m���ЍT�Z@��sc�.?6�Т�'���'*��']r�'Vr�'5�'�X�j�K�:��0�!i�����'���'X��'ir�'���q�R���O P @T��L�X&��;0m�H8�!�@yB�'��)�3?�A�is�d���],?��e	gf��F�>��6����Āզ��?��<� ���'�W�,P6��$R�8Kٟ��I�I�an�Y~>��h�Sd�	�?�E�U~�|Ց��*q�1O~���<)���Ѱ<���)7eN���pCF��z�oZu��b�4����yw�F�K^Ε�s�ɻ$�h9үV=��'r�Ħ>�|�'��M��'9�蓖EB�Wlj�H���樜��'U�V͟�q�i>��I|OT�p"��2�ѹ�	�}�\�JyR�|�nӸ�;��d݄Z�aU'X5<���h�G�g��㟨�O��$�O��	G}"eW"q�eؓ�
���ɷE������O�cv)��s�1��k�s����)5�, 8@���}�2&�������O?�IƬ�J��߯T�-K��I�s h牦�M{�&�t~ңb�6��SW�&��Gk"���!�C fA^���`��۟P9vb�Ӧa�'c���?ś �ؑV,~!#��I�XE��yA�J��'C�i>e������	�����]Y|�	���J[D%[De� +�y�'�V7-Ċ��D�O��$7�9Ox9�C�1\h ��R!�&͈���r}"�'6�O1�d��2,�q�hqX���*)f,A0H�a3���<���Ǡf"F�dܳ����V9hf� �'@"#!���a��\�d�Of���ON�4���#Ǜ��_����S��D�3��u��$0VP=�yblmӂ⟘r�O^���O�d�:�ڴ+��c�nJW!�5�=�2	l�b�d�0���.�'��#G�^�5m>����@��v����A�<Q���?���?����?A��D��/�@�b��	6���+���N��':B�z��+�9���
��&�8���O�y��0��Fp�8��c�I�8�i>��i�̦��'�.-胋Q4�:�Q)��Am��"Hʱ8�5�����$�O����Ol�D	$Q�d0��Gfj�I;`&�Zw���O0�4���żv,��'�RP>��$��'��B�P0��& -?��U���	�'��#�� ��߇x�
m����fH^<)���H��w����4�L���BP$�O�\��g
�c�(C���}!ԃ�O$���O��$�O1�
�:i���2>�D���?av�	sgN�����S�h�ߴ��'z�듒?�r%�z����'T�NF^=�4 U��?��L^j�4��d^+��!����S[@�X o��.�DIs�ڻ$����Dy�'��'"�'N�[>�2pcz0}�0�\�r�M���!�M�,G&�?���?�M~Γ9U��w�p9��l@Pƹ��#ؠ*7|HS��'���|���	C�>&�<OZ�� Q�/��ir��^l�u<O5�C�ަ�~�|_��S��i2!@�0�v��A�9kz)BR!�ҟ��Iǟ��	my��k���;�%�<	��h�.�qC�N>9np��C�C g����⪳>q��?�K>2�tQ>��p��&�0��O}~b��:���i�1�,5`�'C�V�I���d�4}<���n�*_�'B�'�r�SƟ(���B2U�Eo[`�(�����ȣܴLbti�(O��n~�Ӽ��k&S�8�o��d^$5	�$U�<1���?i�p'R�hߴ���aM�(a���ʁH�ϑ�(�b8�u�TB`|�"u�<��<�'�?���?����?�c�ë>%4i��E�+� �;" 4���٦�*���П���ݟ�'?��ɣT�``�D.NR�B�, d�c�O���0�)�S68���vF
�r�|����\ڸ�QJlb���'�r��(蟜ɒ�|�X�p!��-J��a���O�}��|�2Xџ��	�������SjyR�xӮ���Oq��a֊SѦ���[\K8�8���O��lZT�\+��ߟ�'܊	�*+�D�i��^���ť�1Y
�֕�|Y����cD���
o����� ~�qU���eJ qҷ�Q��A4Oj�$�O��D�O����O��?�{$��;]B� ��D@+>�x��iA����	ß|ڴC�)X/O�Pog�
DD�۾,:�2ƅ)mȩ'�������#l��o�E~��+��`wj�7 R���Њ̻_����#X͟T2�|�S�����IǟP�aO
	L��8cǯ�%?t \�Bƛ��	tyb�m�dЫ5��<����GY>��`fƃ!^x��"`������d�O���+��?� ��[#}����f���أ�ɗ
P�m�pn�ۦ���t�y?yJ>9�!_�S���g�L�0��t�" �.�?����?q��?�|�*O,�l� ��d�0�@/��ᘱ�p���wM�fyB�fӮ�И�Oh��������#
d��	��v����O*��gkӤ�N�J�(�V�O��i��I��hB�e� =џ'��IٟL�I�|�I����f�de�&G��̒"�.]x��?@g*6-�4qS���O���+�I�O`oz�I8��a���0��Ƣ��@�J��X��N�)�+dF�lZ�<�C�K�8�Pt���Z�(i"�m��<����L�ē������Ol�DT:@������"�l��^�9Rt���O��d�O��SU�� MO��'�b�V�z�d���V�6U����k��O���'�����'a�X��'�;_�����5"��	�w��)%��kA�U&?�9u�'D�q�	�]v�(n���5�Jp؄�I��d�������y�O��\�V��M+����ht��F��2�B*|���<q�i��O��X�M[;{���K���10o���O��NQ|� ޴��D\�?�+��X,Ph�
��8h���ƙ��u�S�+�Ħ<����?	���?y���?9Ro
	y/�D��ؔW�&< ����ɦ]#ę�������\&?��I�]��- �bW1q?�r�(�=��O����O�O1�ʝ��M�v�:81E�_�	�0��$��:w��<	� �Rz����=������'y��h  ͍�Z���C���|!*��O����O��4���6ԛ�*/�¡�4iR��˔,Պr�Mz�I��#{ӂ�x�O����O,�$��!��r����qP��� �,�8B�lӘ�
��\�1o矮�>��]1�P�B$M�o��� �D��7���I���	ߟ��	�|�Ia���N�k K�	W�pÔ�J/5PH��)O0�d��)�t�u>����MKM>�1#gi��$� �\�@�U"uS�$�t�I���d=RmZi~rcƅk�j�	�,���Ie'ۙa��LP�^?M>�,O���Od���O��Kp�(`�v��H�S���@�O��$�<��ij �1A�'�b�'X�S���톷]���j6�F�D���_��I���I\�)�\�E���+��T7)���8��Q�^�@�B�� �M��Q��ӐX�d*�$K�H��!6-��!�.�V�� �"�d�O2���O
���<A�i�*�	���逐C(��C��� ���'\*60�	����O|�!��ΖW#�#a ļK6x5�w��O����/|y 6�'?�����@�}y�+K�(�ȑ/��ڔo�h��$�<���?���?���?�+�Jp�ui��\T��J^�D�.�����m{��Jy��'&�O�rO��.����s��N����b�ҀY�����OX�O1��\*p�v��	�z[F��1��Nbu���ƃ<���/ ���O��O�ʓ�?��C6����Q���25J\Y� ����?Q��?�/O^�l��;t-�������z����3|R�K��
	#Zy�?ArQ�������'��B7N�z�`��ӵ?C,(�c�0?���'Cp�@ݴǘO����?�giL9`^ސ�5h��p
��(b�G
�?����?����?Q����O����"fj�Y�QI��H�Y�gb�O~�nڀud(��'n�7�'�i�5�1F������Z���w�X�Iȟ4�� >��lZh~Zw ���g�OiT�1 ��%E*���GΈ]��I��J��Iy��'�2�'1��'=�;NR���ϔ�h*��6`�
@T�	3�M��%�5����O�����$�~:p��QDC"&D�h�I�dj�d�'Z"�'�ɧ�O�B�	S�+Q^t�X�E��Bk�X�#ݹ(A�J�OԈ��F��?a��+�Ħ<�Ab�\�:1�b��8`���%�_�?���?����?�'��צ�ɴ��ϟ�"�=:���	�W����R(|�`:ش��'���?���?	4�_0�У �VDv�M^ږ�"ֲi���6!x9��ONq���k��Y�FN?0E�D�e����Ot�d�Ox���O��$!�MDz���l�x�iuϗ48�������4�I��M��+�0���L��}%�l�4�ͫT�X�#A�@�H�Q��t�ޟT�i>UP�e��%�'�&�sc�2B�yJ� �>7,�;��M4U�2$������4�^��O��$�/&jL�#�
^�R
���Fʚ1�:���O�˓1U���̓5�B�'�RU>��D@I���e�v��+Ͷ��׭$?ɓ]�$�I��&��'q\0&�ť3u����hl,�a� 32r��ڴ��4����'��'�NK3j�0�	Ѧl�30SF(@ �'�R�'�R�O��	��Mb��1�J�k�&Ÿ]���Se���0�+O��nZj��[����� ��-�/N�BXR���7���BA����pr� mZ|~��Ӿ� �SO�� ���*�8�C�B �)1<O0��?����?	���?y����iF�n�()�'Ʌ%�`�FH���mZ6]�0�Iٟ���O�S؟H���� zr�`R��		^}�$��O��?����Şxa$m�ش�yb➎}�>4 5�#dlD�S#�y�CP> ��䓃��Or�d�
�)����c~���Ē���D�O���O˓e����� �r�'tҰ�`'�1��`ǖ�D@jfY�1�O8�'G��'��'�����$�-��pGI�/HS~rm�w���I�!���O����I#�Be�F���IA�k���1�B�r��'���'e��ԟȺ�Dwl�����"��S�W�޴[��or�B�D�����?ͻ+�>Mj���Tᮕ��-�V��̓�?I��?�P̉�M��O�u�JT���4�<�R���F&2��`@�B�'�i>-��ܟ���ş��I`[^ �/%P�Ʊc#�Eȍ�'�<7�י���O�D2�9O��� ��	r�����"��X�G]}R�'e|����	��TÔ$�^����v��	w�$J��ɷ���ұ�pi��j���O�ʓd�6�ʔP.2d��S��)����?I��?)��|
,O
MoZ5�4�I��`�2�9T�R|��텿]vԡ�ɰ�Mk�2ʼ>����щ|����o�Qz�S��'l�=��do���:�ܑ;T���.��K~Z��T�찒$�;!���Df�PȂ5ϓ�?����?���?Y����O#N�)#�MK��`
УލP���#vR������M[DRq��n��O�4ٗ�4By�\�ЄH_��8����O.�d�n���4���J��MsE-�	H���+I%&��q+�0V���L�py�'i��'���jsrA�$�"x>��G�6lN��$�O
˓E�Ɓ��B�'�"[>��H��g������	ּ��so&?9�Y������P$��'u�lA �!�1�@�CW�](�qX����e�GӦ�-O�I���~��|��Z;VHt$9׃�hJ�r����P��'"B�'���Q��X�4�u0'nT;��ڀ��"y�<r�����N����?��]�8��'$2h��LB/�V�)��%� }��ן�#��֦y�'\�h����?���8IK���-&�t� ��/5vUct5O�ʓ�?����?)���?Q���i���L$���ϛ$Ҳ�� �K	X�l�T���I��X�IN���� ����1����\�9�B&?r�#�\��?���t��;Q��f4O�5�2އc^��2pd�&��ܰ�8O�}��e���?Ib�'�$�<���?	�a�)��@I��P4����L��?����?Y����H��d��ӟ(��������D1�t+4�6��O���'�R�'8�'t�P��0D$�⤌�E2	��OL���IQ�ndB@�'��ӗ�?@��O����U	�j�iTJ�8�J�!��O�۴�?����?I��i�O�M��ƛ4�`<���S���Tc�ODm�<ԕ'��6- �i�}a��B�Dd#c��5���F(`���I��I�.f�mZG~RDM�l��,M��r�-��YH˖p��Uqǔ|B[����������۟�� �M�1,b̫7̀A�\�����Py"ly��5��B�O����O䓟��M3z�X�HѵM���`���l� �'
��',ɧ�O�yeټod�y{6�9v\P�����ou~��'-���������� )���rAկ܀�k�c8e�"���O��$�O��4���tٛ���_
R-B�-W��b�*�-`F�jqň5�y�y�D�li�O0���O����� ;�=C��W�	���0����,��hZ��zӤ�S�PB������>��]�+��Ȱ!�$�0��$ $o�Iȟ����h������f��>h�Q��0|
��r6B�>Mߚ�����?���{�f�-p�	��M�O>y�o^2X���_�:���Z��?�,O�H�d���G����f��0Btq��OR.,�[�)��n<��D�������O$���OX��-*�i�Ȗ>gO�` &�_�J�(���O��g/�F�H�\���'cr_>@7dK4��X�A#�5L�$P�$5?�QS�$�I��L'��'.��<�FٸF�R�� ���F[��)�#�6q��45P�i>���O2�O`aR�a-�l�"��SCU 8�P��O��D�O����O1�D˓@����?!��j�-�!\�e늣t���_�Đ�4��'Q���?�UO�����б�J�H��]�₍�?Y�A�JTI�4����z�p�)꟰]�(O�L���̩8��K�ʔTuLU+�2O�ʓ�?����?���?�����I[�G�ɑg�"^mf�Q���mlZ&Q�1�	�L�	v�s�����#An�"���3/��+
]���?Q���ŞVa�	rٴ�y��Z��BȠ�c�ZMbQ��O�yR/
0�������4������V�K�c�-�����B�O6��d�O���O��%ě���K\��'�������T��O4E�9�� -}�O�0�'6����4�xh P�!�����	�u>p��B�p��$?I���'����P�~p���TV�#��C�M���	̟\�I�����I�O��,r� "�M�F�\
0K�WCk�4�Q��<١�i7�O�.�6&��e	"-� b{���!u��O"���O��
�Ev���/�nx�V������ x�!�L߬$����F?	����'��<ͧ�?a���?Y���?1�b�0m.�m�q�U����9^L��������I���$?��sU���&���e���s��O��=�Ot�$�O2�O1��"�#�#0�tvU<hgXm��E�
7M#?i�e�M2�	U�IKy 
1���J!h�&��l�r/�*$��'�R�'��O��	=�M�KY�?�� �\�t��r�:h,j�r�ˉ�?�f�iU�Oj�'�2�y�nM�C�¬٠�]&6.z�[��؋��y�i�IcoV�S�ןĒ���nKaPRّ�)�%u_:��B/�8���OP���O ��O�D9�S?1B�`� ��L��2t���	����I	�MR��|��
-�&�|��B	^\���@�q0�t�b��'�\�PC ���'�,L��c��&P$-k��a�nQ�ń��&72�����'6�	���	şD�I'I{�Z0	�)��	(�Ó5~�����'�7���F�$�O�Ļ|�!�ڰwP���D���B�Hm~���>����?iO>�OV�JѡیEK섊D�.5�`��qe����QE�i���|b7l��'����%N�d�/��% D۟$��ߟ��	ןb>�'K 6�C��(A�F�uUN�C�/ԍ 0����<a"�i��OX��'X���W�Dus�҇��Ç����U�0�n�|~RK�:gD$i��?|@�(�89�S�_7f\�Q��,z���cyb�'�b�'���'��Y>�O:h��gE�[�͢����Mt,A��?y���?J~b��i���wq�E4M�d�D޾f��ZUm��?A���S�'-���Sߴ�y��E�O�8I�P��>�P��3���y���4R���䓨�d�OF�D
�]f4�p�RS\����EӢME����O���O˓s��J�.n��ҟh)�#P�r�N)Z����)��H���FV��I�(��m�mR8d�3�t�.��oF�u�N�A�] �#�2��|���O&�X�RLL���&[��V�=��E(���?���?����h�N��JFÈ��eİkM�,r����ď��b@�ISyR�b����5t��'E1<z�<bK3E����������%GU�a�'Ƃ`R6l�g2��?6`� V�9�TiR톩�䓺�4�����O����O��䟔~`���%&�ق�E@h˓@�����;�'Ґ��' �I�r�5'r@��D�^%G����Ľ>������O*TP�Ì8KV8�4�	X��[�NM�]�8��3P��wo�84 2C�R��yyG "a�v�׋!
\��#��*B b�']��'8�OK���M��]��?ٗbն�4�Hɜ/&L�AJ�<A�i"�OP��'�'�r�̹M6<��	ƫ�|(�Y:YJ"��7�i��I0g�d!3C����񆩖:g�(`�� �j��H���r���IΟl��ܟ����,�R  ��h�+S��,�����Ë�?!���?�!�i��q�O R j�z�O�a���0�]�b�+U˚��q!=���O��4����qDqӚ�uXƬa���(9N�9ҁ^�Zᶴ����]ܘ��C�	ny��'�2�'�"��iF����M�C�y@�#�#NwR�'	�	��M�F�������O�h s�
=m�%��l�&�����O4�'�'�ɧ��e��X)B�Л4a ْ&�OM�(Ф�W���������+�FMd�ɶ{�b4P�Њ��łaG2�@��ǟ����)�jy�.yӼ�A��f����eފ/�쩳��v�x�d�O>�l�S��+�������l�;H��xg?=]H�q��ԟ����/H��n�A~b).�����U�IB~��|a��Ъ������GIk�<���?����?Q��?�(�
���ł���K�i���;3��Ʀy�tG�ٟ�	��8&?��:�MϻQ5���c���8��m[��+Dݘ���?�K>�|brhٹ�Mß'���s��G;�S�@�y�p��'�N9z$��~?�M>�)O�	�O����W;N�񤎚AT<�N�O`�d�O��$�<	 �i�lq��'l��'��8â]/5O��(a	��~1�$�n}��'��O4��G�و6k,\z "�*A>�A�\��D,$52�8҂�t�/%0����0���аE8� ���ñ2���'`G�h�I��x�I��TG���'^4X�bH�6�������'Զ�Q�'�6�DU�����4��Is�߀@@��CxA���;O<���O�����6�9?I��[ob���2
lH���I4�v���Ǚ[,'����ڟ�����	Ɵ@������o�]>d����U"r�ع���Gy��i�t@�"��O:���O^�IĆ���O"@B��*N��K�&�6ڈչ���<I���?a.OD�'�?��t�&z&<~*u�fhhHnp�5��L�'ѐ�fK�ğ����|B[���Cɚ$[\2��eǌ�3�
���ş���ϟ|����ny�"k�vq����O�\��� ~"�y���� G`��7K�O�lZv�M�	ޟ��i��z��Ի4����D�X��a�Ƙ����nC~��c��0���,�O�7/��L���ؑ(F:*茹��ƨ�y�'�R�'���'�b�	L�VjXT�f�7-3QZ@�T�2M����O������i>�����M�M>)Q�'���sw#�c8Z�%JI����?���|�6�?�M+�OHT#�� ���m�<rl9�C�'�&�8�ǌ.�?�#�6�d�<�'�?���?�u3�>=��2U��]3q�ژ�?����BҦe@��Yȟ4�I蟌�O}� C����P�j�UE�-#ġ�O���'c��'�ɧ���@����7��#%�Z8`�N))C��z��;]J�7m1?�'�r�	K�I#=�|:��"*�ڐ!�H����I�\��՟��)�^yo�Da{@�:UN=�E!58#�F�4%�����O|n�E�o���ܟ rgʸ	�a�H(}o*�z�!����	�)5��o�G~��?nMl��SY��ָ/�:�ˣN�(Ю��� ��3�ģ<����?	��?!��?�(�6U�S7h�4p��b�7)P(!��O�ʦ����Ɵ�	�p&?�	��M�;n�~��6��PͰ�̙:84������?I>�|z7���M�'>墣��@tn���K��!��Q��'h �
4�F��Pr�|V��֟���Ɍ� �	3�k�h,����^Ο����`��oyrmg�d�'J�<��N�N	��͈!j�.u�C�$�����>���?�K>�0��6jc�4�Q8R��E��M~B�6����Ҏ���O閩�I�m>��p��+�:��rL�B�'���'���S��H3B�&M�R�0��_�Jݢ4r2e����"�4t������?�5�i��O��S�M�L��㚁L�F�X��]�f���On�$�O¹[Ǐy���P.�a��'�?q�$�
IA"-`P�Ψbʀ+%�@e�hyB�'y��'�b�'�"�
C ��9�cG2T������yd�ɂ�M#`Kۘ�?9��?��t�?_�Ir��$�%�!ϸlwdꓳ?����ŞX�q����������\���H�0�M�V����nD�GքU��ȟt33�v���i>i�f�ǫͲ�Q�)1T�d1�gVȟ��I�:a��R�����l����3�uG	M��yg�17����6!
6[��슅d�4'iT�4�'�'��P�R�'��w���GIO��e
���Xސ��BÍB�V9O~�$�/Z �|����;{�D�����9g�5������̓�?���?	���?����O�&��Q� o�I��
L?B5j�'�B�'0�7� z,�˓W���|��1/�]��o�.)���v��ޘ'!rV��a5�V�e�'~���r�Kf���TJA'ʁ��%�^��0�I�N��'��I��$��ß��	�.'(,	�b�,@O����OT3:��Iٟ��'��6͙1��d�Ol��|7�u�U���F��=��K�o~�a�>���?O>�OM�Հ,	2#)��%I��M�\͊�D] x�<��'���4��}��]�&�O��
6a�1�d,�Ҫ�2?y������O��O����O1�r�2����^�Y\v`�s(�Y���q�V�{/
p���'��Mp����:�O��dIiި���b��|TB�U�J�V���O K�j��+��8�?��'w	%���n4���B�L�
�'��	��4�	͟��I�8�	k�4�_�HR�*��V.Lf��t��#Y��7K�~d����O4�D6��=�M�;"8�TPƭ�<{LNa
Ď��l�� "��?�O>�|�r�U�M�'Ķ�2B�$�Z�I"e�2髛'�[��ޟ�Q��|�[�l�	���@'	�l���*�Ǔ�]lL���ϟ������IMy��|�Ε��	�O`�D�Oh|S�JJ�"�8(��v`0YǤ'�	���D�O���%�D�&�r)� ��r������9���63��=>9db>Uc�'3d��I��UVČ2���� �&5�0d"��'���'��'��>����<��p��Ȳ4�(�2G��-t���I�M��iЀ�?��A|��4��	t	�.D\��2 �[�64O����O��$�NK>7�3?�w�K���ӕ{K2px�*N���3�˕�bx$��'2�'Q��'��e�9�xEJ���3=��<9� ����������I��`��Ο<%?�	8?0�!��@Z!)r���ĝ-nz� ګO��D�Od�O1�P�[��̨~H�y��V�>��m��W�jHr�*Q�����&�*.��Ni��jyB�ѥyg-�`HN;lJ�����PI��'�r�'y�O\剑�M��,K��?���Q^b��'*��$9>E �o�?�v�i��O`��')B�'������l�5�"�)�O �2��ӻi���>TV4�$՟������}�2P�g�B$n�`�T.B��O����O���O��$(�S:O"���Bȁ����Y�ܭ����,�ɷ�M#4'л��Pn�u�I8F� I�CCv���'��A#ڕ'������ӛi~�6�>?ǈ Bă`Xlg�����C*:@Tىd��O�U�N>�,O���Ov���Oz=�C�Ƀ>��06 �PU
�E�O���<ɴ�i�~A���'�R�'��S�k��p+Aɾq����Q`8V�M��I�����w�)�"�Z�=�Z�@cJͿ;Z �fK�*�(��pn͔�M��V��S so�$��B�1���S�끘F�bQ�GFW�V���O`��O���i�<)1�i ���Ύ�m>A�p�ث+lH��$X��Ɏ�MK��Ÿ>�@'�Jү��x�( �e����?y�F�M��O��k�����L?1��͚�tb���K�4!���+�~���'���'�b�'���'���bK �H�۳`w��bW�]�g����4"��uc.O�� �)�O�(oz��$$�[����4-X)w���U�џ`�I\�)�S";Vmo��<� ze�������I�*�+ˈ���2O�� h��~R�|R]�������U�N���c�B�(6Q�Q�Dn��p���(�IJy�ft�F0�2��O^���O��vN��y!Ԡ�1H�*e����PN/�����D�O���Q,߳6�ۅn��]8�1F8?�����`�L���'�$L2�?�m�^��Vc�`�� ���?���?����?!��	�O��	��x�X�G�T62�@����O` o�,�ʀ�Iȟ��ٴ���y� ���*��V�V��F��y��'a��(}vb�m�L~�o�n�T��S�P��pB�L�k���:���5RmʨZ��|�T�`�I�������Iן��P7�a.����Z���My�Ev�n�
�g�Oj�d�OȒ���E�IJf���R�z���晑0����'.���)L�OgeB���"�t��@O�0X�i�V�\�6En˓uc�`ц!�O��O>�.O<���҉#�x"���&B����O��D�O����O�I�<Iֶip����'��ܐ)���qf̏ME�M�'5�7�>�I����O
���O�
�+�/~����v�&"��+���6�4?Y�R�����>�S��Y$l�h��{�CW��6�d���	��t�Iɟ8�	ß���!,��4D������,oe�x��/��$�O�mmZi�~�>����|R�Zd�����<C�nP�a�M�'����� $%�֘�����5�*0IG��%��)l�(�Q�'�t�%�������'��'��Xa�D�.,�r
�b���r��'�^�t޴}~&����?Y����I�=L��r�B_?OQ��Rn�h��&��d�O��=��?�A��+�J��@��ۖ�S�/$�)�든i2��|"0��Od�H>��%)z�(h���a�>�����r<A�i�4]��-��|HVGO�5`\��I�Z���'�6�-�I����O��
��V���j��R"q�0���k�O$����6�>?�Ĭݯq�R�TyR,��Y��AQj�@���@8�y�U�X���P��ޟ��	̟�O����1���(� �JN�_��i�e�y�V�:"�<����'�?�f��y�'�0,Ԩ0p�U"-�~���]�T<��'?ɧ�OF��b�i��$�G� ���A�%t��z�.�p��$Ъk?0y��RﰒO��|
�\Zeh�gL�4�d�9�aG��Jl����?����?�*OmZ+:q����֟D�I�����
���y��תs+��?Y&^���	˟�%� 䌒�@4MpD-�.4@Z=�C)?��H_/*1+۴��OU>X���?���v�����So�b�RK	�?!��?����?���	�O�T�$aMZ�Uy��:w}���� �O�l��,*b��'�6M+�i��86 &Y�.����C�Z6��a�Ea���	����(q``m�N~«� 1z�p�S����E���8aS�!� 
ӑ|BV��SڟT�Iԟ\�Iʟ�3�\ +G��0VOF�9�t�:R�zyB �R*���O����On�����%a��T��CX\:x��F��:�`I�'���'�ɧ�O����F㊼�y�#��9�1��
Ѣ4X��©<���A%\���A�Ioy"KJ�	\��ɕE��~l��+�'8�"�'���'��Oy剺�M��[��?y5O�jbL\�̻R��a3��<�u�i��O���'%��'�"�Q�j�놈�d�Q�c�V�ˬQB�i���[[f4�T�����憋��<�Gg�9m_��%f��������Iß���Ο$��C Ϣ}j�3T��/�ڬF���?����?q�iÂ-��O?bf�ޒO���w�O��(e��a<������O��I���ش��$	b��`b���m%���FAI" N�}0Ď���?�V�'�Ĩ<����?����?A��Y7n冤�U�	�]����f�?�����D�Ԧ��É[}yb�'Y哂/�6��%���8Ek�L!$�	!������	a�)Z��*=��4� G�-��	����d���*��[=f(�(O���
�?ɡ@+��811:)���U
T�0�� `���Ol�$�O���ɶ<���ie��3*R@����L�]*�dk�(�$`��I�MC���>i��Ml�zPH��_���5��R�l�(O��c�cӎ��h̫E+�1�+OL���-�oNQ�p�P83;���6O�ʓ�?!���?Q��?����	)1HD,�b#>��*W��L�in�3[�����$��v�㟐����ç"����w�\:}�����?1���ŞKT��1�4�yb�޽;��' �eib���V��yߪq�<���!�'��ğ�I�C���9��e�@�WM��"��\�	Пh�Iԟ�'q27M��P�����O4������aB�9���	d��4C]��0��O���O�O ��nͥai��g'�9��TI������N�9v	�2�R�ӥ8q��^���)S�M/rw���`��o�TݩDKԟ�	�����ןE���'^�hY���[LJ�� �"��[U�'6�!h��~���4��|��+K�*68 U�� ���s8Or�d�<q���7�M��O���C.����V�W�@p��b :i��7֋���O�˓�?���?Y���?i��o�nY3r��l
(��QR����I.O��lڠ�X����4�	w�s�8QѠv.� �^� �p�:�����d�O��b>!J�.=� ���SǆM_�����@���'	�?8�ʓJs\ ��+�O�x�I>�+O(�zQ��J���� �ET�eH���O���O��D�O�<�c�ibL�Sc�'R�d{Vk�r� ,� ML����@�'�<7�1�I���D�O*���O����"�QO�<c3���>������kz�6�(?Y7��1���	5���Y�b�&0�v�i�+�)od�i0�r�d��ӟ��I՟������Q�Atׂ�0����bk���?a���?I��i%�5{�S���4��,6�M���>�2��Q�X�2��M�J>����?ͧ~�fLQ�4����rS&��3dCy����ǜr �}�����~B�|�Y���ğd��ퟠZ��Q�A�f��uY�B! B�h�Iny��b�JX����O~�$�OR�'C��L!��f2z�ȱ)ЍTG���'�nꓴ?1���S��(��Б	�, Q�,أ��j�bE���P�o���Z�Q��S�C�"kT�I�%������W��]I5H�KA������P�	ϟd�)��[y��n���!M_|M��QV�L�zt���냮c����O lZn�6��ן K�$������!6��tS��⟘�Ʉz�V�oZ_~r�E0b&h%�}z��<�0�S	9~",�B���<q)O����On�$�O$�D�Oʧx��h겢����cˏ�?r�8�i�����'zB�'��O{��n��.ż��X�b)U�e�>%�`a�7���4�)�=d^�@m��<�UO�1O�^��v�^0�z�R�i	�<��*o��������D�O4��O�e6�H��5Z��j��Qx��d�O�$�OD�A���[<u��'d"-^G��d(R�nLB����ĵ.��O���'qb�'D�'x��'.وY�\���K�~��Ob9��2@��������2�?�.�O�bU���/Ǣ,[��1,�:�(�,�O���O��D�Od�}λ/��3�*�	ma��}�n��
�����1m"��'IT6�"����(R���3�&��Ea�ά��<����?��)�*���4��$v�ШQ�O��A�k�.�ƅ�ՈL>b�$tԙ|�X��S����������0s��ϻg�`�¡8b�	�owy�`������O��d�OP���䐙r�\`�T�@���ȫ���X0΍�'�r�'|ɧ�O���E�D$眓Sx��!l�HH�O�8�ベ�?��=���<$�Y#[��5YuH��c��@D_@�س޴)�6(�x��պ$e֯'D�ʁ(�8i4H`���}W�6�d�T}��'R2�'}�h�2�	g���K��^,�2���7�V��0���T&��=����R�x�o� �!Hو%���:Ol��DP����0���xn��+P54%�d�O�D���E+��$r��i��'p���!��,�lH 茥P���"�|"�'k�O�Q!�i�I�;�@p�NK'E���pܪv�^� �F�_���1��<i�2�H�\*�l�"�f��Ma���O��oڀ[�p���˟,��\�dN�.��L��!!JZpl�?���a}r�'�b�|ʟD�0p�HPe�$h̤[���j#�yȢfg�����4�CW?	K>9�P�6p�Ĩ��)�W��x<��iʊ��dA>��-���0y� =H&(�8L�ɠ�M�2�>��mq(��B��&{$Tjt�ʴFiV����?�Ԉ���M��O���,y*��˴��t����2Yʌ���V d=���'}��S��l�S��,�Mzae�1�t]q��:�MS@�֣��D�O��?�X�����U<�@$Z�k���Pl:�?!���Ş&[�X�ܴ�yr,J�@�lu� ����`�'-�0�yB��1O������'�fy2�T�z�H��FͤG�ĉ��0<���i#�	s�\�8�ɹ��Q���ǫ:���OO�����?i�S����ß�&�!� �B������rрu�,;?�go�R��Q�4n����'X���$�4�?�e�C (y!��	*�5�2Wq�<yVi��y����g��X�"�h�J���?q��i2�8@�'L�
rӄ��]�}m���g�ʖd@עƨG8j���l�I��4An���'е�q�O�$�>��A�t���|j:X`�H�*����d�O����O����O�$J c���#OW�P�����*ȖʓE/��P���'`��'���Pg��@����2��JNԨ	��>���?QJ>�|���,V��(SM�o�@Q��\�mu�8�f�M~�h�<��P��d�'��I8jTYT�=�b4��JM���������I����i>9�'�Z7��\�����z�n���A���ۆ�.pv�dK��5�?��_���I����I+JUK%a �F�x��Ѱw�@�7�Ԧ��'�������?a�}��;a*6�j��EA�:�r�+)���?���?y���?�����O�����
B.d��L��I�)Ik��'���')�6�N�V˓hH�ƒ|��ڴBB�P�gQ<]��*����V9�'������H?������6(�3'��A�6�0&x�e��*uPe{��'�N'�h���D�'��'�^���n�d=���L�~"�ȳ��'�BR�L�48�a���?����	*�& �����P(���	����O���"��?� �M��'A~:LAh�t���"܄1|(�B�E�4��i>���' �%�|)Đ26��c�'� ,��2��ҟ\�I��(�I�b>A�'n�6��4��	��> "�@h��
�M ���<qQ�i��O�@�'R��[+Zh1E�v���1�`۝@e��'��('�i��I�
L����Ok�'LAr+@M�9�i�����������OV�$�O8�D�O���|jB�T�	:F���[��d�/�>���A1����?q����<п�y�Џ8�~a�OÏ^~��ن"]�N�'�ɧ�O20�i:�$̙z�ܹ�g��r�F :��H�$˝s}L ��&�>�ON��|R��K���&�xH�kR�ζ D`X��?i��?�*O�\mZ\���'�2 �2ͺ�s`��2������C�Ob��'�b�'��'��8Q@!;^�=Ac��u�V`��O�D{���T�b6mz�S�B��$�O��ѧ��K���	�nO��~��5f�O����O����OҢ}R��t���ڤa��QfdE��gׯw�j�)�S$����4hs��'�B7M5�i���0�=o�e��bU�RZQ8�#w���I֟\�I���n�}~b��V L��'&�6ujW�E�M�~�GI��hH)H>�/O�d�Ot��O��D�O:|����:��Ȑp���Vh�ԙs��<�°i�|1K��'?�'b�O<���LJ�A��R$~��Y��n�s(�듎?����S�'"x�9;B'�#Ṵj0I�og�\� fö�M��P�|;���0��(�$�<17-̺8��҂ꌖ)���ի��?1���?��?�'��D����iBb���l`d$@ mnJ��7·�$?
m��FƟ��޴��'����?��ӼCWF.�n���P:ư���� Z�
p�޴����F����OZ�O��NO�y�*��\�o�%�GO�&�y��'u2�'�"�'�����Vx���"�@��iH��Ȑ����O��ɦ=�w>I���M+O>��A_��� R�Aw�wbY����?���|R���M��O�T~;Э	�gܹ)��}�t��5��B]��?IwN#��<����?����?Iq���L@,��5W��b4����?Q����WӦ��e�ӟ���ٟ<�O���x���^)��S���M� @��'��G�>y���?�L>�O�}�R��T�h����i�hy��^!+�2(c��4?��i>1���'��@'��3儐'xòĐub�N�(DKA����Iݟ��	�b>��'�07-��U,����ɆxT�5����1)��H��"�O��D⦵'�<�ɰ��$�ON$�tO
a�1�fY��0 ��O��dY	3�`6m??�;L�89��'\��:v��ڲ��)e��܁���<zb����$�O`�D�O<���O��D�|�V��U��{E/<8� ϖ�q뛶�Lbj�'�����'G�7=�T��g�b垡�"d�!V^�H�"O�O���9���a�7-��#�AW C �y�6k��F���C�{� 2�ْm��d!�D�<Q��?ц���פ��7��#Ɉ����B�?��?���$J��њ�$�����	�!��N�b��6,�y��c Y��՟<��O��D�O��OJ̐�AЖ}L�	s�"�~�BX����"�6�R�lھ��'!l��	ɟ4�1/�p�D9OZ��SR��ҟ���ş��I�LD��w����L �'6�"q�S eOf�!t�'�x6��	r%����O�n��ӟ���$���ԲH�4�d(��=�:���,���P�Q�ަe�u�-��<��TJd���C��>��M��a��$�T�''b�'�"�'�'bX��@��"�����ZO�`�W��޴vv�|����?�����<I�H�R�`�W�. �Bb�ʸ���П��?�|R��N�J�@c Σ��6)�E{�PC`���$ؤv����R7ҒO ˓WW�YY'�#f�cr�ccr����?���?��|�)O��m��a@Ĭ��)G�T�I� W�9�Q!c���^������M��'�>������9���b�"o��}�b	N�I^r�BClsӺ�8yJyiQ.埰X�I~*�;��,S*�-���*�۟q*͓�?���?����?�����O��a�S��6Iv`�;3&\)!�'�B�'>j7M�-$��O2yn�M�I�'���+Wޜw�  �@�h "�&���IƟ�ӿK�p�o�F~Zw�؄�獏.
$� y:�e܍~�B��B�IMy��'A"�' �MB�jͲ�y1ʆ�h���c���'��ɳ�Mk�
5�?9���?�/�"I���NR�9cU$�yf��ך�Z�O��$�O��O�S�M����⚽uZ��W�M�~4mلi������_y�Ov��I6�'����D�*������:wk�`K1�'a��'����O��I��M��VE�H�,��`%���q�\��p���?a�i<�O���'8�lȼ]�&�Z�Z���@�*�<BNb�'�A�i��i��[�O��?)@7^����	�Gmd��4k�w7搊(o�(�'=�'���'���'�哱|
�ph��
�H%*Xh�$�$00�;�4xp8X����?I�����<!Ǵ�y��=
7�����+ U�A*c/ʨXIr�']ɧ�O�2�i��$$�^ٚA�@"A�p��eˀbA󤕭4$$L��.[$�O ʓ�?!��Z�y�'aNɸ��(f^A���?��M����ߦ�Aeo�韜�	㟰k&�C�*�!�t'@�`	WjXz���I� ��B�)� �(9�a]>r#�|R�B

xęXp�������%7���1��K��!6����ٟ8��+�([���w/T5z\^��KFџD��͟������D���'����'Z/�&���Ә�ش��'D�7�z�nÛ�4����ъ�dU �*��_�K��-�34O���O��S,�6�4?��`�%g����F+s�^EC"�K;%'N���M$15�8O>�)O���O����O���O���ۣ.(�D���Qe@�<�A�iz�i��',�'��y2Ň�
��%I�0��j��F�3v��?1����Ş*9.1%��_��ei���&8��a�B�5"�T�'q�5òe3TE��h�̜��pY�!(0�a㕅H�����F��cDb�3�+�;7$�õ���z`����E>�z��#Ɵ'j�"�
ġ�W,�4rc,�%v�)6���N����4N�i������dMz��3[�l�;F`M">�#HT�m���Uϖ�a�́�b���lU:�i6S��E:Ӡ�X���  ��0Z^�9B�A�[�(�b���%{P��"0T%Y��&����S��&dV@1\��bb�N�B�R����G�k�@#5�/,��K��H�a���E�)n��#��Eڌ��4C�΁�&�
�4Q�h�K	" l�hֵi������$�������R�/r?Q�� �hF*!�2�Ϭ:J���c�Q}R�'DB�'�I�Uqd\���4�� �n���SjL�����j�,E� Yo�ԟ�&�D��ԟ��'	�RܓIR����P�H������=l;x�nZ����CyB [�A�맅?���J��4I�q��o�!�h,K�����'	��'����' ��It,.�B�S�P��e�>[f��^�x��(E��M[���?����f\��ثW?�t32��<y�A�E�%8�7��O$�������}"Ccڰ|3�ԋ�i�	&�U�AD����M�>�M����?����Q_���'�M��3R�T�Kpk�2
�2Qn�԰���O��Ox�?�	 `�΀.m¤S�K�F�yx�j��Y�Iٟp�	�>�Pͩ�O�ʓ�?��'��$)ԩBkHU ��q'@	A�4��_i��[���T�'���'E"����"�F| q�M�w�Y�b�"���%���'*�Iӟ�'��X�
a�@��EZ:����!�ǘ<f��X��Iy����$�O���O�˓t�6�
�{��C�fҊ|�:Y���� p�I{yR�'9�'�B�'p] �܎G\ Y�
y��JG�D2��'�B�'��U�PY�	?��T"C�E�B��N�1 ����C(�.�M�-O��*���O��d�"p��L��%B�Ar�v�T&J�Y��?Y���?�(O2��PN�$�'��0�E,���ӓJ� Dh&�i�fj���9�d�O �I�=B�"}2�ӗ�*�jض[یEꣁ���Ms��?�.O^���A���'�r�O���M«LJ]P2�Y(_ގ�`�.�D�O��$�-/M��T�'^�t�cӔ$�<��͇"Q�j9n�Tyb���m�7m�O��$�O\�Ɉb}Zc����g@�(N،	�G�)BCd���4�?�  �*��i	�8�j!q�DђPGݵ5��,ӄ#�H7m�O����O����i}�^� ѷ	D#d%�9;@��cx�Z����M� ų��'��D��2u�FXz� ����4�G��f�PmZ͟`�	ߟ�(��̢���|2��~*W�2C��f&O ?�<�H� 	�M�������s���p�	�2�J}q��ε#�^�xc�0:$�ܴ�?9$m��hl���t�'��'^�'�^#T�b�n߱G6�l�ǌ$�$�O6��?!���?�(OD�����]V\�Fl֣Ws\����d$���	ɟ%����u��P�sd�;�Ǝ�I�Œ��0�M������O��O�˓P��QQ�?��t��L��y�`$�B�2Em\�rUX���IƟ$&�̗��$�'Ԑ%h�`�2^)�1���D
�y�td�>���?A����I� =v�%>5��l�1k�V�BE�^�Rl`jI�M3�����4���&���.(
�A�?���e���Ms���?�/O>�t�K��ܟ<�s�� �MĄ>��]!�_w�P8�%��<����?�L~�Ӻ��E�%Ä�	q�ùV,� ���¦��'�k��`�&,�O@��Oe�Q�jQQ"J4X�����"kʕnmy��'P��4��;��i��ґ(D>�4�3�,�0Xrrٱ�4\���h0�i�"�'w��O�@O�	�8U�D�p	�	pFȢ�J�,G�mZܟ��	l%���<���,Q0�J�a�%D?�K�&c����i���'#b��2x�O���OR�I� @��d�`�.�����1R�7m�On�O�!���d�O���*9 �s ,d�$���+D�7-�O�)��<FX?9�?���"�p�@	��{~R�[�N@��'Y��O��D�ON�D�<�"��'�����$
�3��tbш[�&alT:��x��'B�|�R��ݚC��y0	\�+ ��җ.��2T�6��Op�O��ĸ<	��U����O��XƤ�CZ�(Z�)԰Iifm�ߴ�?!����'e�\��ZPa�T����h������F�.�Xij�x��'k�	�d�v��T�t�'���p�ÿ U<�Ze���|��``Ke������]y�/A�ē\����˟-���XF$��gOb�l�۟��'�G�[_�S۟8�I�?�X�"X�C��3�+��Ls�HOd�D�<��.�`��uWD�8'&4�7o�}b~����Q�M/OڼIዎզmQ������8U�'���H�&��u��Y 0[��ͩٴ���O���KM�SE�s�� t��R��bl(c`]���t�i��Ca�'#�'���O�)�D���KA-�	%�zPS���8h:���>�#<E��_�����v�Z�A1�@{&��Gfp6��O:�=��<:+O��N���Y(h<2���+�楩�kПo� Fx"#��O���Of�ȅ��Q��� *Or�Cvc�����I�{� [M<ͧ�?N>I��X�:�1�NY/.��K��:ǉ'rB�|��'<�	ݟ����,���각U�-��nY�S[�D�'���'��O��$��`Z��cm��0&��=V�<���dq�������	ԟ��	[yRk�����Nd9�2i��xFi���K�1���?������4���d��m.�]�čh�d�����k.2�&��	ty��'���7[>�ɿK�&�Ґ&g�J�"r��?".�I0�4��'�^�Dمh(�$
n8���̞
b��R����H �F�'�BQ� �����ħ�?������-\� W-�
9�HaǠ�a�	^y��'L2����ugB�_�>�ڑ���K�O) ��'�§F�D��'���'��TP���9|:0c6H8N��r�"K�e��6m�O�k��DxJ|B�i��`
Jup�F�h6U����Ԧ��#j��M���?�����Q�l�'�<H*��0U0�i�0��&Ip��eb�0��19Od�D�<�����'|�$ٗ��j1�E"����#��d��gb�:�$�O8�DZ}s
A�'1���X��BA��E�z����3��L�R�nZ� �'�h@������O����O@A���%;J5�`dϡQ.��J�����9�I��"�O���?�,O���ƺbNQ�Ti Q��A�H�^|�sP����d�X�	ܟT��۟|��eyB�&J8�:Y�yy�@��8���޾J������O�˓�?q���?��	I:�	�f�#\�Ā�@(��{�L�<���?	���D8U�>��'���R�|�
;3��hr�5oyB�'�I��D�I������~j�B՛W�tq9�+�47��@g����	����	؟|�'�}��#�~���To
=S��i�@q��_ r�@�#�i�\���I韨�ɕ��������J���E"G�Ԓw�m��hl�ܟ$��@yǏ=B�꧅?I��ZR ̵��y�.�+ ���0`͇�K�	�����x`#"q����@yBٟ\0#��O <�u�@��5	��=�ie��x�M3ݴ�?i���?y����i��W��^9�)�6�Ϸ;���+!ol����O�Q�0O���y��׼l h91�^�O �\1A.��g����R�-�@7��OZ���O���h}bR��amF�7�( P��ٶGhݩ���M�#��<�����6�S�� z�ܓv4\[���C��As`� �M����?Y��(ۓZ�\�'y��OZ�q�g�2I��[�:t�sP�0�'ޚ A�O�I�O����O���]<�XD����(hA��DǦ��	�w u	�O\ʓ�?q*O^���J�x0n��f��;�@���L}�^��90�v�p��̟��Iן��IGyr㐍d7�t�F��/M7��ACeT:}!�UA���>�)O����<����?	��D�~(85�@"�A�C��T;�%a���<����?����?�,��$B#XHH�Χ<���@��`���"F'O�,���nCy2�'j�Ißt���l���,p�g5��-锃#Z6֤��M���?���?�+O���R��m���'�X(g ӱc�4D��b9:�x1B~����<���?1������465pi�e����q�`��5�m�����	xy� �P��'�?���B���!�����B#^��} �4h�Iԟ��I��x�w�b�d�Ox�֟ ���TLp��iO'Ct���i�����I�ݦ	��������?���O�nG<|f�yH�Jɪ.{E�e�,��'�g���y��'��Wܧe��X�,U�eH}a�G���nڰ%(��Qߴ�?���?���B���|y��a���)&��)2�pYeCJ.
U 6MS�!��$�Ohʓ��Olb
ο{yEr�j8�4`��ń6�OJ�d�OIq`B}�Z���	|?��K��3�/�~��| �i�����I�������6�)����?���4oB��B�*5��т�JW�l�0�S�i�"�گZ(P���d�Ovʓ�?��B�����,_�C�,5�q�N��Ό�'�l���O����O(���O��cI60�G�%E�N�J��I
��9O���I`yb�'�	�����ٟ`���=J'�D�R!�n�*0h߆KD�	��	���Im��'��7a>AAq�^����# <m$��&-b����?�+O����O��D�V����b���A��0-�5��Tn�7��O@���O��<	�C����ٟP�c�%=� �	�JM	C̆�#���M�����O,���Oшc3O�����$���.p����m�3f�Б��x�X���O�˓g�T�:TS?U�	�\����`�v ف-l~��"#U0��s�O�d�O����~T�d�|���DI��)8�)"�jM#'��A�`G��M�-O��D��Ʀy���,�	�?˨O��ך��� P'�>�����x���'"�O�>5%V;��{1��j�����"sӤTq��ئ���ퟤ���?��O~˓5�b���DˑT����#j��@��vlW��y��'�R�'��.�D��Z�Z��%�	~Cbv�N�r+ xoݟ��	̟��dH���$�<a���~r��=�~�����Z�qe��M�����$B�|��?�I՟x�g�? �lpn�+,���!��!��*��iO� ɧ~�������O���?�1�Ph�c���*hy���@���'�<Ez�'���'_��'B�]�x�#-��N,�ɗE� 24y�whƼ8� l�O���?A(O����O&�D��y� �w/���]㲂D�Xt&kD;Oʓ�?	��?(O�P�Wg_�|�򁘼0��À�ߝs�x3��i}�'�|�'��ȗ?�yLc�0�X��(<�d��&_�_j듞?����?�*O��Z��V�S=L���* ��[�ܑ�A�ѩo����4�?�I>���?�C ӵ�?1M��h����q�޴��AE+nh�Dgnӂ��O0ʓ�0����4�'���|�0�7B�@�`�s���i��O����O�82�,�ON�O��Ӥ(Z�5 ȍ
�4�k5NA6-�7m�<1wf�	�f�~���*������%�
���5��%/���nӺ���OFu�F�O�Od�>�C�̅�R~�#�lZ�[��@�~� MiC��u��֟ �	�?]�M<)��d.�1q��?,[ր�����5�ſil����'y�''�j�$�9>@�)E*S�GG:�
��Q��* m؟`�I�܂ƅP����?���~��٩w z�*_Gx05ɷ/\��MM>A��<�OL2�'!b��4}I�����
2����"I�}��6M�OP$Sf]�	ҟ$��Z�i�e(-��-���b�P)�4"�h�>i��<A)O����O����`�F>Vɦɘ��H7R�|i��çj��>������?���_������Jj�G5J��!y���<A(O"�D�O��$�<a�-W�cc�ɇ z�� ���;Z��Cg��N'�Iٟ\�I~�	ٟX�ɮw9>t���B��l��F�~,J-SBE_�oV(�O���O��d�<����I�O��03�I��3��d��5���ѵ�'�ґ|��'��,��y��>I��H�AZ*MPw�ݯ|[ H���ۦ%�	蟴�'�V r��/�)�OR��J�B��a�����ұł3�"�%����ş ���8&�@��V�"���;0)P}b�<8�mDy�I��C��6-JY��'��.?�u.!�ʜ����>�ѐoHئ��	ٟ�u\ǟ%�<�}r�+��}X�֩��w���{R�����O��Ms��?�����@�Ę
�zH��ӹ`�[r+A�a��o��5�p�Ia�	O�'�?p`�'Hh�RR�A%d��^+���mߟ,��ӟ,���R��ē�?Q��~�V��
�ɂ���>ܼ5���M�O>��g�<�OR�'a�]�x���B�u��0�)�W��6-�OE`�.b��?H>��\6T�2,��A��i��.9�=�'8����'�֟��	Ɵ0�	��l�s�Y-y����*����g�]3?u�����������m�����ź0� �V�����Z3��m�'����?i���?1(ON��M��|�c���t �����h�Ƅ�#(i}��'G�'0�O�d��_?e[t�@q�q&n5�Ɛ��K�>y���?����?1�G�<���?���"�5���ɠF���W�K:I,��P�i>��|r�'?�I �,Oh����.rmh\��k�%+�D���i���'����0JIw�ҟ���,o~zÇ,O*�E����m�9H<����?��Ko�'m���$#���fB�;~� [) �vT��"��X��M�P?a���?E��Oh���K�8��Q�B�:"|.�1A�i��'�}���*v�lY@����s4z�b��@�1D.6m	�)=lʟ|�IџL���'��v��.y�� ���>7��'�צ��2 '���O6B/-hA�	��B�N�k�D��+\7��O:�d�O�AJee\k�I����|?�	�P}8�J�O�m�*����c�M�Z�<Q��?��&��$b�L,`�i��1��40иi�Lߪ55<b����I�i���F��V� �:�MݴP��{E��>qDÔ^��?���?�*O8�Àdj��A)AI9n��؃̌�IF�$�������&������(�!U�a嬌��mǺob��P�-^c���ן��Hy�C�,���=|V��U�V��Cs����ꓱ?a�����?i��Y���'�j �&2D�8m��j]�j��T�O�$�O:���<�!aV�9҉OHY�4����dX�R5P�4��o�$��<�$�O&����x^�O�,"eB�R��M��'?4��ķi���'2�'.�QdZ>U�'��D��,#��]`�a��-А�AF6.$�O"���<���T��u'��l|�1*�mТ9$ps�I��M�(O��� O��	ß ���?�r�OkLN�	���HU��[д�(�Α��'�B�'�>�q�A�j*V6D�l �hݴz�\����?����?��'�?���򉎓q�̭�#�N�z���:���2qʰ<�'��)@���i�OF��c��m�L������$�!��Ʀ-�I����>RrX���I�O�ia���VN�'��#�:-�� ���O��'>=�������#$K��L'/����C��C�2���4�y�n?np�'&��'�ɧ5�/Ԏ'��Srg^*E���S�N���On���O0��<ٲՐq̶���=6�Q�[�9��	���D�O�O��d��<�mԶYyVy�-&F�(thtc1���������'V�`�q>� 䵙ר�!+#DQ{�K� z%&U�L��۟$�H��۟0Xg�>��G�� ��h"���d����GUl}��'qr�'��	]j&p�N|�b#�	���c���N��1+�#Z��&�'_�'�2�'�� }�&��A��}궬T�s�AH�n��M+���?����?QՉ��)�<Q�'Q��}"��%H�N�w�3�Z��Аx"�'#�ɾAS�"<��K,�S&̆�.Rn!c .V&A�LnZay�ǝ�qn47��d�T�'��d)3?�g�Q
k�e1�D-0�6���cIZ��,C�Ri�?�g�9,~@i�]�"Ҧm��`IV�6�51�H�D�Oʓ��-O�.?� ��,Y�`�����D�PX�T�4��3�Ş�?)��@;P<�q�(1`���� �:��F�'32�'�H���(1�I��x������ A9J%!��C+tVU�>��&�I̓�?A���?�®��$��M�LC�>$��ЅچH���'ۦ� �'���'��X#!q@�طv�8�����g�%V��?����?���?��ƚ�*��l�u�Q m@5����Dȭ9*O����O���*���O����z�pe��Pq��rE�h=$��4q����'Z��'�bU�P�Q(���HK�K��T�W�N  �4�A�י����O����O���{7b�~ZDK_*-�01���hp�'�A}��'d��'q��'N�zQW>���<{��p�!�?:�}8�O�\�.�m�͟d'�X��Myb��ēs�6]�I�	dM:�	%�1em��h�	gy��0cs(���D��] �K&K���U,�J� �`'I�L�	���	*5��"<�O��4�h��Y͑a��=��9�4��d�Llښ��i�O��iD~� K>n� 9���G ؚ��%�M����?1�L�'�q�TՈq$�)7�؉�t.	��4a��i��Y8%iy�t�D�Ov�$�� '���	�#%j�3!����ԂcON�t�t���44-"�Fx����O��j�Qj]� `ծJ#"��`l���	ퟠ�I�81��M<Q��?��'�KS�ʳk������[�'z��B�}�l��':��'�",�tg��c򯁳�-2�i��wL<7��O�\J���b��?!J>��~�0�K��d���WfY��:��'|�T�y��'h�'��	=+�)��튫u�j���)PX�ß����?���䓐?���6��������I�xZp�Lc.�����H��?A��?�,O�䃵���|�Uj�*a��qCe�94Π����\}��'rr�|��'s2������C�
��`��D��٨�끵C��֟t��؟�'�8I��>�7X�q��o׭IV�� άk�.�n러&�X�I� jd#'�ɎY+���ȟd:���7z:7M�OV�d�<��b��aF�̟��	�?�(���?A��
���faZȡ$[�����O��d�O�H!��vrJ��eNa����j�0�ʴ.Dݦ-�'�����t��d�OL�$��B�֧u�	�
x�za2g�����UeR5�M[���?ɂ$��<�����d<4٢��V�.*���D�/�6���j���n����ퟴ�����ĩ<a����a�܄(Wƍ�5�Xd���y���	�y��'�	p�'�?Q���'`:�*�A��(�n]\���'.2�'ݴ�B�>))Ox�d���b�h�*foZqW���֝�����<9T�V�<�O���'a�h�����эH
��ƪɺ:��6�OR�xI{}"Z� �Ixy2��5��F�O��4˳GZ'q�d�BC���M#�&P�i��?a���?1��?I(OR�ȗeՐ+�cZ5sI����'�PX� �'��	�� �'���'RBM�0�N�qCkɂbɂ)��.c��y��'���'���'��'�ᘢc����8�lCKۻ`�j�K�N�B\�7��<������?�/OF����i�f�	̔n�lB��	�t��O����O��d�<�Ϝ�9K�O�F�:��a�%�Fh����K1Iy���D�O
㟐��8���k�*��AK�N L0Z��۱ &�7�O����M���s:�X�.��d�O��Y%Ę�#���N�ҕP���0D���'���	_y2c���O��M�	�ֽ��蟚W3�c�Ɂ/ț&Q�\He"��M[�\?A���?���Op����3}�x�䡃.F5��Ӵ�ib�'Z�T����)�?.4c�����Jl�%v����f36-�O����O �iYB�I����
��O9F����YR�:BdĖ�M����F���6�ߧ;J��T����Q���ꆶi3r�'nr�K1%�O����Oj�i3�`�F��f��H��Z��"��>y�e�b��?����?���Ȏ/�6Ik�`�$<���R�7���'�$q�k"���Oh�4���Hm�ӎ�y af�[?z��v_�|c7�1�ɤ �LY�?i���2��`c�5rV8I�Ꝺ�yr��G�l � �Z�z�ϛ=��O$��@����QP+ԨP���#C�ϻ��ڀ$]�Tpa�F��D<-)��ȥ|��逇a p��@ї(�V�!V�4���Ň�p���q�ǻ+e(�&Z<rz<��M��g����T�*[�uCf�ö���L�gX�ZR�+]%и���ߑT�x�"��٠���g=/<�0s6��9䭪���O���O
<��d�M,��C��<Јzu�����@�n��@�D�R���N_�(OT�S!ͣ~
��R*�D��8c׮��4J� $�Ò�a����LQ|�����	!Xmj���O��?���a��+�����B����sw�Ї�I�r549���;5dqÀv ���Td�I)+�ܙgg_����*V�qG�I�m?��h�O�D�|Jdˆ:�?I���?��л]��1A��J9T�L�9!.��!�m���
�j6HY�$�*��b>�d�?qx��PI�������ކxԆ�j�ڣ:�N�ɰl�*�2��)��ԣ���"�z�R5�M����N�iNl��	៬��'��f�@��sK^� c��^*q�ȓn�a��P|�hĄo�N�Dxb$�S��bXCк����T��$�1�y��')��ɏ��'���'��ם�����S�B�#���NCth	���(1��p�:.�=��BC��:௣?�=�V�P	�nq�G+�.��9�I�["�Mێё��JQ�l��g�'�@k�G��v����%^v֌�Z�'Eʵ����?9����<��� �cڔ�!�Ly��I}�<�Q�
I�mK5���|��ei�A�dꑞ����ˊ|��PnZ:l� �%�3+D̲w���<f����(�����Snv>����ȒeiE��f��	�Pv8���K��4B3F��d��*'�4昕w��MA�Ävq�P⑃1fJ��Y�oU&Q�L�$�'��1���?ɶ��'W��a�#Ms���"%O��?q�����O<��<;��2��5J\ "��+6�蹅ȓ]��Uz -�=oMzT���D*-�r�x��'eўP$��6�p���A4D(6]a�� D�\#�Aܸ>|����=O��+D�(I�.Ŏ_0<��B$�:��d/D�H[I�����W�zh�kѩ�;�yb���^t��+�m�u]��@��Œ�yB`T�:x2�` �?f"Z3%��ybɞ�g�ju�%�D [.�����J��y���\DB�6Y��H�+=�y��K���ԎڵO0R�����y�C��MP`E��CD�[B���U��y�S�K�t閍Hbw�����ܝ�y�֚}:8h)S��jwX�B�G��y�I�+`A8�JU[� =8�R��y��74�x�J�0^2@}�T�X��yR�Yzަ��IP�WwP=h$�&�y�,��FܘI�4,MݔMX��4�y����.�y���ѫB�)�G���y���~��s����F@�	Ѓ�V��y�H��|��M��ǔ�:{�L�b�]��yR�5h�؈ l+}�؋���yb(����f�x�5����y��9f��G�@�<U��90e=�y�$��h�8���A��E�j�j0�yrV8S02��4
�&?�D`p���+�yR�Ջ#���6DF3bJ��6gC8�ye͜'�U�s䖡p
�}�Ձ��yBd�j� Prg��j=<�*�h��yR�L}8t���� x��J4� 7�y�j����Iw�Ē%{�|qD�R��yRݒP�
4��͇�KA�!�D��yb�ɝ	�´ �ō�J��\�c��y��ϛ{˾��sj��r16� ϔ:�y��K�sY��T.� ��TQ ! �y�͉�Hj�u�3!�.|���&��yO�/�<8�Ǭ�[T)6�/�yn�(t��j� ~�x\��[,�y��){��`(�!u"I{�F^��yB&U�*�䩡��r�r�����yLޜC>����+�$��r�b���y����4�p�$�՞|�H{�1�y�K�,/1\�S��;=�>�z�A8��O�X �"�3}RM�4baP��(��3���	2�����x�7R㰽8��ZOܚ�b�8U��Yc��I؟� PP�i��C[��b�����c��'S􀺕b�J�I�u�I���?(���j4�B�2�P�t�צ����@cիo;d�A/M�����|�/L���=�}B�
L�e������X3d���$	3 �����8�g?���ؑ{:�ͱ���s�U���*;EqO����`4�s���ٓ:�^$��
4��)���tn ����&�Lk8�$���E�����=bn���k'�|@�������4fs��8sW>U�*R�Sn2�Ӽzb��&<O~1rUҾ��h�u#��O.JF݊T�H�cr�x�ywb1��W�~O����1��<�՟��3� y!����S=mq�Y���|BR?iy�y�=�|څ/�?Z�������|�\�3�H�y�J\2
l�I�gȷ;��D0/�=���ҫ8 7�Eb�!��h��@ht�	1�z�zg�Z�D�B_��ԟ�!�'DV�_��)
��-9: v,�{Jtչ���D)����I%W���Y�	pH �ƅ|��E��_���B <>��?��@?���Y�|z��N>�إ�bgW��@``��Nx����g	S��'���٦�!
�������T�E��'�q`Ee_%:�6��+bo���@=@��r>!I��S�5a`��#���_rx`r��$�䎏[zh@2�{��d��*L�@{v�3Qy��beAR�k��$
�c�nS�-R4�����.D���^=_�@`d���;�R<�W���3����O��8�_��'��)�O�<��ϖ,,�`aↇfB(`���L�	�x\��	$$fh &�Dx�|�1\�輩�DӦ`q�H ��P�p�D�|�T�����O����'�{x�ޥUcd�r��I�^�|*ac6K���RbE�1HA2�b`[p�'-|➜C�`Z�|��Jɓ,x�`�Ȣ5>��u�myB�H�O>�.9a5���_�^Š��v��<Q�����t���?�I&H�#���q�TD�t���Q1ODd����:*1O��1�=��D8B@��3<��K3OP��c�OF���H j�,5q.$A1i�O�4dp�	Jv�5��9F� V&�"��1B�Y@=��E�Y��(���j1 �����'KM?
C�	�b���a'�$P�qX`C�H�ʓS�P�Gx����l��1����uNh��N��|���� �g}�䃇��=���ȵ-k2D��
���)c��4Y�'4�!B��_9Dh�5���Bbm�#�Ti��<�x#i_�l�n�Rwʧ�yu�B��Op�I?�va&?�^<�띄=q ���ވc�<�$���v7t	9�Bh��Fyr�Ϫ�(��,{�LJ�W-i���ȠI�H�GȰA���'�lh��T�}�ɋV4��ߴ���P���g�89�Ӂ�2<$�zwǫ<�ddNE��u�4"��'U�t�gb\�:a(�AMF���Z���S1~��	lZ#��dj$n:�f#�ɮ&�@$��AL�i/<t��K�]B(�O,Tm��'�,U�b�[����	�9��Qm�2�l��揪p�b�]�PUfl"���������O���R1>�T��d�*e*��P������<�T��?; ����[*ʆ�V�Z�ɐ{"<$x�
S�l{ ]�`\u���#�S�w,�X
t�$�':}B��p
,*!�e ���2V����/��M'����O&A���F{����l0k,�=9�hY�k_�(H
��o�1�xq�'�� i���6@z�2́�&�"��ddSe6b�E{���Dèq$��H�0ېO���~rGQ�^�hYP�G�6�3�����&�'� Ҷ���\�*MZc7J}�)H��I����DK��`�wƊw\�D̏4��Tb�?w`�z��2�O�=�!�6ZM�D���D�l(�YL?9�m��LS[K��Î��P�u�k�֦i�`oi�'6�����pP��<_�f*fў�*�Fx�bZ'�(����gG�!�\Ш���F).D÷IѪJ�v���y�AD}��R<��j}�dJc�^��T12�ޱ$剟gh#<��S�ͳq �3"0*�Jg٭;�>	�WG�v���:6@�E�'���[r�^����S��M=%���'���ׄh�P��t�L��K>&�tk���"��x��L�Pi�(!�yC��<k��e��h��K.H�K��Q&�?Q�F�~���E�D�d�d�c�a�'t�Ya��'S�
L��#
?Y�H�+�}k�}1���Z�"�3핤n0r�ٳ�Z
M��+��I'����m�����m��"�I.zψ�Ӓ��=)a�#<�V�@��x�Q�D�(�����0,e%ؓ��
t��0)	/!yQ�����м���<U2śS���g�<�p���M�<����U���
�j�) ��u�B�#.3Z��ag�R�I�3�
�鴍��f�r��Z���ɡ|Q��Iqb�3}T��s	*��#<�Fi��#9"頕�ܒ:��XA�HԆ�9�'�I7t���1Rx쁐6 
]� ���
�!��()�"��q�/	�t�>�����#B���m����V���{�lq÷B�B4�����Q�,U
Y���%Xc��!F���-=���'p� �U��C�z�!�!B�!� /�l���)� @!@��=q�dq9T�	>t�f��1"Tq���L�g}�Bun88��O��o`�5�3�&֭J�#�%\t�����<�O.��.@,��w��p��S�D��H*"�Y��$,JJ��DY	~�`M3���2TE���	����Sg�hSM�u��E($/O�*���*R��<o^-�� �(+�D�T@N���iŐo�8,�q�X���a��*O=��ӂ_��$�5�9F�����kհ��O�Z���	��p ��Kc�T`4ٜE�ܽ!�;g� y�2�]%��X�O\9�ۅ��D=L�2���o�2.�0�ABV76~l���#�J~�~bg�C��,@ �z��X��L#�Y2�H���B"�,�P" ?AZ4��ɒO��;�\Q�.̿9ͤ2P������I=*��u��F�7TX|b���v'�M�rG85!��[���'��D�=\aԅZn�"v����ͩ1��X}�#!�v�aRaE�-f�Y)�E��0<	���j��O�@C�!l`(�����0vFt��"OR0����T`��ߺ	W�y�&����`!ʏ�qO>� ��Y�o,�x*�MQ�!� ���$D��
��}L��Pul��@N��)�B$扈 �L�+��'���+ܻx��3%N�(���'��ł�s>xͱ��N��J��!�
P�,��j�|� "�5c  4�M�c(����	0y@�@��$
�!ܸ�9�)T�)e��A!������ЭˈR\�Pv���m2�Q������	E�{�n�jE鐜W�H�pd"��!�DҸG�!�!�ϢF�ӄԀk�qO�h@�� ڡ�ΠB�0�H�`"��T��Z� 4?�����4D�p�����V�xQ��5�Q�6�/}r�C5Dc2��m�]>ջuGǐ7�٢C옋gH�����!D������K�v��U���e�>�)Ag@�y�~�'ð]
ӂ�B�g�4� 3fǞ��4��1o�"�C�I	W�����0�l��w'NjR�Ô��UelJ�'�$�tfA�,�L�B �P>%ʖ`�˓FQ๚ ��xB�I"G�:E��֊L�ޙAQ͆�9R�C�ɡj�Q�Dn�_X��A���<)�C�3��@AUd��Rx"C$TVlC�	?0ȔC� w�����_a�B�ɛ(���@Kdj�!Q���V��C��5d��ڲOC�0��'��$p�C�I�E3�x�A��?���A�[w^B�+$f���:4��eKĎ\>:^C�I�r<$���i��}^=h�� �B�ɗ~hس�7L�tq�D��(Z��$8"�L�p<QF$�.�,!��'�)�dR g]b(<a��'!B����g6tG�Y `��#%.]R�
O@@�P�íY�m����TJ!���'�ND�6�+�K�<%s�(@��L��r�vB�	�H��M�6�F4�����Ȟ;���'` EA�0�)�S>�jlp3o�7f��[7�ޏ��B�	2HW�|�R*�N�r��W#�A����m���p<�' � ?Gڨh��ݮ�v��c�n(<Q�M��IP
�)�ӎ9^t�QG�U�Ajbi؄
O"�{���Oa@ gkȼv�Py��'W,�A� =�"i�$mӀ,1h��&lLn<C�	�$� �� ������r��X�'�mK��?�)�	$G����M׀�	D$J&}JC�Ɋ1�X;$IT36Z0�ʲbǽv 
c������0<��A�[���L	?m��� H�<����I8u�C���s/�tXRC�<y��P�>ЄPB�Dt� V'�I�<�IL>;�~ :F�K"$9ӏ�<�W"AP+�3t'Z&sN����Ra�<�`ԙd|�i�	�)`�ȪT�MU�<9�aOTq������]Q�4PX�<����A��`�+��Z�RR�<����= �h��$C���� `LP�<�1'���h����	b�`p�'��p�<i�)C�^��e���1�^���a�l�<� ��v.�:Bw�-{��p炉�3"OR����1�|������CǢ�ۓ"On8� �@�
��[A��{���&"O�%�r����A���Y��LБ�"O�	�׫Ȃp�:����t��2 "O�ٱ�y�~$�� JL�h!��"O$@��a� 4z,���ʓ }�)�W"O����DRn/����*\h�� �"O��Xt�����
�N[�1b�@ "O�x��
6�|�!�ڟ8���g"O��g"�%p7���|:��>D��
͋�F����8K��@��(�t�<�G�/I-�4`��Ϟ=�!�S��u�<��k�	Aw6ei!��47ƽ����H�<���͗tȢ�Ё�8h�(�0��JM�<��j�.+���	����K�b���!�M�<��"�2x�ֱC�&O0 0"�(���o�<�!n4o���(X!�~M*���n�<��$ߜ�j�'�b��lb�&V�<��-5�T�:���+�:��l�<Q��a��F�D|����t@�e�<)TBL�q8y�uN��O����c�<1��՞9�dP+`_#x�j�K��I�<Y���!�t`����(��`ˆIR_�<����y-���[�G���e)\^�<a��p���
 ��'b|C�E�[�<�VT$V��r�	�$c�m�~�<�#�E
xUC�e�#T_�����p�<��G�1w�4Q`!�B���Am�<Y�JA?%���KR&M�!9�Wg�<Ş5w�� �)R���\k��]�<���h�\�Zr���Y�����W�<�"ȃ�ԋ2jR�\j	�OX�<a�j��(�Z����\�Sϸ}3���R�<��!�2�( �2C��8k�L�<�6�3)��
Ǎ�4�๺Af�F�<S��f�8��'F�ͫRPD�<)����P_��;P�ˣ6-V`#�J_D�<�� ������Ĝ���(J@�<ab[=u��}��T���X�f/
D�<Q�J�#5bD�XAE�%� =�e��y�<��d���Hb�Fɛe�Sk�<���D�7�T���Iܨ�p�R�<����$(	���).�����|�<��&U�L�d�2�h��V�%0q�P�<�5 E/d.�d��Eš<�#�E�V�<q���/�D��bs�Uj��M�<9�d��JD�Q��.P����VF�<����QtD����?k2t"���g�<9�
]	Yǚa�,ս�ơ��i�a�<��N.�|��D�Ӕ2n�I��!U�<���T2�t]� ��p!��㉞T�<v���\�؇BގSEd
���D�<� ��2���I��ɇ_5����B�<���N�����UOҪ ��a'�X�<�`g��z_<1 )ΨtN�tq��R�<�QV O�v��7F�9�t�G-�Y�<q�� ]r���6 ��1��银� N�<ie�S�o�d��D.�0<�R)���Dn�<i�Z8tk��Q�Z�`�)�l�<1��,rӲ��D��"ff̸u&T�<��	ws�����3��l�!�e�<9D��9Z`�3�پM��S�Qg�<	�$ψD{*-J���P�jгӀNJ�<� &<�#�|��p�[0V\��"O��bG�er������
��0w"O��u�KL��z����M
�"O��q$H�$f��i1BԭV��4"O|\�پjM��*�#.�)��"ON�g�(S x�Ad�2϶%�U"OLqa��`Й�v�M9a�R�h�"O�ĺv�9AR�Q2!M�0o^D�S"O���mH=R�.�`@G�J�Q��"Old�� �3Ғ,��pyɒ�"Od=s�e�e���b�̌{��嫧"O�q��#Q��j�$Ѿu�h\��"ON��c7}\fБ���:��l�"O�h	��H0X���o�>L��q"Ox��^�f�t}9ǭR�|�N9@�"O�m�ԍӉ ��LtBB��,�k�"O�ô�
-
��թR�=��4��g�<�RM�k���˂x��2og�<��A@�bb��NiΎɛ�,b�<��ܗX�ѐÒM5f@2�Z�<���^W�����i`t��ǋ�Z�<�%�M�� ��S�-ڍ� S�<Y7ꊨqɦA�&*��| ���%��H�<ɡ�m��h3�΀���%#Z[�<��؏G�T���R'G�&A� hE\����<a�爚_�`� -�&Z���m�Z�<�&=l\��iB≤>�X���a�<�Wo!�b豖HK�z�<�ѣG�Z�<)��\8	8� a��*b ����U�<��nζa�B����k<<��b��|�<���6Pv��p�)U�S����� ^�<��%�V%��"^�1Hxѩ�X�<�C�B�)���(�ρ�WC
-:"�
S�<١ �~���Q��A��q��e�I�<�Q�1 ���rg�(]
� �`�<��T'e@!�E�[��h���a�<S`'��i)��P�����t�<Yb���f���iC
�"R��`A��p�<!���5w"Г�螢.�f��wjUA�<q��F7%�Ԡ�W�J�b��}�<q@)�4e�x|:�	�Pt�C!�v�<�8�������`�_~K^<��'�l)��W��x}���W%a�Fqp
�')�Q4S�3 �([@��0�$���d �)��Y�	\��#@Lޫb���ȓn�[�f�M7�ջ7˂�w�x�ȓ'�p9[w�I�_�[@��7ZX�ȓy�% %ߒ=�|�l
���A��e؂sM����ъŎ� 0����rߔ�H����0k��	�D�H���]����=r��p�/Z���
fvJV�F5_5�T�Āԟ_�2l��g�.	�e�/
(��k��DTټ݅�=`0��b��/k'ܕTg��X�d݅ȓ^��8���"H����+�b���b9��M@aFx��l�,�� ��2uB����o^����f��+�PI�ȓ5�� R���T�6$z�/�h�����|QJ)��Z*O�|)��e��$� p�ȓ�px��%�X�v��K.�ȓ!�z�Q6��0d�<_�X"�W�<) �@���ayѨ�&/�`Ɉ�(Sz�<�� ��`ig���+%�H��!}�<��+̮Y\�4����#L]�	q�$O�<� ��:�m��;�Jd���ưl�<ٚV"O�� e]�e�7�.-�܈"O��J�E_����
�n�`�04`0"O��٢iI5���ꆤ��̖͒!"O��#Aڤ%�4-�$d	�'��"�"OȤ��	@^*���qÚo�00
�"O�(�m�Q�H�4�V'p�h(6"O��$�/�:�#s �7k4 ��"O������xL�@F�dc�A3"O���� �`��)C�[&��	""O������5�p+�'>�S@"O�|C�Ʌ6'��\3c��&�}�F"Ote�훑B�J��E�e��9S"O �3��*�^��'Р��J�"ONhءI��p^�mI0R:lh䢁"Oj�z��2I����R�L6QA1"O������fR=�*�8\	E�"O���a��Ȱ�'��Pl�6"O0pA�b�" �e�W&�vs�� "O`8��*���2�/�ag��x�"O�����E2/k^t�֯K�vfl��"O 8��jX8l��(�D�E:uŘ��'"O�,�b�&Z��\r�a�钖"O\�	�Iі4U0Y�%�_�9�ի�"O�ث"���d�+�LU����x"O�L9d��h�ZGn"�-)e"O�1��*5zq��Mʨ3w^j�"OIyI
*�����X�F�sc"Oz(�V�C~	n�3�V-j�B�W"O�=���`S����
@�T"O�j#d�|4���0�v0��"O��*����ڈ�5F��tv��Z$"O��b�����k$D�;��%h�"Ob$����|��q1�bEjDj�X3�':�ɬ,���@��[�e�d���,��B�	E(�̡��Y.17�]3G��B�I������A��"Lh��'��!+�C�I>�J���iԁv�rQBFj� o�C�I�Jp����ϑV}����2x.�C�I�u��(�f���ڸ �IS)�C�ɐ�:h�à��!���#�L*�C䉏'���P&ˉ:@�8�u�����C�I�{�H�`��3A"�Əx��C�w�j��4D^�NDP��f�C�	$��t��N�4��  �>�JB䉢&�<� F�;%�=�K�>�zC��$S%�(�� ��8�<�.��H8vC�j�XcV ��R8)�U�9LXC�ɒ�慪��.U� =2aB���C��N�h�V����L{�f���C�I5"�h@U��
7��d�Ӫ�v��C䉆(N��N�+��[�� 6!|��%�ɲa㴐Zda�E�(J���'3CB�	�Gu�uW��2��"��
B+B�I�*=��f��+�^0)6�[�w�C䉯;}n<Q͈�	�Bp:� �\�vC䉨A
PLZt�ɝ�tB���aƴC��K��\JDl�
�ʝa��Q�5�TB�	���1IL�H+��YC*Z�=KRB�ɏ>��er����3���ԧ��_�xB�;5@؄���"P�^d;�@uC�I"6>j�I��ԉ=YD��Q�|��B�I�D||Fŉ�@ \��p��C�ɍ(�XLb�Rn�M�Eυ�.w�B�)� ��v%3�,�!-��p-��1`"O�XI��%V<0���u䨛�"O.ܱ���/y!
��W��M����"OjY@�*��`@� �R��ȍ��"O�T#�˕#Graj��j��U(�"O��3rd;[�F�FAV�2tk�"O�4�AF����� ���i�j�iP"O��[4���0�Ĩӌ��p�JS�"O��� ���H��T(�l	���h@"O�d �fX����b�,c�z8)�"O�m�WA�]MH`�˚���a4"O�a��O�V����G��8�$z�!�_0��Mؗ�hk3'�3k�!�ˮm�`j�d�z�Tv�9�!�� Wv&4��J_I����BfI	i~!���b�,J`#%�r�r'�ȄS�!��H0�ܱ�
�)��mk�ς��!���rQL�"5h��w�d�P`� �M!�$-���e�������x�'z&j޺+Yb!�����
���'����&��4\bŅ�%)T�
�'�8�b�iʝN� 1�(N�3C.4��'��,)�c\�J����K�,e8��':�`Z�">=�1#�[VY�X�'�L���,��g¾�"F�H��	�',���-܍n�S�� .�x�
�'�\Iɢ@��7ji�	��)i|)�
�'��|i�j��M�|���R.����	�'��;d�/5�
d�C߃����	�'����B딢R��x�7��X�"	�'ш�҆��g<6<�6�ƚ#HL��'<�˅CߞOxH���L��'���b�/ɒ���*��F�bh�'�d�S�B�}p!�F�1GZ�(�'�83a^����bb�߳(a&�P�'���tN�T:�L[A-R(��١�'9&���({��p�P�;b�}s�'I~��*�K3``H���&#VX�'��4J��� N����S�Ƭ
S�@	�'��X�daF�8ʔ�	��k��$R�'��(��H�|!�� B̞.b 
E��'���c��c|٩��9����'�\�퐪i�D�
l)g�RM�'� �9#���(ؑR�ג	�YR�'�H���#
�r,���qN݈z��D
�'��� �ּ ���YK�_���	�'�XC�Ř0��Da
��R��=X	�'=�|����\�����˃�K0�z�'5(�o
���D�5=��'�l��Ď�F�X@"�
�f۪�	�'e4�c�R�pzppקONĠ�)�'�p���Ҍ/g�r�%�7<�z�	�',��a�Z-]Z�Us$K74Ƒ��'<�����	0+I�)wmə'� ��
�'¾hE�K'\�h&�]-$a��'l���eh�u���|����'׬� ��;J~H���sz%��'S�� ��8(��E��cE9p�3�'贴	�
׈`��r5�ix�x�';hp�q�Y�@���(�ְ�	�'�i��۴��(�EƥP
�'���&�H|��7+��
�'�P1�cH�R���K���`��
�'����d��R��	:@=b��
���  Tۧ��9@pRD�G>]o<;�"O� (p��.�*��'�l���"O��a����A�/�;`d�G"O4ȓ5��mQ�e@���8E��s�"O�A��Y�?���1���7�hȚ�"O�ͻ��O���(Ĭ��"O���D)]���9F,D��$��"O��G�1tGT�A#*�SbP�ї"O�ܪ7�	�X�� ��^�]!"c"O&p���&o_�-k�L)i��"O�Hys��CǄ��� �UI m1`"O�Ț��e�й �T8��)"O�I+���!�����Z)3�"Ox,u�(mGTي2 �;u��j�"Of(Ro_�V�^� ��sj��"OL�肎��e��7�*���"Ol�W�
2����v�9�~!�"Oh���h�:.����]"	V��9�"O250�W�0bU)G䗸?M���"O�U��N�N"��fR
��B"O\��u#]�~Y���<'��a� "O:��nV�(1�2�B7L�z ("O�%�ɑ��@�V�L��u@D"O�h����~=BH�V	��F"z0��"O�<P��ϒ0��i�iݼH:V\1"O4��֎ܟz��=xq�W%v*�|��"O~�X�a̻Q�B�u�H�"4ȩ�"O&�� ��*��5�S)Q�zf4I��"OV���3'��Т� G.�{�"O�Q*�cF>����φ4E��a�"Ov]9��Ùh�����8����$�!��PG�Ua��O�q�I��A�+}!�˪�C$cN/MZY���K�Ud!�$N7K�h���G\KD�(hf�%c:!�$Q��a���)�i`A��"*!�D�.<L�2�)W�O�z�hg�7�!��=F��A�ʄ?l�I�iJ�U<!��H/Q�V�p�g�LԒL#�(��l$!��X4,ੌ�^������J�G�!��޿<��9���4T��;%���!��)ee�a���V?=E��&��!�D���R1��u5�A�G��2�!��Ɠ �� b�Z�@�P��$�: �!�DL�p\8�-nj���jW�!�d�>f9�L�W�	X9���$Q�!���;�*հr�pe���)�!�$������I�<��m�`M��Py2�x�F-�T�̺$ʠ����y�K����f+�ye���yb�]�[���qf� ORՃqO�8�yb�݂]���<jzT� �O�-p�
ņȓ=��d`��D9˘���]-M����ȓm�VD�W뇱�,�{ÌJ�W�n�ȓu���X�N�5�\ۑ�(zT歅��
���՞d���V���=�<��.���J('����J_'"��ej�
3��&P�r���%�g�8��=���j� �>] \ŃPAɆȓ]�ʔK���"QO*�����чȓ} U:%+ܤk y��|C�݅ȓX� �׎PG{X��i��G%���ȓb���u�Ő\� ���L��9�ȓ-v��Z��D�/lNՊ�Gʧ|R�\��m���M-�!z��Y�2d���S�? P��R.S�(������~�|Y�"O��[E������A�h�NLV�a"O���qk R�� N�x�+"O^U��`��~T�z���aت�r�"OڌIFD��V��S��g�> B"O�� �,ǃ7�\7'�z�I3B"OlxE*H#�V��f��3�p�w"O`iO�B-��1�Nެ��"O ����<c���+T�U��h�CS"O6pI�E?[^��Ѣ��`�I "O��K6�I/2#�i�!,�:k�8q"OP �E 5)�BͰ �A�&�a�"O���(�#n��	ޛ/��,��"O8�"*[
��iG
=+�X��"O䙁��V	P*�`��52b��@"O:٠��Q/H�<P��1M��=8�"O
ź��M�j��1�3�[K���	�"O�	`��Ԑ3ڱ��H���y�"OTɃc��̖� 7�7���X�"OV�N�*�\u'��E� "O̽���^O�t��E_9K، "O\�&�/w*�J1c�Stm1�"O� ��Y�^,�5�7�H�[j41�'�!��QS��`�A�� $x�n��!!�U�[��G\�����M�lj!�B�P�(���F ���b�F AF!�䛬޲!cbC��i�S��ɘ@!�D�=�����i�
��]�|�D��'�4l�B�\�}�"AS�c�*��	�'Y��?���a��.�|m��'`5R��`�hӗ��,{��O>a���I�(���R}�>��p�ZM!�䍀M< ��5��8����ܓXg!��Kw����_<ug�	(tM�:t�!��BM�)��fȏAl���ӛH!��[~��+C�g�z���&��IA��|y��� �T����J�zq�I�f�T�~�C�ɳ�^M�e�C5�� J"���/���gCzR��ƛ��`C��P�n�b�'��P�bA����K��S�B&����'&D�w�X:W.,-�Bb2B�@-��' �P�� �j��  ��R�8���p�'��8�e�P2$�V�a!��{���.O��=E���D�&�-J����H�ٶ	
=�䓡0>A�(BfؼYIS�h|�Z�CvyR��%�!��$�A�7Ƃ��F�-j��5���3���=�Ћ���I�e�ȓ"��!z���&� �6LS����ȓ�\i�B�T;<j��;b'�z����Z�rr@�@�>ŋBl�A�Dd�?!
ϓG���QF%.���f��й��Il̓O�͐p�W�u���6��$F{"�O\�؋�W� ,J�џa4�e*�'���7�̾T=\�)�a	VH�E��'ʾ�1��6�r��k��|]~�
�'��@R6�N�'��A1��BG&x�
�'Ғ�Q�`|���0KʭG$���'����3Eu2���!�&3xh��'i�i��_�Y����CW�����'j�����έ*�X�+"j��
��ܟ����i�Y1!C"%+������LJT��!�!�0nH�5��(�/ޚ{vq���`��j�0q98qS OM+�ޝ��Z�ܻ��D7iB�)�.ٽM��`��S�? �� �	E/r���	�&�6b��&"O��d:��0�yq��0�-��g���ʗ��J���Oӭp�:���#H I����P���TiW�L9�݄��:q9%�'D�T�2�e���U��Z*h�� -X����&�J0��W=ʵq�g�;*g�d�U�S:@l05'����(j'	�q�M����ϥA��C��n�����K�<)��\��HZPS ���.�	�0Y y3�N�
0�X��&�'��O~��� '��qz7f��i"V#�D��$�!�B �@r&oٜ}���!!�D�+G}B�j1+ݘD\�X�R�	!��}�x0�G�>_6E���B���'!a|ªJ8��ْ�\9V��N��?�
�'�JA*墕�<�l�P��֩��
K>y����'j1O��Wh\W�x@[�"'#�R"O���D�mM�,����>L0]J1"O
���R��y�vW�\� �P"O�,��,��C��\`�b[�\�
��"O�X�t�Т0�T��@۹*�~4��"O~� ��0x]�UAP�Ҿ{�fy{1"Ox��h�	 ���Be�Θ@���"Oޔ��" ;1��) 	<�"���"O��2`�^]�Ԋ҂ղ�t�7"O��tg+K�0ɓa�f����2"O�i��I������DKҧBä="O�I���0��Ł����H;t�D�O���̮qR�IƋ-�.)��+L�\9!�$�&f�0Xa.�u���م�[�!�D��p��y+�3%��1�F�#0!��~�n��Ԯ�kq�e���&x!���x�A���)ζ=�&�ޓqr!�D�D����X1�H|@(z�!�ʄF���0� y�`!B��٬E��y�I���af�H�ZG81���ɼIQ�C�	�����Sl�R4T�a��3{9J��D�O����O	9�4�9��4�q(���O��=E���Z*hT����K�;Wb��W��!���L�4�j�E�p$qB�i�5:�!�$_ %�\+4�]�/�@l�!jV��!��]b}x���y�\Tӕ��2o��	\x���'�<�*&��T��v�.�D)
�'|6�qr�@�j@�q��l�Uy��(O���$r�����3�9����P_�)��n D��cG��#Iu��HY1���6���y�ւ?M8�A��Q�D<!�B��yO� S�M�&I��m��%
S��	�y�cЁ @j�x���l2�m�b���=I���D��k���[�N7W���WD	9+�!�D�AG
�{bn��1�D�Xb�m@���'���Bg�(I��=(�'ޙ �XS�'�!�2r�Ξ4W�b��/'h!�$ȅq�II�%�	�6�A�&|!��8�B��&�ѯ>�0�����".c!�dɛ1�1�F��$6�x�y���PX!��J'��'&�*b�X��B�$nO�OҢ=��8�)&HM�0�Q�E�-LB|��%"O.�j���	/ւP�05b*�K�"O�P��U�8�ѩCJ�M�B �"OR���D� YvHaǁ �|E1'"OPa���L"~�V���S����"Op�d�G�6�d,�
e�:Ղ"OhE��Bƞkl������>��"O�  ���l_-Mr����Ǿ0�u��"O�u"�V�OP�p�`�Lc(¸KP�Ip����1}��Y �E�T p�H5D�(��˅�F^�e�	+�.ȱ�3D�p����4�-�m/5β��n<D��� ��"pꨚ�Ś�7�M*Ѝ-��0<����o�ȕ���U�;��"��}�<іM��D�p����2Θ�t�Iy�<	���R�A���VRr��"EHr���D;�l��d���˿YY�t�a%��%-� �ȓM.�����n{��p�H^�TQ��X�<MC�]:И@U��Q����M
"̹��, >�+��%kⶬ��#ܠ�z�j���L���֚xm��	�'h�Y�AO�Wb�j�-��i��q
�'�@s�Ƣ5M�9ڶ���b�*��'�j0鴫L�;�)鵍�:.C�A��'��p���-\{�4�E���l�s�'т���I&�(!P��CO.���'7��Q�� �v-�.�h*�����'u| b�R5_���
�aϖhX��J���'�a����1D��ReA�31�(�EH_(�y�K%����#C^<w��y����yҮP�-��)�f%I�Q|��8�ybE�)"]�yc�>���H3.���y�o�l`���P4y(�#ӯą�y�K߉K��CF�_�I'`@G�K=���0>2�0]�����@�\� Y�jUph<1�!��LV�i��*چG�Q�h���d3�O����IE�DH�Qr'�Ӿ��E�f"OJ}hq.���'�,p &da�"O���è�m�Z�
�dǏYx��C"O�%� ��ppG��Y#�HdO��#���l��+�,�,_�,ȸ5d2ړ��' �I�*��|8ţ��d���t!V��C�I1s������%T��QぴP��C�I{�Y�wJ�9`�ܽIs��&�$,�$�<E�T]
4%�#�B�!ʲ(°N˶w�!�d�)$���	�h��5��n�F�!�$�H�|��"��N�F�1��y����0����6�8"�I�1!��U*�y��ʄX �U�,�Y�!�J�S<m��A��� L�k�!�$�=��Ŧ��R��)3j؂+�!�䘁g>2�Ce�ƈqxT�[�G�(k{!��3=d��V��xvx�j2G��#x!�ʣ4� ���]q.x�T�T�gY!�$O-g����<Wg6�1A v�!�\�kH� ԄM�VtĠ���Zr!��_�T��Ȕ�22](!9��_!�d
d����v֝�ԏŇO!��
Z��E2Dջ*XD���_�?!�$Y��v��씀4b��A��L1 3!�3F�����O�9P�n�yTM�{!�$��j���P�"�4y����Г��O ����_ b9�s	^�+�QJ�)"�!�ҡO��0����$��m�q)N!��N�:�����.S� �A��=@U!�/7��x�TLL����KQ�0}9!�d��wd0�n���k ̚ %!�D[?)$=0 �f�l�4bC�h!���/;Еj�V">60`��v�ў���S� p��@�l�H`�D�ΘFx�C�)?�\�؀D�,n
vH�%�L�/��C�)� ��0OO-=Kp�r�F\H���Q"O>��f�c^`,�tCD22���d"Od�K7e�
~] �c�"��=���"O�$XR�<"T4} �`- �J��'��	� �dh���u��j���4%zB� `�Ȍb$�=H��(qL^:C�I&{�@de����$c#�"�B�ɭQg
�����;h�X�+c�L��B�ɼ%x@-�� ��s���s�˒R�vB�	 pI4����L%��`�ݭlC�	3[�2�"FV��U�3%Χn��C�ɧeJn�3�M��N�z�"��-b`��OD����*gW��XB�9*t$���!�䞴i1�)]32�>0�E����!���5�� ���9$��́�J�([!� 0L5�y���	+ͼ���)�'�!��Z�we��t���	�칃�Ķ{2!�N*k�4A�bj�.vI4Ha�#1�!�D2P�B<Z ��x�rI�sg��@�!���P�³�<��sc�Z�"O�
���H�:Ě�q`ֶ7�	D��D !˔�Rf�vK4ݞ��S�$D��0�Aʦ2���}��u�A&D�`؀Z���*�M�&lݰ� !D�H����B�n����W%k&�$�`b=D��bsI����Z`"B2bxlR'%!D�|��C
�64�7G՞|/^��($D�,�2��	
�$	f!X�ru�(b�'5D��
0�'��mK�H�!t��	C�8D�,Qd��
{�y�	���pzGH5D��B'� --5t�"��)B3Q2D�H4��"r�8|�ȅ�W54��23D�$Pb �U:����@�4$�\g,�O��=�|��&��c�-ەF� �R%*����y��^��(�
�G�q� w.���y�	�;�z�H��6Y�^�9'"���y��[*nkh�b�,U�b02�ǋ�T�<��L�{$�}��aU�_�����!�X�<	��Wb�0���Ʃ� D�W�<!�Mz.��! ��	�9� TR�<�p��Vv\Q;���T�E�+DN�<i�5LG��(r���m���a��SJ�<i�b �F` �P�J�E��͉��E�<iFf�=Մ5��L����taB�<��#T�I�ؙ$k�Q��
%�V�<!���f:Vq���d��Is���Ph<i��B>3�l,��hC9De(�7N�7�?щ��h<I`I���bm�g�36��ȓD�U�B�G�LvH�4F�s�θ��O5������,�����הC7���ȓ
�����/N<}�>�I�]�gd!�ȓujX(S�oSha�����lhR�ȓZ�n(Y!)�3b9bO_	�t���V��)��mТ)��TaQ(M�������(!���5(�`����,��ȓ5I�*�l&X�����%ٔOi�Ն�oo֘����@T���7M�7����c��@�֩x�j���`�X�<W�"���a&�^�5��U[���I�<YTB��y��(q�*�1�r�rd��Z�<!��
%�(�����j2̺a��[�'iaxb�;-�����T:G�\j�ե�y�ʕ�Pd�6%�:[�,�P���y��A<Ok���Bܮ.G�4#0�ζ�y
� �aRԊ�.`���0c�H�lj'"O���TOJ�sL
��sO�a�Ȓ""O��;��ɦCRRH��Y�Tazw"O�)��>y�&ku*���t�"O�� ���*/@�gܠGC�Tc�"OV����i�.I1S��$8-��a�"O��ƆL',�-BFm��kﾜ�c"Or�
M02��±�S2И1ڇ"O���F�|�J��6��p�haa`"O�h��L�(��m�ԩDh���)GO��k���6L���LQ� ��B:D��S��j�~�rRP�6�\��ǃ8D�r���6��=��� �R$K�N4D��b������@��޵y.�h)��'D����Mm�ji�g�!c(�|���:D��P��L~�J��uT�"��6D��Q��4<?��{e��N0�y��1l�d|��F��c�2Eh�E�y�'�ذ��B6W^��0�y���+�hy�Ç�$_�uRt�y2͎^�\h	�$"l	���y��msR\J�N߫hIh@�J�yr��"M�:1�!�%�u��g��y�cN()���Y�e�5n��Z e��yb����cSD$Ha�� J��y"+�{����F
4;n�`	@mW��y2�
"5��  �b�D "b�Q �yB��#|�Y2��_�%��N%�y����N;��('�C�C�/�y��=U��JBF�5H!Q����y��]6J��`��͒[��2��A%�y2 �!cX�́5��:
�HB$aK1��<a���ۉwh�(Y/��:��[$N�7f�!��T�Eh:uQp��0a��Lܑa�!�DL�%z��D��C�j�1��-�!�>CU�]0c���&��r)�Lx!�J���Xa1c�w��A೥U&;!�k�ÀM���L�օ3[w(`J	�'|�4��Ӣ>Mz�(�H�	C��{�'� ���A=l��e2���}Xz�
�'ר]���(TQa)A�J�@I
�'��6aN>"y��m�6@��e 
�'91[Y�2�+�'��x��K;D�(���пeSʩP�n�dSҜ���%D���MDE�"kj�pKq�6D�l+4�۹-�t@�ML3�xS�b:D�J�j�
/~���dF2}�8�N<��N����H� ��%��[p4$��	8D�� ���1m���d���(i.�qG)D�$�Jњ-ppa�E�ߪj+H�a��%D��zW/Ρ|O�˥��2���J�a'D����)ПgsZ`	��'�ʜ�A)%D��9�J\��X�l�r��B�(D�\A�j��,�	]�g�J ��$D�(ҕCJ�-N��@d���s�qx��>�$5�O�x�Ea�߬��!J��o`,�G"O����/K[<9˄C\�Qr�sp"O.���D��O�I;�CܸA���c
�'TƝ��ª~(�����F�@�'��xa�&؟7���b��C"����'�n��d�
e�<�3D�'^�Y�'RQ�g�Ę�^,(3�5ezMa	�'�41�
H7�~<q��e�F��	�'Sj=`pl���̲p�p��w��C�<� z���i.ڡ8����0��"Oz���-�/k&:�:P�#5îz�"O��c�����@�m�Q��&V�<F{ʟ&�]L�$�I<	aEO�8,T%����	1%��=9	 ".p�a �"5%.��2�I�J�J#|�''J�#����u����g爐Wܬ��	�'��E����W���@*�JKd�	�'��m
��~(�	�Qd�R�A
�'�n�Iw�R+8��\xq"}Z�*
�'�FM��뇉[if��h�6u΂X���hO?E@1��4~��C�(�5_�6 HbO�ɟ�F{��i�$s`�PUX�L�0�eИ�C�ɚ �H�j�H�&^$�3�$�8B�I�
Wz���Hצ�b(�
�w(B��.Y��$��ȭIe�wH>|JC�	��JH"�
�N2⨩瑣+�C�s]N`�����R$j����C�	�Ab��)E�&c\��%�]k�B��](���mұ3xs�G.O��B�.qRöIc��r�ٹW��B�I=^��T��Z/G���AY* aB��2JQ��Ж�,h~�4��t��B�I�T�{��M�9�L���ա�xB�h��Š��-�b��栖�O��B䉸{ꀰ���>M
B}��-��U�B��6?�FI22 ���ӳ�w�XB䉽f>T4ڦ���y�B���@B�I bJ���(Q���|�Tm��/��C�ɨ< �"F�G#iނ�AgM��U��C��G@t�5�ߐ���R���bi�C�	�ڴ!�r�S�?�|�!EN���C�I=/��P%j	�X.\�3�$v��C�ɰ!X�A��D�+@E���,8�C�	47�u1%*Y#�xH:��)@�C�	�,ڼ�ZШ_&����*�)+�B�	�<o0D�u/�A��S�=H��B�I�g�t�iP�G�C<�3�I�-hTC�I�zl��d�N7�6D�Ӎ�8_z�C�I-Ny �Y�*� ��3�⟄��ɾ~P\}�R�G�E US!���B�ɶ!~���lG!u��eִj@�C��$ �������EU�ɓ'(I��\C��7Vc��HD�V�V<VH�6Jj&C�	�E�^1��ёe�Z���c߸B�I��F���Qu^����X��B�I�=��4Pa�6Y,.��s"�i5\B�I�SN���,iTI<mʎC�I?13��@a�4T�S��ޣn��C��W�P�Q�ߘ'��e��;�LB��(1$��#k�+hx����ڎD�FB�I�7?�����\�n���1���u�BB�3bA��e�9~.<c%�C�>"��d�O�b�쪷��Z0E���B1^l
 $� D����/J5���q���%w��%���3D��7GNx��	Z �Ѵ�h�O�<����Ӓ&��T�W�b����X"��B�(�`���3K��!Ȕ�J��B�Ɉt��:1.��*M���d��r��B�I�N� -��ǱBDZ�R�=2����j�XI���
\)��&R#@~L�Цg)��0|r!��(n������wYm��l�O�<a!�݌	H|���\�b�ji�ÖM�'c��&D����!���M��N���:B�E�̵��]6�J��j��o B�)� ��G	����$�u��7� ��"O�x���O�R���4�&	�pp�"O�#��Z�3BM9S$}6���E"O@xh��B�1Ȕ��cU�{�,)�v"O`{��ƨH܂4R���)g����'��I/$I�-Ċ*��@;r�աWcB�I������ަ4eoG�#z�C�I��>E�@Am��0�� -I��C�	S���11,�Rn�l��Ż-�C�I1C��Dp6�[:�� @ϧ8B�C䉅k�A�C����U�C�ɪ�T h4Y�a{�	�`I�l�J)$���?A���nI.-�'��&p�[�e��!�DϪ�����2/�!�F7�!�dڦJ�P�ڱa�b*���2)�C�!��K6�@�����)rx�X8�HZ�!�N1G��)9�A�V���@G��cq�y2ቐy�^p{��B"0GDm����Q��B䉌v�����N:oTl�A�n�;���Ov��d��1�f����P)��% V!��	�&7�9��@Sy4�G$�He!�D2�̀��GC�,��c�N�!�\4���#�m�o������«�BO|,���K�F.L1@��N�<ɸ�P�|��)�ӊ6�v�����
��Oڲ"F�?����.Z�x��ǎ1Sy�2k�0�!򤞽K�,�Qp���e���P����'����N��F�z�C#�(64�l��'[X�ũ��P$T��Ar���'2�� #��tXG��8ָpRU�
o�<YP��0|�Ÿ�%S�t��	��	IT���hO�u�D�j��_3��*\%�Խ�?�+O�#~rgϹE=^C���V6V���c�<9v�F�V'�1iw
]�Fш�p��`�'ax��G0<�E�&�H)
���w��y�%
2T)��aT�Z�'��Ї[�y���^�N�z � ��
�;s/�y�n�z��ez �ț�lH��hV����hO1�<q�6 v/&�Y�A�w�V$�5
/D����"\&���b��P1�!�a-������y�Q!ܭ���� ��(���,LO8���ُH�0�e�_b��&"O~	�A�΀:`d�1J�}Kd"Of��&���t.Q@dNx7��"O��CU�L�(nX���C�'N6u@6"O�t�@柩lfXrÎ�m��eaf"O:a��d����xP�lV��>���"Oh��p�֫P�m+!��/ �<-hW"Or����^9��(x׊;R�qK6"O��#�ԩ�檎�6���t"O����鏜z.z�B&K���|�p"O4�9%Ib2 �"�9,�(��"O�`s�JVO.�s1�3��E�'�!�� \���[%+�~� ���<n�!�D�a~z�q@E��4cU��;~�!�$���8��S_�b�(lcu`U�=d!�DE�n�!�f?��D!�N�&!�dF3ʲ	0t��!z��d���[S�O|�=���I��W�t�|r3���LAt"O���Qo�"y�&�9$�^DH�
�"O���ҊL6���d�
�
�4"O,�qn�0f�ʤ[��	]��"O$��s�	�Y�X�H�@͜u��萱"O�<���'*΂8�d�H��ag"O� ƨ�d��&ad����.ʴ^��!���8LO�YE$�hKT����A8]���2�|��)�u]>mA���3`L�2�@0r�C�ɛho� "�=Z�0�F�ў8��C�I�`Q5CS M�.%�$�M!h�C䉰VO�h�D�z`(�bP��97�hC�I�	�Ԩ��i@�֮xN�T�FC�	�Y�����*).�ځH��CH��3�<��/�9)�d��Fyj'��O�C�Ij�d{�⎽7�}�f*��˓�hO�"<`�{���BL�d圐A�B�\�<�W*Z����k1�ɐl+T�`W�ĸ9�B}�P�A)� �ؤ�=D����8��(�A��CM"�S��:D������=Y�d�����D�J�8�i5���O��d�	0�	�E�Y���45@!� /KM�<�� ���1U�E!��d���@�B�N���K1��gZ!�3�4e�C�Z2do�$�)2X!��Pp���YhRX��N�,B!�$�w�Č���N`�(0!�d�' 4!�������z����cK�w��3O��s�-L��R!Z�R�j �qY�"O�4K��r��8�R�"D6�`�I|��kY�Y��8a�#V2l�J.D�0��h��/�.5s"I�@�x0k!D�(��!0������/vFS�j?D�
�o�>+4 �J�g�<p�^�c*D��+�@�V�氩U��&G �2b3D��a�eWNڮ�%��D-
08�g+�IU���� �ؐ�H�C�$�x�J	$|@�B�Ɏe���3���8+��r�RB�ɳ\ʖ�����Cy����F�
��B�I�b�9Q��Te�Ѡ��E %"�B�Ʉs����Q��%FB��8�G	6CC�ɼg՞��ˡwV���$��/F�ڌ%���'Jў�Ӟ1>�\��B��Vrh)�`���ֈB䉶��r��
7S�q)��MYZB�ɕAZFqpG���D�8ePva��,B�	�]d�	Q�9d����ڠX*B��9'�*pu��6_��d;�l91�B�ɊR=�"�M
�a@�GY+/��B�ɮ:�I���3�<��"ۢw�\�LG{J?E�43I�I�sh[/C�����α<���Z���)[�2��U�2;dU���s~�IPkԵ de�*�	i����y�˚e��7.�6hv!�Կ���'��THa��t���)�F��PH
�'�pq0dbؾS�z5q�L��K�.E
�'����(,���I�/ãl��)O���$\�(C � Ń�7��Epaߚ*/!���N�ђ��ȉF���p �I8<�4O�V��P�p��-\��"O���m�㾔�''"~5��"Or�┪V�s��yu1%jƘ�R"ONY�S��qA6�ѳ���|�>�"O<AZWl��rQ��V(N]Q���"O��raY�{�pXy���k�x5�`"O��;a	�!u��ܠ���E�,����'��O�=�'\>�cWHU�F���g�. ވ��ȓ�|���*A�����ҫ�a��x"M��nӚ7��q�4�M� �h��ȓQJ�u�R�SI�)+��#}�<��-ri��J�:�޽�f�ʹ~fQ��	p�S�? L(���:Np��yv�K-8��m9��'<��xe`�8{�V=��NW=&JA��&<D��[���[�t8�D�S��My��>��0<���U�krfI��=`��"L�<�C`U�h&<Y�%E��'��� @��p�<S��L�%UO�:���Kp�<ٖ�'H�X\P�^2=V��:CE�qy�X��$�PGx�W�d��$�������K�"��<�Oꘙ���<kI���4��4^�Q��`�On!�WΔ�2���
� ��|�zt�K>��H��x#�W� �����&v�8�ȓP;�A��P"�}�a'-W�Іȓ4F�}Hwƅ�6ș���I�L,�ȓe��yaR�2[V����!M"S@*�'��D{���EB�x�ї��$�h0h����Py)GtC�� �
"�q�ty��)ʧN?�0B`�?��y(���3 ���ȓef��3K� =m|豣(Ş&�t��c/���j@�L��T�BӜs�H��P~�=`�d�/���Sc'�)b���W$QQ��D�p�Ұk�FV3�fp�ȓn��H���506� ��aWW^�ĄƓa�Z ��B�q��8�įϕ9�X��-�yWT�q㨅�t�m���,i��u�ȓG��C�Z,�l)���@�6����@�rx��N������(�&z��ȓ1�@A�+  y�T(c�ўW��	��j�-å��� �;�*]3�Y��U3~%�aN�'�80�C̑�KFf=�ȓl��a��܈D��p�YL�<����`�3t�D���c�F�j����ȓR9P������#���j'�U�G��ćȓed��Q���n��a�3S�Q��-��${��L8q�I�AE��z��M�ȓyD��	�邠�΀��I͖0_.p�ȓS�z�1���jF�s@�+��ȓ@��	D)-TbG�$Ct��|wjI��~�|Qק��Q�y�ȓn�J��F?6�:�Qa�7+��Ն��$�{慃�4��(YQ�ȓI� �b �/�T�w�ڠSS����ܭ"�6!��+�ٝ00�����!�5S��{E��sV���ȓC���Е�Ɓ:�dԓ�(W�)�ʜ�ȓ0I\Dᐪ��8��0�`8Z�� ��. �Pk���v\Va��L7h��	��-&L�ه*.X��T��ѫe�h�ȓS���hћ*I*�3q�(L�
x��CY��c-C�����v��
 �`��H�f\J��}X�]�bkZ�9.N���*�(���Үay�QDχ�5��ȓ�
��H�����Ӿ]"x�ȓg�1 ���qC�'N�*6��ȓ&����J��^xZ"��:&��1��ܭ��f�NRN��]��=K�B3D�!ϛp�4
s�GG	T�T��'�P0�f�M3Z���H�7}O����'� ����hr�lz$��|�J`K�'0Ƀv�6H;�d��@� �'�x��c���ĵ���>�
��'��E��cO�[40Q�� <�lm
�'���8!���h�����ѵ,j�	�'�d��5�'ݪA��j^. N�-�'�x��E���%�4�9�	e���
��� x��G��)�h��ګ<f���"O�����Щ)pT ��ܾB�d)�"O��+5"ו2i�y��QMZ���"O�hIr`Èr��*��q�~���"O]k@*�?��	��烡Cz��4"O��R�.Y't��!d�"����"O�=������P��\.b[��"O�U���WA�d���d]�o���B@"OB���(f ����I'Kw%��"Ov�2EO�+���igE
wpAZd"O�zʸC�"��S��} c"OT��4�zB�K�	DH�"O�|���(�p�IcQ�|MP�"OH@{�`��f�@�2�茭eo2�e"O��H�Ζ--�^��T�ҏ$z<��"O0�0"��f�b�Cp�wv�h2�"O0�Ce(M�s�4�#�F,Y8���"O�Y�GF�1ub����'[N���c"O�L����+?��T���!J�)�"O�hy䯈��]x�KY:-.�i2"O�ܘ�L���F���
H!&^,P0"O4!����G�	��ψ'�Z�#"O����NELBx�O�w���"O�BGJ� ,�f��>][0�q"O�%a��E�W�,8���	1	Y���f"O�xb'��|��l�Cˁu�X]�$"O��kY���qY�l�(���"O��8�*��PA�ď7��hC"Of1B� 8�&���O��r!��"O�-`�,�V��!�-�2"O@,�%C��b4k�$�<�2�"O�-r�Ƃ�B:z���G�@Ht*"O�њգC�_��-IUD��{$ñ"O
�T� �}w�1�f#R;{�jU�"ON�!��j�䈸�4Ėe�'"O�����:<�4���;P��q�1"O��g��9`�ly#�V�l҄	#�"O�X��WE��LC�4XV��"O��� !T������!PhP��"O�MS���C�>��G� ێ��E"Or�J�蝀w�vy�� ��*,�6"O��s�Wx�^��V��$q��m�t"O$$(t�\a4��y4)��$���3"O��Pw��n��G��[��Y�p"O���+��.T�SE�6$�T�p"O8�I� 
�2����U�	�.���"O�S�ɉ�3�\,x�fZ�X���R�"O�4�l�;0����CL*n6�R"O���b)	�$�� �tQ֐�"O�Q")Q�dQ���\2��"OzH3 �	~�r8�`��	9�)�Q"O\�j"�P!����-M�t$�E��"O�Y�Rˊ z���c�K�/b��6"O�!w�7.��f��J\�"O�iy�*N7�q#-�v<��"O�4���H�.ݓC�ub$@s"OZMȆ��-
a� �
�.C���d"Ot�����X!��%�V3A�>|�'"O,\D���2q� ��T��!�f"O���V��*Hx�C�n�4!�`	3"On0�P�ȗ5�*�c�Ǜs(rP"O����cί>�{CAP�l���"O�|jV�A;������\�
R��"O�9"(_>Zh>��4jA�S�>��"O� �uPӤC�VY�YQ�!rL�#�"O�rp.EZ��9��E2iVD)�"Oڥ#3M�"99<zT˓1UN��s"O�!��� N��k ��sa�E"O��D�A����U�@�X"�= 2"O���3��')�98��@�H�|Z�"O�p�ƀ��;PX�A�f�>z�:��a"O�uh��^�exՃ!ė�>��!�3"O�T��X��-Ӥ%W�P���"O��g� `�x�%͏wo
e"O�AH����d��F$XD���C"O�Y�I�8.�be�a�1̒�
!"O2���E�
e�xP ��z\<���"Ox�{�n�> }�L�2	�>eX��E"O�P`�a5d��Šr�0REJ�p�"O@��%G�D��x��I��!,�"O����
w�l���H<&�Z"O�|  ȑu�(-���I)�5Z�"O�(�A�Q��tLTș�<"�14"O*Y��$�`��ͳV�4d��"O��Ռ�Z9R�8��d�Y��"OR�"�́KP�)�r�L�1"Of`���ʨ�����iҠ_�~�9�"O�!�c�ĉa�L�uh�'U�2���"O4�d�ֱl(�`0�-�d��A��"O��3%X; �� �#*u,(C�"OS��'o)haCAL��t�A�"O�DC�3p��pĄ/YdNi�"O��ɲFS�nb�t;@��*Z���D"Ol��"׼s1�#ǩI��QY�"O�P
�k�H̞�3�b�+�"��"O��I�k&�i��ҩ�Hb"O���&Ǐ��d@�d͞U�d��A"O(H� �Lt���.�[�m�Q"Op]�c�-{Y@�3tk	U�����"O�1sl�b?jM�z�B�'"O��aǵ*���2���'wP���"Obд�I�=�.�Q`e��h}�d�A"Or$������pM�`�XTe�:F"OVh�cK�v���+����n=��"O`D���,W0�l��27e���5"O���Q� n�2	I� ƥ`IX�C"O����ϼj�(�!`��i� <��"O✸uI��8P��n�"�kq"O<]3�DχE$��wM(7p���r"OVs���Z>4��7b�5vN���"Ob8ˢ#2Z0!尅ek���G"O���N������8~���J"O�<�SŚ*)��CnN�qw�99�"OȜb�#
�%�xcs
Z��~��"Oj�۷�Ǆ^�V'i�D���{�"O��G`� fEV��Vʐ�]o�p�"OpmQD���'�v�:4�'U��X�"O��ᦣ�#1&�8��(D"O��i�,l5yEك#2�{�"O�4����J��:���*��J"O*�� @ܩ7�f�1!��)vJ��"Oh}�i�" X�)�h٩~��0b"O,�Kň��:Ef��Ն�R�*�p"O,ū�)��?�a� 3���H�"O6ّC$��y��`Ã͡׀=��"Oz4�K�-
�.y� (/o�\8p"O�xbV�ƊD�
�:5���{���(a"O��;u'	<ti���fj�-s��С�"O� 581���S�~Y:��P._��y�"O��Yu�ܵ,i�\;�G�0$f }��"O>���>l x
gĖ�ddLHi�"O��"��E�n��<�#��Q�D�HF"Oܬ���'dW�<�5IҐ�,���"O��C��8��x��_>j�D���"O&A��!c��؁F��$4yp���"O[�R�, v@��4aVEzf���"O)���F�{*zŮH6m�p|y�"O$��!��4�aW@�5�NY3"OD�S��53��DŇ�?X�ٳ"O0БMS�B
���Ĥ��L��bd��P�'��>�I�J󍃮`���r/'$��C�*m����C�	b7NAA��a���Y��p1���'zL��� R3YڼTk�"<��hO�R�t����M)E�Q�	H:l�TC�+O�T��X=6��bt"��"7�1�S��M�Ș����S/^�5�T�е`�f�<�-�5� ��էL,\t���b�a�<ea0y\A�l��K�������i��hO��<�s���Ze�I]�g/&p�hKl�u8��Q�!���Ee!ݜ4�@�2D��17 ��!���g�J��6�q�(24�����7�b<0� �T/��+����!��T�f��3LE�v.詁��^�2��y2�j ��h'�Ek���& Ю$��#<���;�S�D���r��X��5�PH��Ł���"�
�<�}z�/P480��3�� �R-�u�Ot��0=y�lC# �p��zl�	�կ�n�'Q����ZhR�鵯³`3��Mʆ"���G�p��%�C�Cd�HG�Ѷd�LAob��Gz������P�Ȃ/����ӂS&
�&B�	S�|�tLs��)S6`�kT�'��#=�Z�,�z�n�H���q�Z!hb�Id̓d��<%?� ѭU�=�|���bP*`L`
�l`�<Y�	?g�0#E� NW|
��V\x�D�=!ܴ8[�E`�2N�T�k�D�2i��A	�'�(q(`�ĳ(���ѳ,�[����Ќ�N~b�)�Ӯ"j�8�D�X�i2l_)@xC�ɔHK�I���,�Ե��^�<�C�I�c�,�q�j�D�T)X��ݮ|
C��h�����@J�rA4E+����0mN�����)�H�!�ڝ3%�[e@��
B�-ꓧȟ:PKC��VR��ļc�%`�'x��G�:�A7�+��|��t��Ĥ>�y���
(r�zK�,�Œ|��$��=�џ�F��؃sz(LP3C�N���ѱ����'�z�CS+WnZ���'Ai�Y{�'����1�S��M�Q��B��"$��b�"5Z6+�q�<Yc�����S�P\^�l!��R��hO?�IEu�T�_��td)�ܓQGxC��ݟā�%����L�x⍩�:D�,������vl³5��!r�.9D���V��+PD��R	@�}�@��s�5D�(q�Kӕ�dhR��C�.&Ѻ8?y��ᓺ`�`u@^b���fA,�C�I�(�y1	\%��Q�]cF�E{J~bq�;7&�`�oO= d(*��H<���2�vE�"�	��iӃgW:|���Dy��'�j���X�m�~���G�f����'$�j&�̟cJ�M2�ϗc��R O���ka������^���u��hG{���Gy��`�!��+ �y�]X�}��6�	M���'#����h�&~Q �:��J(H�=�pV�T����~� �5Bχ08 Z�ɇ&N0ؙ!�B�'��F�*;L58�jΠ<>h�A@F��'@ўb>��Ư�v�]�Q�3�H"3D�xat���f8�qslP��T�ק/D����"�<2ՐA�	̙E�ژptb.?	���?9�'�~�js
�=h �!ַC[�=�(OX�=E����C?%:��<8���@�O�)�HO��D���ӠAχz�� 0끢 L�04�|R�'��Z���\�F<S��"eA_(�?��'`�'ב?7-�"Xu�f�hY���Ǻ�?��'9����.�<S�� ��O����'�2����'��������iB�	zy�$�vEp��	E�NU�4�Ҙ�������=�}��4\��)��cهSp�bv �"nk�D����$7�S�'+@�UkU��,�h��%��C`<Ѕ�T6��`ǔ�UȔ����-sɎm�ȓ$��R2	g��]K J�"rcVa��hO?���.{�Ԉ1f��ʃC�?�yr`G2���
srA�Rf��:S��D�i(b��v� _�~�!��E�O��zr���Wp�\�q��&�*�ksѥnt�	^��H���{d��w���(֢Z�#X�x�e�|�g0�Sܧv���Nh��4.��w��X��+D�� �"� A�TU��/�}�Ɓ�A%lO���y�KP?V'ē�o@�����>$��-V�6�A�Kߍr�؜h�fX���'Zў��4��̙{E.�����)]����"O�#�L�|��ppQ�Ӡ��a*P[��D{���;1<�A�]�|�
a�`O?v@�{�̗~h�5�i?x.���DD�$P�'a|j� M�v	�W.ޤB6��tF���'��G{J?幓��.��D�e+7�h�q ,���Y4v�)K4��e�()v ���!��ܴ?}�1{�P�=T�AȥT��!�-.�T�*cC&�f�:%�[�_3XM��S�nA�BɅ49+��2o"@� ��.�z����l�a4�M%�H�ZA�YB&D��8Ҕ@٦D)�H�e�O%%�<��&��S.\�V#@]�=p�ē$�Y*���|=D��$�A�Ѵ%�"O(U�åO0k�\ecGV�Qb�ص�'��-����5l�7��X�4�9U �ˉ��s�+�G�I�F� ��ةh��-��h0D����%@�Vz�k �9M�z����3D�@k�5�l��*���'K34�H��iC�O�9����CY(���\�<�䌎*1��c�.÷p@BL2V��R�<q��=E�V�S��O�K��8'�O��F{mFW�ĨP�L0#��Q�oQ�y��\/X����G
p��oW���':�z��ʀD|�E�@����|z�
��yR
�9C�<S�NT:J�ӄ�Q%�yҬI��.̩���-���1�y"/&A���Ƒ+��P�~�����>ɘ'�J~�<qF͖4'j�Q�Z:W�C,M~X��O��A���a&�7�	�R��"O��a�l� �,ӡf	4{�e��"OJ�)�NN�.���ߊx��2�"Oz�#!	�2���C����� "O�l��ړa��k��ͅX�NxV"O��hT��NU�����=A�6��"Oj(�G��Ws)��m�g���!��D#�S���X͈c�#-�����S0=�C��*��X�De
2j!`� �"z�C�	 G�h 
�"\�5�Ph�0c�<C�	�#C�  9@�ģ���T�D�kv�R6O�=E��`�,G��8F��c2���̛�p<QH<�,O���1ς8n����Nj���"On������YC�|�eǛ#��%�T�>�K.�S�'c�1��߬
y|�
�-ϡ�2؆�*i��c�d�"e�d��r`�(7�������?�D�V�8Ɗ� Q�%Qv`AZ�GH<��'D,�J���/-{ܐw�˭~F�?9C�,�)��qõ��3��Y�*'IaJ\��Xy���.�1J����W '�5�' ў"|���/N�����N�t�l8�tk�<�f�
=
�<ʷ ׄ�X����JQ̓��=I�(�L_Z�xo��r��(��'�J؟�j��'��q���"$i�HZ.r�s�'^�y��U�D��0˶�S�}Z��`�'��p h�*Y��,��Kڤ�;�'�֐x�V�ޜ#��5<9��
�'Z�)�O�B�V�.�ƥ#��B��yRᇞ"�) f�ɼ+�u @���yJ V��y˵ތC!^	�W(@�ybşs���7��:24"2�\6�y��*߀x $�G=-�8����yb�؞����|� �m���y"�ԅ�B��f���=�N��y��ȨB� �t�L9���"�_��y�B�T��0۠�ѥ|��LZQ��	�y2i�+)|U
��W�|v�5Z� ���y�J�@:��Ar�Y�e��A���E��yR�ޘj�1��X�mg�	��L��y�$�;fC|<��O��a�~)R� 1�y� B�\�\����	]{NI���1�yR�ƀE�qy�$֟W�����G5�yBd�X��S��:V�����B��y�N�b�"�"�$�I�@`���=�y��
�B\I)���P�L��`�D�y2\t ��� jXS�����E2�y��N�T� 8[�CݨL��w����y�3n��8ځ�=J�L�j�KH#�y���+P�L��k+� ��e����y�-�c�"�Y$�X9,�^�i�'��y�Gն_�$��N
3�"�8�"ݪ�y��"E���#L�)�,<�Q�$�y��R�=�z�c�L�X*��(ѭ���y��?/���G�X�DP 瓿�y�C1"�^���g� C�h<�@P��y��ٳ((����ט<]��#��ؕ�y�g�!�r��8�BYД��yɀ)SX�.R�gh՚7	J�yr
�5	��	3�r�� ���̈OP]���S >n�@ʱі'�⽚e9O���!��RZґ�$X?R�`�K$"O��H�FŠ_/@`C3(	��l�"OL�*���/-�Ȅ�j�*���X"O���� [�t��։��|�hh1"O�m!S�2E�V��iEA|�]��"O�I��`R�M=䱲����Q`�Q��"OU�n=a,��#�Va�-�y"mϋsl�"��J!
������y��܆K+J�edX�iz� e�C��y2��+;N�8B@��1|�XX����yB��?�)F��vU��$h��y�U;T:.��@��i�T�S�=�y"� -;I��0�
�8a.RTR3���y+^�JĨ�/Ubr`��E8�yB�*S�P:�'!j�|,c"��y
� ��@�ʫi)�)Z�L� N�0Zq"O��z��)R��v
96��� "OvL��d���nA��!:��S6"O�MaS�'K�Ƞq��+$���*O` x�gǨ7����h��Z\��'39AQ�ȌoȐUප��qAIT�<�#mX�s���qժ��=Y
�s!~�<Ip/���8̀�oO�1Ƕ� ��M~�<Iv 
�T�¬��D�WL�����<d��r-PP���T#\�����x�<�$6R�����A���@�{�<��d�#_֌d(�K�;~D��w��r�<��h�ʨ����V�_�|X�#A�Q�<a�EN�K�n����_�C�.HQA��S�<�醠*�:H�6B��7(e�P�O�<��-B�Tr^�����>����I�<���Vu��|Sq�Y�8!���@�<��^k>�KwaY��T<0EC�<�M��@ئ��g�bM3B�̓g�fE#b�=OB(��ƭ@$��3��*8�tcG�'�F8��� JRmsff�6�c�JЄ���'!��#��-�I"k\[#� _�5�Ɇ�j�"?QêX�
���)���%&�c*�-j��lR(Ӑ!'1O�d;��#"�iQ���BB�y�HM�yȺ�"F  (�IDlj�v-�3 �S�O/��J���9G��P(Ԅߩ*�Dq��/W���{,O��Kr%1�3}�EJ�@��eӧFծ3(9JR�Գ9^�\bˎ�"�\!�K|�=T��+RW&(!�?>:�-�"����r�%7�4���{4�!X�Դo54��¥ёlNpd!�$�&%Te�3ʓl24����iBhTAcdT�$'��D�V�p�@39vM`U�U/���r ���x�ᑛ����%F��g�����T�gc �~R-ؽ)h~�V�ۼ�� E�c�tLε4�'A�� ��2b#���޴�V��'E�Kȉ�@�ŤOq�@ �'(^����LW�|�`8aeM������hIb�p�ڇ�F2QڀaA�I)\���3�Q4� ��=@�`�('�E��� M��@!)� 5�Ywj�K��!S7T��	!BK`���)zF\�2VbS'>���"�$o�Z���,f/"U��� ,O�8���+G�X}3��͞N=Y!�6lh��#�I�6rH���T#��bp��C�ZECG$LM8E Q�7om��ϧ!Ӧ�3i�0D2����%y��F~"��(K��=���T`��)�L``Kɝi��`�0�ĽS�����$����F�	�X�C���
(��&&_.<J���#�yǉ��2�D���!w�|�h�lP���F���M�q�)���t�&#�����tnu2E��Ct���c��?ٞqBߴO��5c��Tr(�j�g[3O鑞�k��Ư���B����&^�@Y��??i�fA)O���h�Oz���"��P`�r�(���Sw���uB�ϙ�y���"��/� 0��1�O�u������¯5���bUh�Z�"������U	��|�wV0�?a'AW	xR�`��+��\d�B��אd��I�˙o��#=i�O��1H9q�K(�ӫN�dz��X�1��ր�*3��Wق��`�[-d@�bsA �i�[ɉ'{^��2�F_δ"l�
M��xشyX���B���@��ӧ�
,�sb��t}8�e@�Q�L�� I�@j�kp�׆�~r�H�4��I�9�\�J��B�R�=ȓ�΋#���m�� m�/rZ�	*V��t�P(Ui�Ӻ�̔f�68�&�}���TNKTX����/P��ZPʏ?=C,REŘ8H0�3
�]��I�+.��i�Y�)ʧA ��5D0b�h����H��RFz�
�%^�JR��q�'>x4H��'��h�ԁ�� �ц1�<��C�� ӄ��DIO]pKo�{�j�����	Kk��=��B��s�,�k���}��p�C��V��(�"O:���lFY�9B�B|���C�E��#.�2�����'���J�8P1��� �4��	�@6�I:� �g� ��-��k�`qPq�\�[��C�	��vX&��X�P���=;�#=ё,H�j�4���!�S��$�!]�V\p�3s�^�'r����G���!�'�d�Zɨ�nB�O�����O0�i�
Ս8�$�Oq�p���L�>�p��C��chv�ɗ���tV�@+t%'4�0SO�7m����b�:6��a�)?	��N%vn�Ig����MS�qX�S.������0X��%����39�B�	�]Ҭ5أol�x�e��#7c���Z�>���@@f����)�'k��@�G�/(I���\8e����� �Q��ȝYY�	Z���:��Hs�O��ڢ�P�y"8�1�:,O,9��5l H����a,�U�'�� 3�F�l���TE�9k �oɭ0\�Q���P�B�.zZbx���1P��:����[	�㟐#"���^����j >a��\�b�H4>-,IA�G�6���;�"O �k@��  �SԣH,�$�Kv�и�.�@�@�3A;�,���h��d�S�DaZơL!��p�4x!�8CbE���	�.��Ca�z��H���=�4@��'fMP1+��jd�xq7K��ܥh�vƾ��K�5c]x!n]*��q²��V���\*U�ܵ���'�|:s�*`�s�n%�<�� ]�"z�5�FT-5Z��(�l�Sl�4��P�
�J�=i�,*\��B�	�N<&MY�*�(k�Yb�kP�z�Q�D#S�P�N��vH's�
E[�8�g?��J�e�ae��$v�)���So�<I�?r�tyDo$	��P��G#6���cqǈD�*T�P�8Gh(�3�C����a���������=�l��	�8��Q�'`�N��)WFF�H�x9B��4��e�-�=j|,�$�7�O�x҃j�<YH�3D^L,�D�����UB#G�W��̩���"�����w�ɟg��T��\8����"O��WC�j���wi�G ,ؖg�;|9*`�F��y��0Ԁl}Q>)�'���A�Ӽ9��Q!���x:@��'��B�,�1��MH���?����W��b�̕�7��e� D�*p>AR�k!�m�6!�q��q�H��)/X�*���8ԅY5J3l�bƩX��b-��oإ2�Hx��/,��� ���;�����Y3#`�V'WH!
x�R�I�g��' t�2.I-c��k� �bsx���)_�,f��N /%~,%L��!���~əT�K�ds���;y��K�h��O��V��9 n\����-?!5F�=AdaiR�ҵ�QSęvh<�W��j�ցjd�*�a"d�Y6 t�f,ܪ@4�b� A�%G�\�Ó4�F����H=5U��jG1�ft��	�4Q��[�
F2�zDSmՏ!�Չ��[�{L;d���z=� 3r]<�/*h��qw��OQ��Z�Bo�ɔNU��`hC,8�H�!�L�u�L�|b��MƎ�YwEȾy��AZa/�|�<�cÔ-�Ă�j�'���k�!�??X����.��`�q�?GX0���O���ÅZ>�0�E'Z7EK�=3TO���d�C�~���g��>2�����M��q��-w�l�s�I���'uj8l\�<�ВS|e#�N�7�&̐�ɚh���	�J`t��m2s��L(� [2p�8"s�+]|j́�k��a
�1$�ȑ���cq���[��qÇ�LĦM���؁��b�H��FX ������2t��T�
R���[�c���çI��Ψ�KI<F:l�	���<��GԘ2�2����ړb~"��!(O�K{J����
�§�O�&̦H�8D��$�_}�?!����@F��q�Qi��y2Q�16��s�� �8Ur�lȱ,�Q!��Y:��8 �� Ĝ4�b1}R�&KM�	�OW�����/g�I�� �F]�	ד;F�Kp�.RlP�g1�֞M����*�5&�R8ɒn�2ak���L��X�e܁����	.i��a�掃I�ةh4�5��<2r���dU�O����թb�˥}>t������i�f)l�l�G�ǎ��>)���,"u�L�4
�mk��K�V��b2�J��䁖��)B�R�T��p�[���Ă�`,�����bJ8Ʌ�ܰn^!򄀨VA���ee(H��Ƒ2�zE�N�,V
U@���R�b �qÀh�$%擡4�H1�g�ٲq(�3/|fd���gq�U¥ײַ�y��?g���!Q�Ӥah�"�+e��'��2��&�g~���r�fp*'�0GH�J�c����'�T���/�
���G�T���s�y�!X>t,��'J�	%���GN�0?aG �f�>�1u�F!��X,�T!���b�6��O�H���Y� �(��f���!�#.+�q3�J&D� (R�Ǌ���J��2��A���# t��`�(7�d����LJQ	w��(��T�?��zrb!6��b%KO�<��+Q�.�	0�ȑ+c���"*e�<���23�"٨�
�=�~H)e��e�I6Kyn��JM���@N�����|�����F����I C ^�P#	J��LR��4~Z5��X�~�8K�(S/
ݚ�!�mɧ�/?�u��+�����
<��Q�vbD�8.�2�xBч 7�q��i
�H�iHt���|wH$��$æTIЄ[G���'�r؞� 6�)2,������;�\Y<O�M!p�Jp��K��Ot����K�A�>�m�@Pm�@�����c�e.�B�IV��iڲ �4�=��a1԰�h����c
�Q�J�OY��X�rǕ�n�`��S���m�>��QfL�҆y�/&�O�R��>tޔ;��1v�؍�v��>#����͹|6-3'.]x�D	p$�@��p��'%��a��Ib�i���7Uk���g�3�>����ɍ���>)�A��	V����!e�2C>�T��O��PUˋ,_%k�#}���Z7�0z���$M
�7�:-yUdV�J4PA�G	��y��RIx�4��d�T>]��
S=O�����i��В�e<k��i��ًr�*��N���N���M�%�'�h�B�!f�;�f�=	�Ph�OF���17q�����F��O�8X3AY ,�DqVC�=���s/� 2�c�jԖd0@����V��Ӂ�\-Ko|�ã��0��`	b+Y�n��͂�f9>��O�͊��V�;�
k��>�E�͓x��ysM�z
�q2 c3�8">q2/ܐ?h�1xbo!�S+>���z�	��C~�m�͎	*E�	;M�l%��,�mt�w��*��8擆)^�E{���!L��M�3-:2���q��� ��x�)ڧV����gι_�+P�LژܧO�	e֢��!��e�� ��\�t�j��C�~��'��0aǜs����.6GȀ��
�E� ӳ�Q3`��q��I�!��	.�>����8_��
�i�?Ku��,8��E$����}�VlA'l�����h�x���A /�^�<�� Ƭp�%/d�}�3f�Ty�U�"���=E��B�U���
���Z#L>�yr�,2x ���%/m�4r�a�,�yb쓑;�hrR#ǝl(>ɫҀ���y��C�}4��ͿY��x�R(X��y��9��9���W�]�Ti:C�/�y�m�m�������<D��i2���y®X0�E����;��,x���yr*_?g5�1Dʯ6b��vf��y"�H,#�2�%k�"Q2\٧h�;�ybƔ3"����JB�S����՟�y��ч �B�k����^�V�p!燑�ybaې]î��ц�0b�P����y��`jF�JZm�`�`	B�yG�.%M����nz��(�(�0�y��W���T:v �+3:ʤ(���'�yR/>@�~�K��K;�0h����y"�Tp���߈2#� 6	�+�y���Q)��*��Gcd�ڒ�I>�y�d� ṕ���$:e*,����y�NX0s�r�*î���	�	���y�N��Lu����a�ڭ�ԃY>�y�-�����&Y
dp2���A��y�l�~�Zu��O f|@�fܷ�y�Ε�l����"�֎*?��#��yb��!<"cb�2W�jl!����yRLƷ]�$ y7��<S��`�L6�yBW�`6��n��(�$ѸWLE�y�/T�9s2,*3CQ�(cLD�C��y�kK.��e  ��)�pM��yR\��d\P��8"_� y�(�yb�O�.,<��`i-�|�g�P3�y��ڛ�.Qq��� ���b��?�yR�Ҹ"�NP:�A�Gq� �b���y���~0��=�Y@�Σ�yҁ�>F{��ւX�|'8 ���U	�yrȂ�M9d����t��h���ycU 1�6��a��[4XC �W=�yrdI�j�}�T�@W�D�y�(ظ�y"ݯ?�젠�E�UCh�2����y��W�M ������(B�M���y��UH4(��!}f���R<�yRN�.��,�W��<'h��;�nۋ�y��#ob�zՠ��F�a8��E&�y
� \|��T1���	q@�'s���+�"O��z�KΊ1W��:�/�06��Q�t"O�I���O`<�H�`8����"O<92!�Fa��@��$Dd��V"O�]�gb�~_np� >�4i""O�\"��]�2"��'�OL��S�"O�dH�a��T~xPf�u�j"v"O��ж ���  Z�_;%B^���"OQSA�V
Ԛh��-A�C/*�i3"O��B �Z�)�j�b\�T�T"O�C"$N�>�b�S[�<@�"O�٘r+�,s�4r�\�2J���"O�4�F�V��4a�!*y�T"OZh	�d��j��04@ӽSM "O0E�g�*ucp9Q�K�P��ĐR"O���P̛;e���3����|��w"O~�8+ȼbo�a&@T�
���J"OTU��ȍ�ΔC�펰��E�c"O��Yb��F?����O
}���p"OrT�RB���(�0��6J�.�Q�"O�i*P��+א ��l߾�J%c""O�ͨ"�ZP�ŭ�c�БQ�"O�!�o!�V�� �	�q�!�W󄉉s�)�ǓX)b���f��
��� �F����	�Y-h��1�.ZiN�7��80��]P��
���㉸;��CW�c}���-&H�)��K�9=�ؚpe���Ol�!j� |Z���I~B6I6I$�rsd��%�}`	�m�%�iHE��,f��~Z�Ҩ\?J�H�E���+!/�@}r�ē(h�8���I��/k�,�2����[��	���"vT�F)�A�8ʓl���i��L� C��Z�W�^4��H#�����p��]#^�Y"�Z�3�	5'n��K�l�p����%�@@Q���1Ē�*`g�OX����D̼�����H�f�!�T�'s���>�Q�䣱��h�c�nU�!y鲟Of�Ԁe,�3.����o�GӲ�Y���F�`+��-_���'*C�U��	���l����7pE��~J(���u����a��"��	�hy�Q#�?����H)b\����e��*��>�j�Sc� �0e6}��d��A������ B�H+T�+%]FTi��[�X���# �4@��j�ń�����8��P�#n�>,�No9)e���V��e�D��qX��UMܺ�˟r���GO�OjE#��t��D��I� �f�aQm�<���QC̕|�0HZm��ay���/�<%���ݸ ������n��Љ��˰[	օ��N戕���ݟ�� \�&� ���.�m��ȡ��k>]��A�=	X"�3ĨI4f�`���o&�p�Q�b�DO���j]X2��,��x�Ah�s%Pقe��O^��*I���q�"T.Y&bUP*�bbDG]
R�n��;E3P��f���xxPF�pf@ŕ'K��{�AAɧ�'Qt� ����l��IR��&�z��@�hMT���h��Yk��S4��!�	
�哌�N'f���EP�0�p���<�I<��8q�~x⌞�1T&d���
ӟ��秂�K��cҪ�35��g� ��6���C��'�ڠ�7|�Q�S@M����Qx��J���v}"dU��l�C�F�ҟ�9�fMGP�Z��)�tv.�� Űbx,z��R>Q������C��8�f{��)ӈ�"j���
�N�#E0�ٜ'm�͉6�H*2�2���\ⓐVf�OB0S�D�S�Jآ�[�F'��[зi��Ѫ�]}�O>%�s� !YV���T5/�	0i�d�)3e�*S��d �I�`(ϓCP��0�F	�y�4�B�i�	<��'HB�eH� �c-�ybjީ	��ҧu�jɦ��X2��6N��I������>��`A/ @���ق[����4�L�mؙSW������9dZ�@�N:��S�O�D1�G�5'�
!p#MO�'u@�Ќ�ǧI�����ڒ��O��E��.2������#�屋y��"���ɳ$���J�/D�MÜ�A��i��6�V�Tc�H�ؒ��)��!�^�( sP��m
*Pi��;T�!�DD$yz�=Pӡ%g��d�0G�!Ae�	*<	�f�;��y�-Q�O,L���X�t_���#���ܰ>q�=t��Z��������c�?{:����Ɔ+7�\C�ɅIaD�jl�1"DH��U #=I IB%3%H-+��8�S� 8:Ժ�� 4Z<Qq%�	u�' l�h��
n���!�Θ`b`l��)��h9)!��O�)v��.��Oq���0 
Nr(ȩ��N��dS �ԉ:���
��"4�� ��(�GD�v���]�P�ԑ�@��躓Eڻ��Ҝ���C.���?Y"'��
tJ\d8��ܸ:�(���*O �:�VgI��\�c�'@x�ӡAP�es���O?	I��Q��i�
���Kg��b�<��C;>�,Z+K�8����D?��%��[��h"e����<�� �v�CE�d [�-�{�Ԩ`���o[�5�����& hAǟC	v����<o�}��'aD�&IU�T	|���9U���R�����Y��(�6͓�U���~�%N���(@����@�Je�V�IC�<��o;��}�B�0M�P����I��c��],N8�$�O��}��S��04�=z��I� 0�B���8��AC i�_'�Z���z��P����򜑵"�)F�LL�'kME�d���BլK��a���!|Ou��(�5> p��H){>(���O3]��x���G#�����Ba�����
S���`�aY�ؽ�W�;��;u�~HC�V��b!y�����O�n���ĻJ9~�A��C�s���A�'��A[�픽�=�5���s�x�:e��P�Z�A�ڱ\��X
7�G��h��$�o�fp�Ԩ�3�x�1 �3=?!�D�+��M�UAЮt�
��S��I��i�����^
�zG	�<;�$AȔ�ϨO�l�t`P�xPy�6�Y.��H���'��m���hj�p���ҥ
�l���k���9w��-fE4m� mq؟d9����p��Ъ�N0k;��pt�)�I?� ����u�������bԉO�И���Ռ0�~�S�!&qj��
�'�.%�ІR��Ab�N-w��P�qҀ6GE��&3Z��B�-�h����8���
0FS�]9byɀ�A-!�Ω@QY��ݻT,P�ca!k	�
ġє u����=����ϨOD ���[(&s"Ȃ%a@53����'Ls#��8(�L(�*ojzQ`�F�:(=����hDІ�7�O�U�!� �x�9�U�-N�#D��A�|�渓��H�� �c��>擞5}�(@�Yf�����h��r@�B�ɼC��,�� ]
�:Ļ��ſ-W �+�늳lԡ$�"~ΓXG�
��/h@ޝ���P;Z��Ȇ�&K6Es���%J1%�5j@�O�`�WhD�0>�W�۴�8�I���Z�� 3
Dn�<qam=��IH�j��[����P��h�<	��,u����>H[� لRX�<QDK˰:0̰tD�BVeJ6�[�<�B(�*�����+m
BX��hR�<�t��3b� ����@�._��з#t�<5HIO�@�� Z��	����� ��d���� Zݬ��=%?�(2l�":���M�{����7lO���2����X�	�|V��IE#��^�=Z�n�H�j��'EZX��I�`#|�'��y�Ȅ<k�8-���˿	�d8z�{¥��K5!�p��S�ON>5∝M���ɂ��A�!���"��e�Tm]X���M' ���A�Aj²ȂԆǂװQ2�@*}")�N�$�xS��d}�Oj�>��`��~�@�b�#�y2GD5����Ăm�b�	�_ 's@0iӁJ.JG"�&�V�vL�-HbG$}��.p��LY0˛�Ej��[1×�*�z��Q=�H��U �<ise­4~�����I�b�p�@�&O1[2�b×>Ѯ͜����ɷN��$G.��E�F|��E���B���R�Љi��iB�S��~l�%O��d=�7�%~U���5vV�A�'��R���@i�R�ն( ��0��.Pq��{H��SR>=�eJR�?��]!�_��2���-T^�i�]��Xpq"D������CS��:z��P�uR _�ʩs�iڰ6�l�����$_a*�M���|r��,��1�q	I+A�N0@��d؞$-K�D$9`������O�v��!�3�0
w��3͝;��%%��#Cm=�g~r+��*�f���Q��b���'�|M`Ak��Xd�QE�$�@�q4|a3qg�H<ٱ�+�;iR
V ������"]FN!��Π������6\�T�Ť�<���'��D�,O���k�5��eN�j�lh��"O��+e쓃W�xa��g^�"�6��a`�=P�*	%��|a|¢�)j���
u"N�fʈ���ŭ�p=��A0d�~�z!k��[�D]<u8��gDU&eyXA!��/�h�Q�:7&�1����&��'oH�c0덡@����4}����� `(
��[%�\�Ar��S&�����'�8a��7eo�����=-,��3A����FF�.(ٖ���O@���-��<�ĝG��
0M׽R�L�Y�s�'c����(��Y���}���] ,��@8!�E4>p�	�&ۮ���r��5RP��'#h���O%-�<J�T3"���[�'��I�B�M�`nH=�O���elLs��H�V'l6�S�p�\��wIP8m��H�p��B�I�<<
�Z�1�E����~���#>l���A<���iRgB�Ac�}�3d�NR�Ph��ٗn�Vɉq%�o���E*�O)RËK��	YB��:=����;�<�Y���!�t18�Qc�d��#H��*��G�F]�'I��(��"̚ !��ޘX�-�/�`�5"� ؑ#�>�RGa�;v�X!	�ݹ@ n�P�K�O¨SG���Б3$�6}��("-��7��)S/G��I8��
 0t|Bej@��y�Y�fa�0@q�Gg�T>����(V	*\���i:���"�
SC��p�N9[�z�
I��#�	�w����5�'������88���7GY�J�����O�����Z�A4~�\�O>��SÁm�&�b�I�R�����a���a���� ���0x���)�>0�0qACD�U+8(;C�(���33�S6F�O��;I�3H |q��>�'��E*�SK� T&l�����?>q�#>)�H�$ddQ9��$�/,�\��c�U�\_J���\n��	�8��݊��]�"��=t^��Յ4�S�S'Lx�O�0wT5hT��=����}~t����c�)ڧ!:@H2 �/Flh��iz�$ �\�����G�7�0<� L�Ql,Dx@̫$A��`6/M�I�VK����q18��B<�h��f��:F4��3ģ�c$���O���m
� ����eE�W�L����	�nW���}ܧ	("x@��?kG��q�J ],�Q��`��5�p,M�c�ޕAs���S|͕'ĊkwF�E�S�O�4�u���A���y�V܅�2���JE%����%�ɿ:�h!�ȓd��CWh�Y1��$j��#=���ȓ<~��@��
Bཨ��2D�p�ȓ�P�F=�t��%�'T�~I��*�} Љ,1��� �Σ.r���+�P��-J �ܬ J\L�y���"4)�mIl����w+��U�ܕ�ȓp+��a��I���@2�X	��X��z������Ap�8� ]%| �ȓ�<=����(R@��4e)D��G���Kۂ}��].d��$D��("��4MN�o�d�^�;(%D�`!�lG"8���c$씢�����%%D�����=����k�c�]�&.D�ę�.�0��鸅�)w�mТ�@�<��E[�~��9��G��zŉw�<9$�߰(�@#���Qm�S��w�<A�R����h�I1v� C�j�<!P�G� .���!bԥ���p �Ed�<��|�E3�H#t��$���~�<I�gQ0g$%+�*�U�̒��t�<�ƠS7!�J���^�s�<9�ֆG}�<yg�ْv6��uA�YܜAy��Yf�<��3�������y�H�kv@`�<q�L$K�>���E]6S��B�I,���	��*R�������L>tB�	�o��yu����u��匂��C�	�Q���&J�`|��W
L�8B�	-	V2�P̞	gD,q�0���=��C䉀�4T{���� �LE�F��K-�B�ɤ0 li*��!�(�P�B*`Wb">���A�J�|�I�aҦ'l0���<�AQ�D�Ly�c�6���r�CXu�<)���u�ͣ"Z"����gc"T�D��@��/p�@�� N�:��P�9D�`9�R�d�`E�͡K���K8D�X�vC&NI����JL#ZP���� D�X�#���ZVpةQ�)Uv�{E�!D�� �ˁgrzq2!^�AFiu�>D�� �h��K�2�P���)3��(���2�HO�/-�4tp�+G�_�,�����ڲm�Op�l%tX<�AS>�)7�J�H�L�QWAZ��� ��Nr2������u����L*�F"~*�'R/21h��֘1ְ	�Avy���A)��B@K��j� �شm�0���	R��=H1瘔V��ز�I�%�(��Cyr�V�$0�h(�O(�>��0���d>����� I��e��^����\�n=M���a�4��(!�h@)��M;�U �Γ �yҨFrܰ��`�>�S�O��!"�O	4��ѐ �"���A�Y�R��H��^�	a��S>��R��Xfv�y�lS<tzZ��#�>-����uF����X0���Ē?�{�%	�(� Z�З�����!}��U!/�O�d�D�)D��h�_��9�^�$�$e;�S�OJM	"痚bU2�&�L�^����	�g���f��6"@��e��0V5�B�	5PS>���C�o�r�ɞ^�2B�	#w=�$)�障Q��m�TfȰ#��C�I�pqsFмH1�e
t.C���C�	4ivA��,)Ӟ9���AO_�C�	%f�FA�v�bBҴ�-*��C�ɞi�m٧�\����C&��)Z��B�IA�>Q��֍^��4! I�<[f�B�IK�>��q�Q�S��␣��D�XC䉗m78���<$��a����B䉆.R�ىR㍆@X�U)�nS&�B䉸A�DY0�a��a��qC4"Q��.B䉳�v傒'�_�N��s.��6��C�	�UU�ZS��W�taP��K)1uB�ɵuT]�"M��X�P19EN�7�C�	G�\-	�FFI�� 9#&ˡn��C�s��p�SNW�Sg�����@�PC��)
�~, ��_�G~��
n��<��B�I	J}��pq)>b�*��U�	�2��B�ɫVUF$i��!�X���a)HO�B�I=u��Pߚ]�xXj4ٮXs�B�Iz́+p��xif�P��ہGzB�;K�y�̗�Ujݹ6̚?CޢB�	�A����ւ
�rj-C�*��B�I�V�ց[�k:L�*W���*,B�I�l&r�����S1d�a�_�1��C䉐=`Pe��՘0LY�6��/1��B� Q��K�ލ!}0Mc��)�B�I��N���94�M�6��O��C�ɞ@�}�҉+6i�q"���C�	5a�Pt�t�YZ։�Bm�C�I4=R��G�9+Qv��G�۳X�B�	d������1P#�`�"�5cw�C�I8O$�Cp�%1�(3G�Q� �tC��:U�ᓵ��?2d�@&Q^^C�I?j���r�ِg�HX�ő!: ZC�I>"~��T�[.\��T�OsD�B��;�\i�A�O�BfIG��%,�C�,R��'��Q�~�`�j��C�I�N��@��?.Bn@��̈Y�C�'"HшE�ŏh��)gk�f�C䉡	'��*b홲�a��
�:p�C�I�9�@�!�w�jy���#{�C䉉`1z pƂӺ$`jK�ܫbRC䉚�T3cN�3R,��.�v>�B�� ��i�v*� ��p���4Jm�B�ɾ����o̗H���؍2	�C��9`l@ASgG�1���b�
շ:��B䉽Yͨ��I�W���qSL���B�	c�N�`��Y6�Ј�#�O<�PC�'va*�D�����.�ZC�	�K��zeI��ʒ���� g^$C�)� ��G��&8Kl�G�̣gl����"O��AمJ.hI9'�ڰ6Nf`�"O��!����[]�H�����3�"OZ���:pԠ�2M�:"~��rS"O̬Ʌl̠��)8��Odº��Q"ON�`sG�@�4�x0�7T�$Q�'"Ol��''̟xe��ؔ*��NQF"O��!���d�b��Ĩەl�z�h�"O:a����ZpH6���Q����"Oi��<����b�K�D)4��"Ob�[���9aOc��"Or��0$�u�l](��'�:�B`"O�iJe���<Ta(g`X�x�jA�"O��ѣǸ*���qg���(x`�"O����iޒ1 ��U�8��Y(0"O�L�d��#�"E��K��Qk"OdM*�˜�q�l �G�P)�*�"O*�ۅ���A{PyR��	1-����"OJE��R�,c%K��b�
"O��#I� (��!�덽'<h���"O`#��7dƵ�fP#pI���!�D�6sf�ypgF���v�Т�P�!��:����s���zkU�� R�!�\�?)|sq��w}�D����V�!��!oln$ȶ�T>f�Ъ�*���!�DJ���R�I%����3Ƀ�F�!��rvy��CG  � ��� g!��Qf�D)S�G�t<b�o�3_�!�-���S����`�A�"��h�!�UmZ`rU%�>0������ϋ0<!�D�ho*�Ô'Bd�H:RIQ (8!�$ڂb�z�#	�*kpe���͈V�!��Σ �3N�^~���!� �s,�p�+ݮL�˒/��!�d(J��z��@$N`Д��-͢x~!�Ĝ�[#`�QT/?B<�Q�+ȀU!��7�%F�$12Rap�O�*@E@��Jـ�v�Q6�y�R"^�!�=�ȓ��Y��A+j��%�?+"B���<�Џ�� FD��/�=jQ�C�Ʉ��(��(pbNQp�]�n�C�I��h�0g�(4��B( �n�C�I-w�:�y�Mغ`�	 ��=6�DB�I gr���� P���Q,�yTC�ɀ"��E9
�)������n�C䉯~��ɓ��L�t:*0)\B�I2Q�̭�&��/u��1ǮGB�&��8W���0}�pN��Wġ�,;*���5�R�Q�`���h.
p!�ʔ;��ə!h�(����,f!��Žo�T��%I-N���Zqn�1`G!�$Y	^��H@F���x�L	�G3!�d��k5��Q	�az49쟌 )!�$ǴI��8i.Ԭ}yRբ�h�%OD!��G�x�8�ED�WB�URG��yU!�-D��Tڑ�Ώ{�N:�E۾u3!��#{��R��պ ��U�'NS�!��OZz�$e�H���Y�*�Yx!�$H�Q�4���L0J�<P;��Ɖ�!�e��m�b�p�� �瘖q�!�$�Hߘ�ZO U.8u*�H�K�!�DU	@|�� �X�~�|�:�EϛG�!�$�8DN�����2M�D|�sE� &�!�J$%!� �¡vj�IB�C2@!�� h! ᚓ$�J$j4 �
(
ɊA"O�@ $G�-Dm8H���)fr��!"O��6�ܤX�0�(Q�8S"O\��� r�j)���-C��(�"O�E	�5t��S���8?3갻�"O�2!��$�X�ar�H�;�h�A�"O
h�&��<_��{��V�'y�E "OdAAV`�2֞U1  �=Ƙ���"OvA��oK37��4�UD��b���6"O�y�!�@0��D#4�A�/���"OP���iǧ�NA�cmӅC��-�"O4e�&úW��0�]?{��T�"OFiy#K�Jj�Pkr��3���b�"O�r��E�E��0��m�_�$�"Ov���ʝb*��UM��ctPH��"O���Ee��p���jJ��\o��K�"O�I#4J��p趈(L�eZ""O���C�"L
��p�!O?��c"Oʀr�N���@Ej��-<TA&"O|;�$�o�peA��P�R"OTl��	�`xZ�����k�<U�'"O2�´�,6�"��-��ge��ya"O �!1f��B:B`!�NG�aH��KC"Ot9"mY�Q8$���,��"OTQ�!ˆ�($ ��/�53k��C "Oܝ�W��}����/�122����"O*��k��5+<�7O�>B���"Od��É��R�`���*R`9�!"O$A�t�^(�y�V� #Q���"O�!� �ʩng�U�T��dB�p"O��Ru�L�xQ�̛b��G�̜D"O\]�To��.H�	���/=�*�k "O���m�,ݴ�v̑F�����"Ox@RÏZ�,Bb��C���9R<��"Ojdi�G=]��XQ��^�(5F9z"O~U�&��*f�<����ǟ:X���"O�T��(�R��B����R�"O��8��P��扪Պ]� 5�Q�"OY[�,CNޠ����_�N�A"O�-��E>_)VU(����S~��#�"O�	ц�{T�E8#�E�/�d��v"O0�l/�Q �$�-a���h�"O��R�Y��%xQ�M��fXCa"O�!�D�(.d����	����3"OXX�����A�#"�2�j��"O�T�U._dIN]��+�t;JѲS"O�|��GL!�
�
���#2:��"O���ۮt �#�jӨ" q"P"O;�J�>�|�D0b	z@b�"O8j�Q(�0�����_b(""O���Ť$D�6��.�� `�"OD�Ș5k�p�Y׍��7�H��$"O��XqCy�p8��M�~Ųeʰ"O�Y4G̸D
C�k�.��=G"O�й�c�
�[
дH�6,0�"O�=P`��\�
�2�&�62�x��"O9xfi
�aI�m1��Z�Rxj5�"O�p��FI��hSVnۑ~Tv���"O�8J�$j���!MU8>��ɉ5"O4���G�gnA���x�H�{t"O���F�˻
�dY�!֧�8��4"Ot��C�iq � ���z5� "O�����&	��f`�Ȭ�"O���vhC�G
	��U����R"O� �a��E��n|���_"���A�"O����.	z�2�! �Av���˧"O",c�%Z>���rlN�<�N9"O����
�aF�4!�5��"O6��E���*�.�R0낖lp�1�Q"On��0@UG������ݡT΀8�"O2�rS*^%���	�X:M���C�"O����'�葑g<%��V"O�J���2V��&�H����4"O–�M29^JP8��C�+ɲ��G"O�ِB�"�&�Y$�o��Hyf"O�u'�5hfLt��Bْ �R�ɣ"O�Q��H��\1� �|��x��yr�Ʋ�a���(.��rT��5�yRE�H�m07j�%#sv}s�鏼�y�	�9uR���V��Q��4#Ӯ���y҂�&��DصO4B�T ���@�ybCA�:�=+GAMc���H����y�eZ�Z�
� sn�[�~4��eV��y��2 ��S�іZd����y�F�!S���[�,A9zG�i6)�9�y�k9dAl,*���q��I���y�3t P  ��   �  P  �  �  r*  �5  A  �L  �W  Xc  o  8z  h�  �  y�  (�  ,�  l�  ǲ  	�  J�  ��  �  ��  %�  ��  �  w�  ��  7�  x�  � ; � � c  �* �3 \: _D �L �S �Y (` e  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&�-�S��y+ʼ#�hU!�68w,�6nW��y�X E�V4�!#%*�v��o�9Fh��1�$k� G~
�  	Y"*�7r\�烖 �P)��'a�'~���RȈ!vˀ!��o_.OŮ�	
�'=:X:࢘/x.`Z'�'Z�|Z�'�I��*Ԯ�\J�M��O��L��' �'	��UzMKX�(�'<��A�ڧ=� ���J$h�@�'��2��UoP��'O[�w�Ft�M��3v�'P
%�Q�׿����P�ӓ��'8F�P�!J�ttp[��+S8���'^|�" �6C]<�!P#�"�"-��',:�!��D(:9�4���`��'���1�G�"9�.Ҏ�Ih�'�~�{�˅�zt��D�J��=��'�2-��F�j��!�s!ƠnV���'��0UL^>D����7`�^���'�0��Y�'�(��֤��x*���'���j�g�47�������
_kx�Q�'�>�6�,wB�0�
�4IQR`��'��9��-�7}i6���><�B�z
�'Y�02�!�>b�&U�҈ͮ5�f���'X�ͫ�gB�xmc��L� �@Y�'Ua�OM�A�rdj"��oU40���9�y�Δ3��U� 
����H��y�d�#X�&�� �A�Z���(��ǖ�yBl��P
I�L����`��,�yMQ8$������+�F(����y�F\��+G�@I�� H^e�<� �Y\Ȉ�;uK\�.�Y�@�P�<���C�l�.P�j�	���L�<��e_��`x��A7�Y���XE�<i%�T�t���u@�D�^x
��}�<A��348h���=0����#Qw�<��mY�A���BG�:В��D��q�<Wm�.P�ج��I&F>(��5g]u�<���8VȤ�w
!yzM�f�
o�<Q.A/iD�	p�,�L��m8�Dj�<i3��<����S�A�|��[g�<�&�3Nf=릁�!nD��,�{�<Q�QXC��p$�Y�ޝ�"�{�<��ŝ�F�D	q�֙#���`t�q�<!7�.�ν �n�l�ЙWBp�<�P�Y�Q���Z�fO�N��}��Cq�<��g��<��'�H?`���L�m�<A�#�*)���`�#T��00��u�<dH�}��B!��l�>HcפOi�<1�gO>Ax�VG��F�2��Uσh�<9#%���@���b~�T	�GZ[�<����9{|0�d�R�+���e�U�<�@,ȥlHְ��!�:�6<��π}�<im�J���P�9�8�9���u�<�픎!{��x�kٽ��݂*�Y�<I���,Pt�m��%�9M��˰�Xa�<!("~�����D���)�d�[�<2�Jg̎]�	��O��i����V�<! �-F��`!��ի�ش�Q��U�<q�Hx��  J���ԣ��@O�<��BP)2�pJ�٤t����I�<)�ю��<��
�ր��	O_�<i�b۳m-d0���ۧ y�\�&"@_�<B�>VV��:G��m���{0�@�<��M��m>�	�d�*s��]c�{�<�@�By���� ��~��Rs�Gz�<	�!�`X`��c0:Ͱ��vKs�<�1E�S6��ÄW,s,�q���n�<� �,@���8:�$�
����j���"O0֣�>g�2h2ǋ�'d���`"OQ#	�SQ����D�NJU�%"Ou3��>i�h�E '[�]�u"O�t
��� ��$�7ePF3t�'R�'�R�' �'��'Z��'
��	���T���\+#FP��D�'��'k2�'J��'�b�'L��'�$5
�F�>������&��=��'2�'��'9��'���'��'�H�P��J"`��t�ջ��I���'j��'P��'��'4�'�b�'d��
0�ޥK)���O��I����t�'B�'���'P��'_��'���'��r$J6b�:i��� {%� a�'���'��'Q��'���'/��'��$bW$���x,�%T
��8��'zr�'���'���'��' "�'t^`J����;B.���)����'T��'��'��'Tb�'R�'Z
pg�V�K��]���?#B,JQ�'9��'r�'R��'���'�2�'7l1� P���qGI�4�2X�'�b�'�2�'9��'�r�',B�'���@��:u|�	�h
o^��;�'5��'���'��'C��'T��';��)�!��? L�L���!���' ��'�B�'�R�'b�'�r�'��BD�R�{��� G,ݒ�ֱ�#�'���'�"�'%��'l�}��d�O����*��ɱ��L�AS�ip��Qy2�',�)�3?�P�i�0��E�`�B$���مv쁋ULA����D��9�?��<)�7Xrٗ/0<x��;V\Pr��?���A��M3�O�瓁��I?��$a��F����\!r,)��0�I�(�'1�>uB�,��[�I�<2h@ԫ��P��MI�q���O�7=�N����̏D�h4p���2������OL�$d�dԧ�OR���i'���yʩ(�A�a��B`.B�o_�$}�T0��� �=ͧ�?��,��$�V�s"Im�dXC/��<A*O��O��i#jq��yR��?S:\��.T�$��͐��u��O���'��'���>I!BE:<c�If���Y��+�U~��'�N��-�0�O�L��0f(�F��ԦE�!��E����gcj��xy������Ȭ�H���(E�CP��Z�K%��˦��$-*?��i��O��T�	pv���d�WAb�jel�64�d�O����O�!�bw�t�������$���Nۼt0ҩЁ�M�49R������4�����OZ���O��$Òs-Xu��Ð2T yq!�� ?
r�o��&�G�1��'�����'˰p)�� �P��IH����GO�>Y��i:�b�b>i����z� .�"���ڒd�숼�I-KH0�aJܭ/A���;"��'�j�dr�9�̼"%u�e�2zH���?����?1��|-O�m���1�ɵ�����`�*��0�d鑫3�8�	��MC��k�>a�i�6�Ϧ%h���s̠{�$M3�H�!婐JL6�o�<�a�4����r	�M?Y:��w���$&՞X�2вң�J$� �'c��' ��'�b�'��0�u�R+�v�0ф�-�,����<��
�nM"��T�'�B6�&�dWi����G�p6JaX�&4NrY$���شDћ�O�ȩ��i|���
���p�&��"�`��'sf�H+GVjrB�^yr�|�lʓ�?Q���?�:��YKWH�
��D'��Ɯ�P���?q(O�Pn�F��m�	���M�dKM�KH�NX��2pDN� Jf=�'��@K�fgmӔ4%��'8yj��nL2�x���4^�N���g�:�@��%����޺ワ�O�P�(O�2p5DA#	N/&�`PD˜<[,�d�O��d�O���<i��iC������v�����YFC�a�wd�H�I��M#����>9��iy��
��떉E�n������p�XTm��z�T�n�e~Ң�����n��	�]�m�vD��QV��)���Vh&%�ٴ���ON���O����O����|�æ��Z��\�RCɲQ�Tc�(8>��	U��'gr���'S:7=��ٗ�γ�F�(FlR��~D�6g�ަ�r޴;���OhLp+űi9��Y%T	�Db� �rH>��I��$m `��n���,��&P������,Bi�^)x�a�H�D�H@���՟`��؟���Cy�}���Rp$�O���O���b4	=��&e1bw�y��,��;��dL��U�ݴǉ'-L�y�E�I����N�$M)��O���cШ�^8zԫ�<9$�����E�X�$J�'̬1��	~���R�O1a���d�Oh�$�O���)ڧ�?���YJh B�҈�Y����;���0���'j�6m.�i��p�o]X�M`�	d�x�A+q�T�ݴ) �Vby����Ib�B�˼񈣦������?]�E*4�҇9T�04D������ŕ'���'�"�'���'"j�NДv. E���J�B>��y�S�ؑ޴s6���?Y�����<q3�\�_} ����'璩���(���/�M{f�i�O1��(�G�{�\�	�,�~H�0�O�g,2T��*�<�1�� ;۔��+��ćԦѕ'h2}c�	C*%��̌q�\(���'��'4�����Z���ٴzN"@`�
l p�Q��\f`�"e۰J4������DGay2�'K�V�m�����qx��@�\=3��pH�NY�Cg 7Mf����_н���O��\�'_:����� �uYM�~����kW�7R.�z�=O&���O���O6���Ot�?����k�bh�7��T�ׁf�`���b۴;���'�$7�0��@@�h�{p,��D�J�ƏWW�OJ���O��O�|������a�ѡZs�LBϓ&�.%�5.ܺ1��U�O��OH��|���?��>ծUK�^�tLhB�g�<u^T[��?�.OB�lږ|��Y������I_��)ھ �>�ѧMTGך Hw�Z���lyB�'ӛ��#�T>�ū�"7��*��X�;^�����Y ��{ �R�b���|j� �OT1�I>�3��~�PfB[�Y}�t�WH��?����?!��?�|r-OR�m��x�r��3�V$�F�'H���ۄ���8��>�MˌR�<��4L1M�!/��C\������<a�	��i=�7-/cur77?�owӾ8�Sy��ɡ:`�0�<p��4#ݣF�p�IIy�'�r�'"�'�\>Iq��S�=9 L�+����"���Mk�����?A��?�J~Z�K��w%n�I�K���=��&8[���W�v�|dm)��S�'E����4�y�#��C�F��b�M�`��ykE�Ϧ�y�o��)����������O�d��m�b�ԣڳ��-�	��y�t���O(���Oh�kU���]�"�'3򤇨>��!; �D_����IJ�O�Y�'�r�i�O��z�a���x$�1��0,ZT�����H�n�x���lZ��;�H�I��`їΌ&E�H�*�@tqA+�@�ٟl�I�P����dD���'���j�3�F�07iJ�o���'�26�K��.�Ck���4����X�u��)�g	 r�� �7O��mڗ�M�V�i��L��i �$�Oʕ�$ǚ��T���Vt�T�ӫa�P���O���'��Iß��IΟ�	��4�����1�@�$K���6��$L�}�'I66�@h�"�D�O���#�i�O��dFQ
2.�1j#���\娙�1��[}�qӺ�l�5��Ş��@ ��%��(	+�	����2��	(O,��0����?	F)���<a�*Tg�I�u/S�f=�| 5H��?Q���?����?�'��D�ۦ���,ɤ��;����8T��;֣�ҟ�X�4��'r�P��v�xӐln��h��4���Pj,�u��!��AaBæ=�'6�8@�H��?Y)���d�w�JA�ːDh�U	�/�7�4�C�'�2�'���'�b�'0�="`�vX�a
w�c05�G!�OT�$�OH�m��*��ꟈSܴ��_������RX�*�*K)b�4�U�|��'��O�� x��i���.Rz�apE��c��up��ݍMe"���K��W��KG�Ay�OB�'-�hȦq̴�EY;�r��h��}��'��	��M��Ƙ8���O
�'��i8��ŀS���ۡ-^�Nr�'�J�>�&�q�`%��'s�P�pN^/��к�y^�W�R�T1�E��j�~�O�`���V�'2�QS�ʫS0~��Q0,�U9W�'%��'.���On�ɐ�M{ Mٷ/��4 G	"z�P`��!¹3�"y�*O��nZO�������Zd&B_��i�e�(
Ό��T'�Ayb�):��Ɛ�`�Ŭ$Z�����ny�Ա@[
�!�+F�l�Dq�օ��y�U����П ��џ��	�p�O�* cS%-w@tt��íav����h��az���O����O蓟��$Iۦ�]+r��`�k0Uv\h��@�=���Ip�ŞY88��ش�y"/.yp�q�t���h^ q`�N��y'�*L��I?�'�ϟ��I?8yQI��'t �@A�P��ן��IƟ��'�6m�>�:���O����i����`��
qIfL�����|`�O���5�	V @ �[
T4a�5Đ1^����zh"�O�1y�~	`I~Z���Ot	(�ii,���4ߔ��oG&N}F}Q��?��?!���h����¶K�J ����ߌɊ�ݥE<�ď��bÛ��	��M��wv a���R���FKX)3-,�c�'nr�i��7m�� b�6�$?�5����NBX��@hʚ	�P6aK�*�
�$��'<b�';"�'��'8D��3IJ�p$p]Ӗ@�,#0}��V��Qߴ4������?����'�?qRA�&["`<k��Ѩ��A+�nZ�8�I��M;��'ꉧ�O{h�Ru/֐6�R؋ �E|"� �DEܢV�b19�\��X,�s�2��a�ISy�N�~�DrD^4x����b�4}���'d��'�O:�ɸ�ME��>�?���A�4|�`d��h�����<���i�O��'�:6-�Ӧ�P�4=Zܘ��+�`� �i�͝������,�?�M#�O$��n��������wSj� ��6X7$MQ��ηe����'#��'���'w��'�̤ɐ_7P�3gϻR(lp@�<	����6�^����'��7$���2�P�&���G`�H� �4��4&�L��Ǧ�S�ڤqn�J~���-y�V ��i��Xu�9"Z��R`�)5�T������Ox�D�OX�Ě�F��� ��߀3� ��iM�y<����O�˓#���(Z���'	�V>�$C�4e��A���"z:�`�:?�Y�iݴ��f
-�?9�A�ʥg�Np�t�D�e�"L����֬T�t-O٦��+O�)��~|	�A�"�"d�^C8��Bɠ�B�'
��'���W�$�4�(�g�3N��-��[�U�@d�%��?���Û���Cty�i�&���C3"i����(�#>���Ob�vm�mz<�n�M~�c�"p�������  9pw.�&������M7aJ*�8OX��?q��?���?�����	�P3�#į�[������+*Сl�o��e����P��l�s���������>t�r�B%nC�G_P�8��
�բQ���O<�|*`A�M�'�HAY�솂s���#��:�B�x�'�n`;'�Zq?�N>�,O����O�09���"R=��`��R(eJ��c�O����OX�$�<���ia
ۂ�'���'����BQ�L-�lr� �3j��C���I}�hq��m��ē�M�7-N�'ǌ�9�	�v�$�'J�Q�#��ћ6d)�I�#�~"�'�>��Fe�84������,0���'e2�'�B�'��>A�	+Ju�����IB(��E��I�M�7�(��d�ᦁ�?ͻ6��C��-H���N
|
�ϓ����O�6�T5B�6�1?!��_�p �Ɂ�(���b�ؾG���!/\�:���J>�)O����Or���O����O�y E,P.>�꽃�	�R����̿<iջi�&���'���'���y� [HVք���cUy�NV�1�l�P�O����O��O1�e��/2�X�u/�>L����j:P��7-4?	�B�*[�L�IW�	ly�H�^��8�6��G�0!���%R�'?��'��O��I,�Ms%ō�<a$GB�V�0�Q$��+ �����<��i��OH��'��'�"�[2H�<tMQ0V��(��$\�Q,�m"q�i��	�pFE����߱a�'�,!�(Zg��>)n�1Ɖr����꟬��џ����x����F���!!C,[4�)�����?���?1g�i��̟��l�{�	]Tx�cq�ؙNk�1�ň�0� ��M<a�i�6=�V��jy�~����q�[�v��㵆ڵm�lP�CK֨��\�����4���d�Ob��|����"�R��^T�E�2&u^��O��������C�b�'$�V>�ѕ�N=�)�#K�{D���5o.?��V�|��q�S�����%��YI��ܿG�iaC��-)��X�L�3����P���2\�/�Q�I%�B���j]3׸|*�mί}�<�IϦQ����b>�'̈́6-���J�@���?`��"ǂ	j���C+�O�� ݦu�?�aV�D�I/��!�'5	�,)B��ْ^����'[�����i���O�y� �O��'�f����n4�����/bv��'��ǟ���ퟤ��ȟ���@��bZ<V������Nﲘ�*ө`t7M�{q����OB��$���O*-nz�-��ԟG�8-��M�א)[����?�|�%���Mc�'�aY��E���,���S_˒Y��'�X�IQ��ӟ����d�O���{$lX�v�K>�貄�̥y��D�O���O��ě�c��y��'S���*V>lCQ� �.���d��O�(�'�R�'��'�X�F�%8�x��VD )��Ov��%�K��6"擎-����O&�B��Ñ-�TC�� 4�ּS"O�O��D�O��D�O��}���z]D]�Q��������)9Br�����5g��	���D�Ӧ��?ͻVG��F. x��.��RM��ԟ ��՟x3����)�'T��f�	C����|�Ĵ`�A�9Q�%�n����4�P��O����O@�$\+�Y�]oټ���΀O�˓[����yR�'Y����'�vT���̰�5� )F�Pw+�>i��?iJ>�|u�X}�e����6h�&̒,��ߴ��ě0x�`���'w�'5剩w@ɳ$���ܤ��&֩`��u����L��ԟ@�i>!�'
�6��;U�D��آ�3���rZ��S��EZ����\����?�v\���ߴ<�VLqӮ(4�٣m����@?^�ҭp�)P�D7M0?a���''���n������/2�d���Ǳa�:���q���Iǟ������������BB�@ ��B�ɋnC:�!�"�?���?a�i`�K̟�lZa�	�h|L"�A:R
���ퟄt(�N<�ֳi��7=��4a�'tӞ�`Ѧ����$5��zfG̀!*��Q$Q�r����a�	xyr�'R�'��n�pӈ�+��O�[�ß�H�b�'��	�MS@�8�?��?�)�� g�:Zf��qh�"{��uCU��0�/O���f�>�'�ʧT�,���˶	�:I���D�%`��X�6����4L��i>��`�O��O�͒��:�,Z��K�nvI�'`�OL�D�OB�$�O1�0�Wᛦ#	p��̱ �S�k�d%��	{n�%_�`ݴ��'�d�W�������潳����]	DD8"�,(86M����{W�Ц5�'����4��tR-O���Q?:AD��*�?V��e9O��?����?����?y���i
%ft8� ۊ5�V��P���~�o�>p���0�	V�s�������Q ӟ3vLE�g�&eX�+�-]"�?9��O r�'���{�i��d��+�֙)d�̸4\��&��D��Yvބc��*��O���?a�@l%(JW�x�6ѩ�'=5>V�q��?���?1)O�oڛM���Iɟ��1"�.�B&..%&�� yI��8�I���D�Op�D����C*P�
�,žf�����!?�H_�?�HepP�ő��'8�B�$��?i7&�\w(Ii�L1���s�P	�?���?i���?!��)�OR�����ks	�R�� �����OtmZ�Vv(����X��4���y��	*c��]�1 -O�d�ᦌ\��y��}ӆ%oZ��MC�E�Mc�O �X�mZ���� x�;e/̐"�D���9�$A3��.�$�<���?Y��?����?9��ؚ�ДB�eM6��u��ɴ��Næ!a'����	̟�$?�ɝs�
Uk�
Η>凞
i�3'�� ��O��mZ�Mc��x��)H�`����q����|��5�����B�i~^�;�D$p�e���%�<�'��j��a@H��D�_�F����"�'�R�':����$Z��a�4jN`���1��)�����7X�"�%��f�@}�3	�V�$�F}Bbk�Z`�������+ )l|� C���f����&fĪ���n]~⧛�-t���i�O0�CL8�ka�.v H� M����p��ן��I؟��	Z�'x�~M���W6��\A��2�dH����?�9f�V�қ��d�'Sr7M/���^���d�Ņ&P�T�0*�(+�'�l�޴X���O#`-3E�i�	!}& ��,�ۊ\�4�G,<DDq(�4_��e�uy�O���'���73�����B�eӆ�Pt�T*B�'O�ɫ�MS�F��<I��?�/�@��V�_1{֮��ʓ�x�li�Ә��y�O,��O�O� M/�8).T�~W���v�ۺ/��Дd��>r��od~�O�����P�%A�#5��j@J�M��4@���?q��?��Ş���禍�ׄ:?wB}�B� 
Z�X!"Ā���6�$E}2�'� �a�6���E�1n�xh��'pҩS���2O��	
^\p#O?�ɠEĈѣr�A�D������-Y���|yR�'�r�'���'�"Y>]"��Y![TL`aCDڊ��)��3�Mk0G��<y��?�L~�>���w�j�3����o7�$���\�7ά< ��'|��D����8O�m�p�� 6��x�UoQ\�S�;O��d�O��~�|�W��S�Đ�*ӂU^�L+�kS?0<<�0%ğ�����T�	iy�'��§9OF�$�O�1��O�`
p� ��3�8�	-����O ��!��ɌҜ�w�][d�<�Sh�
J����6�ȸ����Ǧ�|Zp���0�	N�\,���=����T#w�����ʟ���蟨�IM�O�!�p�����ꃿ*�d͚��Ҡ,��r�Be�E����4���y7�Z5B��ZT�Z�#���P��"�y"�'U�'�hb�i ��,hQ���؟f@k���L���;5�H#}K��sL&�d�<ͧ�?i��?)��?�Q�7^F!bQ�Ρs�PB(bA�'t�7m7��d�OB�d%�9O�UÃH@�4Pœ����4
�$�q}��'<�|��d�7}�9��#֐/�1U	7"�H1��i\��$��+A�Or�O�˓9!�)JŅP�n���(+�̤���?	���?���|,O
xo�
 P�IYb�=ʁ��/���B�C���I��M�b(�>9���?1�4�<BԴv��b��T�HA2LӴު�M��O$�3m�:�(���nM�$��iK+@�7���u ��&��d�O2��Ob���O���"�ӗ"�����
1ѫ��W�
m�	П��ɫ�M{���|
��
p�ƚ|�o[�	�"�gL�Y������'��_���-��E�'����`O��< h��2��	�eʚ*���I�V��'��I����Iӟ����A���\�p�K�78z��I��'��6�{���On���|jd����C�S�U�a�ޯN����'<�꓾?i�ʟи� !�<y:B=��C�H�W"��lij�ߣMvt��|�	�O<ٙK>9uG�r�eن�M�qԠP���?!��?)���?�|*)O��l�V�՛Ra�<~M���V 2kv`hP������Ms�R�>!4�i+B��B�Y84��QA����p���O�6��,<�6-)?$F������ ����4El<4�r@H+���[&:���<q���?����?���?9/��0�t�mFP��Ԩ�4Hi�O�צ�F�H����Iğ�%?��I	�Mϻa��c�?@�����f��6�}�:���x�)�S�:���n��<y)�qT��&�
(�#���<yGD�`��	������O��dU�j	���41&1���Ta�f��O��D�Ot�dЛ��ߏ���'��?|I�A�FA���$A�!K%�OD��'�6m¦�K<I��_09��$3vI�Nܲ��n�d~"�|D����	��OY����l���B��r�r�,IꝾ^���'�'�������D���i�L� f�YS�f�ҟ��4Y'-���?�C�i��O�R��6H���ʄI���'B"��d���ՐشF�f(Y2͛f��$Xj(:�'�0|i�/��zY���2�@+~׺X��m*���<���?����?Y���?���.d�B4�2���0ݓ�+���$@覝�6̞������h%?���2&�BFT;B;�,󧃒 ����OZ�d!�i>��	�d��#.s���+ehL�R����d�>A�37(Ply��><����@��'>�	4V���H�%pd$ږ�M���	��<����i>Q�'�7m��@���	� :�ȓ�?#��
󊙬^��D�]�?�0X�h�	Cy�g�9Q��*F��6?adE�,
x��yĴi���M�(�I4�O���$?���H�� ����t��G�[&`��ɟ���䟔�	ޟ��IM��i쨘����5s����� ��Ը��?	� \�����I��M+J>ٶ钀;H���m���l�DlYO̓�?�*O�!���c�0�m�B	� �Y1.�\�X�J�,T�7i �?���%��<i��?Q���?Ag�{L �(��W�x�p���%�?�����ĒΦ�SӣQ͟x����O���B�k�1@����"F��vd��ObU�'8��i���O��Z�$}��D�;��9��@K��UEҡd뀘�#�6?ͧO����\���'n�y��C�~S�|
�/Q�J�|����?I��?��S�'���Ϧ���E�2��ex�ɓ q�	�$dM�v�,�F��@}��'C���gD9^��x���(<�4%�2�'sBk�io�&���1�W�<�q���;@FT,^��Aw胱D�p� 4OH��?	��?����?i����D�Qaji�#��U���7�3(��nZ�o0�������I�s�D����� ��Tc���2@NMJ��؀�?9����S�'/��Rߴ�y��Q��
�@B��_R,�Ԩ��yr��86���䓃�4����ܗL���
y�@���)���O����O�d��v_�g��'��N!B[����+kf�q�*��u��O(�'��6�A¦��M<�Ջ@�dՀpS.%N"�� �-}R��<$_P%qS�g��OBV9��g�b���"k�%�"�.M�Ԭ���ˈ1�b�';��'���៨�W
ُ]��L���р\0&�)�)�韰Iߴ1Ev5
���?�$�ig�O��šu~�P�.�"S�pI���$TΦ�K�4G=��璝yK�F��(�A�2����Jٜx����DV@���X�$�L�'r�',��'���'��YgאM�����en���S�Kܴh^�)c���?Q���'�?�NƱ�l��FO�H�8�j�'�0t�����M���i��O1�(%!%�Z
π�h�)�;Xi�س���3oWd��PH�<�b�IͲ�DC�����$�Bx���HS'p;Ru���ײ5����O���@̏(a2�4���d���=����̓u�4��
8,�L0��Nq�F\̓Λ��Dw}"�'"B�'�ʩ[�L�a���S"P��}����>���8O&�d��\ڑcO?�	�?5���M���.>���3�*��bG�������	����������a��G6B�`2�K�[/�x�r��M�j���?��E��lJ����'�z6� ���E�S��|X(Z���xs8�$�0Y�4m��O,��b�i6�����4�ҁ� ���dS�sW��)t�4-"k
r��ty��'��'�bNZ��l̓�D��Bvr�!��&+���'~�� �M�f��?����?�.���Hբ��P���0(H
�V��D���حO֡nZ#�?�N<�O������C6�5b?���e�3�B���f�2A��i>#��'�	'��O
�.޲���Ďu\�����	�����ҟb>y�'�Z7MջPo$I���	Ae��	#$ڊ�|�x���O��d�ܦI�?�V�xk�4�n@k5���[	���W,�J����'��v��>L��f���
T͞+��d�Ewy�+�~h�ȑ��Hm�������y�V�\�Iß\�Iҟ�I��O���i��h^���^�:̉��	uӠ���Ov���O���t�����]�t��g"X�>d������,%��A�4���/��	o�7�d���ìT/{�bHY���56�L��Lg��� �492�	f�	Sy��'}���,8�y����0���x�'��2�'R�'<�ɞ�M+�X~b<O`KGLHpD�(ҫ\7"qZ�:����o}�'�b�|r
9�R܋��0\Va�������_�R�Ҵ�m��b>���OL�$���>�#��J�NHA(�
���'���'a��'��>��I�&A8̓��8X,����R�p����*�M#WGT~b�k�V��]�-�Q���)���#���:5�L�	՟��	���
t�æq�'�H���ljz�	�b���Zs��-t�8:�Y'����4����O����O���U�2���eD�8���Վ����˓=��6�9v6��'�����'C�R���+U 0(��N���jƧ�<����Mkǔ|J~��G�H��QÉ= v�q@]�.}B0�7l�X~���B����1 �'C�-��X�t�^�P�4�W�-1p��I֟�����i>�'��7��?�d��A0HN���s+Õu�a�vdL�F���Oݦi�?rV�$�شq�2�i��0��ˠx;n՚ǡ@�R�z��Tɒ�A�������u�.w��(�\��߽Rd��6
��mДkU�Ӡap�l�Iޟ,�	����	���*�n������b�U��	W*��?Q��?�����P]�i�O��l�|�ɇ8�h�$DFC3��S҆RH||�K<���i�$��O<��i��Ɇ84h�S�.?cU����t��q� ����%�z�xy��',�'��e0ZR����

9�<�S��E{��'��I3�M��!F��?���?�,��� ��������B�*?@���⑟�Q�On�m��M{��xʟA��t+`�8�TZ�B�,�ǥ�0`�7��Jy�O�����B�*h�`���;����$�O?���c��?����?�Ş�����J\ \��E-@�Q��c7�1=����럨�ݴ��'F˓�M+pI��.D^�	��8K�"1���^�����h�TU.��7� ?�Rd�?����0��l����&���U�F���y�^���Iҟ��I� �I��(�O�ћ�j�(H�,\��*]-�Vp谪s�v]���O^�$�O��?��������XE����o��C$�9ׇL���h�~�'���?��4XPn��<� <��@`K�PbV<ؠ"�o�)a�2O�� &���?���:���<ͧ�?Y�"\Q����G�-K�����!H��?i��?��������9�r�V�����X
�<�X�RrD����
��J�FS��7�M��i�|O^=�SC��s�t{')ձ-�tl�󚟐�6E���9�T�<擈����,b�mN-@2"�LQe�:�#��\ퟤ�I���	�\F���'4���O^�0�� ϳw,��;��'�@7MW."����MC��ww�Q+�)�,b�r��N�^6�(�'��'�b��_����@���@8�	@�mw�y���-
f�Z�N�+��Oj��|*���?���?	��T����qN*���RE�mU�B,O�o��p�������T�s�Ph���3R�໐� 	�2��׊���O8�>�󩒸~�.���m�(�d=�t��	����)l�*�_L�X.���%���'ɖ�Av �@��pd�!`M��'d��'����4T�p�ߴPL*qΓ_vaB��מ�Z)�vDË,��o����$f}r�'��'{~��eJ=eY�dz�	;�;���*���4�7��Q>���}���2�O�<*@�{�A;r������h�����ן��	n��[���R��82��`��6]ʍ��?i����H�(��dæ�$�؃F�V�ry�� 1i@��)�"O�I����i>`E@UЦ%�'��	�EB���QEA7b�`Q�B����O��O��|����?A�pu���F�7J���ϋ9S�@����?	+OTl$,�B��Iٟ`�I\��c�9��at���I���gU����q})uӲ�lZ<��S�T�G���M�%+܇z.٫1�Ě8!x����4t�-��O�	1�?��g/����Nz�I�X�U�&�ـ�^�s�n���O���Oz��i�<�B�iv��[���T�R�s�S4��c *u82�'7m<��
�������� �HTbB�h_�ݙn�M���i��K�i���O�=�	�"��r��<�����1$�? �u;1���<(O����O��d�O��D�O�ʧC܊= ��X��B3	�4 Ȱ��i�*4�'l��'��Om�a��.�2DS�dN>8�-3s��P��E�	����O>%?�ـ�æy�,�Uy���;h��h��'%�J�͓E�>�/���$§�����O��ė$td qFXX����uG� kN�d�O����Oʓ)V��$�?FX��'�B,��2��`rqCӎ���!�4��OH,�'ڰ6�
�D%�����?b{dlCb�H�~KR�"?��ćW�@�ȕD��Z�^�� ��?in�% ��
�k�D�d��i�-�?i��?!���?��I�O\	���%�̠Ztk\������O�n��d�l�����D�ڴ���ywd^����b,�c~�J�.���yb�'!�ɮl���lZm~�	�D�=����q��Q�-m"	��D�7A�B��|�T�`�Iɟ��Iٟ��	�����
4x��`[p'ч{��	p�My(k��\�W̠<�����O8��X�"�U'�d�`CS�'t�p@�>9�����O�T�D��{f�4ȕ�A.0�i���3��\��R�Ġs��)GO"��Y�Ihy��zs֍���^���ia��,'`��'E"�'/�Od��M{����<����%��I���I�I�8�d���<�3�i9�O��'��'zr�[x�z��t��`)_�'$N���i��ɤ|/�P	����+&)N5����];;��ɛ�k���	ɟ����x�	ȟ����f�(��J� _-q���C��?���?�u�i�V�k�ORb�c�t�O�����0��v)W[�q�Q#��I*�M#����dT,�M��O�����!�=�vW8v��b��Fx�c�i�Oz��?i��?��s�Z��D�{�&��U�S�n_&i����?q/O
5l�5
c �������Iv����"<̍�a�7V�ɛ\\x��'$"�]����O�O�SH���ւ>�N8	N��E��� ,b6�)���Ay�Oc���ɿ6O�'���D՜�2tjrˋ,+z2$���'gR�'�����O��	;�M��d-���D��s��p�`�o�*��'�72��;����O6��G(	jz]۶��MI0�"�O���[�'��6m`���I2����֝~Γn�Rq�&I������
Xdt̓����O���O2���O����|��w�lS�=*��`0A% S�f!Um�2�'-����'�6=�(q�����%t�(J��W��צ�����S�'X�0ٴ�y�<��A��`	t���ջ�y"��>t�}���OX�'��I֟l�	2pu�̪�a z�~q���f�0d�	�D��ҟܔ'��6-^�H����O��ĒT�:DQ0�]*9�ܷ6&�(�8�OzAm��MS7�x������e&ߝ_-~�0d`
���DL�e�����J��1��Բ����d%*�X�xFY����C�S�I����OB���O�$0ڧ�?�
z$�����Ö�9C"��?9e�iM&,J�'f�o~�X�杁.�����.��Q�PոsJ��1� �I��M3!�i1�6�4@7�3?�ag�b��	�� �4���\Fp�������H>�)O�)�O^�d�O���O� ���i
�Z��ͲYE�Y��<٦�ik�#�'\�'���y"C�-��@��ў�`�k�k�a��?Y���S�'@L5� ♱E���hM�A�̅A�\��nӼ�v��cᯟ�$���'j4�ƽC�@�*Ӎ�$E`���'���'�b����_����4�6i���K?Q1���:�<Y��M�2>�ѳ��j�f�D�}B!{���l��M�'�-V�P9�j�h�*���F�Zٴ��$�2H�����CZ����N�60� |)��_��T�t��Z9�$�O��$�OP�$�O^��9���,{���J�������v=v����H�ɪ�M�pŏ�|2��P����|����J��a!�E�I���!(N>J�O
}m�8�M�'AۮpQ޴���I7d�d����k���#�G�e ~��4�ŉ�?��0���<	���?���?4��6d~(�!�B�[o�,���\/�?����Qצ�4H����I�t�O5|��K1�=j!��C)��O�E�'�7�ϟ�%����:�m��i�4��x�@T1͏*~�~�XD����4��i��t(�O��a�c�Hq�-"H[V\�b��O����O��$�O1���oq��
Ȋv�.I�@eH�e��ʂ��� �aw[��Bߴ��'���4��楘y"1h� ӭR(��Pro����dr�P味Nt� �����	��`(�-OB�9�H2�ՓE/\�(���9OV��?���?��?Y����E+A�Ri2F��t�����I<f5��oZ!-�J�����IJ��������1\�S��^��'KA���'3ɧ�'���׀�M;�'�\�2�I����� �[0
F<\ʘ'��Xj�� �8��|�\�8�I��E��}�D����c fA���A����d��cy�io��-(C��<q��L����7b��ecZ�#���'
 �����<	���?�O<Y�E������F�ʐ4i���@~r���fx��kb�($c�O`���I+$*!O%ߨI����)(�e� �& �'hb�'@��ş@[��hx8&I/P�*H�g������4s8\ ����?y��ir�O���>�(�	��� �T�SC��|6�ۦ ���M��N��M;�O�\�Wc���ӌɒU��q�gi��ڑ���݅�����Oj���O��$�Op��X�V[�K�8R�]:��F$���V��iU4��'V����'@��x7��9Rc�u�v��{�`4����>��i*7�L�)擒bJ�5B�I��j�8k�7If�MؕE� $Y�'�$�� �ןp��|�P��@�$�#k��9�
SP3�q�&�(�	̟������ly�B~�(C�O��XAhĚ����A�4��\��@�O �mZq��k�I��M{a�i�b6M�"��ߑ~�D�F	P	F�h
o{�T�B%,�# e�n��M~���3�4́��Ǔ`�����ɞNTv5̓�?����?a���?����Oi�T�`�T�H�.u8�+��'
��'��7��)S��i�Oal�m�I� ��8���0��A�?1�܌H<�&�i��6=�6�"�Du�V�rn40SG�6����e���>]�E̂=vz�d܏�����O��O��d�=(d4���G�w��@��Ӭvz�D�O��b�֎� �'b�Y>�Qǫ�yL��3.�90B5)�),?A�V�4 ޴�&%'�?��_ h,��(��0 (�ri���-��EV��)���dIBן #�|�B�)Gܚ�AQF5
����2�'tB�'~���S���۴7"Z!ۆ��g�B	+��Le�8{��]��?y�����$�o}�sӠ���L�E~�ܪ���"�x �F�!��4^ς��ڴ�����~�В�� ��ʓ�l�yA�7n*��4G��B������2|O�YB�.��'�ȧdM�,�|P�M���bB�O����O��?�i�����' fC8�Af`��5��4Z~��Hh�@�%�b>�j�g�aΓUX�yC���&$���@B�A�"�de����iʣ�?Q��!�Ī<y(O(�F?:p4��o�#T$"��'�d6ݸX���$�O���N5���Ӡ��0�$�H��L�㟄p�O �nZ��M���x�˙>T@ͩ�n�`���X�ᒈ��$�8b����Jq���'?A���Op��S^� 0����^Mi���~�!��*'9a�;�D��S����(�D�ş\�	�OX���i�?ͻ��l�GLU����sON4yGTdϓ;ś�iw���oZd�<�nZD~���h숴�S�-�>����"-l����X'u������|�R�l��ҟ��	ܟ��I���S�߰\0�R�cȪq��1dGyk���r>O>�D�Oz���$	2"��%EK"<��H#������':��'uɧ�OQrqR��?C�<�jr"�Y=�r��K�%�Ɯ���Ε�/�$;��<�D���;/��u�K�/�Y��A��?���?!���?ͧ��秊:�f�X!�D�� 42D�f�q:�Fi�lYٴ��'dr��?����?�4�E	�j�p�(]�}�������E�J�H�4���§4�d	P��I��Ԡa�O�Y��Gϲc���qa8O�$�O��d�O��D�O��?���)�)=j�܂��U(�@���iy��'�7�3$���O	o�G�+�6��C�>m��(�#N2_Bر�J>����Mϧ!�¡۴��D�'x)�`������@�uj�i���f��'����<�	֟������@�)�D�e�$k߮UR��Iʟ$�'��7-B�S�Z���O$��|�7i7`��C�i�vU����a~�k�>�������� t�i��з<W�P��L�G-Iqeי}N��b%)�\��|zg�O�,;K>�V	NP�8+v)� ��� c��?���?���?�|�*OoZ�K��]�$Ȁ�A_�pc��_�f�V��g�ğ��	:�M��r��>)�w|&,0saX,D�Z���ҏ$\R�q*ON����t���3����"�(O���%Aa����A�7"�i�C5Oʓ�?a���?Q��?�����+$�萋���	=Nj9�c.�~_��o)B�t@��ퟨ�	k�s�x3���+Z��� I�(38|�U�м�?I���t��	o#��;Ol�"��H�I�v� �)��ך�q2<O����5����5�䓘��O$�$J9:(1��	=d��IG�S�X���O���OT�<�f�Ҥr���'jRgQ#��i6�g� ����X2}�OdU�'g2�dͪ9�z��cŽ1��X;U��9,D�I�{Ujɉ��s]�$?陳�'X��	�a��ȇ�L/L�,	�E���8�I����4�I{�O��Ӻ$���`�Q�>��	��H8��GtӬ��G�<���i|�O�nI

ĳ6��-+w 죧��L��O�+f��4��$�>a�\���� 
��1D�$�*-s�C�h�49 -&��<���?!��?���?a
��L{�����8P|DҦG�������Qџ����t$?�I��)�"�[��r��c��X*�O�$9�)�S�sa8�Q� M3��̒��<P�*�;	D�'� �@u���0��|RZ���ЄP]�z@�C�\,��:�՟��IȟP�I��Sy�Lh���Ǡ�O4��2�O(06���q��)A���bo�O��n�\�;��I˟�'�jX�&&�;�݁ &K�ITP�/��Z��֓�P!�������v�S�ߥI�Ň�Y6h���?�D��ic����ϟ����P��柜��w��A~p�6Dz!"�[.�?9���?!c�i��ÝO��cr�ؒO^��q#!\�QM�!-~��e���	ោmz>��"&�צi�'����!��J4�����n~,���Nۘy^|����䓭�D�O��D�O���Xd�$mᴭƈ6g2��7hØ+���D�Oʓ!1��GI9���'�Q>��Ӯ�t�8G��6;� �u�6?�PU���ݴ,ԛ��&�?1{$爙���1fΤ0�Ĩ��G�G��L�wB�֦��.O�I"/�@<��ܔ"4��I�dT�+���`J��OZJк�";3rȐS�1�Z�&�m:��c��EG��Ї�+8a9�����F0|q�j�Bۊ"���6"�v�a�X����i��D��c� q����d@�R�åyjr5a�E�^{v�ꔂ�#?���cAYx�4�K���XpiRS��?
��!��N�r#Ʊ+��9�v]Q�GVD��@x��G�y�������'�P誰��i�$9FK�!m��Xٲ�����8���T���C�Ĉ͘|���E�\7�����%��`Ā�vr���i��k��ꓢ�$�O �O���O��#�Z'i�0`�>��h��]..���O��$�O$�ĸ<a�n���IB�İQL�1,��j�
��vP����t��ȟ����(�.���d�$����*t�`c��V�}�]ҭO��d�O��Ĳ<�'�E���䟼��LC	%	Z=!a�Lg=��&���M#����OF���O�1Z��|�'�H	��3���j,,��A�ݴ�?������s�T��O��'��$�N1��ia�ǎ�Qc8�
 �Q5�`O��d�O��a��	b�1��^PTtj��J?��Zt� ʦ�'ޖ ��u�2�D�OV����.�֧5V���J<)RD�\>t��
P ���M����?qE�����'�q���ʠ@S�J��p�`덲N�N��i�x	ub�R�$�O��$�����'��	
�Y� 9`�o<Z��8�4�8 ш"���O,�+P�Bh՛C�����rEᦍ�	�<���(:�Oj��?I�'9��B҉GY?�X ƸP�
@:�}2c 5��'f"�'��
	��4������a�lq�ρmH6��Of��%B}�V����L�i�Y׈�11���"���h
`�C��>)҉Q����?)���?I+Oj�%eW�=V�U��ݵS0��q+Z�wS���'��	ԟ@%�d�Iԟd���	��+VI��,�A
%����%���I����Ipy��Nl$�ӐZ"��:�t�^8���T�j��7�<������?��N6$�'��P���`�TIF�Y�\�(�Ol�$�O��Ħ<�qǉ�^���̟�0�%S��I�=<���t�L��M������?��q+���{�@�1mR|ܰ�hZ(4(�e:$`�M#���?-O8��2�Ev�D�'�B�O洙��C�"��D"ccK�l�֬ �!���O~��ڽ_�v���Q��0�N�l~�9E��OS2�o�Xyb#Ƥ(�6�����'��c!?I`)����b��i�(aP�lড�'�y+��'X ������J��T
�]�|! ����(�M�Ǌ�.v�'"�'?�D+8�4�K9(Gx���R9�Ι"�HтI_�6��O���O�O�s�x�	^�t�C���m�֢_�E&H��4�?���?	�'�=�����'y�$_?m��Q ��&��E�S�
<Y��'�'T���<y��?���m��hA��e�T���@J8l��i���!l}�O�i�O��O�E���j�qhf�9N������B�䟰�''bY>��'�������.v����!�&����94FO����On�O��Ӻ#�
�(��<)��D6^�ƌ������IX��=��9OL�d�=��3� ���aMT	:�"<S�A"0Jеi%��'��O��D�<�'JFզ�#���:V�����.\s`�&l6�D�O�ʓ�?� ���	�O�p{�
&qN���O��C�ة�Q��ҦU�?����L<r�'e�L��31b	#��3��Q۴�?�/O��dG%@$˧�?��������ZH�&�c\@XH�l_\�	ڟ��'f+�����
ނv�����e9�JǦ����OR�`��OV�D�O��$��Ӻ3�k�4]��<b4��?+���������Yy�
;�O�O�x̡�r�X �2�_�v�*-�޴C��{��?Y��?��'��?ɡ�c�9V��\SO)��Yw
����'=�"|Z�
N�d3ܕ@R.HN� RƎߖ}r���'R�'��MӢ_�����72�Z`Y��g�� @J&�:�،�D�X�'�?��'2��!+8O;ͨ��E:��]۴�?����#��X���DW�9�.]"�ȆO
� 6�B败'��S��1?���?������C�l���	P��f]�s		�cʈ�jT��^�Iҟ��I�	RyZw�̹��AN'Zzh�ȵ��# ��4�?�-O��O ��<9 �H�`���Xa+�Y�)ϞAP�	94����L�IJ�ay�OF��.Xz�!��ry���&x듆?i���?�+Oy����n�Ӟ@�� rd1N �b��G8U��4�?9N>�,O�i�O6�O����}���ިj۴�?�����U�$�$>��	�?������B�Z�~�0%A�_�O���?�����<�;�i�fk�Z1�ĸ6�U�B	�m�py�n� y`�7MBQ��''���??���E������A�	��'	�Ħ��'!��'U&�B���FI�%ib%��,ď�L��󠅳�Mc��,+ٛV�'���'D��K;�4�(��A	n�2�N �/_�����Ҧ=�	韼��|�)��?Q��W =ʘH2L�q�ޝ�m�<9�F�'Hb�'^ݓI'�4�>�D�O��H%�4��Xۣώ�"`�@3��Ԧ���ݟܕ'��g~2�'Vrڭ(�ڹ2VŖPs�,�$��.�6M�O:�y j_�i>q�I��'��1�Lǟx�2����K/'�}3��kӐ��?IN>y���?A.O�����\&!!���8���1-TVQ0�%�t�I��l&�p��uwIӺi�ΐ�ciΥ/�49��_��M;������Oh���O�˓b����C6���h�Y24.�za��/'!B@U����۟4%�������'��X�T�#H�ĥ@ 炭#9�X��-�D�O���?IV�@���)�O�| fN��XFE&e��b��٦)�?�����Ùr��'=�h@�I�z��8�2I���ڴ�?�l!)O�Hsg�C����s��rf�#B�L�B���\��R�c����?����?������<��#h�̺Abr�e�f(�;z�mZVy�f١Cs^7�\���'����5?iaU�`��pu)����z��ߦ��'�Л��'K������V�Z�EQ���a�_>Q��Xz���Mc��A09��'��'���O�>�,O-���{���kg�Ì.p�P��@�Ѧ-A�z�T�'b�i�O����JB%g������
Ywe�N�Ц!��ӟp�I�6����O���?I�'�4�Ȥ���r'�\衰1�����Iʟ����5�d�)Z��?����j�*��&�ҩ��C^�0�`�iD�hx꓎��O���?�1RB��p��ʤAsH�8���[̜�'���'�B�'A��'��s��0���<�:H�uOB�.�Y2j�4m",(�O�˓�?�(O���Od��O]�ك�j��R�0`8�a��X����T4OB�D�O����O���<�%�3H��IT�e�ll2�E�E�a���|̛6\���	yy"�''��'h6�r����s	�Q~���34�E��irb�'�2�'��ɟrc�l�����dΥB4��gB$!���
DXK.t�v���<���?��xY}�O����~PJ�) 0_�H�Ʉ�����'��[���0&P�����O0����A��`�)DJ�0)���)����n�Z}�'���'��ܓ�'G�s�`��|�@`x�nԈO@1Ƀ!ϡm�N�mZHy�_��7-�OR�D�O����a}Zw����CE2o�U
я^k��Q�۴�?A��0BQϓ��˸O\��8�LY�U2ڌ�c�M�_��u�ٴ-�"-Ӈ�iA��'���OV듪�DÙ2��A+!��p1x<P��G�l���l��ogX�	Ο��'�����4��+3�]�k����D�7�4�l�ޟ����������8����<����~""ؽ}�h=Y�$�(E��-���M�����2�?i�������} �����[$����-d�5K��q�`�$�"i����'��	��D�'�ZcŞ�:�F�7)���� Y�X(�O6P�79O
���O���O���<�7/�7Fr�xH�;B@L�r��}}j}�W�@�'�rV�D��՟l�	#. t�1��0QX �1ǀ%��J�s�,������ៈ��By2�_�yM��'ʔs��[�|}�RLZ�C�r7�<����$�O���O&� P9O:��S'ʩc�l� th	�]y�4���ѦA��쟸��͟��'��@34j5��^8)�G�:(�D��!��INŨ�i��|B�'����yr�>1D���^~&�JsO�Oj��R妵�I�L�'��I�Р,�	�O����Y�? &4S5o��2w�����z�<4s�x2�'����m�b�|"֟���l<2b���ʖ.	b�鳵ib�ɧk�vٚش[�؟|�������q���1�N ���c�^� C�&�''�b���y�|��I�(h�"� �Y
2�tI�Ǭ�)$4�V�Z�f6-�O��$�Oj�	L�j���� ��,� 
E�=Ȫ8)W�i�T ��"������bt��S�FA�VD�HG��M���?���(������O����!v�p��*��tz��)?�^c��B��-���I�X��+��8�9�� @ T��c
+�M3��r�דx2�'oR�|Zcپp3�f����pq�(���i�O>�!�6O$ʓ�?���?�(O�y�me� ř.Nj]�fL�Z�6�>����?��x�Z��U :#�L9[�N�(�����<!*Ob���O���<-n��(�O�&4��+"��dN#��y��O��d�O8�Ok�iJRO�g_�, 
���a�KBD�:�;a�><��?����?�(O:��h�g��*v^�r�I�(�x� 3��D^�k�4�?�L>����?�!��<YK��A��މ_�+ϒ�Yt^D��MK���?�/O��K��}�Sџ��ӛ{RԈ)b��b�� %#S�9I���I<Q��?)�&�<AL>��O| p� �����G�̘5D��Yڴ��H�g:�mڋ����O*���Z~�ڢ9\�2a��x��<@ҟ(��쟠���ß8%��}jc'K8)[��3�K�j���%��⦽!�C�7�M����?)���2���K8�%X0o��`��@�q�%�X�o���|���X�Ic�V���I�0f8Yq��S�0�D.e��4�?���?�����P��O����Dx3(��5�Ju�fR/�pv�`��OD��ǍA�ٟ��I�
�L�l��&��A#b@:w�j�(ߴ�?�����$k�O��+����w�
t�x����ؙmۚ%A0]��X4!���|�'�r�'��]�l�gY 픱BqǙ5>%	�6[+��H<a���?AM>i��?)&�@&N�|Xg�Rw�Ҽ9 �D�[������$�O����O�˓_����<�nt�"�E=D֬��ʈ&l>( eX�(�	h�'�R闇�rFȚ����5�Q�ag^�`2���?���?�)O�zt�a�ӹ:0^�����3�����D�{�`�R�4�hOF�dF�A����!}��;�`\��A.�\k�H�&�M����?���?�g*��?����?	���bG͑@S�-��%.:�+D1��']B�'sB��ᇕ����I�<\hAQpBW�-�]B�
_���P��	����M��?1���AS�֘L�\d���lv��߂rX<OH�R�G$���?��OƥYu�7��U��#����i¶����'�"�'"��O_�Q�4�/��	i�cU#}" ��'{�0�i�b8�3���ܘ�����V�_���c2�!w���kC�_8���o����I�<I��Sڟ�Im���'y�$%mȹ*�C,�I1�ٗJ̬�<�b+5��O#��'E��Nta�#f�2Ht�hh��V�4��7��O�p���X�i>���矠�O*, s�L�w��{�E�,9C���E_���#4�Iȟ��	П��	� X��b�ؘ$���xv|�aE"wf|X��͟��	矠��A�I矤�I�^M$�0���g���a�)bҬ
���,���?q���?���?!���?ɖ, *���CծR?"�ˌ*4B��'B�'��'R�'1����O�0bt�з��Ѓ��r���T�x��Ο��	�4�ɟ�@��I��T���;�D� ��?�މ���Z3I�Z,��4�?1J>Q���?���NJH�$�d�7'�E9���5N�	-3a�d���O��_ ��$����'�4&<B�@@j P�DM�dP�(6�'�I:d�."~n��.���� dP;�a��H��*�86m�O��DC�pҘ�D�O��?y�����"��C��1F��A*��{�N6��O����4v���������Y�*�%�v�v�k���`u��g�V��6m�OX�D�O$�)NW�	�̣��M#�d*��k�����KѸ�M�BNDI���F�䇑Nap���v��0�n�0'�\l���IڟL+4�T=�ē�?����~b���+ �4� $��S_����E���'��y��'P��'[��Xs��1`d��0�TY���	�a�H�Q���&���I���%��X,�X�#��D�u%i������	�<���?�����dʺI�:�qaS�,�l�1��jp��&�Y�����I]������	���T�w��b�h����*&1HƂ,�	ٟ �IǟĔ'����DNy>-bUJU�/o�x�æӥr
ֱ�q��>i���?�H>a��?��G�\}�C[�Ju���:����o����O����O�ʓJ�
��w����ácF���f�5rϬ �V�y��7��O��Ol���O���!����J����cT1IJzi��k�,뛶�'12�'}��3������?�ud��|�F�������G���ē�?!�U��Ib w�S�T�3�΄C� E���`UIמ�M{.O�t;���릡�������L��'��n9Հ���i�%u`18��(�M����h�3�@6-^��@G��!�`�s@H�0l8��Gڭ�B�'�=O���'E�P>i�
� B}���K4*djW�A9op
@Xr�iX�����Z�����$��5Tb[�iU&nL:$#�bމ@Lh�l�����	Ɵ�y�	���?Q���?17�F
��dgV�/���d!�y�O*)���Op���Ov(g�"GJhS��>&;��
�ݦE�I/I�`U�O<���?!����j�J�;BŤ�X%֕O�$	�\��k��*�	�.�>݃���ڐ[q�\�n�!r#�"L���"O�� ���(u?j5�q(�����ɓ�L�z�CV��T��m$`n���ы_�,��`��z^�9�2g�7*N�1P��	j!���$�$&o�,��s]tLUe��N6�ña�)6`ё���f�v�T�	��Qӌ���Aȧ��W�$�!С[;�  y����j����-�8k�x��
)�6�D�[�D+���3iWH�ʕL@��r�k�O
���OT y��2���*R�L�YWBE��k������$v�ኁD�)W��ͽ�(O|`:0a4aⓂ^�)-��.@�9�Y��mJ	�A��E9D�j��ڴ�(O�A���'��������$m��U8�E��ʄ@�'��rҀ�64TLE�"�6� �0>�x薇]��dj���A6�q�G�?�y­�<�|ꓞ?�-��w!�O��$�Od(W���z�����R]Nu�4H��G!*�لH�3PE�m�F!���ʧ��?��e�3���Q�_�orp��_�4�0ѕK5Z2p��J8�6���O�����2(@�3COH�)d<<y0���IȢ�D�O��S�Q�	�%�Z�zP�7(M mZ�hI�+�C�	1*�� F^�o��|{s�ȵ�#<A��)Rf႞\���Q��>k@]ؠ�S�?I�Tȴ-��˅�?���?����N�O����)l���T,X�L괪�%S���I$ٜ鱁�G�^��;vݟў�4�Ѽu�n�� 
&W��H
�jX��?ٕi��`��C��ļ7͆�3�_R��"��V:ZYX �C�g��|����M�	џ�G{�_�px^y���+�=��� A���y Ÿ^��c	L�_>t�p0,�h��#=�O��	�T|H�4y�r�y�lE���I��)Ml6����?Y��?Q D��?i������ޘ0bI�����\yv��
�v(�n_�;��Z�H�Qc�y�(��[3�	5՘�AW�÷_��q�7�W)O�A�P��B��yB�W)�?�g�i)���|�
��̠Ofz4
��a�"�{��9O�@Yv&E.U�F	Z7��t"OFu�5�.f���PN�,�4O�EmZ񟼕'�p�ׯ�~*����Z>q�@��3�Z�|���Y�u5���-�O����O��)�C=��xòe�Jô5��|
��ڑ|&��13j> �A���L�'[�AVd�K@�� �W$)G�O��A��:yL<(Q��H���+��I����'~�8Z�fG;4z��Jl�6p��5!8Op���KOb����`BGN�Hqa|��/�D��c����aJ�.��ahG&/��D��rp.�'<�\>[�̑柸�����D;ʱP%��3M��d�4#2�fPqڍ��G��ʧ���?U��.v��9q�ӗ?\�q���QWrT;�*
����P#�n?E��cj0,�1����v�Jʖ���1�fò�?)6�i�F�S�S�?)�'"v4k�)��8f��⥨
9�[��Up
�3}��!���,&Vf�� h-瑞�K�O
�!�5rw4�k"N������O���X�*q	���O���Oj��XӺS���?	�oSu�T�k���j;Р���N?9��	s�����O�P����>	2$�ePP!�D�%{,�
�@ţ��׋t-�5����v��,��>�^��I��'���	럌�'���4�	w"Dr��:2�P��'J1��可G�ܭ�ïݾ'�[�O+�S��$?�D�Q�]�q��;B��$D�!�d��ndH�$R*gM���TV:�!��$'FY��#M�p# ��!�ʤ�!��jٴL{щ�	 0r1(���O!���R���
[�A�d��O���#
�'X���H��=�ݐa�M�Y���
�'9(��7�E��5�ЭŏQ�f�8
�'���rm	2y;r�8 ��N�=`�'�- PA��^&���&�$?X�E�'4��K�"zY��iO�V!��'��I�%V�<�C�h@���	�'�<�rQ
]�l\�(�j\>9jl\9
�'��Q�f�����	Ʉݠh�	�
�'Z��R��b>�8����:cK��	�'��DE�'iE k6�����,[��� �ɓ�
��i:�)���(%��"O�۠) UFD=d�S���	�"O2����1��<颫\'4���2"O����J1��W@/4y~�*�"O�t♤2|tZ�L�-&Zz�z�"O�H
UH��HkPa��
�#eU��HG"O���F2��xЋG2/�:<��"O<Rg֖n�Y� j@�i�9�"O6U��&�1���1�(��m%h�"O��@	�M�pD��T
~�p"O���cY5I�D8�W�ɞ3NS"O�U3������ނl j�y�"O�� �3s��8	�l*V"O,}R���a��<!d��P� T��"O:eyA�9 ���)�Ɓ-SE\���"O��F��:[�Tq3��4d��#"O@V�3{����b��Bzn1��"Or���DV�~�H���S�����"O�XIBC��a-�Q�p.�%��� �"O�����ȻvE�iPЍ
9;"�۵"OD�҅'�S+�!t�ѷc���""O�<�q��[�8
@����rr"O�c�!��E,(�����1��"O*|�Ɗ�$و�f��\�V��&"O��J�L
����Y��t�"O�e1�""$�C�	�h6	�v"O�,�!�������3`C\��E"OL��U��j�H�Hpb�6}�B�(�"O)HgHP�"��St�O�S���"u"O�HA�F��DHrS��>m�9�"Op(K�K�Q3�A�KF<Խ�"ODٲ�n�0&�p�㜣_��p1�"OL�j �cgb][S�@�(.H"W"O&�D&��J�j�G��t�Ph���d
�] ���Z؋�Lʙ�$����3%���*6"OδӤ�Ψi��%�lHkTt�3�My��
{��|�'�j��؉y��T%�(�����'1��֢�+{�0� A��Sh���@�h%���$�"[�D(3��-i��t��8qA�z�nJG��'FZD;@D���dRQ�	� o.��	�'��}��/H�$un(��HC�r��҉{"�W�_L�O�O����^�t���@ f���!�'{T�X��<J^��Cvl�K4�i2G$�� ?EQ>��:Ih6�C������w�d�ȓV,���֌�Zܭru�O^s�alZ֊��$�&]���3/��`�Y���.# !��/�h�c��=U��sGir�z�'��9�섲��i{R�5y�!`�'�$���dZ�n���a"\vY
X��'��)``�)��i�ڗq��)8�'5����MuE$��w�_Sx�]��'�hQ�'�!.�Lh��:Hy*0�'�2)��E��<����)�82�H�'�x`���	YtQ��ʍ1$èP�	�'�乕��#I�E#eQ��''F}[�5pa@�h�,L+Dl��'���س��7Iʪ������tl9�'a"�� "������R
-R�Ax�'�`�dB&M�n�)SD�,2$�'���#i���#4�5�5z����#2�#~��"�%q�]Ia�J/�D� ��R]�<��E�X��B�����"�) ݟ$��
�S�S�O���(Ӊ�6�~ȓԄ7'����"O�}q�׸]XT�2�����fZ�@�`�J�� ����h��$d�Yg�ů0g�Lʶ�'o�l�68OhCPoӥ#.�8�_G�c�"O��!�RoZ�����A�(
��	=<bd�D��s��)�꛲c��)ЍY���5a=֤��4bU���{Q>E�V�S�"m�".��v��FE1D��j�(�'���� � �������R��\"A)Ɍ^��IR�����>�O�8`e�;}�41��u��lic
Ob<�b�הx^��R��>qp�M�A�hm����,-zm���0=�����<��t���3P�U	�M�_8��*S�V2b��`y�%4w:�*'EX�x���Ԡ�N�.9����3g!���.,:l�+et������}G�'���y�!r��=�6ˁ2&��!G���`}ܔ�S@��9�D��yba		TDh
S��4bm��!�\��yʐ�(+P=��C�����#N�.|�B�%/`@yd�P�G������7�B�	�v���z�/�3D߸����ٻ,G�B䉻L	���dO��\�Iu�YQ�JB�I.;�((h�+U�c��<����j�NC�I�@�X+4�߄r}��0ƅO8�C��>In�k����zi�"G��y�B�ɭ�ģ���m�x��P/CϐB�	��"��$5خQ� �N�P�^B�ɣoZ8����ُy���R�D� v��B�ɓu������<kڨ�b0��9?�
B�%�VL�W	@�!�����Γ�7LDC�	/bhQ��[o���E�:�nC�I}&��<##l�p��V�"I8C�>>�6x���0Z~��0�,6ZC�I�Z?
q�UF�;#�����[g��O�<�6��_o�x��
�m����.�T}�*٦��?I���y�?f]��ݚ:�H�!���x�B�'e�����C,'�#�l���O�ٺ�.
i��b>��.4>�ꀙ�9���7D��h��K�H���Ú^(Ⰼ�<aQ�:
cjaH>E�TE݌)�l���_���)P�9�y�� @�$��3?���2 ����;���r����0<���Ez\X���>d) �3��Lg��T�Q�	�48�y�cF$F@t×H�=_��#�\ܓos℃@��H�	�Qτ<n��r�\<��iu�'.�Q�$/�1ۘ'�d�)6 ^!_� g֥�D ZRA�"���q�@m��s���0T�-�%pp���<w�Չ��$�O�ԋ��
J�@�G)��k/z!�c�N�Y�����Ϡ=����y&����'0�;��^>,�JݫCИ3�je��$�Eܼ��'�1%�T�%`�945�q��̩-��ՙЮ�Vb�	�Ǌ����ȓ �	$��6oYt,q���=j�&�l�d	tU�b%��aVԻCE�W�,q@Vg���3��.��z�'э}�H݉D��D�<��J�^	�&��/{�lU[ǯ��+4����h
z��c�G�1|*x�O�AQ����0
$�$h�O2(��@&ma}b%�R��=لn=�*����פD~�Z��G�V��`҇�ҫI�~L8D�G���z�@ޣJ���Tfߠ�1Y�
�=�HO�8+��@��,h�g�*Jp�-k�玱FrT��lހtξ$ 4BkA����Ww�<��MƮd�`;���Qb��a���Ba�G��-V��9��E֎$#|���k��ck��`�&ϑ�y�
V'*�p����.Fi��˕��\*`t�V���?a�.Y�\	(��ɟ0�ى{�dP0~�@�� G�sH,*@���=�q���hu��ـ |���f�,?�nU1E^�j��Q�B�L�>�����F�P����	�.+���L��)���	�%ݿK��b���-͟�越I�AHD	��!�O�'*.�)��	;�fAئ�G0i��ąȓ7K�,�MA�N<��kŒa�"-{���-PU�D�ԣ	<V-��R�OC D���^̀E�޺(�a�N��W�Ԅȓ5���Y�������@D�
�n�!�I�E?�*��(����B� �u	��>�IG*T|T ��֝��Ya)d���S�^)AI����¨��YCcWu�̺�e=`���a�i�t�@`sQ_���"��d8���	���hD�f+�	k���5�:��)+L��	1�
9 i��V�+6��T>I�� B�#G��=|��rK*R舔{/�Px2A��F�0�Z��E�Dhc�bЯ/�48h��e�\�r�E�&���ݟ0�V�\��i�O?ѷES�dϊ#B�<R�R�"�F�}�'`T��7E2�'G�	��P ��Q!A/�'�Ƌ�Kg�	 lx���
��ɔ$�H�I��kI�PV^�i�k�.���!�A͠4���ԙr��c��'"��pYGN���i��ڋw��$@�mʒ��M�D [ͺ����AtX�-��`ʴ,��A�S�;k�%F}b�ވV�@Z7��,t�-Jc�Uv�������qK��F΂tXt"c�ΨH��a��1���qѸ��%��
�)Wg�%fl�����;��˓O����O�k���ϼh��P�!r������F6�@�u�Z�v

ĤO찀4f���3@ް����V>'L�ҪĐzi*�yF�"�`#=�+]����c<�r�O�L)�눳#��q���
C����挾��%�U���WJW'Gt���q�ɱ:�SC@�e�tq�'�Ă���a
���$�S�QA��*B0.`�
��p��Y]&2%�������L;"�ø_u�����L^�m��Ĥ"8��Q�G0:�����&=��M9��$5;�^t2�o=�"�Js&̵KC2q��D�<�%�t��]��,{x^u0�gc~reQ
�p<���A�V9"E9��,��e�#?��1�'���["*Ed,�TAϛ85ҌqC
�a*B�B� ���' �	W �bp�T��*^�t�\�n�".�H���Ečo��Te�]%b������*O�:1�'�6��ꈆ~�|���iN ^&�3�OZ�3��ˬ �<M0K�"|*bGR�:
x�fM�OAj��B&	L�<�"¨~�v]���
M����!��~��'5 ��%�P�g�\��ك �;2�,�➥o�C䉺{l��V���-��!
��t,B��!=�h̪��?���f�1[�PC�	�U���#��V����oРk��B��^�(,�Vo�X��˶ȍ�BY�B�	�)5��2�� ňW ,f�퉀"O��J$h@��dt[A,�"HxՃ�"O<Q�*n[r�x�I �����C"OT{`���V�pIyc��4��|s"O��R��<@��3$�=ȵ"Or,����%���C� U���Ys�"O�rĪ%)��H��Rpܐ4"O�e�c�WYk
�HBmA�HdЩ��"O܍���U̈�uN�?Ur����"O2- �ˏ�}(�)�mPnU��B3"O2`�B��xOj\u��@"ɫ�"O���aB� _v�E��'�;�"O�)�@FY��cʓ@�y�"O��[�m�_�L!IU��p�0�J"O~�jflD�>�2K�$U���Q0f"O��H��q?������2A���:�"O�%� �89����J���"O4]�a@2�H��dd�|�|i!�"O�Q�(ݚG#0�k�m̽\QPi��"O.t���U�k�
�BN�Nȕ"O\��ՇS"?r�ĈW�P�T�+f"O\h҄�2�x`�ŉ��4���"O�L� �L�D��zEȢj���It"O�!��6A�����W�Е"O�}ڴ�"��)4��&Y�e�V"O�0���lX�ɰ)A��t��"O�`�㔆s���p%��$ўt�A"OhP� <�<Ug�*W��ݨ�"O���K�S�Ѣ�E˨�p�#S"O��y���08�,��$ڵy6^A�a"O�	�ɇ)=(h
1NK,(|�K@"O����N��D+��]�F����"O:Y0��X�vL!
�-��1�F"O����nP�i$���t.U�D��"Oؕ�:�m 5n�hz���"O�tPv�Q��q:�O\�(mH\�"O�`�"1�$�(W�ͣ>@y�t"O֥�1c�ޞT�G/6�5d"OX� I�H�8�d��GSށ�"O� ����H�O�Z�f�4<D�;�"OPJ�,��B���@���xK� �"O4prW@C&�K���i2��c"O����q�9`�.�l�|D8�"Ox%��-N1l�X��7����C*O�р0�F� ���c+.���'�:|��#m�2t���D��b"O�	���ԁt��)���@��`7"O��b�G�J�r!@6�.d@���"O2�z"��+$���+�$F�00�,2"O)�S�R���!�R~�b�"O�	zs�B$c��s�S  �N\��"O�jBhW�<���a������"O*� ��Ă2K%�g�7e-:!��"O�����olJ�y%�ÇNLDC�"OT\a�G�nX�p�f� m���"OPśRA�{�������}�	�#"O"u4 9�գ���wԀxF"O�	h�,<���GŏQ�T��W"O`5�S�^6��:#�l8�Q"OL�`a'��,W�1���%}� hf"O�qp򇐓)d�|������T�� "OVx��<�xRf`[a��h"ObPЃn�@<Z��%�-MP���"O*��*I,(z���OK
Yݖ��"O�4yv��s�]X��M�9ø�A"O��)���?;)���'� P�T�"O�-��C,{�0�c�� *�܉�"Ou���8�ډ8�EX"~^L��"O4����J�lF� d�#�p�*O����H�^`q����r��)	�'͜	i��A*c�zy)ԆZe��p��'��C%L�-#�Ҡ����b2�k�'0x��$���Rm�* �]&�y��'�b��G��u���N,
D ���y�C�;�
q ����d� ���yB��u�)Ag��7@�d�k���yr�ė^�F�:k5d����y��:/��t�r�Z5R��iC��΋�y+M�	at����=x"�h��H��yR���P>�A��>̄�eA���yr�v$�g0
��o��y���U���� h %>�a��S�y�Y N*^L9RG�O��Q�F�S��y򄗦@J��%#M�����P+�y���5IZb��?Ը�ʚ��y���}Z� :�F�-�`�C�y%Q�L����� Q�+r�q�A��y�hH(nht���#�Z���|q��~Q��!�C��P�8pb`���ȓf�Ƒ���J:i�.T������v�ȓJI���!%g_��D�N4�Z�� Ĵ�4��"s�1IcĔq�*��Ɠh�L1��T�6x��qH��(�*���'ONu10�NX~� -�:�{�'��[������j�%����'�DY���;[H������찄�N��ԓ��>c�ި����?`��ȓ& ���f��v����O�o��P��K^���E)̀s� ��2P7�l�ȓ(�QD�;Z�t�3�A�	0��``���-Ɔ;��頄�=xRU��Ў�R�K
�1�aB�z
d�ȓA
*�qc�ő,3��YR�Z�s�݅�S�? ��B�dqb���nڨa���t"O������9��G`P�.�� �"OL :禃,wd,!�����a"O�HZ�o�'Y�N���-�W�fՂF"O
4�E�7�LT2�-� Vj�Cp"O�I�#	�XP�|z�-��0O���"O���T�
i�.tZ'S:���St"O>H*񣒈?$����H�H�zU�"O���Ǡ�&i|��S��үg�R,0�"O(|��/�V�B,Ɛ��H1��'{ў"~0,��:���x��L�R�A�4�֣��'�a{B�N�k�(r�ښ���!Ä�y��UɚY"sJ�`��u�EC�,�y�M��b� Đ��L�KH�#�M�8�y�X�F�1p��Fz���1D��y2-��u�8Ao��廱B���yD`�
Y���׎\�.�J�8�y��BW��	���	W���s ����y�JD���,�i����rg�y2JM--�\���E�=�>�ۂG���y�.��n"��&��Y�Q�e�yk��b B� "
�9>d�%1�g��y򯜾$�|��ք5DT�r��:�y�ǖ!��ỡ�5�I󔠊��yB¶x>�ѦC]7R@%1qf�%�y��*j$�WF:2�����%���y�V���\12�a� ��/�y2�5��� A�v�\h3�V"�y���z��A�F�i��	8��
��y2�Z sl��g҈fɼ]A�͎�'�ўb>�`��N6!ft�w��\Q6�"D�Ȱ�A��u�d!pw!R�_y8iPR)>D�P�QI�2#��ځ��X`��<D�l@4G� 
�<y��L[�a n�1�M.D� ��o"w���'�'�2��"7O�=9gMD�5�^Y*�ݞ6���3jj�<�q�K
��WA�B�� P.�o�<��[c�v"��v�Э��oW�<y��*ZtfT���ǧD5:�!)R�<�a�֒ik�G}���H3/%D���	�3�<�q'K�=mr��Dg7D��/�>>r1R@�� ��65D�t/ۋ[q>�F���Lb:}���2D��Z0�@Q���c%� `R'$D�$���0�8i񡧍�V�cp�#D�`�fR$r㺩Xc��;1��ò�"D���G\�c�f"\�R�Z`B�	by������2���J���C�I�{nZ�!"�τ_ٖ�
�N�,b����hO�>�Ī�*��4!%��*a��45D�ڣ%V��d����X����+2D��zV�ӜUM~8�#E�!�D��*1D�|���T�e�S�<m�Բ�.D�t0e#��JbR�Š�P�U�,D�<�Aąd���@�ɕiq��W�(D����N:Xذ1s�Q
k*�P
��"D� ��K|����吧UOX���!D�D ��]�;�,e
�� 2N��v"D��ʗ��F�$I�TN;_�*�I� D� ��'�+b dTz�mO�IF��4�?D�$x��@)@�Z$�#�	T'&��S�"LO��0��뙴 ��B^�Uv��&D��4�D�E8��T��x�Ա�@#D�l�WŹ���#�e��P�UC&D�� �$�ӭ�Sc�v�@l;�Y��"O:
`	�1&)J6��	v��%"O�fAD��j� s�=��"O� S�mH?"e�A��!�(#`yi�"O����m�&-����K�]�� �"O�D�s&�9�����*��q�$C�"O)�c֬w��1��+A�(�H��"Ob�#�R=��=�pJ��
)�"O�|����r����˕e��B"O"�p%J@�`d((���$*R"O:m��Z
�:$(^�7Β��1"O�e$�R6v��ɠ�%r�Z�a�"Oƥu-�֦���EP�Q`��D"O�8�	�7��A���8��h"O��R1�>�p�$@�-qz��T"O����&�O����"� (;��-�"O�0�S톭��А'#[�T��Q�B"OlT���lP@�C#)��h�>�0�"Olt;Ƀ�1q,Q�� 4?���S�"O�Ђ��ͤ-�\����P��P��"O��7�&�d-�`�(��$� "On�"�� ��L�(�L��BB"O8=���<N���7��J%"O�D��an%Uc�5s="O�0�t�^xdH;��X 1�U"O����V�s
�xsR�:r�N4Ȗ"OP���߶��4�PC�|hb��"O��(T��KM�� �
M|�yT"OF<���ĸ9���2Q$���"O�5P�
\�vh��C����"Ot�pf��(OLMY�cP�\���
�'
��*�:z4mQ*̿h���'�T�r��O"�Sp�I|�=��'_��&ݚ#�EJDK�I��'�Խ;����K��a0q��CnL��'/�E�3��03�eH`A��4A���'7����q9��9��D$-Zq��'0���t`߉}�
��w��Ts�'<|���?�4p���r���Q <D���&lE�T!�	���˾
jl�PF�<D�� u-_B�9p�ʇV����4�7D��i�GI�Rk� ��H�J��L a!0D� p��'M�Q�[�b}|�� �/D�$��_1���엷y��$3D�$�'!�3�9[�lS��@,�Vg=D�`Q �@#��r6*����A:sd;D��C�G��	�*5Pf$Ie���8D��{1��E%x�P��T [�Z��4D���-L�]����s� )Z��4D�0
�
�^�xI2�(B[P<(Ss3D�LK���4`�᱒`	@����!�D�f� ���\;�,C�NT*m!�%U��	�B��,H�+�G�cN!�䘤5ep�Xt! ?��yo]:.B!�D_4�2�X����8�.�+{	!�Q90�bM����e���B�$
�!���` �SC	@�2�����}!�[�n:����VK��L+��	�%I!��ވ�ND3�܆Y������q#!򤙋
pP�,߿�BuAD�p�!�H�6Lز�ʖQ�2�b���.y9!�$Z1%������A��٠4��6 X!�D��ޕJS͈�=�T�w����!��&��l���M*HxT۠��2\�!�� N�k���S"�DYa��!S�:!�"O|0����A�%mԡ2ʸ��q"OpH@�����
���A"OV5��C�
��)�Ah�v�LE@"O�'c�!P��s�%_��ųs"O��h��L��$8�7݊��"O�A��_�_$��dA*lz�S4"O�=���]b�N-B����	4"O�A�M�&Ԍ�p��06��5"OBЩ�l�)Z��;2	��T.�*v"OX 9D��-�����)7��%�2D��ѣV�u����-�4@�����$D��iEۚj�L�Y�M[�c�޵�l$D��Z3��� u*`4Qzt�Hw
#D��b�@�l�����/����a�&D� �oY38�a�!'G~�� �&D���p�I�lꍳ@!B�.FmA�h0D��`@ L-�h(�
�6�⼊'/D�D��n-zpuSrm�8u�Ҙ2��*D��c�GVj��,Ò bi�x��h(D�R���L�\���߯�08"&2D���Ȟ!�X�S�N�!-�lK&�=D��0��]OB^䨶��3 ��`Q �5D�$¥`��g#���M"p�V�H �3D���g�{�	�)ݐMi���U�N�!�$]�a$A8��VX� ��Wh!��_��hp嫜".8�q*��:!�D_�"O)���
���� O\�q�!��� &��u��c�t��kȬ@�!��ԩdTlM��W>�`�i���!�W<2w����̢�8T`e ��!��ǥ9v�	��FP�Y��5��9�!�ƹ<9����$F�'X�i��ϳU�!�"a�N�ʲ��/V>i{Cӥ_�!�^u�"��!�/"�J����!�d:Q$��}\��)��CP!�D<X�8�`3fT� X��)�<!��M/_�ɘ���1�J����?4!���b4��A���bY���U�!�0��G/)�"9@���c�!�Ъ{�~5qb��E]� (�M8�!򤀬^�,�ԪAc���df�<�!��\�D�d��ѧ��t�:��$E�5e�!�dC�HE�В��M�$u���M�!���DZ!��	nt�g���]�!�d��bg�Z��i�D#�*y�!򤍌e�J�z�M��P�&ES֣��w|!��W-
kl�c�F�<�"b�bP�{!��� �Mc k�Y䤨 ��i!�k�<��t�F�8�ڀ	�b�!�D?3Hj��G�;u�F�[3�L�x>!�d@
�HD��v!���ҪH&@�rńȓ>>�E���C�'J��ЧQ� ��5*d(ڧ��?�IJ�MY		h`��H��,cA�B0GP��� �L�Z?~l��n�-�P�Ea� �q��^��ȓi��@��Q����g����$��ȓ$��RU�ͽm�=�Ǎ>�����޶�¯� =L���&[�G�ćȓ9|1X�ҁ_�8���/q�B��>� �r��ҢY얁���X+i��0��52�dy�Ƅ"/_�*Q㝒aQ�ц�eK~������Q*�ȋS��D�ȓhI:,!�&����� es���S�? ��s�g�64������#f��X�"O���BL�2ֺ��%kS�8���s"O�%.��	�tm����0H�"Obt��ڛQf�I�B !$�M˥"O�
�뎵&��$�d����|��"O�� �@s΅�aD�u�g"OD�����(�6�z]��Q�%v!�$�
�P�0�=Z:�u�0NC,�!�D�z+z%�竜�@�^ Sӭ�1_�!��%M��F*I�jt�9!�ۧ1�!��ׄ���rI3_��z4'�:EE!�Z�$	��г_D�Rb��lV!�Dܻv�b�9@	02�mc�Gͼi�!�DΦ)�%R �J"sj�
��L��!�Ď�X�p̻�^U��yW$�=<�!�Ď�bj�<KB�I�n��$ �P�`$��dW��^�i�b�"D�� s��y���Sy��e�!�B%�"cΒ�y���Z���xE)�6 dth�!���y2(�"$PP�a*�8 ֚HqB���y⥄ut$�륅ѾHb!Hqn	4�y�G٪U(��s1 ����d����y�mӖ;b�)�U�SN�����yBd��oJ\�D+T�I��tKga��yb��>O�u -�A\�����'�y�O��T�t��T�k4 8w�_�yb���f����c�R���o��y��U+=�&t 2/�Y��(A����y���
�)���@)#ß�y��Q���r���o�zPr%,
)�yR�G<�����[6�I�́��y�DžR�M�Ҍ�N�T���y���:g�\�,�\�<X�����yb�X�#�X92�#X|p+���yb�R�y}�p�w�ܤ&+�a� ��y2�2�\\*"nL��rUp7Aۛ�y"˞�2������_�hʀ��<�y2m��i��x�R�ݑb��FK��y�'�=3)h9�&@/T�@� A�?�yZ�
��82�����#=�d ��'���U��)#�°�ѕ8A4��'���C����@W��v�B�)^|ԃ
�'q��������Ix���5�΄�	�'��at�
�+���J���+�P���'��a���2��!H�Ȟ#M�\k�'y�]�#�cI���Wg�s� 1
	�'���S�͐"N���Ȕ�j�&I�'������z`�(����F���=�ଣ2�ӓa<���Fڡ;��,�ȓ��Ē�\�EĮ)�	]�b��v����b�ka��-N�� �FFw�a�<D�83C��	Z�l�
�1*������:D�D����x�d9ж��$$�Α�3��0|ʤ�� "�J��a��	�a�}�<D�E-��e�6��:lL0��#^�<�ԏP$6�P��0�V y�0�h�H�`�<�5*S�|a`D)��q�hboǟ�F{��)�8�:�Z��!r|�se;l.,B��(&,9:C��-)T|��c\ M*B�I���p�\�,�r�r�4@�ģ=��'{F�< �0�l��eĨ9����mi��r�,�?�J�h�n%x]�ȓ�I8�mõj�IآėS���ȓQ��s���-EI(�[�*E8�����S�? v��]!^�4���1)�y�q"O4��K�rg��q�@�I�I1w"OxQ�A�C;�$D�U�y��b�"Oj�� ��=G�B��f@���"O�Y���-4�,q�^�{�4�*�"O� �(L0����֣�#�Z,�"OV�:0����9;�$�=./f�3�|��)�*F��7EA?�b�*ê�c��C�	+�R8P�K�2X�B\KP��P��C䉂.=&UF�V8
�D�W`�JL�C䉮a@���LY��"�+a ��C䉁t�ʨ�#El�|���z�B��>^X0�r!P�I��[6/J@¢B䉳z"a��	G�F떀r�,̕Q�ʓ�hOQ>C�@WB�[@�5to^U�$D���� ǖ=�U��!s�8���!D��B�Ɲ�2�:OSj*"!�ƥ!D�H���Ԍ*/����)߫9�шŠ"D�8��F8.��4�q ���Ѐ��?D��!��R�(������8D��0�ꕟl�f9� m�=��@kFH�O����S�O���7�,mk���f�Ҟ X�y��D.LO(� ��������c�{�"O*M��hq�4�����+Z�R�a�"O�	#�P�Z��Q2��N.`n4x1"O6��Rh��G\D��E�{�4,Z$"O�Q �A98���]�8}�a'"OrP���{��h�
d�ఢY��D{��i��Z�Q(���N<�3$&K��O\��$C�gN�20뜀m}��KׁU�dl!�$�dEn��W�'�q���~k!�N�ZT0I�b)/z&���+C� W!��M����IW�1 .N=�A��cE!�dS�e�@$@�dT���;H�!�D���`"��_'��9W�	�R���)�U�
���+"T��-�wmZZ��H�r�'�|d��(D�
8\sw�
�m�~���'��L���	I*���'e��c��]��'=�YP�`��a
��k�JؔM�R�';�ԂE�;P�"�k��pu6�+�'�V�Z�J��׾(9a6<��%�
�'�XŚ6�V��d�����-c�4���$(O�D`���)
��)gǄ%G���%"O|�I"OF�A�l�c7bD2��|"�)�S�8k��xD��ZR5��hE�M�B�IgP걢I�_P=iU(G��B䉄L(�8 ��R�F�t`H)A�B䉉N���A��ܷt�&�ɕ�ǿ<�B�I"B퓓��=I���F�d��B��vr�tfl���L�5`V~B�	�?c�<R�씍$�.���M�'�`B�ɱ���1��C��;OM�p*^B�7<y�陦c
�'ج�UH��r�0B�#��48�\0O��Pe����6B����ȖJ�N���Š,�$B�Ɉ]��D�7��=/��@r�
�^���)?iS�ʏ��d�x�t��<������ :'�b�g�Wy���0= J(V �$�c��a����l�`�<�F���R�~+ug��T5L�rd`�\�<��
V�*�fia��Y�,9��Y�<� �3J��БoFn�"D+q��j�<qbʒ?�0@ C�E*�-K�D�l�'�ax��K)�4�1�����<��F���y
� <<����/j�Rm���#��aX�h��Hyb�|�W�L�V?F����46��@�M��92 '����:5z �F�R�8�fj�z��C䉐0>�iKj��Z!�W�<B�	%����g2:��dUFʾC��8(��4# cV(-7d��U�C䉣 ~^���B�?z��cV��=#m�C�I�"�����*nĹ�LǴŎ�O����O�㟬���<�Rf!Uxy��N��� #���S�p�H�AI���т7nеR�
]c�'D��^��l�ƨL�+45�D�1D�����K /�����,
h]ј��$D�<�!�CDp|�7��"ҸE!)#D���ҋX2;�z �w@Ō��z�� �O��䖧J٠�?� Y���!L߬����W�8��n�F?Ȕ�'"E�*R�Js�+D��C�&ݨ;��}K�H�)W�>HHi7��X���S�@n�m����:	C����`C�I%k<�0�W�^�-�P���ݫ�B�	�nmt�0��Xz�L�E��C�ɮc4ڄ����5�f��k���B䉩^D��p$�?]T��΄	�4C�i��K�HW�*�L�z0��`�
C�I�a
3���r�2�A;� �=��'���V(W�f%�٘��
$*�^e�ȓvOv%92h�m�,��FGϠR�Q�ȓ8�ޝp7��8xe���#u+JH�ȓv�5yRΟ�6�N��ON@�ŇȓH�`��jBkg�MP1�U"]�}��!��5�SCY<)~�ͩƈ�9w�C�I�M�J���3{ʌp�MA��RC��$�^����˅kHL��/�*�C��g�4��� �6; �1��s& C�� (<%� lؽHy\<�V�;6����;�S�O��uK[?P�1�"N<:q�G�'���'�S�"~�6�V�JA�1� ɺ����$�y�+�8Ì�Q);��R��я�?y���0?�D��qu�8�"U�)��b��m�<	4M��"�yQ��Of��d
�Fr�<���ԁ1�0�	 ��#X���"p�<�a�a@N����Kj��b��q�<yVd�Ft�TaRlDE'�i��u�<�Z77���J�|�R�0���V�'y�?ڲ�������b�M���0���Q�<y�Ր/�@uP�Z�\���)a�CK�<y"�@���)e� ����bJ�<ɵ�+��+%���!��z�<٤�]�9�L(��J(Ӑ$��~yb�)�'$G(�y�G�v9���Ǚ&����I^~�Z�X���j�'kc>`�Ѥ��<���O #~:c�л_����сN�
��%���q�<Q���$(S��9���pR�k�<Ye�S����"�,D��8u�V}�<�SƇ1|$VL!!�R�#����+]Q�<!э�'!\!�u g�&q���R�<٠�@���\��D��愛����'ɧ�)�O4�w�����2hpiڣOF�cW��?��,��6��=^�l0���L'hW���'�ў"|*Eͱu����Q=���/Ğ�y�'[VUQa x���0;�<�4�9D����a�S%���f6r���CD6D�С�$�9t�h�W<M�x��*6D�Ġ�`R0(s�tqG�ޝR�VD�U%�<�����-��=6.PD���E�D�X�C�)� �i�	7[;��p�:=A�0G�'�"��$;�� ��芢kP&Q�'	�^�,�	V���� �#�%܂,g��6��Z�]:'.D�LP�"	�]���
V�ոh���bA�&D���#��\|B)R ҷ?�0tѠ�1D���`�]B(P��:  ��-D��õGR	`̞u�2�� x*�P� D��Ċ�]��M��N��wf���y҄ٶv�(H���	&�D�A�(�y�� -J-,�RBl��G�(�yR��3pDy���u��&j� �y�f�Y����<o$�;��՛�y������񖎘�a�8t!jU��yүʕ�jI��E�X�.ău�m	�ȓ
0  EǤcU��#�<��Xl|�3��ȡ+y������=�ȓD���J���T�PEh�Q)����ȓp���@��0{mb�&юl��m�Eb���n�걱��ƌQ�T���:�>dr�0fO�|��U�@�}��S<�����@0ayRȐ�'�l<�ȓ%|j����;��h��ܼ;Φh��Dl�$j�B�V�f񊡡�R>l�ȓ+���	��@2Z(ղ&�yk�ȅȓ�N�����~�
��/_ V����f>���3A��^ }�B"xj�xh)O��d7?Y�JA#|�<-QF)B�����W�B/!�$�?�:<R�U�:UD���ݵH�!�D�$ ��Yy��K'`@qqi�/5�!�$Ҳ4�R���+a:�Pi5C!�dK�}?�!b���:�h��a!���q:��B�I�;)�LZcʌ3J]!�,�J�%���ɧ�̼VK!�$�:(�����T�2&��>!�,1���sI_0X���i���(!��-w���{��R�0�Q�&!���q�LQ�ۡ3�&q����P!�Dt����;��Ԙa���z�!���x1��:�OȤ"��P���~���ȓ�����( ?v\B�&��
je�ȓn�r�SF��/ۤ}�c�Л�fX��$M8y���Ǧam� ʰ暖	�h��ȓ\b�ݢ2�	n�F�1t��E׼i��3�&!��i��p����*�:�Xq�ȓ3�h�z��%Q�0���˧��y�ȓ��|ä&��5��D��9k���)T�;�j�B8�X�㩐�@g<`��m*|]l�s�F���N�c���Ia<9dn��m����qG�'>9@�	��@�<�c _1IL��� B?C��dqЭ�c�<1t�_h��@��K%4�ZYy�Nv�<��$�8�V�0b�E���R���s�<٥b'�i;�"X���
fA�x�<��W򪰀&%@�I�x�h���wyb�'�a|��VG��fU�6k�L;��J��y�D��d�5Sqa�#\8�d��,D��y�O�5+rM2& ��A�qbM,�y2��8-�})ef� 4KF���kW��y�)����w"��/I���ŇȓaF0�AL\2'��Y�u�]�]z���Q�8�q��'I<�r�2�H��a	8�[�0Z{�;��p�28��;k�d���H�e�m���˂~����_�&��cϝ%o�v��@�A�-2<��S�? ir'��-�cp/ӎ�$�"O,��!�Me���@�%* �1:�"O��2mD�*�1W�C�o���X�"Od|�g�P�~S��;�扅$G�Ma�|b�d�|2�O��� ̢F�<����
YR� )�"Ob4g���z���ʷh;��x��"Op�yVBG?*�Фqh�s߶$
�"O> ҧ��2�)A.ܚ�9�"Ob @��ǂf���¥(P͚��"O��۱�P����%�['K�\���"O:	[�, �;�� ��gz���O�p�T텾Z#�DQ���l���Ӵ.)��9�O�܀s���M�aP�ڲW�� �U"O4��!9��&���>8x@"O�H�ݥd�
��T �;pђ�hv"ỎCG�ˇQ�t��H�V@�j"O(T�e�Wd�� ��B�k0)�V"O�@�P�+M ��dcσJ�B����'7�7Ob5(1�w�vt��2T�d"���3�����m��	Үn�4���*R�}��	n��(�`�0V�؞W�,��ҥՏG=�=��"Oh�$�כC�t��u�'T1ց�R"O���g�'+��SP� C�X�2"OLI���#
��FA.$�T@"O��VI
BX�s��� nkԱ��"O�e!ׂ_�/X�e(��5:T��'"O��3A u�0��A*(��"O�Q���<Ⱦy����)�����"O<����?u�(XuA?�Qc"OTI9�n�9����E@��|���p�"O�(z� �D�)oц>�ڸ �"OR�x$�9����N��j�lmze"O���C�#L�qi�,@V��p�'�2�����45
Ty�
��,uru��O^㟴D��X��M�g���$F��B���6�!��ښ`ڀ�4˖�F��!Tc�!�d@3�h+�-I�4h��LN�OS!��ևf�L�)&-�¨�t.�D!���2����9oF(�`n� A/!򄑅O�ls�HY�c���V��D!�$Y-�e�㧐~K$ո ��++��K��(����KTw�q��^n�S"O���Ï*oR�I����0��mن"O�ld�F�؀�D���:�"O@$bw&�6F�$�� ��x(k"O6!#�����P V�j�R� W"O"�{P��7c��%�����"O���� �+K�\a�QdP"���"O~j0�RJ��Y�#ӪS��!A@"O������4	�$���	`t����"O@��Q�Z8TN}{PC	(Un��2B"O��"T	݁]阡*�(�%)^�8�"O���ʀ�	�EA���\D� �"OhEk�E�3?J�Yb�x��K0�'��ă=.4 I��J	�V"�̔�R�!� ��u�����n `�%��B�!�d��>8�$!H�
��;``�!�dL<U4�83W�����P��2	�!�#���E��wƂ��5�O�!��CC}ʑ@ ��'\T�p#޳8�!�D�$M�l�C'�թ@��� 蝊c>!���6�LL����~I��kD��<E>ў@�'�>���)*8`�D�2�02�o'D�h�e?.��Ȑ��/�"e�3�#D�� ��RQ�o<u��L^2;,��e"O�����
+�`AP�卓D�l%��"O�4��e	�@��8��c�}N�g"O����\0��
)NU,A6"OV0��LZKV �I��:�X1Rr"O�[s�M+3w�1��:fՆ���|R�'ep 8h]>�`�R�JKNl���'�>�
� O�0"O7_Y�!�
�'U�\i�bG�KGx�9�O�Ot�I
�'	FIa�̄V��TšģM�Paa	�'� e�ѬA$]�n� ��%1TBd��'�\@GɅH�(a��(Z�Pؐ�'0<�h$D!b�^��3�UVn���'ܰ����s�Q�dԏD�.i��'��xcY& �R��4����'`�����7'�ԭ ��-X�h
�'�.�0�ۆq��ha��e(:䙉��)�t�q��� !��`���ũ֞�yi.�Ĉ%�H?���+Ś�y�MSH����� y��Z �_���':az�׈_KZa��!�6و=�Q���O(#~�A�J�1&�q  C?n�L+�d�y�<!cG�<�q��c�5?���
ѡWr�<��]�9[�(p'��VT��c���m�<���%΁y�됆u�vi�E��S�<	!�'-��|��E���DZV�<q#Gc��9��^�,�V�SR�}�<� ��}�@� 6Oh�D�+�\z�<��ĄJь6Ǯ,n
�1g��2�y��;v��`;����)G�����ߠ�y�g�;u_FlJ�hL�W����E����hOq�.��`�S(7/�`#��,��)�"O����Η/�TXѩJ���|�ן|��'� ��EA yx���G�R�@��'a�	c
�3KJ�r�&(F�2�.O��=E���&+����s+S8&���4� ��yR���l��g'�(���
��y��U N�iHD�'����?��'�ў�O��y`+�i�����KB�X\��YN>��)9d�$��fUb�85�������S*i+�N�< ��1�U�M&�L��g�m��K�MV�A�.҄3��B�	 z-$�S�kD�J�Ǌѝ&�tB�>��@�gֲ6g���k�lB�I���$
B�)Z/ؑ���v�nB䉌t�X��%P�t�Zʓ�hOQ>	a�FV�N����UoZ#W�ʌ���6ړ�?9����7}<.��.X�'�����;!�4̀MS�)њS��9`C_&R&!��5v�k�eP,$��U���7>!�$��?\�Lb'k�UزqpGˆ!��ϼ�X(ʠݯh�`0��Z!���}��ȡ�{�� ˡ�� !�d�v&>����9��9�JP,S!�X�.���д�K4K�Z�ڰj��S�!��'��[��Џ|w�pZ%@��[�!�ċs�"��,�S<Q��o�<�!�ċ�&�f�Q�1!��dn�-V�!�9��P�$�0�8I[��^m��{���L�T5ٱ���z�d9v��w�!�D˴mA�=X藎+ \��3愮�}��s�6�Y�P �,���0o5D��J��F�X�,���:3,j���&D�Z��LCt5�R+G?W>�9��$D�� x�2d�FC@���A[0P X=��"O���`E�+^ƵPTbȌW�轃��'E�󄟹l6d�jTjC��|٥�Q/��	K����A��Ǭ`!*���-�L.|O��D;?��.?�zh�G�7�2Hr��O�<�QÃ�}��H�	�*dLѹ�ƚN�<	b,o�4I�3iU;;�<��m�A�<��ə��ى g�;C�:��W/�W�<Ђ�3U�tJ���
-ж�k�<��M�.fҲX��7}���FEe�<� F�
�>Pz��L�K���R�M�J�<����"�Y���g�����C�<Y�O�TP�h�P&͌���i��u�<i���9��{�/��� j�G�r�<�� �5k�B�рՃ��Dy��Dq�<��Ⱦ7�6��C� F��=Y��VGh<�֡C�G��C$��qz]X���)�y�֭QU�4�
e�h���+�yE�a�>4����X8�yYb�K��y���`D6Á�R�~l��NS��y��LtuHǌ �X�����[��y��I9� �M�@�,*2@��yr�53<4Z��H�E����y��

m:� �G"�)DZ"�y2Iו_�,�뀃�-�f�ё���y�	J�n{l�j��R\��$�B��y�*��u�Pq�q� �d�Gꃩ�y��"s�(LG���d�2��C(�4�y��@�k.��Bo΅	�\h�+=�y2A��$&�鰳-I���V�͝�y�&�}b�
�C�8�X�w&\��y�(G��^5�c�٨�`�
R3�yB�ۭVT���g��Yhx5A��y�06�@À/�0UR"�0ျ�y�	�$s��*�H۾X#P ��y>����^�R��wI���yr���vl���ReK�M?�uj�����Or#~R�E��V� 4gT9>\�@rC�g�<ѣ�@ Kd>�[b��I�9 P�a�<��D!*B���ǩ����H7/�A�<�����4I�({����S�e�<q���ܘI�%�MR�`Z!L�]�<.	�!� M2�c�^���%RV�<	��]��т0��?�����hT�'a��L�<6r�|
�̱B����&�?�yrmA�D�0qc��(܂�9� ���yr�D,@��L��'"��y���6�y"��2sŴ�K�L> ���u`�2�y�菣k��i[h%�fG��$�J��'5^�J��A$�Цܜu+�'#Hm 2��}��9�T ��'! �N�+{{�`��&�s������X�h�Q����;L��!�,��w��h�p���[�,|�"U	?3ms�C�	9J�`�0O��xm^0b҂� ծC�I=e���bd�^H��:s U�+�bC䉪ŞXZW��+ZA��[V$�0?=C�I�S�v��Qo���s��"DC�I�^�<`D���@�4)R�h	OY�B�I�I�@h4�]\�y��A)���-�� ���uX"�9��G�5�7f,D�X��F�*��DF�K�.Eb}HQ�$D��(C��O{������ a�逕�=D�,��@�b�f٣��MZ��b�-.D�� �ղ�ST� ���DW\���"Oh�s�Ȋ=�>0�5��W�:"O�QWl6��aq��
��ļ��"O:��c��&W�~u9���c�@x�"O��G冎+0��㛯Ҥ���"O�yU�U+%��xw��(��L��"O��S�*��˷cëZ�BU "O��p���$6[���FZ"�"O��5N��cY�eȕe_2��"O@�h�&��I��%A8\��*O~<�r�Q6u�z�0�c=��a2�'�T<2��ωY�����J�>� Y�'�)
PL�	sR�Z�1z �h�'Ϧ��%!Ƚ;����0:/�����'�Q�DD��*��!@PLR�<�a�'�>H;f�*z�P�$%E�J�tM�*O��=E���3F�:�HCn�Cr�B�����y2�5d��en�@���@���6�y�?ڂ�3�k�5	r�@�O\+�yb	����#A�:�!�����y���<@�𡢀�4?h�E
�(�y�&� �B�3��UB���9��y2׋4I�+vK�9f��d�A)�?i���s�+V�R�C�dB��h��츓�+D�Z��F�Ȁ;u(L��B�.*D�p�cl �aEn��U%9|&�$�$D� Z5f]1Vq �Ze��� �<�yҀJ*OۼE�3�jͰ�lϲ�y���X �ip!!T�`iB@������hOq��Q����&wa^ah�+,x�hM���'�c��k���H�M	��Dҕ��1~t��)�'n��1�QHҏ0��=@��]3n<�	�
�'o�l����1�de�Ճ�/��I	�'#����J`��p�����.��M��'�LDIT��"dH4���&R���'�fА��H:Y�d,D�&`��q�'�l`�f��`�I�P&�1"��'�4\��E��%�ɮy�f-9��P��hO?iQ� 0(F��0����2��.�v�<)�N]�*��!���Mq��o�<�%�Q'P��k�Jz��g�<Y#�Շr+��;�N�4���#v��d�<!bE�k5�,�����[{��넫[�'Da���W7i�(ybThTl9Vɚ��H��?y���R�>�b�\-5�Щ���ӹP�>чȓH�ܹ�@aK'YQ��%����<�ȓKu~-yA �Tx��y�C�V����ȓu�4]�vk�&^��1Q#�^}p���>���9P^��p�I�[�X�ȓLD5�pÈDb���`i��y��m�?���~f�)m�8qHC�]&4=V�Om�<y�(ƃ'Y�3���|l8s!h�e�<�4�����)񇙿
���Z �|�<Y2�ͳ3�B,Ӏk�</���FSc�<�"�D�{�r��)��9�i�dDR\�<CL[�w������LN�<B�#Y�<��<Q��To���h=R��ET�<��Ɲ��8��/V4z'B�9a%g�<��IM#5ﬅb�N�A��S�Jh�<	e"�[!x�p�Ăt��{�jc�<s�¢�Nl�EKF'$
�*��V]�<'cp��4ڡ����+�\�<�G���x6�%� ���{0�r�q�<i�(�d��}QsÉ(fD̈#�o�<� ���Ƃכ׈�p#��v�ؚ�"Oz@��#c�D<ӵLU�*�"O�9P �%	q����+Ã��("O i:E铬g@z]�JNJ�T��!"Ot�$$�	con(�'�"�����"O��*sM	��=Ip�8��Ͳ�"O>(c�!�7��P�%�#i�`]��"O:$��O�/Ŋ1�eM�6��-0�"O|l+e	�"C�m8EJ�[��4r�"O����ޑ"���GF�(]�B���"O�*�i2���c�EZ���4��"Ol��o<p��	��F�W|B(٧"O���$h�;J֮���52l��ڡ"O�D�򦔜8��4 d�HY��q�'�1Oni�1��.���8 P"HU���IP>���f�=f\�]ؑ	8O��R$h7D���Q�:S�
�-d��Ј��4D���dC�'vh���*��:�\	��	4D�8r���/
����B�'I�,�Kv�&D�4)w*�tg�h��+�Si�Ģ2�#D��r&�'	䢔r CǍ	E �u�!D�,���;PN5�0h�5��ɠ��3D� j�ȅ�.�촰!��1|���C�-D� ��C��x8\�2�+@��r�5D��b���b �X,<��bwA4D��x��J/ �T�Ů�%��x!�4D���h؞|6�lTȑG�3@7D�@"W�\�9M� ���ւd;#4D���l��.>�s(a�JD 8D���1$9`��-�6�B����A�+D�4# �Ɗ8�y�Dʀ�����@&D���$�5`B�2Ԏ�)� �!A7D��邭U S�t����U���ɰ�9D�T۶#��Aj�Be��Ґ���"D��)�.v��`��%�6+�<D���PlN�a�@py���o?­���9ړ�?O>�˟x 9��W�d*u���B�2(�1"OD�����h���V38s��ѓ"O�2Q���F�݉G�[^x�[�"O@��)ӹ7����e��0^�0�z�"O���B� ��E�S��+@،�7"OQCE��s���c��8���C"Ov!y�kУ/xPh�J�7�՛��IJ�O�ad��$�W曵u�JZ
�'�2u!"�=r�~谴c�����A�'� (N�jX�0���
j3ތ��'^$�V�ܗK7\ q�%�ZB����'�6,�Q呅aP��3��S�����'@x�Q���X�����嘨Y��Y��'{��0b#\
8�*���G'QF��`�'`x	k3?զ��UH�1�Ν�
�'rʘ�b�E��h�R�{
��	�'����S�\�
6��d΁�s���	�'Ԩ���X�I�>`s�;5��`	�'V%crdE�(+j!hQF�4�ޔZ�'k��趢
h���Y܈jj)i�"OluZP����< �V&�*��4"OZ(��LޗK~0� �F�%�81;f"O�Y���ݵ=@i#d�4�lEa'"O\��TbӸ@Y*F�^�*�~	�V"O�$�D�P=JeB�$�M�'GP9C"ON1�`)��}~1����)��ڑ"O&��1�;�ܡ�W)� .�0"O桘4 �(Y����G�|�,83"O� ����F��'7�����1j�h4ȇ"O��I�I�pRJps����|@�"O~@�D+ķ;����DiX�a��%Ke"O�ȊfI<S0�s����hԢA�"O���d�@ "�L���
�hŔM�A"O��`s�JJG�Y���Y�h%"O:��	:;���0���R��&"O��*&����!V�A�dI��"O,�S&Mͭ��a� Z_�N]Q""O�(�b�[8Q�e�dgH)<�r�e"Ob K��ߨ�`I�f׊yPe(�"O�P��Q�oȒ�E��%Ԛ�S"Otq``A�
�^m��A2!c����"O��ѥE2>i�`��BpjA�"O���"M#��ʃ�C�;Szl��"O� 
�S3l7���d�gEt�Ku"O�u�uBW�U���+��Q�|���"O�i)�-8���,�s� 
�"O�����V^N�)�-۲U�0�J"Ohղ�g��T��x+g��?��1�"O�p!aA^�h�,�0ß�N�u{t"O�@9�*	�z�|B�@4Gj��T"O:$Цg���is( �#�:�"O��Ƙ*�v(e��U��)��"OȐP���x���
�����"O �!���N��m"��M��LZe"OΔ��ɼT�6�@�͚$��Y�G"O��k���y��Ѓ�d��T��Q"O���M�5~���É�r�0Q$"O��4�� <�X2�b�8�p�"O2�hb�R��(P�qKBa1H "O�h� �p%� b$˃����"ǑȖ��D���d*�	�a�S"O|�!�EA�₤� �ۦo�l4+�"O���ʝ����V����p�"O�- !��I^xy�e�Tw��*O��!�Ț��PX0�(5�@��	�'�Za����8"2,����(��q�'`.u���K &�΁ ���0]hY��'�$�fU��a����'JFB�'`��KF
WQ0�u��KYjd=�ȓ�|��&C�� �1�D��z��ȓO�D�тɒ�:=P���	P:G� �ȓ
۲��#
>�(A��[�	R��ȓr���0�#�-$jiP��S0r���f1�A ip��/?!�"�ȓ$^��eK_G��}#%�KR�t��](�`F� fYF�$��)�ȅ�B>(�&���l:��;:��4�ȓF8ib� ��A�᝹Gt�1��F�<H9C�D��F�I�eI1w����,�H�($OȚ}����M�U��v:UJ�┏M`���mZ3o��5�ȓ��,H�ɘ�Z-��Q ^]� ���wU���B�4Bv���cA��|��9��=�X`r	�3un-���22\��ȓ;p�YP�OH"+5���.4��e�ȓ�<#��[�k��-3�Nݖg�i�ȓ��=��X�Rp.�+cU���\0A��\�:��ǨW�r���7<X
ĉ�R?\:&ԤN��B�I��X	�"�"���SKŢ}Q�B�	*���A�`AL��`���! ��B�	�y؆yb�����b��33ސB�)� `ԡ��2.b�`� V#p����"OP��πaYDB
Zu�Hk�"O��P����L��{�8h�ȉ�"O�I��K\�ܨq�a�"Nʹ�q"OR��d�I	�x��!�@A�=H"O�lZPfX�J�lu9ޠI)���"O$p"@'!<#�Y� +u@���"O:q��:����M��L�0�v"O�0��nU8
� �!LN�)�u�"O8��7L�>h� Z�mös	6d�'"O���i����@L� c�X�"Om��� WG��� LR��xU"O��۔e�*l��)a��?�r|�"OV��L�
%d���B�e�2�5"O�ш���4�����H�5�r�s�"O����O�^��D"���:�.8g"O����9�F�QC<dӨm��"OB��"�2d�0��0����w"O`|��މ�`���L��X"O�q+�� 5�R�ٖj�%�l{A"O��h#�RO��4���F�1��d3�"O��eO=:1��k�&;~֕zE"O̜�SaF��>H��	͐z���$"OQ!�B�O�|[�HL4%v4�!�"O�Y�$��&x�'R`9:�"O�� �CƳ$�T}a�Y�l|�4��"O�\��*� Cm�a[7�BSθ3R"O|}���9�0� I�CN�;�"O��f+����ãX<6	��"O$����� l�������#8��"O�eP���<q-�)Q�ا4&bt"O\�@hD�+��ȥ�~�0""O�Y��I	k`Y;HY���2�"O��@kķd��5�9�"{&��ȓi�)��V	VA#*��2���*��0TO'U�U���јL��P��E�}"�*G�=���5�ջKE.��?����3�Q�1D����"���ȓm��!���-z�h�!ǥ�S~����5LDЂSM�}+ dX�ҁi׆8�ȓ�^)b�O#y�^ 8�ʴ8�r���P��H�u�\�JA�͛2,��gl�H���)�ԂQ.*<�s��h�Їȓl��㮓L(x"	��T����(��0��݉�'�`�t$�ȓ7�z&��+բ��b,�*8��sz:�C(� #nj��ΪmG ��ȓzJ�+�M�&8�X,Q'4�Z ��[C�h@ǂ�: ���tkH"E�J��ȓ�]%�M-N	�p�u�P�\�\��}^�8e�]��P�N!j�i��A_��^H|���C�# t��"�[�<�$H�(賣Z>zR����r�<��͋�*��!���N
Հ��R�<i�dĶe��D��S;FC�����V�<��E^�K��*a�12��%0��V�<�K�M������y?(�9Q�R�<�ק^2V���-�� i��O�<7.�+tW�%�&�ͩ(@������w�<iF�Y~f���b�\�h$���Yp�<�c�/S�ĤPu�V�����SH�<�7�#K�L|���P)o��-�!�]D�<1e�A,\������eF�C��Qi�<�$ D�gf �J�&C�j[r�;4�L�<� t��B�`T&����]�\b�"OH�H�HQ,Hɳ�EϔJ��Tò"O���
��+t!9E�Q�y��-k�"O�ѐ�*�(<�
�S���\��l�Q"O�h:����ĥ��cZ,,��"Oԡ��f�,4�M
�}JFmٶ"OhlP���hM��b�kqA��
!"O�3�m]�\4Z����}[u"O"�����3���Z��#C��h�g"O�I��G�-SĴ����u�j��"O`���^�	�h72���"O�xIO@�+vV�(d�Nl�\�[�"O��H���;yՄ�cq��۠ũ"OBE�`�4~���k�sB!�W"O�� ^$���h(ǗW�"ɒ�"ONzp�U)z��4�΂P�ˇ��y���}�8z2FH�4�� ����yr`�,N7�r��ά>Ob���]��y2�4Z3�X
G��
|��օ���y�);D�Ĥ#�Ώ�k�d��+'�y�F��4�A���Y#5��)�@���yR��#!*�lJ�I��Z����V9�y���+�<I �j�!e�P	 �͍�y�$&'h4�3��}o����J׫�y��#4̠h�a��v�f�Ȗƾ�y�KYp$���s��ȁ���yr���-�3w��˞4�\�ef*D�X3�)Ez��ѰMF,H���b(D���֫�\��=����AD�!s�e*D�H�FY�ki4]�TgD�l�j�Cp)6D������q�Y做(���"3D�T�d Oܦ!['>����$2D���O漁h�d��/*�Ƀ�/D���@*S0<���Q`���m��U��*O��@�,�9T�6	ȗI_��.��"O�Q�T>Fx�aC�V���3�"O@Ub��k���A'�3�xY��"Oi�3a@�p�4����H�h~H�D"O�,�c�W�=m*�H�!B�b��C"OL��G%Y��kŦB���1i�"O�x��J/2ʐ�#��%��!�#"Oq�_7]��ҵ �.�0�'"O���F G���.n>��:��y2Oރ���b�M9[���Q�OD*�yf�U����@���O�a �ć�y�%$����
ƿ1�> �ViЭ�y�
��S���h�*��,L\�1	��y�b֏!t��'�C>t���V�y�!R $n�9���86��̢�ˆԘ'�ўb>E����4�|�n�>�e�s+1���b�zuI�v:|�6fT��,�>�6�����0lD��S0,�)V���̓�hOq�p�H��9"�]�������$����ȓ
ѐ4O
�1b0h3�Aʤo�������?��(�#B.�`�UQ�9{�}�\�<���Z�!Aܑ���۠F�`� ˙~�I��HO��BN�1Fo��wgF�q!b�,�y�44d�� ����'gB���'|j���	*�fXD���K��B�n�2P��ʓ��D;��Iڌ,/�x��ޖt܀�R��.�pΓ��'�ay
�q3x4"�#׾PC��7H�
��'�d0�g?�T��9�������[��7��K��}R�X14o;6Ulո�� }�j��H)\Oc�U����ACc�=YbvE�$�'D�� ,�G'J�	^���T�0J5!�:�ŞL��0�-�c���V��	߄(�ȓX%H��\.^i2�xg��Y��Y��`Ā���#@���� )6�xBN.��v�'���"�D�?e�Up�ƀM8�'śv��`���)%�/^.���#
�L��'�ўb?�TI�{�N1� ���r]���/������yr��P��T
��ܨV�F8��"O�5XBɸ�p����ڼ�3"O���e`�@���q'42��H{�"OJ�cf�E��6���fG�nYX5ؒ"O���&%A;N��1�ɸ[O%��"O��I��?	�Ⴢ��g80�'��E1��w� ��ZA:l�
�'�"mBo
�:h���~��
�')�ɱ�صu�:ȑc��+�Xа�'���Y�J�#~� �­âM� ��K>9�$r�����>\��� ��]+8)���ȓA㒽(���xQ�E�+��х�d	~-��Ǒ��0���ܪX�ȓ $�e=7c~��O�>�ґ�ȓ6��2����;^(�b�`̷+.؅ȓ	�#sE�:B�扊�( ��� ��<u�}�w鈙m}�p��X�Go$�G{��'v]�w/2
� fė�CƐP��'~8��dL�	xx�THfz��ד�~��p��ᔴI��!z$k�%<�h�)1���z�'�T�����n��vҙ�`K<)��?�S�'#@*�@FG�<x\��$DJ;�*P1�x"��"~�Ɏ(Jv��D�P#���Ve�=����<�I<yS��",EX	�2�ʳy����'��p<�w���d�<���B��Vm9c�O�v�<�c_"C��
�K�+�`ÍPg�<Yd�Ѳ$���TI2C�)2U�Tc�'��IR}���C>x���E�Ĳ�����.�!��̥x~a
�I
c�"$:Ǆ�J��	\}���<��q��� F%1�(�����$4�d�"�Љ���.(�Y`g��{�!�D��D%ΐ���#N|�wL_�:��{R����#bז�&i����}�G��uxC䉯JR �c�2�b`ʖE�&���D.�Iu��� �&��NH�smK&W`�C��'xH��bV����6ɝ�O��D�5���	C��.�E�3A��.�a��O.	�A�<�x
U�[��Փ�"O&`�I�b��x�H�9_� 8G"OɋC�|���;2H^!��"�"O����*���7���V!�<*�!�)�V0����W������>�!��)5*@��7Ƀ���W�{�!�$��P�f� ��E�L�b� �O�9���E�D��	IC��[9��p����yb��c�2GJ�'}*�AK���'�hG{���.Gx�n��?Q�Y9$D�<�xB~�*�����&
�¶�	P_H9�g"Of9�����'�iU��{��'�n"=�����$��nF�{�a��	Bk?�����%P֤�q�ġn�朸���OHC����[�&���q�[�Rlh�'Ya}�`V�R�y�7J��..���������p>1S��8e�LtZ��9�~�Z��EG�<���֔kh��ۅO[�k�2 �� �N�'oay2��(T��j"&��q������y�EC�.�Ip�� 9�jLP©��y
� �	���E��0#g�=��Mj�"OXUq0o#"��\��yҎ!"O��Ҡf�x��xR@̣�T18��O�b�L��Ĩ~
򬝃i0lA1Tп7
@H3��@8�x	M����Fz8�q���$6+�ik�J!?�#�S�Om�ܻ��S3-�q�(
0[_��:���;��U̧E��BCaY7B�0�b͔�Mބ�'�F���	�- �kq�.k�@�ˣ�M�N���HD{�Oo: 4/�0�Ebp���sr�Ef���y����9A MOoJ)���7�ē�p>qB�ܩ
�v�Ȣ)5X�x�R�SUx��'�T9�n ��ɣ�F],0�@�"�>��E�T?E�Ot<$�̫y�`Xs͛9N��,0	�'�LC�Ҡ8-�T��N����'|��j�G�9	����\�K!����'�ڑ�VبQ���1 �?o��LH�'T�}ZE��Z�8��W�Q�ք���'%�ibB�!@��g�O�q?���'o:���G�����I�B:	�Ԣ�'[`�`L�+9����C�����0I<������)��@$�X�_u�y"U��y�O����D�L���[֍PnZ]�T-�!�_B�l�WV?1PX)���V,1!��)? &��7��p��8����f.�����	4Z7Dx��O����O�)F�n��d�>���0d�y�C��)xd�k���F�<9PN�4��x���&T�Xa�a_A�'�R�D���+6f���)D�������yBG֬7�j��dˡ�@A-��yBhM�b��L8s�Ԟm6xqa���9�y��'6�p���Jip��v�اRE�!�	㓘�\�~�Ӭ��?��xq�N�9S���ȓc �e��@�6R,�s����N$�'XQ���?�փ��wK���h���	`%m`8�Dz��L�kh�ҥJ��_�Rd �-�Mc���sӆ	+�-ע�����ID{��a��Q����4����p�q��HJF�Ȼ!��2r�tYbj�D�r	���#1�������|��Ί��X���b��2��C�4Df�T��M�X-yn(^ʸC�I���gL�p�R<J��M�2�\B�	,a���#��eL"\��jN"-2TB�I)z����@?L���xW�C�I�V������=��]P0'`բC�ɖp��]₇�9;墁�s�#+9�B�ɽY���
ubh��a5� u �B�I(iH�뉴G�bmr��ޗ\�B�ɉJӼ�Ȗ�G�n��m�R�@�f�hB�I���P��뉀��yb��G��C�I��H���#]�P"���
dVC�ɅC5̽A��<��t
�F@�o��B�I@���Q���<�|������B�2V(��EdT��J1�E�8Q�|B��q�}�rd!IXT�uEqB��/э)�IfX��t��&F��-�ȓpz'-4<���	Os�)2s��n�<!І̕:��*�GY�?0�����k�<��f: 3S�<�e�T`�h�<�6'ͭ>�\RƟW�4�I��Ta�<Q��4R�f���Ɣ�a�X9�NS�<��P�W�L ���4��p$dM�<i�
�� �R���l�~q�WlXG�<y�Wy���"/�;<2�U��E�<	w)��[��0B%`�F:�����@�<� xH�!�_=*�@�B�s+��:D"O�-��&(h�A�BY�7G��"OV�c�@�Xwje�� �F<u��"O�S�m�c�v 9e@�]7��P&"Oȡr���7Y���w�@�DJ�е"O��K�(��Z�4��%m	$���"Oi �Ԗ!�L�Ĭ��Y�n��T"O��j�)����P��>H�"OȽ�nD�e�@R!�ىp��`"O���_�����s�^8�"O$Ѩ�m� �\�C�JF%���#U"O���C�޺{>v%���;�j ��"O�e�saL�1�ش##��Gpp@I4�'7����@4l5��=�B-�k %���:
�'��Ʃ�9	�W�T�!�lP	�'phH���d���Rb�R�P�,R�'���BY�J�BP���#"�s�'*�$0!���v�x����:���	�'�^@���]]"!`��ڏ�ވz�'�Lq��	!,���`뎋
�Hx��'�v�9�A�0-��i# , < ��1[
�'2")�qd

�<���V{�B��
�'+���0&A+h�\�`얪ew<�	
�'�ȉ�1�O���ph�5d���'[D��%�Qb���Ro�Y���r�'C��q1)�%�͉���U����'Q�8��Kq�2�yr��U��8��'\�	�E�	M�ICqGS�R��5#�'��	c2DW5#��h�+ْR�Q�'i����x�%����{�����'u�r�*X2��QQ�5v�v<��'�8ۓod�JU��wOlR�'�DP���ǯ|u�eT$�b�4�r�'ڙ���C1YST��4"3gk�HJ
�'ɌHe� �����߿$| ��	�'Y��u��$Mm�dH����]��yb���yc�L�C�܄S��A�!�yr��
j����O���tzu慨�y�˂8�ȁ�'�o��c$���yr�2&���і�l�Z���.���y��=�B�K&L�[n�9*[�@	�'$��r �0A�<B��5`DD#	�'��Q��.�+��y`biӔ6�lX�	�'r6 eJR��Q�>-X���':\�B���]4,�`"�1$:X�H
�'��})O��V��m�gC]=* LTk
�'crqc�%��c��ʰi@ u�����'z��ceҀG5#(�t����'��15ʗ Y{@���f���R�'!:H{tO�:<}H��Ԛ@/\���'��	�D�ѝƤh7��3|
�'��(���r�DȲ��7 "�
�'�
yڒ�c(>̃�jĴ))Xq��'��USp��'+�^����*�:�I�'R��h˒3*I�s�("��Y:L<���@QFj�b?!�l�8O�ֱ���^�~Vpk�f,D����,�)�nxCG�� MF�I�����MD�]ТB-�3�E�:��){@#�ZB`,,j�ɢ���?�|J�Χ5*�����8*��ys�ӱ2��b�A�M����X++�4�)�B�V���Xl��'�\�릫�F}�%5L��8���w��^��HbT��m�h�r��{��/ޕ���{#i�9Q`쓭*<zP0@����Ƀ`�te�qc� ��)�'{W���b��=!٘��o� sQd�GB�K�I��t�~�Pe��wX88��B�~ܩU	6P��'�$�K	�Ϙ�� ��p���mx$�
�-̣V��t�DS��J�53�qOq���HF^�v��A{����K�r���ʟ.��	׈\��p?�Q��S�H��C�2��4ÍI��<ܙS�İD9S��P��>)@,W�iN��z#&d$��c�KJ<9p���t,!�lL;K�\�i��Ʈ\�TIX/O(UK�'е�|9BM�"|��nI�5���#)�.*�E�å^{�<Y�Ǐ#:� ����ѽ?ޜԺ�甛vy��'}�!��N+��Ϙ'��� �]1_�4��h��T{��J(Oxa �:�)��#=D8�'��w�`u ���2���I�(\�~���`'�'P2�����H�	a��3Tl9L<���7c��w�*�KT����ēi�5�$	_:M��� i�<��\���h��S��S�Ir�� Ϝ�%�~y���8r?�3I��҄!�)��-��a�p.�A|D���Wh�#?��lRv�T�?�3'�K�l,U1��;BT��ڷ!D��P�.Řr�j2*%B3����@�>�Cđ�T�.�"}��B�+������(l�^t��m[�<���B;*�S�-0�%i"*�V≱Xn|c��'�V�!�0<�4�u���n��0�^�1�Z}Ȍ}K��܌J��h����ybf�k
r0Tƍ�(��K�c܂�yb�V	eֶ!�#�$>:`7�W3�y2Jֽg�493�`G�S�l�^���A7�x�$����%�z��=��[-W�f)��ℏF�Ĺ0�D�c�'Ѿ�bU)<-1�jA����	+���A�*� |��6��*�
h�Ѳ��!�!bjM�I>��hxI�wI�8����٨T�>I2%ǂL�<d���&}����E]U���(�p�%[ҎJ+r���n {�6	���3&ꤠ�0`~ybd�qȱ��]���/M[ZX8@� �9�غfl�eyr�@�c�0h+�𺋔�.IQNthp쀙8	�̂�Ӻ��F��8=�@���j����.
m��8u�5�]�[z����Ɨ]� B���z4h� �J��9���ئ�S����㖍b�:����_n��]	5J�y0l�i�8���Ц�\�P����7,�!�64Ҕ�ۋ2c���t�
U�p)b�ã͸'�a%aХz�J�1���,�9H�D�Y�Ex�
��U�&�iCԱN���e���qr�lS3P1{ADY�}�&�y7�-Udt3����A�I��~�CXH��Xg��� L�)�vv2-�eʚ�?8\z�h���!r: �c�[�9:LU�	AL,Bw�8�Y���|�t�0�O;$��O	:7�I�~6 ��
(�Kʱ<����4},0����)G��e
b��	�4��;����-*��ѐ4��)%��іM=E���ҏ�L�v�B��
h���3n,)���*�y�>�F��%I��\
��@l�Q�u�ªeB�\�$�ΦDh�v*�_>�rDM%I��@Z@DAi�Y�%`+fE,X F��d	Hk'"�:�,8G��d�H�b��d��F"`-c0�غ������������B^�.@���l��x���ɏ�Y-���b$�X����V���UB^�)H���u<���Y�HG�Gr�P�Ԋ��N���[�8�c'R&Ti��`2�>%?���+&�jD�ǉ�-�̽�`�ÉX ���&��D|�l�rN�	"0��U�Ϫm�fP�I&.����p�O"����;O�}7h�l����D���iӐ|��ĭ��yði������}����C7=n.�?��;�`��՚%G?p��A�hϲ��'Ct�+W.�<�Q������03<�F.��2VBl�&�<�DG��q��X��˘u%z˓b��5�D���t@W1;	����y��XKe��(4�p��`�z؟(	�A�-r?���`X�og��p��8�	�nc��X���R�Og�)��Fg&���KCZ(��G �y�dw� x��ɔw��SK�/�\�Ä̙�Vj��dR��<)�Ƀ�K�&�;ǯ�8�rL"a�P�'%��)�<��>e���V?�許'o��>Y��"(D���o^���)@�d�2jG&!O����Y��	J��~R��G*,JT�4!p�rtM�yb�¡Y�r,��̆�"I��"Ƈ�?���ǰ_�x�Ҥ*lODh�6�5	�Q��jKBT� A�'������N`oڏ+��sC�V��i�1�I5�"B�	(*[0A��p��1�DCFT	6����j��WX�|���H��$b��:?đ���D�f�NC�I=Il�E���&�Ꙋ��EN����d�]�	��y�O��G��'��[��/!)������^�)�'��%�DT	9�L����Iz���@JH��#��m(D���Y( ���5��Hɦ,���D)��{�,��
�D����ܦmk�
O�qb!��t�6��#�2D��yA�`B�Xf�U7H�r��$�U����6��䍒�,8��m���&�S���G"ҫp�Xh@��,D�4P�A�
�tR�k7r�2��Q�5��  ?I�F#o4<Rc!:���� P{Gaǲnmv��PN 7�L�e"O)���Qxe`4�
G]5zuFQ�A�V� ��G��Y��~�Mɕ>0D�j�=Yb�l{�
��yR���M��y����	�J=��)�?�Dɞ5~Pzy��jԲ�0=A�eT |b���ʩJ;����C����ă\�Nl���ԠW�vm*6��$P�9P`j���ȓ_ݾ�IhR%,�j|0!�}�"!�?���&B��AA3̐�����۲"3d(N�˃`XSGT��"O�Y��{TQA$/�
4�E���X�T�4��G ԔF��	o��~�"��`���ꄆ��G8"T;����y�M\���m�b3T���9�?��O����q�����0=��M[�T�o�~������WH��X���=+r���E�r���p�J�Onp�d<3�,�=9qe�D����ײJdp��ÖF���$���#�.g��8*���d�� �`$Es��xS!�:�u+B�0
EV�9��w����Z#
!ni��)D�\x�i�	OY�=� �ΉOX�%�PbV\ru���u�ӡ��d(l�����2/hp�#f!!D����C]U�b�+XT�A�nk���!Q�*�\��兟u鲔G��œ�{!x�-��������2�yj#4�^" #Ƨx ���G�D�n Z�'3dl���Lx��p̟�p���i��@6�5P°�X�1�O��@GO������oڮ/f�LcƬ�A�9"�����"�K��Oh�
a�#���x�pL�eL��v9���s�آ=q���!T�eI�(ǠYɢ!Zׇ�~����	>\�P��:����cZU�y���?ظᒈ�	M��	2���D�yf �^�V���8GH�J� [*1�DHba˚�>�X�X�r���HR%_ɨ�J�j�"d��L�E��=K�.]�-O��s��Y�Xr���Ke4���
X�r?�BR��'��@�T&��>���xG�#"��'�(Onq
�F�^�T�"�%y��'떧"g|\���/v\��E|RB7T�t���D��m�(A{���aI0I�g�R1�6蓶C`	��ɰ&�����
,�QoZ�h����X����.	X#=y��m�Jݹ�L	l�ĥ���W���4G��+hz) �n�2�(���۸'�P�C��.>>@i��S�oY�Eyw���,��΃�n�v7K�*��u*�cY�b�U`R��pܰ�}��,�NxJQ�T}3��Ǭ�'����m���\I�S���g�<��ꉀ@p
��W�#0n��(
���(4���}��
��.f����OQ���cA�,� ��3d�T|Y�DfF:<b���M�:K��a���
�J��������#:�Zp ��+a����]���nE�-^#=aѪ3IfH��M;#��%S<���$�3zq���s��H�' H� ��Ji��el�|���Od$�Kʒ%4z�e��2Z9�]��}��Vl���nIh�O
�=h���%_��`�H��X�\ē�<�Lڵ���Y�<��oE���~j�Ab�FQP�)D+%8���%F�`I1V)�����h��D�8.���F��/�ͳd���n͡�b�O�����_=O��ʰ�?#<���
=���_�/s�d)*�`����*<�^�3�N�Lx|��"��~Y* lںp�	ش�G_x���i�;_&�ɻtB�*#�:5#2�&�`�b��%��=I#�"��3 G� ����"�,!*'�g�<Q f�.~����dMu�^�p QbyBG@4Z�cE��A��S���z���B�| x�C�I W��m��O�"�l�ñg[
��У�K-�ax�`^�5�l���tiI�Ŗ$�y2Al}z� .�)���K�Ic�'=H��(�Qn��RЁHI6�P
�'�pR߸/�����ʞ�Io8��'��	��o�&K��庅/��z2j���'���hǩS5T���?�*���'�,Qh#Ҍ	�ڔ#uI�<*�6�8�'&@��p.#�6�3�X%֥��'\h-6jBM��Ћ��jk6h)
�'�j�HP��b�V\�őg�:Q@�'�h�&��1`���c!ĝS,� �'�8Д ��U�h�KcJ��TX�"�'�l�I!�W�&�ң�Y8T�l���'�
 �a#Ѿ2�!�ǅ1p���1�',���,�v���ҧ�DN,@�'�6�Jp�F�肁B^�m�^p:��� v\�d�9�@ԛ�ė��$,i�"O��X0IY�-�����(n � �"O��Q(|ݢ���_8h��H�"O��(�'I��{�,^�rƲ$Hg"Onȓ�$��� �k�K�̒�"O�ѪsO��5;��ވz�B��"Of�떠�/c�L�uӫ'�ʐ��"O.�+�ݭP,���жRt��P"O g��G�-e%�!VtL�""O�"F!M:�l�{��^)W�͂Q"O �$�j\.��Ei�H6^m{�"O����֑r}҈H��c����"OLL� ��,ڝ�Дh[���"O8c��G�A.����O���R�"ON� L4R��`@�xb�T��"Oz����5�xhyĂ�j��3"O.I�V�^0C7,��6C[�e�i˒*Oz]�Uȝ�u^x��Q�͆Ŗ�b�':191B1,��Y*F���$��'h~��ԫje��R�e�����H	�'��#���G@DaQW�T����"�'��}����0�����o� $���'��z�O���t�r�C'.K<Գ�'��kb+-u�mqEˡS����'\�5��/�&zgZP�4��$5�c�'�y��B��E����^)/� Г	�'`b�5��u̑9��"�4�	�'P�%���(T�p�'�'^��'�~i*�/�'9d����ޣ7�9��'<H��D�B�1�Xai�Y�
Y��'ญ���G	C(��do�W �*�'���ہ)ݎ~snh�$��z�E��'((`Eg��R^��� �ː#�I��'4Xɦ�TR� ����kు
�'�P�1埲�&زSE��~��'`z$+��2��qZ��~���'�Z���n���&�#S�?)���i�'j��aȓ$楠b&��݈�'!��� �(9D�����W�T��'�dz�F͒�Yk.ٻF�"T��'H����/~��|S��� ,�$;�'ݔ��3��Y^����7i��X��' �zǧJ t 8�Q�~�d�Z�'�N������ 1��Ȣk�<��
�'fH�����*p���+,�a��
�'��tC���3fn����YZ̴��'fv��vbR	F> �5//N���R�'�n�bʍ	C;���e!I�lLB-��'(b�bmB�ybq�veK*!��)���uB�>�lK�a&�0�ȓc�r1I�'I;LG��7���~�V`��̐:���:Xd��c��x�L�ȓS�IPG��3�,���'2�n��ȓw1F"�Ҟ/rb��@h��'��@���P�>�����	�*�J�'fj�I��F�L�������
�'g�y���33��)���45�]h�'�	s��ٟJ��.�E���s�<�%H98徠SB��' _2Ⱥ �o�	�N�l�e���ÀR�F���ՠb@�v�!�T�;�i{(K��+FN$5�L�&�;�B�7�q��'ͪ�����^}><��aEoL��'̮ �6O�&���a����I��ǜo�-X��[���04k�4A�zݩ4k8M8l\��=O�T�ϧ\�y�I�� Q��)�7W�yi�Œ_�-�b"O�y�6c^%��!��F�l R��՛�D�3��<��"��>E��+$���Kя��rl��b���y����7��	����z��E�&�B�+���Op� �	�R]1�1O�r�I 0,����N�(�J�DO�Jai�;,�Q�n7��=�Ë��X>���C �p?Y���1Ɇh��B��"Xl�"���F��aF�?FH	�B�>!V�
�^9�9�64�_�<���iu:�#U�މH�E�&Bw~b
��$$�V��D��S�k���rfQ<2��i1.[��jC�I]�|3�e������Y�o�.��>)�+�-�n}�|�<a2፝u`��rU圯�R���U}<iA�z�~j%S���*�L�W� D����䗜F�H]!d�V���QB��a:�xbŐ�XP�+��x��'A�(���
:���!��y�挭
��D�Q�T�&�P$�����jO�X��+�)�S�oJ�[f��I_��`3��8*ԖB䉂H4�!�oA+�B��ˌ��B��$bn�2�A*_p̳ѡ�F"DB��=_�ya卟l|#�JW�C�/c�@Y�C�Ux8�g�+z�xC�	iv"���iM4QΚ�0ӦG�E0C�ɯR���BF��g�f8�Cg�
��C��%:�"\A�ć�B�z4C�BT�N�dC�Ʉ{.P�0!(D�i%0����$%6B�I�F�ș���F�;h�Ś�O�>A���'v�̛�F�S⓸9��[ �N"�����]�8� �ƢW�3Q�01r��)�1�|a�����5Cu��9<(M1v#���9> Y&����#�hG�v�X�9K>�;y����O� ��]A�N�-�@�'y� dLJw�Ti�Oq������@�<oܩ����U�ҫvN��a�J@�ȍJ��]W.�b/O�W�%�S�S�u1ӎΨ�Wj�.���1-OH0�2`�(NL�x�_w�e�ARĮ�w*�,�Zwx�a�b)b�#��=/�I�g]}2�U>�Q��({���0�΀?&<3e!�8\�I5��B^x̺�B2W��� ՘Q �z�E-�$0c�]�?�Y���C_xĒq�C1QT��D$q�|�B���:�1�>N�Ug�D߈$�2�S%땠J���X�oԚz������v��8�0�߂�V��w��.k>�j̱
6�p�/�}�����q���@3�(�Bΐ�?ӄ�e��<�����O�顆�/�v�ء�<�|�w͋'TйۇbФQ�M���	�Vh�RCI9x$mj� ߴ%t��τ,6���'�P�W�e����T`�2�i�9�ǔ�,;�mχ������B����$X�t^�J�kF�C��	�
�c���S�r�h���;R���Cq�A/ t��y��I7l�ι�bO�8��2G^�DR�\��j](-����{��z�ڡ���h9,�c��2ۂ83Q㜎$���c=��pq��H29���1bj;,�K��
4ז$q�܏#�yRoY$|~`Z��)'k��rG!ǁ"��u�G�f�|�0�ӣs�F1QK|b�IcwpݣЪ
!b)H�z�O!b���p�W=
�� JF�*d{�J�i�arz��Pj"b%T�:v'��C��ś`�b(*��^)|�h�r�c}Q84�@����s����FB"T�!�C�-Z�0 �Qr�
�NEg1$պuh����O��l�D���,Y� p��?�vD�<�㒿Y������h��+1bQ�j��;"OѦY�w+��9X5`P�;p#F���%~C赲S5{�\yz����g���J2)>�q�ǈu�<j��+&G�F}���>�N�{�H	*��O����	�#; ���O�=g�4�/O����>[b���3d�c�J��ʱ��ŉ(���+ �=1�a�@�8PYrQE�E)t2�j�Θ'(d���O �?�2�&�'�>и���np�1�O^L�q���y�J�T�����ұZq��Q���7��C�{�][���S�}H�y���Ҷv�@��\�@$��{V(D&,��PG�$�L�2þ������htJ�MN,�y�eZ0.Z�҂�	+�h�����.	]��@�/*��'�>��8B�(���G�k�6x�0�٧"z�C���vEh
�.d"�b�� )*���$0R��h���,��=)ac��AF�,�"ă�m^UJ�'Cr����ơT�s&8A�i�v�Hċ��aaXͣQ�=��8j�'��ɓQ�#=�!p�$M�-��(�rE��z-�WDc�O�r ���6m̹�@a��8��'vy*�XR�Z�()k֜E�דq���u�1}"�0j&��L���� �nU���")D�$1v-O���ذ�ņI�^��pg�O��+ �\�V|�ۓ0��r�ը[԰�kb��
_����	�Bd�\���	�� ���G�p����P<w�m��"OLX�Q+�>I�^��N�!RP���I*ye֌��t~r�� U�ư!q��ּ@��OR���Β�>/B%X"OX�@�Z%d|�b��~���;��� 6�]RQ����7�U*4bD����w���ȥe׃?NP	��<;?��	�'�
9�P �}�n�а��1��"	~M�K����D �g?yTe�Hp�l�"�L�6B�D�<dJ֠OޥjB��l$�t�`Pǟ�D�ܨ#؉�&b�W�� �a&E�y��8����:kl(��,|O|<�F��{M�(�1f��1��U��OJ�������B�I�0�Y #�&?��T��	���thAaYm�=�p��j�O���dlƩ4hhrQ��NC��@�'HX�q%�#h�b��8Lahx�ua'[QX"��)��7�g?a�&�:OR5��B�;�Q����|�<aQ��S>�1xv��?��J�kş �#��bMA���k��D� �*G�4i�+�*�$�[��4|O���9V~B]� ���v\%���7N�q�$#&�C�I�uZ{�J��BO�zq.M�n �"<��|��0�5ʧ�N1���m����b�tԆȓC�K�T�s�xT@�%N�=A�,	!D�e�D=*��|���'Ŗd)&��s�4����(<�`ݸ	�'��=H���-k��H���F�Vih	�'���� 	P��G`�<����'�ܔ`�	�-�<���h�0Tp 	�'F<��"7�I�%��5%l��'ҵꡆ qHp�kV��l)�fG��ꡀ��y�i�a����͍�XK�؃c��yR��$"��8c3o�T�>�Z'B���'�ҙ����HF�ԌC��&��'ŷU=0�F�� �y⧄>e� ���� ��%g�?VxD�k� ��
xZ�U�R�|�'��m�R�@�3�ZaxR��]����'���G��b4f\���*H�R���ߜr\H�x�#ǧL����_�sS̔Z�͞)S-"��F�
�N�H}���)�p<�����-�"�BU��M�hJ�"e����-.&�B�&x�9�G��nmt5%�䂲L� M����T<K�Vd)��;�	%Z,�����`�tE�����%��vH9HP.�������Z�s�.]�Ђ¤��)ʧRW�E�ň<���p'�$��8{�E^[�\�H�S�(���<�C���s�z��.�\�hd���<v�2�`� E0��g�)R�uN��i#�Ț�j�<5���2��0X��ʖ���xR�
�S����1oP�>c`����+\�'L��=FC�/a_�pX !�10�vnC"7 �X��J�N�p@��%��O�x@�\�-�4IZH|��	2(]R1`ٿdx� 4(M�^( "#�&$�Z�}c)����8I'H�<�B٫d�^Ky]!`�(�[Q���'on�b�&[��ٰ%)_mTtbЦ�-GC�O�}�� �	"���~�4ġ�oH"}0�+�>�+ߒA �@O~�=)��R\��%�[Tp"�#UX���9���o�&slD�ac �Z���)B/�4�418�L;ܑ�P�O6��C���80�D��ɴa��h�!�^J�	�)m��i"��%V�����,�-�B�I?3s�\�Ư������g�t�B�'6: ����V�S�'(�nP���Y	'N���fI�-�p�ȓ̮�q2�J
�p���L2@ ��;����x"�x�R�Ҁ[Gn�ȓoe�1S�P98d��f�KH����O��@�5ʏ0&�X�Ɇhx�ȓm��"���
|�]���k��ȓe���YiՐ?x���zE��ȓZ��-����g�DaFf@�Y}^A�ȓ< �hst�%b"b1�%��m��@���E�@M=w�Z��ST����=qv����*d��2ˏ�)� �ȓZx��۷Zj�0��%� �N`����u�!`G4C�(�����
V^ (��p�ո2�D�$2g��q6���S�? ��hpP�N�bW��+�8�*�"O��Ic ֞)� ��fh�V�j]Y�"OX�Ql�=3��H5�ЉZ�z|0#"Ov�Z��.<�`c��+�lEȆ"O�ݱ�!��O:YSO΂ ���"O<L��7��5N!Y�&EC�"OJ�Xf�Kd�����,W��	ӡ"O4i�ɮI�m�#A����j5"O�e ����p`o�9��"O���bDA�U�tS�`�]��5	�"O��p��
4�L�/Ґ5qD4�$"O����C� �YS�.ech�s"O���G��*e���I�HF�u(�"OpqPo�+@7F�S�c_1_  %"O�dz2�ԅ�RjV�bk���D"O2�+���<z��_#D��"O$��1G�-.�,`�fDs8��"Ob�in/:40�4��)n�u��"O��a၍R��([ M�0؄�C�"Ox��򏊗��hY�K�;%�0�BW"O �f�3s>��PQjŵ.ȶ�E�'T�����7��y1�S���4��`�d��'���A�Oܞwg~p���^�_�ɻ	�'k�|3���VP�md��#�~�a�'^aI&�*}�CVP�iS�"�'��-� 	A�(��}0��`,Đ�'A�I��DmE��ht--_��$x�'�9���w<���\:V�^\�'Ӿ�K���K�8�A{6¤�
�'\��{�I� 2_���g^�k�̘x
�'�$|�"+4�HqY��B�,��a�'�j!S�+N�$�� (3Ϙ��� �'XP��ЬT�~cPUB�E� !"m��'�d�h���.B�4�AN�&D����'n�C�N�hsl�����D!;�'U�Q`��	�^�����L��z�t	3�'��L���-A搥BR�E	s����>v�U	�Έ��o�U]��`�`���6PP7����I�N����:�0|ꄬ�Q����6�=1��8���[}2D�4q��̀Am��n<���)\ �\��e�7�5#�ɨRT�jq:Qty �R1���?�����}�F�H�#ϏW�b�����8P����H
4?��I/)�����I~�PG9�,����3\qBm��B�t��C�M��8��&)V�$>7�I�Ck����ȯ �J��T����f�9�F٦� )q�(1�0�"q�t푐Z���բ�{����R��9B�վ1�XаsR��	6���S�L�1>T�6߶jӘ�i��=?d�0���kb�io:�'j��D� R�.�rE;.���
8��&w2X�',LOd��r�$<�� �oS�y蠂s"Oj���ҹ^L9�6m̑<\VA�r"O��hG��Z����N��2"O&8*��I%T1��J��N���"O4�7!ې
iV��6)�=Vt����"OȩہI 8$Fn��ը�U?�Xɶ"O$�A¬��Z,*��XRR�a���y��L�99٢�l
bր�����3�y2�9R_�1��]@�Ur���yrB��/��]H��[\�y ����y��±!��l��YXc�1���5�yb�
R�����E{ܭ)e)#�yBO�lgr;T�x�N8�d�V��yR�M? ��e�cg�o�t]��M��y�J̡h�a�j�� �q�ԟ�y��	��� �̼2K�j����yB�Y11��M�q"ņWX��!X�yR �;-�X:2�B�Jo�x6H�;�y
� ji��>s���C ��>�:Ecf"O\�@3�]�=���2��-V�h��6"Oy� /^yr1��D���;@"O��X���A"A(d�\�]����p"O@l#fmu=8diA
�H ԉ�"O�x��Aѡe�2e��䜨=,�Q�4"O�=醌��{�ĳ�$^*L0�3"Oy���N�\r0A�x+F�;�"O�h#kܑ2`��"�D����"O����2 ���ҫ�E�����"Or�R B�&�Pqze�#��$�"O~�S�#ܚ��\B�Ä ��V"O~�`4��8L�~��գ�
Ͳ��"O�)*3D�.%՜��V�Ҋ�(��F"O��@�+"7�� ���ğ3���"O�Y�/A>(�)�m��.�����"O�g"	�l&\X0bЉLJl8��"O�)Q���?�\�#�ȏD?��T"On̹�h[{�zq��F�,&�4C�"Ob�9g��b T�t�߭E��"�"O���d��W	* a@�ܯ~� e��"O����8B������Jb}�e"O���iȯq)�׭�+.>��6"O�&G�w�D  BP9$4iI#"O6<��́�FxH����׃_ZXa�"O� �A�X܉S� ��W�65j'"O�aD�0R��e�*$�B�"O ��G�$u����H��] �"Oz� %G��f�D�q��_5BED�g"O�Ph�C��L��'E�)Gh�3"ON�0�H�҄1�a�^���a�"Oz��4hƁ'l��Շ�s�E��"O��5�DKӄ	rÈW��&0+R"O���uZ�u ��@z``�"O��� jHA��mD�`�2P�E"OZ�yG���W��@k 牡��%R"O�j���2xpD�:����y��@�"Oy��8�p��P������"Ox�Z��%�|��2"�ĹX"O���D�Xm�UI>����B"O�-hR�D9\`�"�Iފ0g\�� "OrpiQ��,�p=i��%Q>����"O*]+�¬x�u��	\�*7��"O�t����c*ƐK��*�H0�p"O���ƚ��Yp�B%;v�X&"O�p�@�A����q� ��A�,�x�"O��ǜ�t�H�hVf���"OD�(䊐�&��STH؟VV���S"Od���)�!$D�9����ډ�P"O*�b�]�\�K��6;�)c"Oj�9���uX�G��Gɴ��"OxX��B7{%hHk@Ä�|Q�0ap"O��S�IV�x�J�croTQ0"O���!�]�R'��+���u��ɫ�"O���G&G^�3U���A�l��"O� [T��#-+A@ �?	8�"O@�ፗ �$D� �5 }X"Od��C+�5n�I ĄTF} "O���\O�l�)CT0j��"O0ك��-oā�Q��';�.ȁ�"Oj��r�Ɉ7�b@���.	�֙ �"Oz+eH�&P��@Cg�����; "O.�"ǟ?e�{AK�\}
��"O�Dh'��$>=n��T�Y	5m��[�"O� �:�$8d~E����vl��C"O<�ɒ��8�!3�a�{]̨�"O�5{�b(N�άr��[G0�c�"O����r�l�'�?���"O��kA��QT.ՉD�Ҩ-��IB!"O��a��X�.`���&�J�m���A�"O��BG��+g��Ac�M�Qnv"OfyBPȉ�2s¡bQ&�K*�z�"O�U#�.H��	�qc�BB�h:3"O��1A_�tK�)���F=7Z���""O��b �4q%���A�6aIna�"O\Mc���/w���(���MDQK�"O*�դ �yɉ�a:�1��"O �@3n�l}Ԅ�ņ�)\����"O�uc��^��i_2��A��"O2IZ�J�2.�F�jE	G�6�r4��'Ĝ��q,�
B�s!K��"S����'4��Cd@�O����w
F7�H�'f�WhX�?)
��B����'~x�Y�EŔ#NIBI۽p`3�'r�e����^�iCZ���5��'�0�B�[�y�P0"����x�'��l
���G�vh��]}�X!�'}�9���� �FP�'�8�
�'�X�1B�4���)��Kv�Y	�'(�\���ٷ�T�3l�=Kr%��'�����U1����2�D< �'-�|�iƿqL���4E.-�D��'�d`��M6��q���[�E��'Z��! �Y�7<�pj��x���yR�sLd�kp�]�Y�cU!�y���_Vb��!EH�u�He��>�y2��? �.1p5gp����*8�ybf_�ؚ�RƉ.���� ���y��"r�$<d�%�|[��X5�yk�81�LĊd��.h�0J3�.�y"�6&�Rb���T�е�3��y
�0f������RUИӁ����y�E ����Gu�YCq&���y�%�z�\Ջg�:�fhhe�O��y�Q7V��]��+}��2�J���yr�[UI��M�&3���W4�y��I(fG�B���F���A۝�ybaL:F�&����S�E�☘I�9�y�#�r�$3�k/S+�遡d 0�y"&�;}>�d&C%@�P!��	�yR톡A"̵h��Ӌ4e��*ao��yr��`�x�Eۅ;u4 !��B��yR�e�:ݛ�ā,�dM2���,�ybI�Q����)W�Pz��B��y2
���R\��.��O���t�8�y�A�p�tr�jJE�Dw��8�yRJϱQlĺt�
i��,!�nR!�yb.ɔx��V��8�T��%⟏�yr��d�p����x���kB�0�y�#@08�^�w��xvj�S�B1�y�#�Q����B�5z�XM��L։�y��̩N��"��*	�F$޳�y�'�!��U�Z'�0��ɘ��y�EO��`I���b����#�y��iª}��ڴ�$I �]�yb��zh�H&��|��hVl�7�y�jòx��K�i�> �ۅ����yi&-�zy�d�~V[��I7�y
� �r䄆�(�؄Q���+�V��"O��P&�>1Tv�:�@�q�x���"OZtZl�]��h���N����!"O�����M�l��|���]<Et���"O�x���^�&��J�-!F� "Oȭq��P� B�<q�a��vQ\�S"OP�KHQ�Z������"QN���"O�U㘹"���F</M�Mav"O�\Q�J�2:Bx7^:�M�$"O�t�H��@[7�K�1*H�"O�둢E|*zx�r�� >&�z�"O����/A扻�*����#�"O`ɐ%��#V�Jpa��(x.\Z�"OX ��Ō��m�%y�ܝ�Q"OV �*֘Y����nԼ�j�*B"O��0u��mpT�펷�6���"O��c�"�,Dp�7΃����V"O��;�l��yxĉ�������E"O�9�!��) �����	U7=�HE��"O�ِ���l6��V��(1��0{D"OLE��F��R(�&��-!��c�"O�!�q��J�jy�E'�FOzi`�"O�X#����7�T��&�G���"O.�0�)�"r�B�*�k�)d�A�"O�mC �Ѱf�����*���b"O�uI�C�'�f��H�#:���V"O��9By�h��#��.;���1�"O���܇?��}�V��+��4"O��BD$KD:�ӑ%#4r� �"O,,�T�Ŗ9��he敵%.a��"O��3�+��1��Bf�D"�D6"O�9	ca[�`> I�a,�X�m��"O\���	Рn?�L�E��#���"O��{��޶z(h �KJ�_��E	"O|tXUcH ��S�[��zl��"O��4i��58b�q��� "bѢ"Oj�J�\4�j��u�p�&"O�K�:R�Ċ�O^2F/T�p"O��
'� 0��a��]���ا"O��$���yb苲Q��E��"O�1p���S�h���� K�"O�yc��+�
�I���x����"O�=�!C)b^u6d7u�Q1�"O�0@ό��r������w�� "O|�(t��=~�����_?<Đ5"O���M�:,��C"�}IF"O�-K�봀Q�.A �{d"O*��6�Q8x���[#-_w���""O�@�եY�x�pX���^\�IB�"O�`�茻Z2�z/A[I:�"O��t   ��     b  �  �  �)  5  X@  �K  �V  �a  �l  qx  ��  �  "�  ��  ��  ��  8�  �  ��  	�  L�  ��  U�  ��  0�  ��  ��  h  � U � � �  �' &. 9 �B �I �S �\ �d ?k q �w Dy  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hģ�%�it"L�B�x�'�6,�pvb�q�ΚO~��Ey��|Z�(��-B$k�-Z:y乲6�	d�<y�+S�
���w�þw�����k�W�<�WO�,�R�"2*ܥu5�@XI�<�2̖8��"�m\�)p�ESG�<YƦ��S�T���m�<`8$��'o�<�q
44���rT�.U�X��k�<�T@),VzH���F0��	�1o
h�'a�DĚ�GJ��aj�(K�f��tO��y�A �GЊ�/����(?N`�J���x��}����b(9����;TI@챗�Jn�<9��6?�]�s�ߟx�r���B�<���4V��ع�V&%���*�v�<�T�D�p��sn��U���`�Jn?��'�a|�n�1Y���#hF�M1�i����$а<Ɉ�DJ�ax��E;z��U �o��!�$��x���He��4v�&���0�!���
b�Y&���V{�.".�yr	$���K�2�e��W�ѰGڌO��C䉋���� �!�dPc�:xB�	�Re�0�ɐ����g�
�u�B�	p�,\rCiA<jS8��� ɮ)�&B�I�U�����ָ&tD���H�xLB�	=���+[�&�����=��B�1L�!��f\V�.���Z��C�	1D��+����n�Pp ��dO�C�	�n8h��ŚT�Hz�왽RjC�	���A�jׁ	o��@2c׸O��B�ɢv�bTbW����as�hUp�B䉙l9�X��A�|�QҠ慂��B�'�41��E�t�B�[#�u�4C�IHc��눫q-4La�j����B�I(4��p�$�{;�!Z�%��fB�)� BI3āW�����Gف[���0"O���A�%|�|@��Y��%�"O>܃��P�_A��r&�Ƽ�ƨ��"O�l�1�ˮ'V��%����r"O�dK�E���^��e^�z}�7"Ox�Tě�%'d�A���|�@�"Oje��Fȥ^ T�8�j� ���f"O����)D�й��iB�mǐh�"O�<g��]����i��SU��"O��ʕO��w46�Cuj��%UJ�(3"O�����-L���F)*VnF��U"O���eX9Sn��2HԳlQ�=�W"O�����ݕ'��[�� �A�ł2"O��G�'�x*��T�c3��9e"Oũ-��lg^�{Di�&p|pc"O�Q�t/
�J����v�+ud����"OR��u%��o�@��p��zP�}��"OLxd�Y��p��t �cL�0��"O���J�_�� a�$��>7��&"O���c�<q��Ѥ�W�X2� �"O�EZ!,�,a~�IA���%K�bx��"O�Ej�IPIl�Ё�&]	
UJ�"O֍a"�W."��('����Q"O4�I=#����� 8$W�(cS"Oʡ	�jػ�}k�d�J��Q��"O4��FgK�,��y)�DQ���X9!򄛼[��2'I=FD��K�Q�!���-�Yʓ��PFQ�f%ܟ�!��V�:l���O�?H,4H����P�!�)Gv��a��0%w����&!�dY�zC�iP��l{��;2��~�!���D^���!�H!Hb�K @��N�!�*��p��BN/VG������k	!�$U��^�Qu��'%)����O�)�!��a|M�n��T$�tB8$�!�d*#%n�S3bV��jD�~�!�Ԁ�`��R�*.��&��R`!�]z�e�c��d5�=*���H!���`�ԭɗB��\}<���Q7�!��%3n$8
��Qr�!C���<�!�$�$�tC����p�NHBs��n�<�BHء9ju�F�Q&>����Tt�<q��\6_|�Q�`E�#W��L�*Ar�<E�P�Pǆh�D@��l�{My�<��mS)w[rqb�V�)Z�D���k�<	q
b��zc�ڌA.�B[d�<9�K]��ăd�^�7N\���x�<iO��C���wd��q}�1z�&Nt�<��ӿO��!�>!׊�����Z�<qQ���Oq1�$�;Y .؀0�o�<��c�.���S��Y��f��e�<��x%�X(R�Uečw�_�<!��<0ny�j��T���/�\�<Q��B"�ǉ]�Ct��!L}�<�r��|�xA�!�Qd�a�m�v�<a����cz p��{�A��K]�<A$��7h�)z1새�Ja1G�c�<Q7cϓ)\��i "jތ\�PQ_�<�	�AI��	"Tu�^�q)g�<� �?O�.Qr�\�X��@�@y�<� ��&� �R'@.[m(@��`�<���Բ�2A@.<���5�]�<f�!E����,�O�Ys���r�<�w���TƢDⳭ��*�@�J%��k�<� �p94/��=����d�V�h�d!�"On����7�:�bfT<rr��3"O&lI�� �|�0ur䤔�1�B�H�"O�l!��ы2��HT�هr�E3g"O	�fC= X!a6DԛJ��'���'8"�'f"�'TR�'��'�.�����] 5B��\�$I���'��'72�'L��'K��'�' ��Ǝ��&� &*�6'z����'^B�'���'���'�B�'pR�'P��rRK��1�-�h�<�uaA�'�2�'�r�'���'�b�'����=Y�l�.W�%� �CQ��5!Vlm�	ɟ��֟H�	ǟ�����I��D�����1˔���ڮx(��E�|9�\�Iß��I��@�	ğ �	̟����t�� ^��E	�>o{�Ē��Ը<4��ԟ���L��ҟX�Iϟ�	ǟ�I[�Ɖ��I:J�f��t�*�	�I����I�L��۟�������	ǟ���<���x��qzb������Aׁ�O&���O��D�O����OJ�D�O����O:M��Nݻ8� Z���?>�=�Ԧ�O����O���O����O����O����O���#��~'Ri�oA!\���O����O`���O����O>���O��D�O�y���P�NAb!�ڎ&g�Pf$�O��D�O���O��D�Ob�$�O�d�O�l��jнkX����P��dP!#�O����Ov���Ol�$�O��������	�����e��WL^����9��yJ�-Ƹ��D�O��S�g~�gn��"bJ9�j�[ֈɟTu!͗�w�	6�M���y��'��QRF@�.~�v�jUĖ6�H]���'R�\Y�&��t�'\��t�~2�K#@���s��7m���%-Q`��?�-O�}���av&�Ȥ�� V)�}�rʍ�*�&�����'񟌁nz�91R�_�:��!�Q� ���#`�ßt�I�<�O1��5��}�z�I�H4b�y@�C���ى��{l\���<�p�'kp�D{�O|�K�-:������ l5�)���y�[��$��c�4 ޮd�<��$�-���P�Kݵ!_4\0�ȏ���'���?Q��y�X���5���=y��!Dڡ��$���"?a��b/�D�r��Z̧b.�����?i`��#�FS��d�r���i���d�<��S��y��
��`-(�ȗ8e�j	B����yb�sӸ�����t�ڴ����Ĉ
<y� 9ѧLS\4�ih­W��y��'��'	l�(1�i��I�|�E�O��Bh�)G�"a!X�ة�)���'��i>M�	ߟ�I�x��<~H��ó�ߒD�P��mNL�'oL6-�"�����O��$%�9O�
1���A���Z����R�`}�'��O1�,��������L-TƦ���ͅ�a�A�Φ<�&�ѷ����@�����D5I�Ty�EY1�t%�t*�C� ���O���O��4���v�6�O�n	�(�K�P��w��=T�B��c��y��u�⟸C�O��d�O��"��c�"L&=B%��h��m*!�dӦ�a�j�C��!�'��c4�^'�~���6�ȱ�<y���?����?���?!���S�o��,ۭ6�}��K�`e��'���}�P�B�<��i3�'\������(�*_�!�R���|��'1�OoJ�0b�i��I5�|<'��T��MH��+B�,A��Z�qv�D+�d�<���?q���?� d��4��[�%�A�eѩ�?�����D��5���ݟ0�IΟЖO��aU.OP��T�3&Ub�K�O"@�'���'�ɧ��^(�FMp��4m!8IQ!�*v셢�T6:jA����<ͧX���Dۗ��W�F!Xd�7Ú ��/ܥo�b3��?1��?��Ş��d�=)�Bۢ8���b���(�R��9k{�%�'j67�������O��T�;o�=�7D�v�^s�,�OB�d�|},6�??��ěiN���<��FځDĴ�CcT�&<�B���y�P���ϟ���ş����ԕO�dXe��	���R�h�;|����c��yjP��O���O�����Ц�R�8e�WO�.=�T���mB���	�I���&�b>A#a��A�\�⠲�-7��ͳ��̾h�F�̓+!D�"����@'�����D�'uޭ���-<�8*L�$[��s��'�'�RV�`��4T�H��.O��$��V�y��"ն$С#�$'<�T��O����O��O��	gH�28n�Q@l� Jp41a���(C��g�hxlJ�' Θ�I���s�˱>3V�� iX�t��a ��ȟ<��ڟ������D�T�'��KG�P�26&�I]F����'\R7-��J �KP���4ﴵ� ߿9��0g�=&�F,3�>Op���O��D�)��7�/?Ig�è��)Z��>�p��Y�}u��9�m\�+��HsI>	(O���Ox�$�O ���O�8�V%��v�`����x��B4+�<᷼i��(���'"�'��OB� �/� 'A�\ 2C&�Ep ��?���d�[}���='�vX)䏄+\3� �SE�!���?�p�h��'�8 &��'����Ȋ�&���TdљZ�&]�f�'���'\����TY�@8ݴw��@[��R6��h�y ��4 Ψf���������S`}��'���W|b%)��Q&�J����&�^�OT����'k�`z��U�?)rԑ���� H��a!F�F���`͏F��$�:O`��OJ���O��$�O��?�S��i�T��A�(z<1;2E����IꟘ��42�L�/Ob�l�K�	����<��VI�,G�$����ܟ�[�z�lZI~B�� z����ou�����YT�|�����Qg�|�V���(�	ӟ �iQ�Q8��G
C�?�R�qĢ�����hy�BtӬ�ۥ�<Q����I��W�JcDᆗ�p�X�H��S&�ɨ��D�O4��%��?���S�R�#M^�h�,����VVHR,��1���A�q?AK>�􊆸^��PK(	�]$-J��Z-�?9��?����?�|r,O�n�7k⍳��Nt||s�J�� ����^xyr$a���Ls�O��D �^5��NV�:��`\�M���d�Ot���|�0�TMƼ3E��O%�] 1!TR���s��+S� Y"�'��4�I̟4�	�h�Iq���P9|.h�S=qR9��פgV7������O���%���O��nzޙ3(>u�$A�I�:&z"}��%�����D�)�S�[�h�l��<�s-ɲ��A��)b8�8����<��6��Č�������Ol����3W*aS�)+n�ܰ4��#;�x���O����O:ʓH��V���72��'��G��T�~�Za
+2l�4D�Ӻau�O�d�'`b�����rC�ȶlvLm`u�@�!����m���ғ㍊
Fny'?����'Cn]�&W�(�f�]�m��ac�̼rW��I��p�	ȟ���H�Or��U븵�B��+!6�2(�7 2
~Ӡrf��<���i��O�N��1R�jV,�7u�vAr2c@�]x�$�O�ʓC��p޴��D$<3\��'1��4EH�H�Y���4N�4sU�!���<i���?!��?A��?頧�p5��P���D&x����N��DJΦ���䟈�I��\$?����'��)"̧'+��q��hDl(@�O~���O,�O1��E���˶�b\�Bf��F�@��ͣ*$�l�+�<YC§?���$E/�䓽�_1k�1a�* gCJ|�A�=.��$�OH���OJ�4�R�%���B���AƇpC~`�	��k�$M1a���g�*�<��O���O(���D�� ه�2�m��N5,$`��ln���;��H�����>��]�$�z(���1BLP�O�7��I�����ӟ��	ԟ��IG��.�1��%I/�:�L�j�`�*O2����0"s>����M[H>���:Ӑ��$!Ʃ ϠX�4萢�䓰?���|�s�'�M��O�a0�YZġs�/5�`E�Ӭ�9Y�\��'��'A�i>E�Iҟ��	!�(y��h�R�P�)E~�Na��ϟ��'Q�7ǺR�t���OP��|�L H�6�𠆤bvth��Sf~�>i��?�L>�O6i0�M�
]I��B 0X|�vC�&��h�iw���|ڇ����&��ԉ���ɒ�N%$�
`C�̍��X���	��b>u�'�\7Ӄo���ٗ_!�F�J���y�����j�O��d���?y1Z� �I�f��X�G,�}���"5eގN"���	՟�ef��5�'U�� J�o�+OȭX����@��i���	�\��5O�ʓ�?A���?!��?�����Й{,*l{��Io�P�Y��@#=�-mZ�n�!�Iʟ,��c�s�LR���[�'B�F����U�N �v�r����?i���Ş]U����4�y�'��a�B S�
�*6�*x(^�}��'�B R�+�k?�K>�-O����O"���#�X���j�Ɣ��l��O��d�O�d�<��i� B��'�2�'��@�ḋ��.	?UAZ��3��d�s�����	}�Ɇ?����C��m*�� �aK-�>��量\��M��/�y?��o�$��q��F�R0��&������?q��?q��h���$��pP4[g��6;�r쐣#S)/(�$M���2sBUOyҨq����]�o��e��K_�P�^���G�0v�IƟ$���h����uWB�1��.ك50���'R�N7T�[�f�� 18%���'G��'��'�'�@ܺ5�V�DO�0fy��MC~��� �Mp����O�����D�>a=0=�e,8{#z b]�;܌��'���'�ɧ�Ob�!13*Gs��M{��ȍ�"h0�@1Q�r���O�E�� [��?��7���<�7&�1>��s �� r���ssL�'�?��?��?ͧ������S�����j�#X�@����J�v�k��l�\�ݴ��'�`듣?)��?���SŌ-��bL��E���=@`�����'	^��%�?1�}���[��c6m��bA�� ֞Y��,Γ�?���?Y��?����O�L�d�"h��' j �:��'DB�'1j7�,@��˓Eo�&�|⁛�T��I��O(�Uj��4�'HR���4��!_����|��)U�Gy�@0 ���'�p����'gɞls��On�O���|���?1�y5�0��o�w�Cu"�)V�ꝲ���?(O��n�+J{1�	����	i�tᔶ�*4 �È\T�]�������F}��'w"�|ʟf��"�
t��"c���[`J����-ؗ�f�R��|� ��&��Ёg�ָ�d�6<�z4��ٟH���`�	��b>a�'o,6�d��� ��6S����H��<���+�<�iS�O��'����W(th�Ą:��1T.l92�'��U3!�i��I
MZ}9��OF�g�? �8Hd�z'��Z�A�y�&A��;O�˓�?Q��?����?Q��� .�TAa,��vw<x+�#?��l�XI���	���IJ��矴��������1B�}8тɔ!�p�Q�
�?����S�'ڰ���4�yb
1z�n�m?�l 3��6w$�B�}Xv���'t�'?�Iݟ��	X��%2S� R,Z�����F B,���L�I��0�'ڔ6m�,��D�O���N�<ڵ6F�i ���"(��⟠j�O��O��O���&ۂ3~m�F�Q��K���� �ıJ�pE!6�-�S3J�����A!��ʴu9Q��!bU�3K�����ޟ,��̟�D�$�'���XǬޟ>���T;d� �3�'��7�+%�l�D�O؜o`�Ӽ�@`dux�	H[�:�����<A���?���f#(y�4���׾Y���y�O�
��Q�]�F�#�d�#��r�|�T�������ܟx������&�y��D���T<$��R0K�Hy����P���O@���O�����%����qDz2h���-A*`@�'�B�'�ɧ�O�Jxȕ�V#�N��5d	��pŨ�nR�O(����?i��9�d�<)��Qm�HasC%%ڨ9jւP��?I���?���?�'������A�V���r�˂�(*�Z�,6SK<�����럔��4��'1���?9.O�(�Ѫ͕PFH�Y��.'�Lt���(�X6'?9��ɋ6�f����䧰�k�E�*��w�R�"�yP���<���?����?����?y��'H�0�U�6�߫Kcje+�LϕWt�	����ܴak���Og���K�	����!��tp���BJ3$�^b�\�IKy2�HyB�Ɵ��!�J�.��.�<<���Bɒ���$�'���$���'<�'��'�"���OM
D�>d�4�P��ِ��'�]�\�4ua�uP-O�D�|j�h^�Z����fC~}ʀC��K~��>���?�M>�O��(�m��=]��*RS�g��%�P�ЛbK0AC�i;z��|⒉���%���jF�G���+v��_H$�r��������������b>��'��6M�	)�iiU� >���7-XL���+` �<!��i��O���'�R#��3:��w��l��1�e���K���'K�@���i��	�p,�M��O��'�^c��.-�P}SA��,Q����d�O���O��$�O�$�|PoL/^ ��j�d ��ֹ���&ٛK��U���'������'LP6=�J���E�$m�h���f
�50�Ӕ��O��b>a�ǦMצ��4��MH�pz����b�0�6�ϓ��K�'�OL�HI>Y/OP���O���)��&����b��jMd����Ot���O���<���iJ�	���'���'�rpCD�C�b�1".��&i�@����@}r�' �|��E�VǪq��\�d���EJ-����>�-��D��_�b���%���Z����(J},l �R)g0�����SE�L���Ot���Of�d%ڧ�?Iq@H3~s���Mô@H����?���'o���,Ozll�Ӽ#p���q�3�ф�����<Q��?���ڑ�4���F4I���P��'�\JR�ݟ Z�!�b��;ꖔ$)�ĳ<�'�?����?����?�bJ
~q*T9�/ �[$󦩝���d��ч�X��������'?��7�D�B�'��-8U��5.�>lJ�O�d�O��O1�"�ȃ����L�4,M�THKgꁕO�7�>?Y!혩W8��I�	@yC�.�4p���Bc�����G<Q(2�'(2�'��O���?�MC��Ԩ�?��j�<<Y�cU��=Y�dڅ���<�i��O�d�'���'4���)SejuE�Rx���t�*�ܵ���i��I	KZ���'�O�q���n�ڊ�Õ�������ȕ�,=��O����On��O���*���~(m��
�,$$mk�:�.������I��M��.�%������]&��
���#��pڴ�P�-T��1a�.�I؟`�'��TZ`�i����@M��6�V�C��5�����t�mbH�l�Iq��RyR�'�r�'}���QXp�3����<5� �c�]����'�剖�M�p ���?!���?�(��Y+'��H)>�IBf@/5�n��F��,��On�d�O��O�Yl<H5,B0�OҸs+V$���ӍQ�Z}n���4�B���'��'v���m�_+�a���S������'�r�'����O���M�G�ĕ}��:1H� l�&g�;9��Xy)O�Hl�p��j���������X��5�?[�U�p�X��h�	&oPj�n�l~Zw�XѸE�OQ�u�'�d�d�7	��岇*ē̮��'D�I�X�I�x�����Ia��	 � ��d�s<����M9Ԩ6mK�"��d�O��d3�9O��mz�e��*j�v�pC��\�J��៨��H�)�?Z��UlZ�<�3�W _nP�y�/�x����`�<�����	m�	Hy�O%b ��c(ʱ�+I�a�L���W�.L��'���'��	��MS���0�?Q���?aRLd�\l[w��h�x��h����'���?Y����| � ��N��n �D`�+���ĝ$�l��<pA����Xߟ(p��'�K�LRZ~������ �BY�`�'���'Wr�'=�>Q�	!aO8ɢnχ�D5��HQ�XM( �I��M� ��(��B�	�?ͻTr���[�>t���gA�$Ե̓�?����?	�/@�M��O�Y���F	���� ��1�/Af�p��D�|�K��;�$�<�'�?���?���?��)[>
a�m`��
~��xC�������Q� � [y��'�O;��+`���H��� ��Cg���Q���?����ŞM������V�VzJ��OW)*~I[C�P��M��O���$�L=�~|BV�@ۡ����<�f��"m1l���@O����柸��ݟ�Suy"�~�n�`���O^��/��T������Qy&!sc��O��l��n.��՟��	˟tR�EC��+..�D�T��OJ��m�G~�S)$�i����Ϳ��?c{�чe#%F	ȴ��<9���?)��?���?ɍ��J��:
d`a�L��j1��-���'�2.c�v5��2���kJ`�|B,v��2bT�
?�]
'�4Abҥ�<	���$��H3�6-=?)���(NmG%K�R@ts3����e@�B�O�dbO>I)O��$�O����O�#�*ޫX!�ł��ڣ(vJ�"�O���<IG�i!nP5�'���'�哆Qα����	(r
Y���;}�8�YW��۟h��k�)�2,��/��!�!N�xGH �uc�8/�����U��M{�[��+}��>��v� $:f�K�N�Ѩ���u�f���O��d�O"��)�<AG�i�������z��E���'b����>{[��>�M{��>���l�����9�<�����<�T��(O�H�p�pӚ�a��X��n�̀)OȄRE��?R�Lq�i�70���4O���?���?���?�������'S����煵t�̍;�`(�nZb���I��P�Ir����0X���T��$]�.�� �F$e1e#�K�.�?�����Ş.bx�M#�'K,���M�����S�:kP;�'ؔX���\?I>�/OF���O��Yt�!n+¤�i�x%JE�b��O����O���<!��i�����_�L������aR������Is.��?!WY���I��%��"��:6q,��#�in�E��2?I	L�2 @<;0�Vz�':J��W:�?17�ܘ�08��I׾	�x؊����?���?!��?�����ON��fbΏ�|���0���2��O|Ll��s���'��6�'�iޥke�ŔW}�m3Ԡ.@X1+�v�L��֟,��+zN��n�T~���VÈ��'-�(��BޞUĥ2s��<��J>+O���O����Ol���O�A��&�V��IQ):.�QRt�<��iA�q3��'�"�'��O��FR�\)̹vڬF�di�-�J�*��?I���)�e������]q�	��
�q*JqI��I�Nc�I�+vƕ8��'�:�$���'%�]�F�)HC�#S�/l'԰�P�'n��'E����4S�$ߴh�y0�#�NȘ叀�g��Q��Պ|��������}��'���'=�ʦ*��E
���̈́�RK K�X󛖗�\K�.��F�Q>��]������ύ*z�8`;�㎹`���ޟ,������h�In�'K���Hg�J��T��@ �����?���,p�f��9����' P7�+�$Q0G��������1�.�k`�[� �O.���O�i�@c�6�;?A�ٳ �Aۥ�=3@�IF,	f���r谟�$�T�'.2�'�b�'�����4z4�`ڋ.~t�2w�'N�S�ȰشXn�`*O�$�|*Q,�D��5 _�s�XY�W���3�O����O�O��8^U e� )�8Xni�!	W~b��U �/Ϊ䂕!9?�'_��dB���G�����MIpH�HCb[�!����?q��?��S�'��D���z��,^�ڠ�vȅ9a<(�	F�R/y+L���ʟ�)�4��'���?�$h+p@��c� >p����9�?��x����۴���P.�8�'���I�\ RǄ�n���C˙g��IcyR�'Bb�'���'��T>��/�]C@���(L2'i��c0'D<�M;�!M��?y��?�M~j��8��w�d�լ�������2MPr����'M��|���Ĝ�h��6O|v�(�L�ŜjdV��D6O���Ί��~��|U��Sɟ�
�\�&�`�ȡ�Q 	iGI������ڟ��I@y�&l�>�P�e�O�$�OH��1�E<r�<�f��;df�{��5�ɉ����O
��2�閦�5� oA�m!܌��=?a��؂T9,%�Ӆ�$��'S;&�$Τ�?��Dڸ1��ݹ����lR����O��?���?��?9����O:8��gJ�8��e��h߳u�Var0��O.�mڢ|��'��6�#�i�eYխ�Hr�p�ۉ~"�'%}���	��.S�rl�|~�FJ�E�'$�
	����%rֶ�¥�F��IJ>�*O���O��D�OP���O�bb�t�*̣��<L��m"�B�<��i�\�J�'�r�'��y'	�Uy���fdB�x#�(�=���?���ŞAL2�k!�_�n�1��c���K���N2�M�'&��F����|bV��� ��\5�M��I�I�����埌�Iǟ$�	͟�jyR�wӀ��ǫ�O����X4^ �%�'Q���V��O�Xo�J��e��I⟸�i�i84͋�o#����J��p��єs�oF~�c�D
Q�S
3;�OGG��9�$�/r�@�x�E��y��'���'s��'"��)�||=��^8?װ���H�H�t���O��$����3�K{>��	�M�H>�v�X�l��1m2o����+�	���?���|*��Ĳ�M��O��W� 4��MȬ_����ٙ6h,EB�?��?���<ͧ�?)���?�6X�&	�s��Z�����?�����V����埈�����O��!��ǌ4&����Ad~	�!E*?��V����\'��>�dEpd�6�P@r��� }H��ËS����s�4��4�pp��'��'%�LҬMX
<��&ύe����'�"�'\��Oq�I��M�CK�/B�Y�(>�L��f�K5ph�I����?!�i��O���'`��\�I�ȋ��D�JY��P��J�'��h�ԳiT�	��"� ��O.��ܱ�(ԧ[��Bw Ο��͓���7m�O����O����O��'c8��W\:7�L���(KFb�PD�i��B��'��'���y��c�����O��J6�[�vY���嚲X3���O��O1�n�6AvӚ��ԺT�GB�#�qG���ɥ~t|0r�'}�$�p���t�'i�#G�F��>�#�@) �[�'��'��U�`��48�Ha/Oz�$â����s�J�y�*��d97i<���O����O"�O���i
/q&�RӬ�o�,=R�D����K���{ 8擃K�� ���`�tL���`�J�(uɀ��%Uڟ�I����	��<D���'q�<�%J$(�X�!���S����'�6�G��ʓrR���4���e(�	  Y��F�f�b��s;O��d�Oh��W�-�6??�ѥQ�R����K~v��/G�=�J"z�Vm$�8�'��'r��'���'2��RH��Z�N츐�H�4q�,�U�d[شd������?I����O�$��琸u�D"��I�����>���?YJ>�|�EP)f>��b@iˮ,�r���F:[�&i!ݴiD�Ɍnpҙ�v�O�OD˓(u����Ug����	 TfZ�����?y��?i��|�-O��nZ;]�~H�	12�R"(&�0 {uc�"7 牊�Mˌ�K�>��?a��#���Z�
~��aU*M%���-��M{�O�`�������w|R��-����gmνc<)p�'Pr�'���'[��'��4��`�ܐ��iTh�W&2AP��O���OmZ6��h�'W�6�1�D�1�%��7��l��U�	�]#�y�'��I1/+�Lo�A~��9n���T�(^����6{�p�׬Fs�"�E��myb�'a��'�`N�b�8)�ۙ+lA�pB[.QS��'����M�J��?	��?1)��R�����RĂ�w�*3љ�xJ�O����O��O�P��geJ�4��ڤIE��E�K�[�8JcA&?ͧ9�@������F\�h���F�x$�� ��4;��?9��?��Ş��$���d[�tJ(�(��@h���"��&c ���'H7M.�	���D�Ob�����l�����F�|_�a'�Ox�Dݻ^a6-$?�,S7q�2��ry�,�l��D!Q)�f|��I�d��y�Y����ڟ$���X��ן,�O�&�P�h����&��I��<�r�gӚHim�O����O�?Q����E�;@I�����0���0��?����S�'[� m��4�yrD>B�Z��g`�����ڢ�y"�Չir���`��'j������I�R E���Q;`�Q�=������O|��Od�d�<���i@��'V��'�r�B!=&�J�d@�1_�(`��d�S}�'�|�F�.aAvʦ��e;N�Rӡ��*���Y�dN%	1�Аq����ȨLȱ���@�Ԇ�:A�щvj����O0�D�O$��-�'�?aB'�f�Z� ����l� �?Y0�i�b��R�'���d���k�ʹ�d�@0C���'G٢|	�㟄�Iџ �`�צm�'D��P�	_C��Y�ȵ���N�4K���K3����$�O����OJ���O|�H1�谘���?W��bR�ې� �9ӛFE��B�'x"���'�4�C��,�\�҇�$��\R��>���?M>�|� A��{r'D����6C�g�|���n�f~�m����I�MN�'��'ZnL@a֠�0��`	L*("4���ߟ��Iٟ��i>��')�6mC�!6�$Oe���ap��� zb%�n��ěܦ��?QRW�\�I���I/�.=x�+F=#_���@G�B��t.�ߦ=�'����t�M~����(M5(��,�&(��4�I�<����?����?����?1���,T&�l�q���
�6<�"Aƞ'��'U��f��c�d�<i6�i��';邱�UmH� N�Q�@�*��|"�'��OF=�ش��$G �L�!�ْ��]<�L��H0B��m�	/	<�'��i>���ԟ��ɰ97��[fF�F�4�)GK�9G�0�I�(�'� 6�� +O���?/�2q@���"XP��8��`��� �O��$�On�O�ӄ_�Q��:+���/Z�H��MP�`��mn���4��[�'�'�ܱc���>R�#3�;L9��R�'/��'�����O��=�M�u�լk� ��w%�;O�I����.��ɪ.O�!m�]�=O�I�����`XB��׮��X%"麵�I͟�@i�ͦ��'7=��?���n�zB���wv\[���'�A0w3Or��?����?���?�����	�"P��U��.K�� ���L�9�H�n����i�'o��d�'�T7=�D9���/��%xuŞ&]��8�L�O���<��I��h�7Mv�� >�%�۴u��u��ܟ_�n<B22O�M+����~b�|�_��ퟌ�I/����H)|�v�B&ʀƟ��Iߟ0�	cy�Gn�J�R�O�$�O^0��=$��T�ã�1M!
��O5�I����O���(t��,Z�+
R6RX��3?�W��\�h G۸��Z���8�?�g�[Bܪ7#�'U}�,�a��.�?1��?����?y��i�OB��Ab�
�Z�S0j�4���L�OzmZ�}�D]����Xٴ���y����")Q���G�j�qG�y�')��$"�]n�V~���wΤ������C!�%L۸�K��4YWX���|�U���I՟ ��ǟ�	�@�a��h�PF��K~4e��S`ybgӬ��O�$�O�����C83�`1HR�[/i�RY�SP�z���'\����:5��T���� u}�QWV�.Z4!�C^s�ʓX��h����Or�qH>�,OU��B	�uh�CA���JH��J7G�O&�d�O��d�O�<9d�'z|�q��R�lQ󶩚*��*���Sr��#���D�f}R�'f�'JZe�錃1$�Q�ҿ���&�֑���B�V\�D�����C3�N�K��,�F+�>O���O���O@���Or�?YXsA�
q����)z_83/XEy��'�7��.l����M[O>)F��%_�X(��&�L<Ô�ʔ���?���|�BE��M+�O��˧��
�H��d�Y�M�l��u핁=k����LF��O���|���?	��������	��
���A�>����?*O��n�  ����Iџ4�	b�$kKsӺ	��j�+�hl��ə��$U}��'2��|ʟހ�"�����w�5�}H���4b<2�Ñ|I�i>p$�'�%� �0�Ն<К��aJ(}7�,��-:���4J�T�0���9jsLiIm�Bք!6d����$���}�?)]��ɟd
 � A�ݴXc���dKG&Ϛ���ɟD�b��Ԧ�'&@aw�Y�.O$pDcI�{
05G%��Z�Mu4O���?9��?I���?1���i�n���v�J=����!Fn�mZ�R�l��'#���'�r6=�9����B��-@|�'��0<
���O��O1��lx�xӄ托������[6xu�6L��eL�Ɉߛ���O��;K>�.O�I�O�҃��g�\x�re��DW��ɠK�Ol���O6���<��i�|ܱ��'6��'A����Ӂ:�6�"�G.%;��x5��}}��'���|�ǥ �"���1�$�â+R�����1#F99�7m3�S�r1�$�O ��׮;Dr|@��:6��]���O����O
���O��}��<����%��Bd��h�cҢC$����x���/W?.�	;�M���w�j|�`�МY�􁈣L��Tq�Œ�'�R�'�b*&D�����Sa#�h��T����5��?k�J$k[.F-$������'d�'#��'Y\e�C�D�fŰE��kߤ`��T�$��4#�3���?����'�?��De}\��3�O�$�"���D��ǟ���q�)�ӯ?�F7�I�6��]���? �qFa����)O��ci�3�~��|bW��dLS	RҎ\��C	�j�:A���l���,�	ן�@yr$�H��PD�Oҕ @c8N-��׬����m�>O(�oZ]�@��I㟐�I��l�a ������	E�s��9���n�m~"#L�r�dD���w]��sf�;0��c*L�3�J�ȝ'f��'�R�'��'v��b�_`�\e���Vd\�a��O����O�%m��*l>�����޴��O�:��D��r��%J_^��<����O�f9R7�;?�tmE�R����4HU(_�|QꐬXh2�iE��O^��O>y-O���O��D�O���WE[�lhC5�KA�O����<���ix���2_�X����.�i��i���2����h���dWn}��'I��|ʟ�iթ��o[d���Xba���̑{�$ k3"��O���| L�Oz<9L>�&O�>:NA���R�8Ć��1l���?����?����?�|j+O6yo�;ڐQ��럲w|�Ȳ�DH���%Ty�k�n��ȪOl�DK�4D�<�5��)<D��#��Y\�˓)��L��4��dʣB�\���?�ʓ>���3�[�b�a��=X���ϓ��d�O���O����O4�$�|�FA�^���IT�%��C�,�6^L��ȃ2���'������'�7=�� ��D�C�a��L�% k���M�OJ�D;��)�/Ru�7�t��`(�L+
����%]���a�z����Щp�"I�N�Iiy��'�B+�f��yjN)9��"�GY���'��'��	 �MSՌޜ�?����?���_D	�&�
cچ�C���'O~��?����v�K��f�Z�9`b>[�|��'���!3���y0��zT���HП�z��'�rp��F�+��-�D�9� �s�'U��'���'��>%�	��c�eO� �(�sgX�m���I/�M����S����?�;9=j���;Av,�/�/��ϓ�?�,O�U�~���o��9�т��`@�$�(Tm�E��h��%}(xq(��䓦��O4���O��D�Od��ȑb^��O�(f����٫!�����Ƹ|��'
����'�n��#ʼ-�N�rR,m���s��>�������O���� ��#�ݖL�x�6��3]_��)��;,J�v�}	S�O�`O>+OR�"�[ ����抆g?�M��(�O����O.�$�O�i�<�b�i�S��'�8ـ7#Y��B��W�b�zh@�'�|7�:�ɏ���O*�D�Ov�Q��%jpt��`Ǉ�$�̩TF܉K�H6�!?�2�X��x��;��ߝ;q�е��AQ��6�|��h�X��ҟ0�Iϟ��	�����!�BO� ��{.y�����?���?�U�i�"�ZW�P��4��J\�e;f�E� N�c�S�Dܖ��L>a���?ͧ|���ݴ����b��m���,N�t�X0nY�
�d��Gl���~��|_����<���� �"9z��I���<B��v.W͟<�	Uy�$~�
)��j�O��$�O�'-�(�شIRu�I�ŰL=i�7?�#P�<���d&��'f��H��[�dMB�PEY8i�j�rf����ҝ�d�1��4�P�r��P�&�O(�)p��a,-cg��:�.����O����O����O1�l�lN�F�~�Z�s���.���f�ICL�����'Hbz�d�Ȼ�O��G��̪�'�@V�@��M��O�����Oyh��y�N�/�����e0�ӤG,�q��&y��L�K�k7d�`y"�'���'�"�'�B[>�p-V'ט�{1�Ljca�"l��MK��J3�?����?iN~��&^��w[�uK����h�(��=�L#��'��O1��X�u�w�t��o=�A'� "ʸ��շ)`�Iqd�0�'�\Y&��'�r�'Y�ٙ��3,S����M�a#J����'�r�'"BS�lZߴo��	���?	�KŎ剐���e�%�P.�0:�5���>����?�H>G+T5~q���C�*=@i�7b�R~�Rd1'gD>��Of!��<��e��^�
�Y�l_�jP���x��'���'y��s��0��=M��9p���nyLj"��̟���4'N�Ub���?a�i��O�Γ�0�z�ۦ
S�pw����N�@��O����O�T�P#bӂ�&�ܤ��J�?]˔����ؔ�P�|��4����u�	Qy�O�2�'��'���bq�@�@ 	
;����U��21O�	�MU	/�?I���?	H~Γ]�d]sG��>��1c
"~�My�\�������'�b>C���Qm�-��ᇩK�����M�h�u&4?�.ӛ?)���M(�����D&-��,�QR�IB��H)a|�w�,���b�Ot�T_(+<��w��4-�F�:O��n�F�z��	����	����ǀC��頰.�c����Q6 ��Hn�k~"ă�GhB=�'�䧾����i^�}��̐$e>J){����<���]X��S�\<|�ءgԫY@�9�-O����򦍃��1b��i��'mbؠ�́:Қ1�S�J����|R�'��O��US�i�	�v��+f.�Vx�P��&�-@��:�M<b���#��<��o�i"|��#�	�;�ܥ��ɉ�O��mګ9_���'�R[>�� /q�����M ~ ��Yw(.?�S�������&��k��@�K=z��h0��Sn�H����H�;�42.�i>5��OΒO&��dF��d�&�ǉ:��h��O�l�:K^����$^���)6>P�K���_yKoӺ㟔�O��D��=�"I�q�4<8�.F�.��d�OH����~�(�ӺKs&���j�.�<��,K�E��I3"d92��C��<I,O����P3Y�̽��������
���o��I�� �'R�i�˦�ݙQc.{@�'���暈MR���П\$�b>�2@���]ϓ(7�@�2��Vll$���.B�D�ϓ+�����&�O��jN>�-O�˓�h��G���z�%�Z�{��!��I�M�Â͍����O*��7Oބ$+\d�bK?��M122�I��D�O�/�䞵!�h\B�I���$�4m�	�5���ʍb&�&?ݠ��'h&��	g��Q�#
4)���@A�F�R�B�I�D}��G�=~d�5瑨i�VT�I�M#��Ì��㦱�?�;iF�	��ϙ�� 2MR�0��Γ�?i��?y�	ҩ�M��O��X�:���S0D$��'��6�8�
de�6/��@$���'��'(��'���'s���t�LeSp��8���V�dSܴG]��9���?a�����<y���$�ڌ	%�G�X�B����m��I��D�Iv�)�әCn�uz�������JC�	�8��X
u�Z��Yq�Q	J�O$�I>,O�!ysh��*���4
�/p����O��d�O���O�i�<! �i (�F�'�8	z�k�+��t)dM
�B�`��'%�7M9�I�����O����O����s��$yE��".���i�u�l7�>?�d��'���O�q�
�NBh4=83
�
J����M�a��d�O����O��$�O�d8�S)������$XM��J�KZ�o�<�Iџx�I��M��`������'����C�%W��3I��GMvʴ��H�ӟ��i>!x5I����'%6��6b�JR��Qw \�U�∸��t4ԙ�	u�'7�i>��IП��I"C�DIIŢxɈ�����5P�I�	ןH�'�7MU�U����Ol�$�|j�F�##<�	1#�%Y0�<��j~R��>����?J>�π �QR@т3��A�.�$=&2�t��.�+��!��i>
�'H.A$�(+q��cs��)0E5$(qBR��\��ڟ���՟b>��'�6��-�|iVkM,g!8D�W�fH����<��i��O!�'���c�`���� |< �B	�!S/r�'��I �i,�I5�~��1�O��}d���̀�b� IF�ǅc�a����O��D�O����O��ļ|�OƶO~��3m�	�^��B폪}ݛV�:_~b�'WB���'Ϧ7=�`b�-�>�Hő�`V.fT}"���Ob�4��	Z�\I<6m|��@��$�d��,�
}�*ܓ�Dp�D��MF��Ҭ�}�	Iy�ONM?l�X��G�sĔ�r#�$6�r�'���'*���M�⌑��?Y���?Gbѡb��-�!��@v�!1�����'���?�����[v䠰�M)6�v�stNB�B���'m��G�B����?�)�~b�'��]���ޜC}�@��ǹM��$�'r�'	r�'��>���{�$!C1����N�I�IPb�TY�I �Ms.���?��g�F�4�*�Ѣi��$���3V��-W��z?O����O����7�<?)�g�`����	n�B��:&��3戏-ƽ%���'n��'��'�'.Z�ITő�8�,����Mضib�P�t��4�l����?���䧇?	
�B��p,�2 ��9�+ٰ*�������IA�)�S�dE ��ۅ1�����E̞vѺ`�#�W즅�*O���ԥ�~b�|�P�,�V�L���M0��|�x2��֟P��̟h�����]yb�g������O����ѯ�ŉ&嗃W�À+�O.�n�t��A�����8��ܟD�¨�y"ĩ��	.MOz!�LY�q��Tm�^~�"eE� ���䧩��D�(�\�r�]=���D�<���?1���?���?a����O(zB*�(�)H���D{P�P����?��rU�֫�����'�6�<��N!p�<q�vB��]����)V�Or���O�X./ 6M.?�;]��5*��L��0�"��V$:͹gj�#�?�t�6�$�<���?	��?���
r:`����$��S���?+O��m�02�V���؟���`���(\\p8!U,�!�>�@��yr�'@,��?Y����S���\`\P�oX�;|�J�!TT�0��̆8[�}J�T��6�R)AA�IR2H-·��eD&B1>5����	$�)�SEyR q�D�S��P�VA:���H��[�� ��I͖M� ���O�eo�Y�	ǟ��OT�$�g�N�B�*��LMi����u�"���O$aUH`���Ӻ�⪘*�:���<9q� D��*��x	T1�eg�<I,O��d�Or���O����OB�')�Ĕ�d'J�H��-�F��2sߌ��i���BY���	T���������q��~q��pR�E�Xh�Xs� ���?����S�'r�ƥ[�4�yR�\>j���p.��
MIq蔀�y�f���y�������O���ǅ9nEaf�Ҡ#1�]۱gĚ`RF�D�O�d�Oz�_}��m�	���˟���ß,B��oΛs*�; �y�	ٟ��O����O̒O��!2w�F�ʑ�J�M(n4�e�����'K$*��Dn���CUh�����҂��w�h��W��F�<��d���D����D�	���F��w"P E�n4��"OO�w�P� �'L6톉Q����OYlZS���]�g�����KG�d|��M��q�6����Iǟ�:eȀ�u�uwH��p���a��#�n1"F-Ӭ@� ��e���4b0�'���'���'�b�'CR�'���X�/���j7F��bD���f[��Kߴ7�����?�����<a@��n�eQ�AѨ ��M�L����8�?�|�J\�0Yb�K� A(�� c�4"Y#*���"��X��F���O��C1j�Q�G�Aj�X5$� ��i����?1���?���|�+O��m�Hi�	���Y��iJ�O�K��:¢�E��M�I�M��)�>)���d|I�CTt��ݪVL��w�u���bӞ�%޲�K&e��d�PO~
��#��a�ՠɁ�@P�3�J�T{�h��?����?���?	���O�5r�\*.KxI� Ġ}������'�b�'A6-V���O��n�Q�]���W�\(XI2r
C9�2�%���IП�S�E�X�n�t~Zw�1#�S0Zz4q2���������2%GSu�TyB�'3��'G�J
�ej,�A�KXQ:Y��#��t���'�剜�M������?Q��?�)���@�K�`�]!��L�nV���㟟X��O^��O��O���mD���l��#���̇�iW���vE�c�E8��Nxy�O6���	0:��'k$k �[��k�1�m���'*��'�����O���ɂ�I
	�pt0�J��9�n��/K�r5+GƟ,����M��̻>i�S��(�c�)]�B�e׿{�b�3���?q�(�-�M�O�.�#_��)ֿ���_�q�Ω�bE�4Hd`�/U�~��<)��?q��?��?�,���(���0�n`�# ��Zi�gȹN��ϖZ3r�'�����'�6=�`�#JÌkh�s�/ZY�(p���Ot��6��i�N�r7Mj�p2U��4��Ta�I5g���1&b�Dӡ��W�2IPH�IPy�'�� T;~�"��%R�A������?����?�-O�Ll��"�m�I���I�L�(��-�/Mdu�"\�'���?)�T���	ʟ|'�� n)BEH��q�ɇ 	9j�t���㖩�b�Llj�(���\�����/0~�����
+��	 �B�HK蠫�O����0��W��R�*��l��hI��?�BI��G�dX�jUJ��*�$ �eШJ��i"��ɭX��QS6G�Ht^]
-�)��*�k>s_l�(fע^ͪ�bA�L�J���sWE��Bb~�Ӡ͆i�z�C��J�kk��A��5�807+ 3j��d�\;hP!΃}�*`�A�G3(eÁ�//���3"C[�� [C
�?��M��j�55��{�#	�+��Q��ٟ|�>	�@^�	 ��2l�����n�n!�(/N���`0�Ȁ�J<z͛��' {��>�/O
��;���J�j��vs*P�rj��a�8"�\�����V�Iߟ|��Ɵ�'�\���e�D�$�#�/*/�A�dLض)�0�����O`�O\���O�`��ۼ0�H�3�,N�XbL��n�*#鰓Oh�d�O����<akۻ-��)\�bZ�	1��SMb$�Ì�u�\�l��P���h�	�zCb��"��cօ��Q9lH�eO�^�8��'��'/�Q���W����)�O��k���O�81zg�(,x1����}��o�I�x�	"%�V,�=	��U
4�Xѡqj�M�T�;��̦�����h�'袜�`D�~����?�'G)|Zr�W|ˆ�K���E�L��x��'�Ҧ
UBҘ|�ӟ�ȱ6dL1m�JD��	�e�ܠ	"�i��Ɇjb|hߴ�?����?���k��i��r�k�a6j\҃��4#Q)�Teu�v���Oұ� �OF�OV�>-豌� ��BE��`���Ƀ�s��<����ئA�������?� �OV�}lLȂR�U3HrNyѵ�C�;�>�jC�i��	Y��'��'S��@�Ax�@��[�\0����>�`m͟���˟�9��Ǯ��d�<i��~"�%*��=��&X(�x��G/��'���c��|�'���'��<�P(�,7(|b&�';���p�/n���ǝ\�4��'����$�֘�~��cg�ݝy��i�pC�Q��W�lA�L>q���?q�����{�áH��
�|�u�[8"y��x�'Uq}�U�h��b�I��l�Itx����'��<޲�n�{��yW)�۟ȗ'���'J2_��c ���)E9C����$[53.��T���M/O��,�d�O�����h�I".k�\T�é/Y�d�RD�
M�듚?	���?a*O�	�%VT���'j���5�X�o�X����+s�Z�Ga�D��2���OF��^+�|�@�to��1�e��(�,p��p@3Mz�H�$�O˓5��|� Z?5�I埌�ӵQ�4��Ċ;H����5 Ɛ~� �N<���?� ���'��)�y���0�e\(]���qtѦӛ6_� ;ǈ��MK7]?��	�?]:�Ov�+��-,����֐6���ґ�i��	��Ʌ��'���i��.4`�� H�6 
��B�wӖ�s���̦Y��`���?�I<ͧ�X��TGC��&0��G!mm ,@�i���'���|ʟ�$�O��A��Q�Oڸ11A�&���8CH˦U�I��H��?13
�{I<ͧ�?��'K0��a[���G��*��!A޴�?�H>1�\?����Iޟ4Óo�ِ�ք`�	���L��M���*I:��'�x�O��|Zw�����	���@;�K����M<�����$�Or���O�˓		BU*`ե��# M?@{�� ����'�B�'�'��i�yQ��.�`��O�#%Z���|�����<����?����DD��r��'&�� �$4c�2As�oM��`��'���'h�'��i>q��	MΩ0B�-Q�b��RI�R��Ol�D�O����<a��kP�O(�̱�%�'dD(���	(x/"��g�8��,�ĵ<ͧ�?H?űFHJ���ŽJ�U�f�0��O�ʓabJ\c���'��\cTi�Ƈ�.�zYӀ��n�&mZI<�.O0���O �����Ԏt*�Ɍ*U��A��i`�	�d2V�1�4���ǟP�����$�%�>-!�a�IqZԃ`�ܷ�?Q*O ���O��� �����-�i"Aƾ2m���d(P��M��`W��?�������\�S��AK3W���e��4���D�E�W�����]Fx����'�R�E�� ZF	�}�z\`w�dӀ��O
��֛!�>�$�����p������@h��n��u�ԧ�yo��m����%��q���I��@�tg0(�S���"QQ%��1F�xm�ş09��dybǫ~j��A�*���o�=	�9[�ȿwdO�݈A�$�O���?�V�='n�� K��sJ�p��_�	z���+O��d�O�⟈��T?�3��*���
�G��m�b
6@��$  1O���<q��(v��h�O��Dk�)�
x�A�G�,�#ش�?�����'3bP�P�W�s�VA�̈́ACd�*��7ni�_��	矴�	sy�/�TM��f�8��0�=�3��D<baI�U�	c�Ry�O��~Zra��S���KѨ	wz�q0ߦ���@y��'XVH� \>A�	�@�s�1A!o]��}#ƣ\�8kʠB�*1��O�ʓD�ExZwpN}cq���x�ٓF��0��i��O���W�6!����O����Ol�ɼ<�;x�� ĝ>$B�%���A�OT �m�ן��'�\�Y�����>�Yص�Е`v��@�<�M�%˵T����'��'��d7�4��9��>8o�1��	r �<���l���O^�d�O��O�3?�/	�f8~���-�|@�i9�ǭt����O��$E�r��S���>� �lz�)n�A`�3�൘vY�',P�\���O����(�85#�#(<�V�¥�~���o��$��B֐���|J���N͖@��h\��+X�z�z��x��' �'��\����oJ	C��>n,�K��	�_0�	9d��Py��'22�d�O�	6$"�9���I3L94E�f�Y*f"�6���x.��ş�	��'n8�k�n>��3M_� W�A�ܦ!��4�>����?�M>�*O���O��sF�
�дPC��Z�<�]���F���̖'V"aP�<���@��b0B�{uEB?b��j�nǳ�M+���'$剀m�Of|�d->*xV�Ҧ�Q3��|�0�i�r�'��I�|��٩����d�O��ɑ�mlJ���G����s�JxD�'C��'1B����I�<��O(vĳs*ȶ&	� ��łK@���4��$�>)�QnZş�����D������ ��I��+���j񥖱HǼi�b�'��*�'�\���}��	V�P��F֛?۸�kKզEb�J��M;��?�����BQ�p�'L@��a�wB2D�&�M>Q��B"�i��e�8O
���<�����'7��ztH�u,i���."_�x��f�d���O����W.���',����|K*t;U�M�;q�,�@���[D@�>IBK��?����?��C�E�
���CŚ\��	b'�/���'z��Rd�>�)O6�D�<���[vL�[Ad���R�`p���Md}�Z�y��'n�'w�Z>牢G{����k H��� q	CKb��y%�K���Ĥ<������O����O�в�˹F��Q���W�$e32U��O�d�O`�d�O��s !��<���o�"	�PC+
�~b�j�:�MK/O���<A���?a��R�uΓu�5�E�
7�8�F�H�Ƀ�i�R�'���'q�	�nÞ�@����$�K��Œ6E�a���;�섬x�rLo��ĕ'&��'��hɽ�yR>7m ���U��oK��xsb�Y*2՛�''�Q�����F4��	�O����Rdq�	�Nk����:V�>�*�(�m}��'T��'HvC�'�s��'q����Cl�'#f|��a
��̦�'���:�f{�"�d�Od���,aקu��A#)d@"&G��X�$����Mc��?�w�PT~�X�|�}��(�Z���P
A5v��1]�AThˉ�M����?I���R��'Ф3��Y�!qDM�5�b�:���r�8=�'0O���<���d�'�� ��؉HS.�k4Ilu*���p�:�d�O$��ӟc��'S�	����Idpp� 	�N9����S�5.\m��� �'��x������O��d�?�w�Q�@���EDݕ_�j!�ǫcӌ�Z��x��'��I쟼�'�ZcN ��� ?�uB���MѤdi�OЁ��=O�d�Or���O��<Ad獷\6���Pl��XC�ړA��}RS�D�'�"U�@�I����	 �\��D� Y�a�q��62���h2�+?���?��?	(O�8�B��|
��҇S��d�%䂃$B����I�y�'vR]�|��ݟ���\9��ɥxT��Ә,p8᷉ X�|A �4�?��?q����D��L��OZc��\��I0%��� �H[�Q� �4�?�.O`��O��ğ  ���@?�0E>��L� ���C��}6�F�'P�(��H0��)�O��D��p�k�fN0*����P�;h��dTL}��'�R�'�ȹ�']2X���'o��H���D����AW(j)oTy�F�w6��O����O��QB}ZwF��;(�;i���$g	}��h�4�?y�f������S埨�}��#�
.N50�Vr�i���Ц!����M���?q����P�h�'0$j�NJ3Rf��ys���&�+q�g�B�5����'��|����F��$CfL�<.fV �݋yb(lʟH��ʟ(��A���D�<!��~r�Z�	�P0ʯy��2�Q1�Mc����ߨH��?������:�#�<�<�%�&n9m����*��d�<�����D�OklO<X�x-;�)��R �k�D>�	ps���,�I⟈�	i��'8J11�Q�,+���NX�L�y㢪F�����d�Op��?i��?	��ƉjC�"d�M0&��2L�:7 ��͓�?q��?i��?1,O������|�w��C�����%.�F��DǦ��'�[������<�������f��!�f�6�Q 4%�Sʲm+ݴ�?y��?����ē!H���O�Zc*�a�\�qRi[�t�P��ٴ�?Q+O��D�O<�D�2��O���"�E��UX��	��$�G�i��'��IgJ ph���d�OZ���{��U���F��a[��B���'d�'��J�y�V>��I|�de�qm���Th6f���3�T��'bdP��u���D�O��D��֧uG˞�>D=�UmZ2U����(�M��?9���<�X?�r�'~rd1�!�g <�4@�X�n� 3&04��4�?A���?Y��z�	@y���<x�~�BE+�R�B�ʓ�U8�6�l��'}�Z���
��~?���w���y���g�R3`
�ٻǿi���'����{����$�O8���)`} ^Y�Ѩ�i�nqHMڴ��&��S��'Q��'`���c#܎�ʶ'�k��B6�d�v���|�i%���I��H&���E�k.�1��Or�!q�H��D��`Y�<A��?����+D�� _�O�b@����J��۫7��'��'~�'��'2V� 8���ז�ٶ&ܚk�t`���C�?!)O��$�Ob����s�R�|rbD	�tE���?n��!pq����%�������sd�\ڟ�(��^�C�4Ad�\�Wr5�����O����O�ʓ6�D������%C���D�N�/rޘA`G0XM�6m�O��O��D�O�ɒ�i�O��'M@�Aï�h+�Xs��%P,5)ڴ�?	����M�!�%>�	�?�m��B�@��Ԥ�-��`qԭ�/9H�'��'8���C�'��'s�郮 !�1�Ȕ����p��[�_*�T��X&a(�M�R?u���?a��O���'  ��@ *�!~����i���'�����'�'�q��� ���+I��3(ig>@PV�i�Fdq�cӚ�d�O������q$�,�	�-CB�*�FU,^���j�ɐ�2��	[�4e`�T���S�O�r�9�(aA3H�z����d��
#d�7-�O��O��s�y��?i�'��]*�mV&v�D�ag�-V��ߦQ&��Q�n��'�?1���?�T��q��}"���1n�@!���t<�f�'d�H3F"�d�O
��&���p�0�CZ� >�c�f��L���S�Y�.S۟|�'`B�'(�Y�X���v<�D�8*f��F �<(�z�}"�'��'{2�'vvD�!�ݯ},����)G%4f��c0n��y�R��������Jybe�����>�] �8zR�`
u�&|:xOf��*�D�Od���R��d��:8b��DnS��T��E��vhd��'���'o2[���$8��'X�``3���eHs�B8�|�i"�|"�' ���x�b�>� �&G�q�T�� +rI��
�ئe��៼�'fL�K�3�i�Ol�	�&e"�łv�)x������x�d�&���Iş�e����|&����e����
#'SD�I�ϓU��tnQyB� 0��6-Kg�D�'��4�)}R�� �	A ����[�7��O"����%Q�+�$ rj��̫m]ʙ;����H�~6M��!C��mğ�����������'j��u�̢~b�I����je>��fӾ��)�Or�Ol�?��I�3lx�P��-<-�hq�!_����޴�?��O�	�'Fb[�0�	x?�AT�@9@`bt䑫)�(�����C��h+I|���?��Q)"��ǘ�ȼ�v�ڬ~|z8P�i��CR=7'O���Oh��?}⋛�G��m�%��!;�P�Z0����$[�0i1O&���O:���O^�Dƀr�XD`��u����4	Ԇ ����0��O����OJ���O\�OH�İ�@jҋYm�m���.V�|�uӄ,�Ԕ�X��̟h�	[y�Bn�V�ӪL��)�"7DEb�*L[NlO��$7���O����|����rq�处1!tNʛB�r��?����?)/OltJp��b��\^D�YԅV"H�d���7��ɓ޴�?�L>���?a��y�c��*ԡ_%#�B�Q@�7z@o���	Hyr#p2x���埔�ʑ�N�H�uM�oATUXU�Aq�Iڟ���;}g�"<q�O������+�ƀ"0B/�P��4��/4��tl����i�O �ɖG~2�V:�������w�dx�p� �M���?���O���O>h�2��h ��l:$�Pݴ\���q�i��' �O�hb� 0D���5��B���ܓ����Mk�`�'���$_L�dL:�n��MY�T � F�knqn˟��۟�h�G͓�ē�?I���~ҮU�~��ӑ�ˠ0�<������'D*��y2�'\B�'��Z�k
�N9�����J.H��AY�o�~�$�=��\%���	П\%���(儍y��X2 �P���/���o?�h�<)��?���򤓞p���mm��	_6Y���@I2SN�\�	����J�I���I6LrH8�E�<o�A�!fS+'���!U�)�	������Iğ4�EH\�%&N?\�,��L�4iJ�Ibf�����	џ��Im�Iџ�'� 8�ܴ&½R3H� ]���"GΘ�4��'��'�R]�����؂��I�Oڽ�`�2�*@+C!T�$�X��Ӧ���͟d�?���	�)=��82/�"JhD82b�A�bW�F�'^R�'G�j[(Sxb�'�"4O��f�Vֶp�rK�{v@��+�<nd�O���<IAj�j��u7�&/~����F� ����܋���O<pqE�Od�d�O@����P�Ӻ[B���|m�EɦA�C�B(��c�ݦ�Iy�V�O�OAn��" 8l\@�H�	�b}��4H��$+1�iR�'���O݀O<�$Y� �(���Ӄߴ��E
O�qRQ��I��Pa%
_R�2DdїW���:A�7-�Ot���OF�5��z��?��'@�:�f^�<!ܼ��kp�D����?	���?!u�Ҩu�`pU�D�Q�ƨ����iƛ��'�z�A�e=���O��)��ư���K��.��� ,$Z U[�m�1O���O��$�<IF�V3���T���^�6�H�b�l�h��x��'�r�|��'��� oY&5C���\����H^�t�<��y��'�r�'��'��pJ7ߟ�Uc���dgDt(Ã-T��೺i���'��|��'�� *T6�ڔ#�f�q�X-.2��#�C��@��	������� �'�(\�E+&��&a��X�o�;����lI��"�o��`��T��E����~� �u(�M�!%��8��Tdk.� �i���']��'����p\>a���<�S5o��鹲�*WRm� �P*6��HqM<����*R��֝�]��W���7�ʠK'�K�i�7��<�m:a^��L�~"���ѕ�̲��Y+�	���Ś/���r��i���$�O���Iw�'C�������Q#��C�tg*m�xj�4�?���?��'3��O>�zb+�,C��,��eK1Y��8y5�Φ��-=���O�n�#&M�k0��P>Z}3"ݛ&�@6-�O�dg�����<,���丟��g�7Ll�������0�ʕ�O��&>M�����ɥ#s m{Ѡŏ;2ҡd&	����4�?9!b:H����t�'�R�>�@�O�Qv���4W�LȐ�XP}�����'<��'aB�'�ҡ�7�x	�M
Y)2�ۅ�*f�zY�������	`������?��%C@!�1���P"��H�%oZ���?����?+O����Ą�|��i�<T$!� j:_]�\
�c�q}�'���|�'��Y���$N�/c�7�.o�JD�&g�%\�	�(�I���'���eC6���B4�MH�.H��05�S&���n�H%���I��a�1�	�Z���Z� 9���� �� 6��OZ���<��-$ȉO���O����&�?�
\��i��uu�yР?���O����=���<�P:�.	9Ֆp��疑�Pm�Ty2��/?K�6�U���'k�4�(?�$Ɔ&c�Pm��� KGBY��B ݦ��I�c��.�S�'zO�ҁ��%/�0Yw 
'n��m��qR Y�4�?���?1�'X��O��Jw.��ef��b�L�pֶ����Φ�qi(���O�b��L�&�	T��p��Z�P�Ib6��O����O�p%)�L��ǟ��I~?���R ���2�7n����!H	E�&6�<����?���KQҠY�N.W�r%��l�# "0-q�i�bk�<�OT���O&�Ok,R&34�`Ƌ�^��!��.��	6Rֈb�0��,�IayBcc����:Tl���s�1*]�M9��8��Ox��=���Oz��?n���W�ʂ����֮E�NN�:%���O���O�ʓn��yx�;�&A��o�~�*u�@I�UY�h�iZ�	����'[��'��N1����g������."�\�Td�=#�������	��'S���Ŋ�~z��g�
�B�����(��'���B�iI�P����ן �ɬg�v�IΟp�J�;����c�Z�S&�����lȟ��	Ky2Κ�%���'�?�������Ŋ5�Q@���C/���5��886�������l�g�+",O��Si��V	�9:\�q�Ł� ���ٴ��V*�	mZ��P�I��������9$� `���XW�ճ;><}ɓ�i��'�6�h�'zBX���}�0�^ �1�h�L��)�FnC��M����?���J%W��'�h�vc�6fH�$���4?g, �Ёw�ji�C<O����O��&��ɟx�',�!d=�-Q�m��`j�U��̅��MK��?���"�(���\�,�'$��O~|���-*�t��jߥJ��z��i?BR��+GBv���?1���?�	��c:��;�nO�X�n` �K[��V<O�j1�'�Rb�~2����c:FAA��دGQ�����xݶ�`3�x�������O4�D�O��H���d2�m�2��$zb���)]�'b�'�����"x\�b owL`so� E^V�2�D�O|��Od��O&8��%�?�"qo�*L%hA�\�dV�he��˓�?1J>!�����&ۛ���[��e�&��vyuӝ��$�O����O�ʓ�V�Д���Ö���V�R>Z�r��>0��6�OʓOH�$�OH,������I��[�'X4��R�<7���'��T� y�"����'�?��'�F�8$"5-ON�Q�	�!u,�r�x"�'B"�փ�O���z*�5���[Rzt��Nm�7m�<�I����V��~R���Ƙ��U4jh��/CP��YP��iӶ�$�O�ʐ�)��=L�Q8ţi�"\8�ϙNLf6��/���l������ӟ����ē�?)��N�O�������j���SH��C��OQ>�Y��\<*˪���MM����vL]%%�p��I*h�sT,��Х�vꐹ94:��INz"����%j��0���G�3�����@�*aTf�l�$�b� b�vDS�+v���`F�@�'�FP�f�E�9�a��.���A�AH�K8A�ǉٸ*!ڀ;A����<�@+d��]S!���,?j&��`
7Zζ�[p��u4�i$�)~K�|c�WvN���'R�'�b�^�k Z�M+�O�m{�i�=7�� �!
/kkXL	BL��=���.�"�U��	�("?Y�ko��P+�"#�|0���$>	´b��n�Z!O�Ql(2���{Gޢ<�G��ß\���:I����Sfz4��gP�b&4�D{�	p$�M��i�=;[.	���Mj�C��V>�S'$���
	Pr�M#$Ȧ�	���d�<�B�����̟��O��Ņ��`;0p��*рk*&J��_M��'����Z�j�6B��DN���G��O�Ӽ���2SI�:Ubp��І�dTr�<����&8�TPK��e�q�K|��G�R~�0��e�D��f�'�i����?Q��� �\��^�c��E8U�_�'BBs�;O���D
�>I
qj�&O.2�>y��(ìa|&<�dK�u�<-���&0�������[���"J�h�'�2P>�aiT����Ο ��׮p4�Xhb�
qK�����Şd�i��g��oM��d��O��E��\��ĵI��1B�.)#��#Bj�*D���۫ h��6�	���'���k�N��n�Hͩ���(K��##��V�r�'K�)�I/�Ċ?&��p�f�{�*����X�Y|!�$�	C���ӱ��;�>0��(ߟ*w� ���?��@�"nz��	@G�I$L�`���ퟸ��-����0�ʟ�����|������O�E�����d(�� @4�m��:O���ʫ�p>��Q<���ŭ��04�=:�H�~
���g�3m�>�s ��	=d$�g�'d�]!&�2F��0E'����V�'�%c��'m����,O���<)�1.��dh2*�\��I�DZh�<Q��p����F�V���!�Z�
ϛV�':ɧ�))�ɳ7���`AꈜÔ��g	�5
wdC䉩�Vi��HܯS�(��@�$.�B�Iy���A􉈧d�T�x�*�g�B�I"OƜ�� %Cj���M =��B�I�K ��aN�,a��-�&2�B�	=�|�p�HȏZS"��Ǜ�q��B䉦>Yi��%S7��+���B��B�IRFX�!U��ծlA�*�!D�JB�	<a�~��e�^�i�������)�DB�	����rΟ��V����4S�"B�	+!��IRT�¬M*�`R�=��C�	!``��'Ճ[�i#��#|ϨC�	�y���򄀠$��ɨ�I�Z�C�I�v�fe9 �/�z��ׯ̈Z��B�I��d��1�!/b���h	4a�C�I�=)v=H�cB���G2g��B�I�%(��P�@���3E�kԐB�	��t�ᡏ6t�4�`��=$tB��\*�lUm��5b@��:�B�	
z���Q�Z=Qa��%M3JB䉳LqTE��}��S���1'�C�8y&��j���p�1�c�V;h(B��P�j�Nh�.���l�4��C�2{������HyN=%��C�' �ѓw�@�g�v��T�4%�C�IZ���uGӾp/�8�g]��\B�I�8� �NC�v��i�� $NB��h��M��݀H�8<H'nÊ/�B�I�Qp��b&���,�4��	A�rwB�I�+�j-#�IV�o�Ę �  6#L�C��
]��$�D����b�1i��C�	 	MB%�0�X�/Qz���Z'�lC䉨f�%X"��g ^�����\2�C�I1�D�Ơ¢0sdJ����X�C䉥3��Ҫ�&j���W��3Fy�C�Ʉj���H���� �<PCJB�	&|�����O)6�ֹ"%�ڬ	�(B�I%P��	k���X�j�1�f�+at�C�	�a�@����
����"rfC�I�
rh�C�ך?�"��Ji�B�	"H}4��O��A�Вԓe~�O��҆�Q�S�'��(����-^��e���"(L��ȓ[�~(��W.�^06��]J�]���,!�>�?�'�E*7�M�I�����O 5�2h:�'��C�C/c	ꁠ&�54ԲHP?`24І�	�8w��`(O���2+@�'J�Ƣ�2����t�'B��F�[�k<�0�	�8<h�Q��$���T��;ޑ?��FӋi��qX�*�"�>���I:�$� �.��{���D�i�p1*�	sS�iItn�YY\t;�����RLJ��M�M~�=���ԗ;�8ͩp�7pTm0@��I�qO&8`@H/�s����U�? ����o���q�f�i�$D!b'nӎ �`�^RX�<��aV	Y��P�sAǊIߘA�7�ϙ+v��E�OFl�F\��SNt>��l�����:��6�̍r�P�X����#4@��ɏv�@��x�B�z輛�C
J��ԣ(�~���:PppЂ����P�?��R�J�(�����yț�<H0���,v��Ohpt��.򸧘OC��)��D Et��	r|,��0O\$���A%)��AaG�*)	��is֟�O��9��,����'�(kH,��%%�X� l��*�z�[�e����#�"�a��@n 8����<����!.C?��Jd���=�e��N����߰i��ِ0%�^R�-Q�寧l�%χF?�'r=H�[�'[20��O2B��HS�ZsH����*}=�ϓ^{X� �3�DVs\���rR��pl�e����ppܰ��GD?�U�]F�ӳY8���'`�h�DcǨH\��q��I���'�20�O4ӧ�d��6횴*�R��L�{.B5���l�h�2.tӈ����D�B�V��qm�w��}beV:Y�I	��A�t�Ф��R���p����<Ic�@���'�^Pz��A�^�\�%�!6�T ��#��u( \O�L;��H-1n�d�%ǞE��#&-c��O��c�-�^��I�E:lRa@Y��<�����?�0I�C�O��d.�.AR�.$TR£���OU�=B�����̋F5�a	RfO9�T�Q	١��$I�9���|Z7a��=�.�0��ϻ0}�,#�H��<�c�d܆.>特*�ţ1�\}
�B3zy��O�B��'kԅ��MF9��؃D	�+(X�J��pcĥ�� ܙe�(l�%e�.i`l������y�F�dsd�H�o��QS��s1F�3��O��с哪%R��1��&�*��� A=�c���@QM�S��v�B�C͈d�����" 0�^�'f�EFxZ�M�c�|¢,O�0��c	�� �Bس��ѥJ�*��?���>���ƓwEb�97��8W0�i�b�`��:�MS�	.=�Z��'-�yY��� 7�9��B�t�
`��ʝ��<t��3A�,5K#��>-ܢ<�S�-~�Щ�W5Va䋂51���P�Dܔp� ��%�Oj����7�&��@�n쳴 ��2l"D��	V�*]	c����(Ex�a�(��<�@�%[���FF�,]�F	�B�$�4]��'J���F
5�  ��iQ��BN��u' �*!ǐ8$E@4x*�q�.ݺ$�����cy2�ȸ�O�iをO�L�I�0�ܴ@C�C�3���U�Ą!��a	Q�E4�:u;gb�|��M�A�pܵB�OK���vhRt�*B�w��'�H�Ƚ%�,Z�4J��'�ز`M�0"�!��T���S
ǬLz�
7c��H�8�z�Qߜ,�	1 -������G0�O��HF�L�C����1�A/CXp���α?�O��P�ڽ#�� �p`C�f<�c� �:�+��?-@��s*w��B�2S��/T��q8�?�� G�4+��$�G�]�3��=�QH�"S3R�Q�?�^t;E��#8�,37'�h��M�s�VeL�u�x�J��[h������-ZʓkU�}Fx����0��l���	�;s"��Щ1ܨ���Ƕ_���)O��q��
���q�޼H+�pb^<W���0\��[��ĶL���B�'CՄ�O��ڒ�i����<;�V���Y�RI��'�f��.���hP�[�N�<ZF�V�1��x���_а����%�n���ɏZ�B�Q���
t��("�nqCGCu�X�B��Ѫb�|X����p�4u�'�����!�c��� �š��
 j�٫")��mҼ���@<��8��C>�'#��2y�*��8M����[(cĀ%�$8%��g��$g���2���T�5��؛0�O�[���VQ��R�o#�S��톎E"�T�ƯC�)[6!xb���
�<8�&͍=_��D{�jڶ��ig��ONƠKwk�7�~��P������+���#�'9�����#�/�tId���h ؽ���I��$��k{�X�eoN�S�8��Y�#��v�;��H��9�'���(OrX�2O:6�pD�N�~I�葆A�DwԡaG W�=��5�l�>)��Hp�'�^! jP�(mr��`c��1�HQ��"b!��IQP��gߘ_Utq�����E�	5|O��j4jީ#%lNP`Ą
x.���֦&�OT�qUl^�v�T�������2L�2�+v^�v�ўX`�Oեt� ��C�Lf�܀���V7V.�,ۇ*�)W:XA����O�A�(*$\-[�E.t��T�'�"P���W��I2�#	8I�l��Cb����8����9@F�8 �7��O�}�6�D�J�B%;�ل 7�x0��(�X��&D�S�L
v둩GC2�T�
i��,ЧW�ʴP�cF�\m���E-AL|x�'���h@o�m����)��Zrp�KA����?��� ���Oj���&u��XЅ��3ݔ�A	N/.�
T�P�6�Ozp�ѨS�>~-�F�T&`����&Ϻb��Q�ƎQ�'���U�'�Ld �̞��)�O�v���s*RIc�%\�w��â��vFxr�oD����[�Lo8y˃M&�?�'7�A#��7�2]
��Y�N�	"�N�s�%ÅP���BE� F���>� �h���93�@��Z�4�Y �}��7k4Qx�BBøe����'}\I+ÃS
�!�m�3q�j��Gą�r�84��1�T�!���A� ��,5(�C8��(Ԉ4ȸ����2l�)ϻJN0�h�MİP��q�I�16̑���
�0���CA�X�Q�ǨK9��Lja�=?�C�I���=�DꎚK�:� ����e�������]8�{2A�t~e#'�ߛB>5A�h��yrFC!�v(��_�h0�IqSM������:Q`���{�����xiW��t�`a�È��!�!��6KX<�W���R;'/�:�1OR9#'�7�p<9�R!e������ը"=����B�e<9�B�v*�pY�&�3;��}bȍ;K*�i�*>���w��~t�LЉ!,�u��e,Oh��ՍPܓ0����m7r����)�~f<��
��ѻ� 3��d!7 �;�l��O`��F�)��d��(y2AM4ɸ�igN (4݀�����#�d�	��ڜ+�ЕC�Q��/n�؆�	D_]@���,x0�	$P4��W�ƹG|�1�'�TZC�	o�"�m��.��"L�KS�' �}j��D���(��(�\Xx!�
m؉q�(�"�B�� 1����2��81�ց���
y�,RS�>}�/	���}&����J��t� *WG&jd�#�0$���#��A�4iy"���V�*<���B�D2b�ZDL���0?YGˋ`5
0�kɨg�0ga�<� C�VI��S1d��14f)���`�<)�"YJN�ۧ��G`%c⮘t�<97�V<;4@q��D ?ۤ|B��@u�<�A#�'}�̘�N�!l�<�G
r�<���YtН۠/�'/��k�	m�<1-�/J��U��*�8r���"�S�<ɲO�; $	[�2,>�����MS�<i6��T�Y��f	�!c�I�*�F���^K�,�>�J��P,�e��$.�V�����z�<I��%l����ˠ^�q�k��B��v�'a���C�W�T;��� �'�vЁG��j���CM�ӌ�EI�*|zC�	 WS����*H�tR���
�,�`�񤛨$U&��=�ƥU�~�\�� B
v�. g�r�<1Qe�f]#Qk4�=I�	Fh��� `"��>��`H�E�
�bA�ڼ(<L��/�M�<�$h�)�f�:��Pi���Uܓp}��@�'���`Ƿ�ABJ<Y��CJ[(<���\0�&��FE,?��:�2)���A�
O�$���Mb�XM��EǶ4��'$$Y�Ec$�)��!���G�gjj)�����~&B�Ɇ��M;��8����)�, _�O�0�KRd�S�'f��2�.7:��x� F����d�
A�B̓rk�)�'�.�����C�8t�NH������ka$Y�ȓG��P�˛h�=Bq��5{R0=��y�peA���k�Hz�L�������}c�H_�i�,=���S�n(��+X�,s�#D�L�v K�j����NeQA�X����$qŸ��w����r��:i4�4Z���w��5��	%Y����d����VC�Z�R �ȓm��J&�ZT��ҷ��#a%0�ȓ><&�����D%�&,�D�l��ȓ0�
���R�0՘���O(D��v$F���EF�'���#�ƖI{���A�D�q�)Ȃ2{�i[łG�P}��n�BӃA!5
��!�U�J6�ȓc�����mE�|J󅕒	c�ɆȓB��	2��U8н8s��$;I�5��S�?  D1F�Y�\8�Sb�5��ظ�"O��r��Ȳ5.[���!t��˶"ON�Rv���#���s�B'nъpK "O4��s�K$~:���5(ұ^�^�t"OtЀ�V�X*d��&ʀU�rK�"O&�Z�l՚�B�Q���Kx�T�U"OܝB� �>X��E�I7Cab���"OF�I0f|j�+��&4M|9�3"O�%tD�E)�!A6$��N�µ`�"O.y[��ܧ|�8��q�=+����"O�4� �$_LbUz�J
>b(qq�"O�}��
(`x���鎱7����"O|ŀWc�9+^�kA+D)�l��w"Ox�cPn�8>ܸD�+6<���c"O"yp5>�๨�HH6H��� "O��!ҡ��yz�m�g9�Ars"O�<����Rp�!'đ*)@��"OvQT,O2E_�i���<���"O	I/��<��lb����a~���"O�Ԡ�N�e�����JN���"0"O��YՏ��t9��(��*
�>�"ON�- .1���s��-RsD�+�"O2h���}m��Q�@Ʈ^S0L�p"OXI��@0nP1t�G�eCY3e"O�-�D�F�Z���q�\9_pa��"O\���(�v(�8[ ̬
�΁��"OzL�� �ii��F)?�܄�V"Ov��.�4�Y`g �G�ZA��"O@A�	8 \�5!�.:א H`"O��c���;e T9f�D��RE��"O����c�x@7 	}�NY��"Ox��(ז^��`C!�w-XY�"O��cr��N�J8���ӉP����"O�S ��!R�8`aѺ^�J�e"O�%��(�;G��`"�ͅ�a�:`�"O8(Q��(_¤h�lA�,Ҡ�Za"O�	�b�R3\�����50�t�	'"Oh�R�	âD���F�1&��l��"O�L1B#%�Ƞ��H�pyh��f"OlJ��>M�!��O�$��"O��Qe@�c�|�8 �z����"O��(Dg�.D$��s�T2
��,��"O4�C�,|��+��
3���"O��ʆO�7n �QǷ%�
A�"O��l	.i�C�
y���"Oܐ�$Mvڬ�ADƏ�P�
ՠ2"OP��ANU�3\(b�MhJ�"O���$�N�FbP�eBMdn���"O"�B7p��pju��6|G���"O �ӆ
�$E�E���F8j7jHc1"OT*���:;{B��1-͚y�rU��"OtTb���%q�Iⶫ�0L��1q"O�!N_�a�pI����3f��PT"O�x	`]8=e�m�� ͠
9ԺV"O`�2�	�T�$-�"��h���"O���S	�,pz4���m����"Ov�sUHM�s�Ht�À	�-|�y�"O����C�c��l��Oל"�zBr"O��6�H���o�k��J"O� 0ʅ�E����r�)&U:���"O
Pէ�5@�`���Q�c=��"O�Rt�R8J��԰�A5@�F�Ц"O�0�tȗTo��B�x,$%2G"O�}��JzJ�dA�jŘ��"O� ����-ƛ4�B8 b�ʢ5�ȣ"O �	�Y,��Y1!��Q�:��"O�`��=Ţ�F)q�^Y&"O&ܻc�V-Oz+T-��b����g"O6��d�ҭ����Dm(��EГ"O����?y��)�킭���;B"Or�X��b�L��£i�[j
�'��ܠӠ
2O�02�B]M���'9�0�/*T�D�dǜS��'X�,C.r����f�`
�y�':��t��%B�\ih6L�]�c�'<Ҹ�p�U@��U�%�=	<P��'Ov��F6~�,){���I�F�S�'U(�Ip��.���h"-�X]�ő�'����4�Y�P]~�4Ǟ#<�i�	�'�����#��h�@������	��'��b%,<,x'� y@\�
�'d�51����čP��8~&���'�$]�`BZ*'�&��a��]c���x� K1d�j��W�`=)f
?�y���+9����dCT�g+>Yu�^��yrkF�b��,Ka�T�|��5H)�y����5��@4h�:��S��E"�y�bU�3}�����Q76�нK  ��y��؏Wl����� 'S�P�ż�y⠗�8���РڀQ6Ib�G7�y���/�*�
�G��S~�`ES��y2iݰNd©3��<\𠂃(�yB�ߵy��;#^�qG��PR%�y�g���%ѕo��B�������'��!C�I]�H��,Ք�����'lԉ��!�:`������0
�'ߐ�{�+
�CR�����C}�$1{�'�0͒�)I}�ܱ�?	l��'vFh�E6̬� cQ!{��T��'�ʍ�3²*Q���3d�6�h�'&\yi�!7I2+�9a�j�	���d�%�Ȼ���Z��D(�+�3a�!�ě8�ړ��+.޲�P�J�&�!�$H�y'P��5�Y󒑐)�Z�!� [�>�ء��2�"|��ɓ%�!�B�j�H��D�߾:���錀S�!��
���-L\2�����~�!�QZ��}!�\"$`���A�!��$OF�(B��R�4�����1	�!򄇇u.	��JG/@���6 ��!���-}�)Y�gU�z-�ܚ2��j�!�dСH��9��Y�4����h�
�!��tp6�rG����%%!�$΢� ��2(�	]i
$Pt��>v!�5t@|�p㈦TU���e�4A!���>C��]��x����.*!��o��f%�H�H�h���>�!�D�4{؁���Q�.(�P��3;�!���a	��֍��>�� ��gK!�C���������0ɰ�h�8D!���H�����!�P�E�"
��L.!�dX2v����[&�)WA!�P�=�QЊ��_�ޱf�)cb!�d����\�R Bc�ь7L!�ą�M�(�)���
`�X���K��!�d�)<R!�ޏsPek�
Y%!�!��	-F۰AӆS�(J��qO�0�!���6,�W��yXB,'ծJ�!�� �®�;1tQpD�,y��[`"O�y�3"��~���s�Ý(��!"OB!���h�0�۳��6�఻u"O�UI�ǰQ[��ZDm��/A*�S�"OLu(� I�(�LÞV4J"Ofܰ����j�&�"␉\�2"O� �s��|uR����I4)�vt�"ON}(2��"V @���?1T\�T"O@��棕�MLh�I�@r)u"OXI�A�&,���Q�A��8 $pr"O�4�'d�*7 ��K6��;S�5G"O��B���J]6�p� M�I:�|3�"O��;$��}>`I���,蘲@"Oލ�@�I#�RճcCI�h����"Od�k�"b���$�-$���"O܁��ML��T�G��9��,z"O���`L^�A�*��b�ȧzT� �e"O�@I��'1�]K��\+F�\( "O`9yr��Ȁ�`%*}Ԣ�q�"O�Myr��|�B�af��x@cg"Ov�a�O�M�B��7嗛	�<XR�"O\�)��L1G���p�I��2"O��'��8�Y
�Jυ����"O��x'�//a�tc���+R�w"O0�)dL��~�&H�!S-R��ݪ�"O�B���&5�@�@�A9P��!��"O�H�t�=xF��p�O wj!�"O����i��p�ޙ�C�).+z�V�>9�Y�4�j��ƫB��@P�,���ȓ��ܛ
�.����5A5�-��%�y���ԧ/�t 3f^5N�p�ȓy����Ȝ�/-��Ғ�گ~��Q�ȓ�$h���O�*���˖gX(�����њ��i����[BH��856��ȓoGHp��P���S�O�5��ȓz�L�Am _T�Akpm�UJ���l�4!pC@Խ|�Y!���?���ȓIbDy�A��,���5N�n�Pͅ�]%"@i���(c����DF�=d�B,�ȓ^%��҇��/jYx�
��Rs�*��ȓ���'�ɮc%2#F�>���ȓ8% |�eN 8t5@G$	�3*)�ȓ9��R�G��)Q+���Kt$!��M�<���l��R��)�R%  ��c��U�I��+-�|�RI���~��h�� F�̑:�H�}8F���O��a��[����r�9jZХ�`"O�	u(�&0 �q�(�WuP�V"O�i`vJ�Rt��ƇƩ�T"O��� ə�H�z�ʹ}�Dr�"O�˶�z��<�� ��A�"O����][�h����<�f�1�"O^A��b�2Ψ�([ vڄ�ȑ"O
�A����^d��H@�;R��}�A"OPʕ�ScG�1�pK��K��]["Oh�(�J[
R���zS랋b˖���"Ol	
�Q�;�,����ʕtb��r�"OJ�X�l�pD !y#h�NL���"O��CC�
��Ѩ�FV�t6� C"ODc�H�FD��dV�*� �A"OR[�&\�D�T!��J�p�6"O�e�� K$2��9�gBǜb���q�"OhpY �d%*TX%���
p9�"OƑ�Ek $@1�i��/5�dMh6"O� @�鏰< 9��~���6"O ���$T"W�� q�N�)��0�b"OVqi��Y�L-�D�Y�4�Vh� "OP�.��t�,ПK���q�"O�(h�`[+N<�̍H�XD�5"OZ�@�0Nm�2$�7�b�;3"O+�kO6{���JeI��o"0؛#"O$H@Х��5ր�A��6=6u��"O��k�j؈=��RiՃX�8��R"O��a�OȎxt��'H��ή�@c"O�����bK�6�Ά�8)6D��遮�2�&hZ�Eѭ(�jth�
4D� ��D����@��u?B��c�/D�B)��I���m�t�X� 1�"D�H�Q��6���p�&ѡv�Vcr,"D�T�Bi	�$݃RA
r�B���@ D�B�.A�L:���G.KDE`��0D�� 	�|䣷���'*uC��0D���4�]&6�N�Z�C�'2f�1�.D����ͥe.��	R�i��å�/D�x�`ӕ���ࣛ"#�闫0D����F'(Txk��x���AQ#r!�dſ<��۲FM0�|�w���/c!��2kR^Ma�N
R���!	�4�!����;�*��d� �!�� �5�!�d��`��*�&�}�2K�,d!���0�:�I�)�Gp��hр�>>M!�䜩q��c�D��Q�>���D?!��ٍ
�� (��e�)c�.�/[!�䐓u�5���B^Zx���ьy!�d6� �`�H>G����LߟO�!�$9�$ ��*��%[ץ3{o!�^,���x��C�lD�A"T4sn!�ƬBGH��$���y���`Ћce!򄑀U��P��\ wpxKa �!Ux!�$S�=�$5��˔|QR�cwE�uj!��W0JJ�kF�Q�\E���C�ދ8!�d�*(�H�c.X������P!��U�`>�i��&����(-I� !�G2N��t���̥j�	���v!�$�+wKn�9ቑr۲Pcׅ
�\�!�$�;.����N��;tu�񃄧!��K ��#�4~:��&��@U!�D]�� ��N�*	*�%`�J?!�ē�2�![$e�<�NY D�Ϣ;!�䆓�|��b�9]�"��4����!�ė�i��,Ғ�; �X����F�[J!�$�\y����U�z͒t%F59;!򤛻x��	�T"�&|���i����!�H�D	<ݘ��ƞ
�P���P>y!�dΚ	`�����u�D�薨<!!�d�y��a�e��+����c��  !�D�Q(��0�e��9�%G!
�!��7e=T�c&�=<���($��'�!���]bHĺ��� \���r�#.�!�$����;�L]��5 ���	�!�� �b.�̰���L߾����	w���D0i�z)PC���(�-M�y2 ߗ϶�:�����HC�9�y2��6!}@Ġ����!�W���y�K;\�r�ְ:Z��g�˰�yr+��L����f���gЌZ'��-�yb&_��I+��R��Y���Z�tC�	(�+�ڏD�q�٧~�RC�)� ����,\Ҭ�1�-o�,�p�"O�P gKL�x�n���� 6$ءU"O�{�GJ.p�@d8�#�`R򄊁"O�+&�� Q{n袄�@C\��"Oe��n���i��K�CB��t"O-��%��)��a�;�6�S�"O��Jt$�Lq2�!A�OH�� "O��iΡQnU��Đ-{�"O�{C��+P�RS�Z;�"O�s������cC�^�d��D"O4`j
l�l-��D��4�0x�"O��`1��kȀ��зcT�"OP�3���/h��ī�I��x*��"Ov 1&LDfP�gɅ�Ac�ѐ�"O�A�8kq�MI�
U{��E�"O$���O�	)ZF}�D`��d�����"On|;'�PQ��W =@��YI�"OR88��"z�x�nZg�Ĭx�"O�ۖA9.Z��K`����x��a"O,;�,��.���gM�;<��TzE"O�#q:B��db��Ά_�΄B "O*��#�X�m(�'���]#�"O��(�C�CQ<�ٗ�pЬt!"O"����m�>�r��rÔH� "O*8(�GY+�������;�����"O<!�����/�`�2��иI8��Cc"O��HңN:p��u �,e
z��"OI�e�+϶��O�f����"O�œ�։n������>]���"O�:��B�)�0ؓ�Z3@�=��"O���f%��zޜ�[��8�F�T"Oh}�`��Y�����,��u"O����
g��`��D�*a��#"OXt���L%��sG�K7i��
 "O$@�⁙�qv�43��8<N�@��"O2��dJ.,�k��+:��Qu"Ox����ń�f���!���p"O��3�K�>IvaP�E")Zցb�"O��JvEԠ1�ni��ŉ?iMLA�"OB�ckN09�VQ�q�$��3�"Ob���� �5j�z��כ���g"Op�i��_�LNͩ��=��`"Ol��D��$�=XADT�|��lk�"O��cH�z̰dG4����"O
l�R(E���� ի�ݲ�Y�"O$	�@�Ē
�	� ].9P�Hq"O�a�/ �$)�a�D�1v���"OX�s�3#���掯 �Hh�"O�P��]-.��T�G�� ��p	�"ODљ�LP����̎;�x��e"O��v�Kr�LڒŚla�tD"O�q��P'3˺�@��EyF(��"O��Q�F��BW&LB�EΩx�2�� "O�		�Q;�=�օY�S�r�"O��2�"זg�Bt�3Nݎl�0`�"OhipG�pdl8���0J�<��""O�A�C��&Um��j�K��D�2E"O��7 �IJ�J��ؙ,�P\iD"O�`��酙m`��z6j!�1��"OؐCl�6��A��Ź��Z"O���u�@@���H@�3J�`��D"O�M�E"�_�Jm�P�N�q;~�F"Olu	�a͖B�d��$�~"���"O͉��J2?�9�	B^���2"O� �XaqfLۤ��4�˄&	""O ����a#I�v��E"O��j�K�H$��W�ؠh�dQ�"O��h���O��I���,X\p7"O ��W��)g�"pHT�ܶaZ9�F"O`�� ���}��ٵ���\/0Pu"Oh�S`GQ�$�iBr!ԑ,б�"O�%i'�Yj����F�~t��""O�q��;`�0%�EZ�c �� "O������n�b�J�	+D��"O�)"�׹MD����K͓3�|��P"O��!�ծƙPB�O#ZH��3"O؝�fO�'Y88" �O5��1g"O�B"d_�x�բb:T� "OP<��E"�a�a-C<{Ī��"OtpjƂ*���#"�)U������g����gݚE�v�i��%!�m{�d1D�,anXטx@rBI��ڂ#D�Ti���������i�V�!l=D��s@ǆ5��rd�.wJV@B��:D����-���h�`�L���%�9D���#O�����NW<�ڠ+Q�%D�Xɵ���qZ4	�V.D�t�a�!D��+��Ee`���K���hؐ�?<O�#<q�'��/n^�᱁~̚�0�f�<�E�7��Tb�ZV;�L�EUg�<��aQX%�V��`4�X�@Uo�<1�DF�e]���CT�=�Xq��(Li�<����r���)��0W��� h�I�'	�'��(�� ��&���=x֨F��(�ȓ4>��Asi�6�1���֪v����?qӓT�p�O\3g���d���L1�?)�[��-$����b�
�_�a�ȓ��Y0`˛�?R8�c�����ʝ���~�1Q([4%-��S7�Z�gf�A�ȓ"*���wOޙda�E���Z9QV�Eb�S\]��1R�E-���˓"�&L����hOQ>Th��
P aA'�!:E���O0���'��IВLwr�hV$P'�|���K�c!���$�nI;��xLӢ�D� p!��v��pT�Џ^�1��*FVZ!��].ۆ��2�XnT)��1n�!�$�*96>l��A�=gb �$M�-��'Eў�>��F�Z4��)�g�K�ߪ�� �!��x����Y|���F(=j��ӓ�OF��D<?1c��,5 x `���X�ĉÅGO�<�S�:�fȑ�kˑ!�Zd���LH�<���iŨ}A�흊����`�h�<1��ȝV>T��� Z�8Fʝ��l�<ɰ.P'�L���-[�%b��Rp��b�<y���B���2��Xj��Õ]�<���)_��Ŋe-��U��0�&�@�<�# NE�i�g�
$��Q:��N[�'axb!�	4���ژ�d�2[uHxP�"O\$��!��QJƆD!=q.�bu"O��N�+M��(V(��h���d"O~��BZ	��q
%j�5��q�"O^PCt��l||)k�i�+K�ܻ�"O�1�҉)�C��p�z�0"O��Q�ݻL��xp'�>f�(��0"O���0���:�����^2��'"O�r�A$2�-�����DJ�"O}#�*�`Q�b.ߘI����"O���កV\��B�-ֺ7�6�9�T��D{��� 0���+��'�u�C�( ����"O0�����;�����?� �"Ox���̨v��t�! �h߈9�A�'`b�)�'3���Dʠn ^u�	̈O��!��v�� �����?�`��JXh"�M��n� ��ˏ*Gm���BOڶm���ȓ@�����zL�����)lX��'vў�|zG��\3"�7�	h�\��oSX�'Eax��	�x�걃�%��,�|��Z��䓙�'u>�c ���|�ԩېfL�'��%�5D�����}�*J����f�2i( #>D����A�)��d�����HObH�<D�8
�d�+E 0�Hv&���^A!��.1�j0�KH�nj�,��H�*Y+!���y�x0� jF1N�E�0f̘|!�d\�MQ�AI�#2 �j�P!>!�d�;3�x���ܢa0�XR��@�!�DK��J���G�#m'6p4AR!�D�&um�L�3��!H
& (�j�5/J!򄍟;�����J�P��
�MD!��Éh��Tq�� B
R�H`�!@��'ub���Y�{���� �T��"E;�&J Hd!�d[�H�sE��+
!�T3�$�%8J!���&�F��F��i&��q��f�!��&���Q3f;��A�g��� p!��[@�3S�]�"p]���A�:!�̧J~�%Lݾ%�,X��޷~!�B?e�Yb��Јk�"��F�'�񤏺��%%���.>�,��4�B��l����%���TIˆ�V�RyNC�IR^,"׆��y�$Q���=�h�O*���On�=��k!��$��t1�E�"MH8I[8Շȓ��بs��.t$���A��4f�1�ȓ��f�0���"a��k�n���C10�2)Q�ݜQ�-�}�����P������B�e!��$e|i���$/��˓�0?��f�amJ`)�j�I~�$P�([���D{����x�j���>X�L4�����8̊�O^���"W>��"	׻�, +���A�!���DY��=w��Xȴ�ȭ4�!�d�/<o���3ƛ�N�&�!b䚳N�!�Dث0��Bwm�I����3�	6�!�$��dA�v�Og�*L���d�R�'\a~B���7>����Y�7q>-�#��y���<]�^}b��# �:}���O����?����0<Q�M��8PJ�3�D��}_��Pc\�<�V�R05xa�'l�`q�gTW�<�`A�,\nQ؄mǫs瀱6c�z�<	�Δ�;w��Ha.�)G	,!h�N�v�<�QgIT
����H`~�s��x����<�������f۞9��CrD�u�<�å��#���4N�I��EH�<1Q�٧(�Y��с5]J��%�A�<)6*
9Yq�,�;&8} Ǖt�<���ӂS�x-�@Ñ�:T���Gy�<����
j:��D-U��D�7�\x�<i�m�\'��@P��50�ܺI�q�<��H	"y-�#���5K��d�ip�<!1)���a���ݲ~PU�Rq��hO�',�b�����ؠ�"F��
[���ȓ %LE��i�6r���
��;r��ȓ[`�"�܊/��̛����1�������1k��/B��]+��6�&��?����~Z&AX�4�u�$j��|�+�(�K�<� ��;Ro[]��)SK��吙k�"O� "C�bЀ���O�����'+�	�<х �D\�$ȑ�I��X�#n
@�<��	���-�_�4
�T�<qG,[�'FL��b-�&a(�y���M�<�g��
{��(Ø�P��)xfB�I�!��a��S �=z�/]8D���p��	�B!��#�8e�����*�lC�I?���C���7��h�7�unC�(rX�yC���1U�5��/��O�^C�I ���deM��L [T�&[�B�0z��豢��n��c��B-��B�ɻ/���抅*ND�\	�/ %O�j�O֢=�}�c��o�@�겣�*�`��P��Q����	p~�f!K0���&'B��f��"�y2���.H����h�!��Ɖ�y¡Y+/�B����[G0��j��y�� B���@O�;�6�2'D���y2�@�K�m�a�@�LZi[1g���yR�šq��P7�Y,Jn�aNۉ��D9�S�O�28�$c�4M?����'O�(��'��rW��ag�h��ގ�<\�������>)ub��#|��Ǐîz�y�4#^�<�P%B�=����C-j����OA�<1if��a��&(�R��z�<AB#��A �!�
e*e@�<��ٓB�	���4^o���Q�F|���hO��;�@�z�+��v��{R	��E��'a~rj?L8;�P�0#"�1b,��y�(_����ȍ�#2�Z��ܚ�hO��O�c>�ɕ��{(p���5���g-D�P"�I�'a����D6y����-D��2�^�c54y�U�=�R��SD'D��B �Q�@8(ړ���"n�yz�2��]���I�	͇.?���2@e��.D��F U�����F��q���+D�t2@aS��4�+�b�_x���T�=D����EB�.8��C�fY
b�;D� ��(D>MI�ʁ�r.$]��:D��`�O	["J��DaZ�|��� (5D��f�ֲ{�p��&�VIҔ"�-D���ĺ+��h��}�q�eH*D���U���̓�k�1��+��J�<�u�O=��P�a��!c($gOJ�<��MG�R��m��ȋMKV��f%WH�<� ��"�*�iRO@�Z8h��b�I�<䮖�G��i�̘��X���MB�<�s�V-Fİd���Y�_�]"��_��R���O��a�Mƛ[J��b�-Lt���'�4<�%K��F�"H#R"D��t{�'Iha��ۗt�(�A��.�ޥp�'�% ���	"����H4����'�؉�r�_>�A���)�X�x�'��H�U�,n;�lq�G[ʴ0�'�N�"1���Oxxm��Q4�������Q�"F�PH���Ce�d��hA�!��[/HTH��%�Ա���<�!��z=�4���rVDj��d!�ě�Nņyrb㓦y�1�%'\~Q!�DÂHG,X�V��p��2���!�d�5# ��L"
�t �ğ-+�!��Y����-	�H��U�S��	x����@�����
���x�`�#D�X3򯆞���a%Ê�x���$$D�� z=�'�
�b�5�Ae�3�YXu"OnI�4n��g@��#� F� �U"O�L`��Y&�h���+C�T2L,`�"O���Y�pH}X�J�\|q�"O*��B^on��!Q��;{ʱY`U��E{��	��u������<�����<l!�dU*|��n���Y��`�G�8S!�d�>P&lx0��Iu��昢S[!�	+{�����09i�	����FK!��ÊUK��� ؏D`4k�b
�J!��!'ز( 
�����jB'U5!��6veH�#LP�M�L�F�!�$,Ou� �v;h�듊M�!�$�1-Pи�扖/�0����(qB�)�'(�g)��%��uG�ĜZcb�p�'W��#a��>e���@�`JzЛ�']�l�� ݣ(�VL����.l��H��'��a9�(B�1�F���lͱvo�Qr�'�L5*Df��<�zi9G��ts>X�'�Rt,ێ@���;u��tS�@�'�n:Ѓ�6,�RY�*��p8����'Z89��Cz�9ub�9ls�h
�'��@����/2�d����:_#,���'T��(�·1~Qz�[vϙQ$�л�'��Qz��¶Xۼt[�L-C�t��'y���g.�"\���Ko;4̲�ϓ�O"�r��8MG���*� D�B �� LO8��bQg��Y �OA�Q�r�ap"O|HA c�_e�x��	O߸!��"O�L�U��Ka$����/'�2ɓ�"OQi�)Xھ�[�
��(���#"O����.E�|�z�AGj[Q#B���"Ov��R.nm��k�H܏[�=X0"O�k��I�;��`���U{�"O��T�Rj�f�ؠF�GN�t��"O�9�5X�Fii�šk(&A�q"O.(��?�ʈ
�M��E��|�t"O�thu��^�Rq�FK��J�z�"Ovq�`�V�4�;#k�:->L�"O@�9'��*gT��ԫ^��آ��$�OĢ=��[���)���<<��QƋ�8?�	�ȓa^��]".��ى�BD�eK����f�Vyi@ ��C���!�V�<�����2,���c�T����4i�&P)�3D�c��B�6D�i��
�_�qڱ�)D��ٕ�0a,��qU�C1��Hȵj$D��
Ң���Ⱥ��A_��s��#D��Q�	`���	,H�,#D�l�$��:NHn��c��>8�A��?D� �ÒR>j-��m:�)�b�/D��j��T�q����/S�Y�ԙ3�,D�\��e�}���Q	+B���7D�"��,3�.t2q�	�v?�{� D���R I0z
\�왳rp��TA:�Iz���T�"t���F��cA�٣؂C�	7f�
,��hȲg|Н��o1e�BB�Ɇr��e��OD�ĚSw���'�B䉝���S⛖_���!�䆎7�*C��+r�|r#ƌ�,f��"�C�-+�B��-w��C6�n� U�g&��^8�B�	�-��	�l^g�H�d  u�B䉫j�8�	RE�%8p��qZ���C�oOּ�CE��A���wrZC䉝=!�٩BE�$v�;0앾8M\B�)� .�T�V�8x�� !�Cp"O䂦��+�N��u G*��hiE"O��jv�;9�N@��dV�
�
%�&"O�2N
mb ����dOf��T��;LO�p0V��G�ȉ".зר�y�"O�]C,:Ze�-Ҳ3��K�"O��������iJ�(����""O�H��G�1�v@`�@�#���'"O���")�@O�3b%* ��"O|�srN��Rڝ��C8CnD1u"O 5s�&ڞ<��	[RZ|��"O���a��}.�Da3*Z�qV4��"O ��t-��2����K
;p�9CF"OI���'�]��|���P"O,a�W�:f'Z��.\�M��y!"O
)�e�$/l$���/%�
q�0"O\t��Mݞ{�<	`QA�4�$��"O�X��C��:����9J( YU"O|)X��F�\�+�EJ z�"O�yCЯB�H�|'D*����t"O��Q��F�L�DjWŀ���	�"O����jU�c:D8z��N�~��`�"O8�yՂ[�?���DÍr�n䱰"O⍲Qi	�B΀��d�E�(�"O��E%�%i}�ت��A<%���O��h����l�"��֋Ĺ*&��qF"D��s�)eԺ�����M�]@D,5D�0�6E�5'qYcD��7\4fu��2D�z���,So�ĳ�G\pHHA�u�/D�8� ��=d�0�h'�ϩxcL2��7D�ta�(��c�,ɓ��7:0	��3D�8z0K�P1N��.K��� *��0D��ҥ��� �{s�K�XƺL��g+D�xQ���)7H(��@���|�<D��"h�}�t�IF���NjАg�>D��jq�ؓa� D;�,��^gh���>D����#��]T��U��]tH�f;D����� M=�D��t�x��7D�4��*:���fAΆ"��K�:D�d�V�xa�i�W���7z��� 9��:�S�'	bx q&�k���r�;�X�ȓ�Bw�.C�m�&�!JT��ȓ�lktI�y��Q��h�5n�d�ȓZvF���H -� 	K�J=9D�ȓ8�2ŐQD��I��P���N j��ȓA�9����f� ��J�'hr����@X�E��c�x��Y>�Ș��mhT�s �˫&9t���aW&���ȓD�����@-x��m�6���K4���ȓ\�٢�� $@L�%Àz���Ol���q	�?kD$�Y"�B:SY\!��7,�x�<_�R�9"CX��i���]��5K���P���,Awf݇ȓŤ0;��:h~֜�1H\�o2���
�����H��Fe�1~� �ȓ&��M;#cE������ʗ�̆ȓ&$��J�#N�q��vǎ8ɚ=��H�.Eˑ�I6H��XŀƋ?t�y�ȓ$ͮɂ�-�3�dI���*D��i��M:ڂy�C����űqf>������*�j��J�x;AIݝ �&�k�]�,D{r�I(����î:��ԡ��
bC䉖s:� �ֆ͸�\��vG�<C\C䉩b�)"��I&*<�@iD(~B�)� 0�+�gb���/�� ���U"O��j���{�,1@o��'�v���"O�h���.NU�4�V+-2�00�]>���j�K0M<AUd�:f`?ړ�0|jw�O!p�ܪ�����B��z�<�� 0�������\�d���w�<٣-��
qZ�e]=Yr�� ��X�<ɑ%ƞs�|(�gH�(�!Ñ�Cl�<Q�,C)OQ~E#7g�"`�ĺd�a�<)�N5�V 0eD�5P�FD�]�<��2��pQ��<�\z��V�<��
;5�ٱ��%5LMR���X�<��$ ��A�����3��Q�)�V�<�R���;�J#ׄ�N��y���]�<	3ϑ5�t@��+�4n�Rt�~�<�J�Z{�e ���Z�2U��o�<����jA`��'�	s;�ᰩ�@�<�6	D�F�98��mZ�e�V��E�<��b�J����b��6Ov\I���D�<�BǪ\K	���9k52�A�<��!�B�yE�;�L� kz�<Y�$�R2����gWRc $Zx�<I7 �:
\��h���9�*U�t�<��I�YA^l�@)�\�֍�%�NZ�<I����MJB�c!^�O(�S��ZW�<��&�E��b��s��R0�O�<!�i�4W�|b��Z�,�C�R�<�bI�x�iǨ�7�
�P�$Cv�<i�( �_��]b�'D+O�"հ�l�k�<����4G�AÃ�L2_�\8�"�M�<�3c-v�,�N��.�XͲ��@J�<�0g��Q����T!9�=1�i�D�II���O�(e�Dk8!|�X� C%r��r�'����@nE*	A`���Z�T	�'��X�S+�;O#
8x'N̋�&L��'?���S�԰yQ����c�F0�	�'���XRBVt���` (��0�,��ȓ7 �ܠ`Q�Q�`Ԉ�f L��`������u���iܸ�WoEB@��ȓy�mrTB��J����Lŋ{(�хȓ{L�k�S(P��t�e�M�G�J��ȓ ۸Iq���ݮiʣ�#�����	W)��^ظJ�)�C"����4��0�t�Iv|L0'��1b�v �ȓh�
Y�d�@'����=�ƓPA��s�#��q|h�G��U=bx��x�㝵%�:h��]3Fb���@���y��ؿ����a-٬0C����`��O�"~�E��N{ɹ��/D����g�<��n�����"M�[������c�<Yc�1Y�>���K�$���zS�_�<�����Jrd� �����`��S@�<ђ�ݾzAH���� �,>���V×e�Q�':�	�?�l9��g�`p�ȣ ��2�"C�I�T��cY���ys2MW"e�����O��	�u%��D�Vj�}�,شy
C�I
%��Z&-O	[h���	u�B�ɺmj�0`�#+�q�­� Z�B�	LB�*U�xm�tJ�<7�PB�I<T���ነ<*yI�-&L��B�	�T����?�� c�~B�	�]+��7eQ$�J@�@f�:�&B�ɂ+-�`rrJ7k�� D疯X���0?�`�ؑ; �=%B�zV�Us�<� ����OӸ<G�������;����"O�,�T��9m4����.]>{��r"O2|� Ɠ����!�A�UIp�9�"O�y�V�G��|u��K��<�|d	�"O��!�H����4��u�T�[$�$:��<���K�8�b��q��ԃ5�ĴM2̇ȓt����L|�YSs��)TxP�����P@��s�(s5@�#^�X�ȓ)�h(k��R���Zw@̝@�Ćȓg��0b	_�(����)Ů_:��Ɠ�N��6�Bx��c3NN�RP0�1�'8Ԅ��3O �X"�O�Do�t�.O&�=E�T�%��P�RcU�@�J/I��y��K\��%<C���!�/���ybfF4=0b�S�U%$��ps4�
�y� J o���RU��f��d��1�hO����ěj$d�JY{��*T�݅*~�y��I�c�B��6(���1sI��pa���a�@��ْЭ-Ȧvr���U�(D���FN	�r"�+��F�
L�rG:D� ������uF�Z���e��8D��a��
t�xس�Ɨ&8�ĕ��+7D�p��⚁/�W͔*{͚����5D��yso@L��R��:�d�e2|O|c������SjJ�	�&6�ܸ1t.6|O˓�yb�	b�\1w&�&w�&��2+��ygB,}�Q7,�o_�5r�� ��'�ў�O�BԒĂ�:>��!���@<=���J�':�}��O�a:�=p�O3.w���'HN�y��5ȩ�� D�3�4A�
�'��9�d@�	kP!��`-Ζ�*
ϓ�O�a�����'Ӫ���┍��c���-LO"5P�-H-�Dt�6�\�7���
c�'�D�
���A��0�S�K�Z7�'�ў�>=e�ΫI��T����<O�u�p?D�����7:u�4� m�T�� ��2D��"B`f�M� �#����5D��ن�,��i�Vfߊ{���t�2D�XQ��#?z`�*�(�k�н�c�#D�ԛ��P�ұ��	
�db����L,D��KU�֕h|i$�ǪE���s�,D��/�/;G����ENx�X� �4D�`�_O��R��Y; k���ď'D�P��$����1�@@���hܑ�%D� ��DЖZ.1�G�}�^ ��#D��jSO��8�A�,�f�-��0<��jU�"p8�ՌXQS�FhS{�<q+�)z���'�5����u�<�o]}�T�Š 7cl�ـ��Qr�<)��z*<����:(>�( gCm�<yU��:FN�����B�wj�m�5)j��|�<�(*X?N�C��U*��%�!Rg�<��?�y�&�\��"�Fb�<��I��o�t/��Y?�4��MG\�<�tʖ�1�e҇ɞ�`i�oBZ�<A-�l-C#�L䤠jTdCJ�<����pf�4��
>��U
"��~�<$�P}��tJ�*�?�`p���{�	@���Od�{������!@�S�� %�ϓ�Oʠ3nԡQf�8�Q?a{Z�0"O�U[��I�P���7!P�J�V��e"O1���9b�4X�UA�*�$e�T"O~��d�TiF�%0fA"N�l|q"O�}���\-{@�DU$L5}��r#"O� 2��@lکAJ���4&��04���	i�( !߳k�`�s�]�.9	�k4ړ�0<A%M��h��hYSF��Uh�䟼F{2�$@�Nh�2�.躥��)ݚ)%���ȓu�D�k��V�Fј5��Y:!��^�a� "�x�톝et�ȓc4��Ð+��@�� ��/psh��ȓ�iӱ��0��<� *06�晔'���Sv�h��UO	>)y�0��7�ZB䉢:T��'��]�m�����XB�	'�Ԅs�ޕJ6�xiuh�7�$B�I:]BЀ&�ޖ�X�Iu�L(�B�I�sz�t�ՠ{v��w�_-c�C�	N �I&3,%�e$/�C䉮&b�Uh�Ɲ1F�C�\;2C�I?l��'��l��a���$bb4�O
��Ā�e���k��73!��x%�ъ9�O��=���0թ�+J��q� �4|XL&"OZə0��D�XI��S�Ph��T"O�dR����,�ك!��\�E"Op
��H#<[���mCk�aSS"O8����L�0#-K�Y��"O���0�ÏMf���&G�uFh�3��'<1OZ��G�K;d4Xe�ұd#~��2"ON��P�]�#x�%�\�r�"t�6"O�x�$M��P|�jT�33 �¡"O�1jG�Q�Xl� "�^*�"�"O���U䘰W��ˡh�Cq�� �"O� �pL׋�F���0+2̺R��'�ɧ�i3?1%ğ�]z 1�P8(����N�<	TB87|��*2���#�6��4�G�<�E��?�v=j5��-dj"����H�<b��"A6@DA B�bR��l�<Q�kB?K�a��i�4{� c��g�<vj�`�x�(K�`I�1�&�`�<��8xؤ���22���@�fO_�� �<AfD��P~��v��P�
�В����hF{��ɝ)}�d��@���i���⭏4F��B�	�p%��;W�A��J�:�$M�,���0?9Q��@��D�*[R)�ekRw�<I�jɮ%$4Z��1�X��AAu�<���=:��U�#H�
�%8�j�<A�oVKDX�z�
�>{i�U��F����F{��)�	0Al��qg�V<J�A ^�2C䉋B�D��&DS�w����t��)uC�	�P��q��C�,�L�xE,�ԒO����қ��H�Eծ ���p�)�h\!�C4��T�� ��;�b�=?!�䋕,k�%�s�[@I��#O�W�!��Bxx�ǥ�}#����ե!�D�8ސ,�R��;i:�Ş�u!�đ=i�>e�6C��u�$��d��ў��?��O���!�Ԓo���" N�F�h��"O�#瑣;E���C�U5|0ѫ�"OBmj ��x����C�=q����"OJ����x�$E��	,<n)�"O,�;u�2yf�K�Ѣ=[����"Ov���e�&gl<�g���W�ʦ�'0���Wg�-��#������ex!�d��yB�c�*:
�bq2�Q$��O��=��2�`m�5��]Z�����"O�"1H��sGp(���T_�v!""Oح(P�b��E2q�G������"O��FW�g���?oܙ�7�'��	c�)�'�� CG'�3P���aK�!/b����'Lў"~�C����<�0
��	�F���?a�'��T@S+�1ӶR��1S�&��-O��=E��E[8S@8��L8sX�xr�@��y�`�>*iK�H�"w5r����y�
֨K-D%O��[���B��|�<�pO��F�g�!2@J��4�@@x��Dx��S$;��ly�ⓖO9h�9�B��y�LH��l3�'�;p2<� L���O0"~�s�ӏ8M����:�mѴ��Z�<�d2g��PG�[�XO�p4.�m�<aÏ�J��q�� S�e��IRUNg�<���VO�\!��ŌeRJu�b�Gd�<��ƃ�F)�@�J� IY�L_�<�vK¦��`�I�!�Ft�R$JZ�<�S\la��;�.Ůz2����O���O�	!
'�(%n�.D�Ac����XB�	��L2 �͸>�0��F��?L:B�	�,{���3&<��L]JS�C�ɺ>o�X� K�l�	���_��C����1A���)������'*�rC�ɞ-�0��I�=Gt��eoRz0<C�	�HSĄy��R�(�|Pc'O�ck\C�ɵ)���
G�T�2'��c�(��?�B�	+,�a����Q령��n�:�"B�	<x
�� U.Ԯ0-���@/dE�C�I�����"o֎��������C��5�p:sѾ[�th�'Q7��C�I07�Z云F�;1	���6��C��0P�l�ҵg�~�P��"�
G��C�Ɏe(L�Q�#?nqԚ�%N�¬B�	=��L"� 7\6A��K	(�DB�	��z�q�,Ґ� \{�d�<�"B��~��҇A��m��&���H�B�+ra�e����%M���Dl� v{�C�I%2?`p��K�j<�@��S4C�ɝGRe��k S�f��'o�4"8&C�,C�D�+�c�6d�u.�;B�,C�IT�d(�El"$��M�+H(
C����ta�C�M� ��?��C�cz��a�B�	&���(јe��C�	l��|����<5fi��΍� ��B䉕W���0�!T�(�y���0m�bC�	+e�q9��T�����kP?>8C��/`}�V�V�B��T���ʮE!�C䉮rF�Q������+I	Ls�B�I�E����d�hjقA��.OvB�4 ����D��?AR�{ahŠ1s~B�	��8p��
�D��դ]�bB�	�70��Q@�tA������n�C�I	�*�D��?g�@8U@�,z��B�I�H����"T+r 5��B��ĩ��鎺9>p�hGC����B�I�p�Kbk�8+F8��KR��B�ɗa���#ɟfR �j���t�vB�ɕN��\ѓϖ�W�6 ��ꐎ-�:B��9	P�д�۶U T9jF�ͤC�B�	/�F�j�D{$��sn�#yy�C�Ʉ:t�.��~f�U���:~�C�	6�&���S���X�˒�xC�	���p�F/:H�#�	>4��C�	:;���xR��*Gv�9"�.� �C�	�o�vH�!�(l��v����"OFU����f^h��a��1%��0"O� �0@�m��P�*c��0��Y!"O6�R��T	N.�e����LӲ"O��&	�+�J��"@�]�
�?�y��R'���8'�D��p��L0�y��A�b9�Thӡ@�-�|%1��3�y���ScH���Ӊ{�j9x����y�x���D� CH�ݹ��y"���DT��Q�߷3���;�A��y2�˼m��icL�z<N���y�J�~󢰳D�nu��mA8�ydڠAp��Q�\)|�Z�8���9�y�X�H����fˬ@D��"�D��y"�4�Ҙ��$Z�9�LlA���yrD�D1v�����r��A#�yr����-"H2��+����y¥�_�:��b�ht�mCB�U��yb%O>�2�fvl�慖��yr@�6kK����J$c��y�(��y�U:��5b�dG`�21y�X��y���n"����S�fX�C#�y2%J	=�������(E琈�"��y�)1c����TfϪB�6�ZP^�yBJ�-%��8B�V�?}�@pG/B#�y����"��ER�6L���c��y�+�T���/�:ex�$�Aa:�y2��)pw��S��4VP�G���y2��ra"����B��%��IG��y�ׁ{����{��0Z�l�y�l��C��a(�C�] �철+�/�y���$�&DY��M�c
��0n��y"�T�7U���We��]��y�%��y����F=zrc��N)N�l�,�y�i��#��;"G�L�<�:sB ;�yr�AZ:���J�	Di6���D��y�
���8҃EĮ< }Y�����y�aL� ��P�RE7ު�{!e��yB�έJ�� �͒F��(c��,�yfB�B��w��t���	�R ��'� #U��s��mC��ܖ�Ҵ�'� ��BO}�	�hܫ'���	�'�h�˂��:n����#WPk~�`	�'����C`ߎ%%�@p<�	�'�T@t�23��5з+�3f9��'F�@Պؘk)�܈�P./I8��'8!y�d�M=��Z"+"Zc@4Q�'v�VS�V��2��8j����d<D��۵+�:+�\@2�AJ^]hR׌8D�t��Kj�j�bc��7�
��g�6D�D3�
���ZŢ�BęI|����>D���uB�n�I����wJj%�D>D�L�!i_�(�Q�A�ǑW� ��&D���Nɔ?D2��3��Q����m:D��C������	Bf&�PBt]��8D�䉷������H&�KA��1D����Lƈ�CG�Q�=7�595j0D�����B�m=@�D�ʽ�X� �-D�pЇLZ�Rp�1�UB�MzH�PO.D��zq�	- �N�5��a�S�9D��PVd�&_Ȑk�Ό�
�f��q4D�D#��1��$8a+� ~H�q�A3D��k'o�"X�NDJ��"<�a0D�� ^QPX�r� ֌%̰��gA��yBjJ�s\�B�*"�J,K�/+�yr��0D�s/�P��QD,@.�y
� ��s$���+lL���h�z���"O�z���9x&��7&�;��0�r"Od�g��]�r�Kf�@�p�HxY"O��{��m]	rd�3� �[�"OZ�"tAC�.�q#[�6����R*O�d�0�3��ؐ��gF`�'Gp��!���d�P��tNp�'p~�ST	� ]��������k�'��UY�&��A1�����?���'��I����x�Q���$Z�\�'��Є횣[�}��k]�=X���'Zf�dM�o���J�@�r!�x�'�4A�1蓳;"!brhWj�&�s�'W<�Y����@��HW?d3V���'����D�}3p���MS\���'�q��NH�p)� HeN�M2,3�'��`cȏ�����@�=��!�
�'_���JQ=���IQǋ�;h
��'!�}���
r���[��)5t漺�'�ʴPU�B4���
&��ty	�'��E��O�L̐�3ů�N#���	�'�@i���:E�~ @��� z!�|�
�'�n��H�?|`�(剖�;沕�	�'�b51vb7j����!K��1���y	�' �����.d������9��	�'A��*V)&�:�kW�D� x�t�
�'��`�� �ɒfe<&e�P
�'>Jk�J��������X�
�'�敘3K��b2đ�E	<_^��	�'|2T�d�[�h��x���^�[�> 	�' �d£�A�D�V�8�텉T����'ϰl�+�v�d��H�Q��'A�}:v���Xn�Ѣs�A,s2ur�'�����93֚XjC%��?�=)�'��5C7$�e�"��O��:J�[�'�:<��+DMh��¦Q%.��̹�'ذX�V�ҝc���b�
�,�����'~`�&�v�B��U�G�N��lc�'[v�1��T!+xl��F��2Q�]h�':�$3� Y�4��Ϝ�R�4�8�'�P�s��k1���7'���漃�'�4���o�?���FU�Olά:�'ZTK�'\�ZZ`��&���o���
�')�[ ���x��#k"�,�
�'?^@�0�2l���V	]?e���S
�'h��dX� 1:���o½:�'�� �f.�Q�yyTG�f4���'���#T-#S;����M�ǒM�' ���F�2��k���@��'���(�eٔg��lqd�.0V�#�'vt��N݋Yo���rA�'	td�J
�'�h4�R��z�`�΂4OF��	�'�d��
΢-�^]I�bW#	MJ ��'a�Ly�G:e2���5��LDFa��'�ִ��E	�&bA8�MءK2��@	�'�i�Ə�(&�M��lÕHHh��'k���W ��V
$�f�'*��iC�'�d�d&�`���H���%�0��'����Q7L0���sM��g4H���'[�%��[�_
=!C'հiVָ��'�D]
`	F;j�:�ˡ%Ю\!��I�'���K0�R�`I�����V#�EZ�'Rn�+!�ȉX��@Qb-]6Vq(I8
�'D��u�C�7&Ĩ�a�:;��{��� ��ʕgL)-�8���Fm#�"O@�r�F��R�b�5>b�lKV"O��s慖6B@j�TJ�aDXyC�"OX�(5Dǜ4�,i��)��_*8�h�"O�[Bg}
1kF� ��0��dɇ�(O�X�2���Z�`�Y �ջ?�bԄ�\�V ���˟q��Y�6hߺ�������s��a�9�6ɸ�ʑ?Ψ��4f"�O��'�����
�dҹX%��2���1�''8�v�ګy��CuȎ�-��s���2�S�4��uR�B+�b0x�'I�y"隆Vo�wH&�&�P�E�=�yb#J6/|8РrH�=��P�/��p=��}RE�
Rk�Q��F�E�t�#"���}���>���$�"?�j�9#�ړ~��K��pJ!��<`~D�1B7 �(E ��ɮr/!�Ϥ�a�s�9Ţ鄫�	o��OuI�v�z|�!�5%�4R�h�#M���ƓW�H�`K�,~�1w��
m4�Y�0��'�~)S0�O�g���S��݈V�1<O�Y0�}�0qu�4�E�	\��Y���-���hOq�� ���5OV�!б��slD({��'��$[�V���)�+�^Y����8�qO����Ʒ"^:�i��a�B���#����T�'3O�"=	!bέI��q�ۼ4 8�ⱃ�k�!�E�^�X;����:dhX�QM��xR�$ʓt��0��29��E��8��(��	�"qO��pF���$Zt9j �$��Hp�D>LO�H��*"qN�8�휋AL@(�O� �C^j͹�Z<�lHh � ��٦���I�ay�U��K��(��q9d�FW�0#<��
2?��$wV2����'M�\[r"�,�!�(�B� �� 7H�����D�'!�D	��(�� ~�0���Q�`{!�$ڙ ��y��]�@��mjP@��-y��o�E����?!A���E H<EP�0�g�N�p?�O�p�f�ފ8^ u��-<�d��"O��Z�q�~X�тG�j�т�|�>�OJc���E=8�p@Bc��?l|�'��5���;O���#���e?��`�s�`0c�x��)��d�X 2�+p�ͩqA�7q���?)��I@%WB�M�)$ٺ*oȧ~wqO����ɭ?@�`�,�
�
u��/@fm��E{ʟʵ�m�|&*! ��F���w"O��B�j�6� H�(݇�u���?|O�p$�'YU������o��]	�"O�4R��g?*�;$�T71�D � "O��C�� ~V�DL_?N��}2��'�ў�[�	݉-�xmæh��	
:ժ��+D��A�I�S��A1�W�5&6=�(\O�c�� ��e> ���7� E�Q�&D�j�G.q��!���-7�R �$�	:�hO�O�Ԭ�TnWj<�2�CŖ�@+�'L��Af.�6�S�c�
��H)���4<O$�r�T�@�)C��,o�ځk��'�ў؃��eA��Wb��𕬞=n��_�t�>ɧńE� ��j�)
s��).�z�N�'����~N�f���PA�\&K�����"��b1O�=%?�B�G#*ތ�҄����5Y�)�	l����'�|�`��ޤ�
@hR*Pe�l��
�'"���o��1P���A`�[l"8
�'c�8*��%|>JE� �!X�p	��hO���') ����O�?���I嚟��>��D�Oc�5��#@�^�PCE���6�X��3}
� 88�ON�g�� ��i��=��W��K����-9*D��"�cj �Q�_/�b�P�'?��1�$�|��"A;��i2n_�h1^�)�Mr�'�ax"!���z͹u�>qJ TA��M��Mc��O��Y�'����ė~n�Q5�|��)R�}и����p\��F�O�㞀[�-��T�D��(L�\�~�R���f̓�M+�S�D���6v���q�艓sL���Fb��}�!���VTNez��n���z���6L�!�֦y.!����2�V�0����XG�e�0B�^�H�\>9�b�1rhÕ�y�f����%��A�8�p��ЭF	�O��dV	pu��R����"�2!y��<i!�d��h�N�2�V:\�R����v[��D|�S9]���7�X�tl2=����l�����i�+������8([��w�E�+L��ȓ	]\<`�c�����w�ة$)�(��0]��%՚V�J4	vJh�m�F(<!��̞;��0 q�Q'tՠ�Z���'�qO�D��sƂ�ӣk&�}�7"O�e�v͂+6�d��1��*Apl�h��	T�O�n����1���:�/�&(����'a��r���-��k@�!�8X����?����j� �)��.��,�>#��'hў�Z̓l<`̠a����	L�p.u����H�ԭ�?l��s�DϷ4K0P�=0�2LOX ��������c�صUyf��"O��s�d��lU��s\X�1��BX��S�O	�#�җ �sNm���2\O�c��vD<d*N�@��B&Y�L!�S�0D�@��K�"4�9�POF� l*E��!-D�D�'׋Ĉ숱瘳i�0��+D�Tpg�J�< �����&����C&=��x����q!��{��ӆ
�1���k҆5D�`�����fȈ7_�^EJ�h�>L��G{ʟ�U�Ʈ�X�謱�@�<���"OH�0�N�jHR�ܵ='j�)G"O^�Xyw�P�Y*݂�Q�c_e�<1�hш<����E�~
�-@��C|���0=�s莣9np�YfD��N
�����Fy�<I�$�>��"ce!,�E��s<���\�\�uIW�2h4�Q��0͆�N/n��w$�(�,�s�Ӽp���$��E{�����8��b �ۉYH���@�<�yb!�4 M�
�ᕋ&-����N��y�J�N�D�3�C\�sx�ƭW��y�D�o���,y�Nq`��1nB���'z��O��d"�!t�yX杣��0���u�&�ȓ+��1BNϤ!�
�2�JEX�e�'�~"�7$-�X���H�$�Ѣ��+�y�h��m�JI��	(W�$	��
^=�y�J"*8V�ɰ�>L��s���y�e��~2(�g�T�Cɠ���b���y��@�,�Ls,\h��M��ybƄ}�h0B!�:z�����p=ɉ}��B�O"ΐ8Ǝ	��t{%(��y�!��!}Nx��L�.��u+X)�y���9E.� )�)*C�,U�);�yR��.C����&�G���⋫��'ǂ���hO�ղ>���2A��l��	�)���y�Jbn��Pz���G�(x�� �����I�Ҵy�G	D�|pb�)A�@#H2*��%�OyKg>g��5���W���y��"O 1+1"�{��e6�dM�W"OJ5K @�F��dCp�ʊ(�@pb��"|O� p�2fl��s�|�V ��K��q�`�����O���dLT�6Ȉ�C��
0 �H�¥G�H�!�+F�f������T��e[/�ax�	�B��і��/1g��t�F;u��C�I, ��y!�_�flYA�)�n~z��hO>��4jN�|v��MS�28$a�70D�l	G,R�y�J��\�="�bO2�D�)��=�'Jȯ7�lyZ�̓�F�1��`�<���lvnx��I�kb�	wK\h�<9ra��1j2����>4J��C��`�<�$�$"�:�f�w9��SŨ�\�<ё���v: V���<��rN�/W!�$Y�<(c�D'�"L�&d��:M!�&r�
Q�	�)4�����W:!�ʴM���IB�<8j�lQP�@ aK!�dW��2%S����9Hv����6<�!���_�N���2v��0��Z�A�!��J �tp˥BԤj���*����!��+�@y��Ο�A���z��ű4!�P6o��M��%��m�#�^3B�!��I�	�"�Qw��`fƸ�E:@!�Ć��L�)�D��EPj��pc�<=!��́4�.��a�� ��1K���K�!�B�[���k�/@�i�G�:p�!���yrԭQ��Z�H�B+���!������ H�(�ȱy�IF�2:!�Q�ڼA�K������!G��!�!�D�?���@��F����ulֱDk!�ق
u��R��=%M��3�-P�7�!��ڸ��|���#Ya��J�k�)av!�3`��D���L�)E:�X���	X!��_ D�| dǝz4֌&(͔WW!�P�@���ϐ�9,h�aG�<@D!�o���[����K(��Q" Q�g(!�Dܡ^�*ّ��ΗV$(l;5��Av!�d�� ,Zwl�8==P5{���!�_�hli�C�?"D�"�MG�c`!�ĝE�޸)2�(.;���[�fY!��3犌24H�f%��[�Fu�!�7;�誐b�4g���Z�LG��!�$�q�{ %Y� �}�����h�!�$�,�(mЕC�>̰5M  �a~r���j��Y�%[;ٖ����ֵ,%����%
��yRc��A�><�GDD&	˄Ts�'�y�GE }��i����������ʪ�ybc�9��X�nV�$Qۊ��y�#�:mKVL(�Z3_��ۥ��y���cՈ�YhC�L�N�(�F��y�jѪ]7��!ᝃBʈaC%靅�y����1�����B�DҪ��T�Ǟ�yr Ɩ�d�Q4�ի=�f���J�<0��=q��SCFE=5X���SP�<���� 7��" c?U:d��
N�<a0�"^�^<�׭U�R��EÂ�
I�<�� �)8�T��n]� �|a���E�<��#ݭ3M䬙 +*^��B�3T�x2�f�&8������II��5D��ACI˥���`nPK��%`�&D���G�T'.m��B�C���@($D�:S�N%7n%��'"ځ�F$$D�\	/nTl	�$O�|�pT��7D�p0�Z�x�Ry1#�=&d|�ō3D�Г�bZ!��u�7���saRP� 1D�PC�"K�<`t`4eH	Z��H��2D�� ��	��Kp*HKC�M�0\x���"OԓwL�<(�)��>+Ӽ4�"O`��P�R*9CLy��DB1f5���"O���k��3�D10#�N0F �#"O����ƅ9$�B��c��%���"O��c��9�` �P�H�ʵ"O�O�\����X#n5D��"O؜�$��?/�~�J'@�,q>Q/�y2�@�xLy���k&D|0��̱�y�*�2p� �4!ӗL2�Cs*͚�yB�6�\\*"�����OE�yb�O�LMvixV�ԎV�;�ޕ���ک�\#�{�����5�&� ��P�V(]�3�~D!�\�y�`$R&A*
��D�!VV�'+��B�� WWax���A�����yh�јr��4s���H�(@h���D9^����D�L��s�"-D�Mp����JKĉ���N12��AfA�.�~�*�+Y���i!
ڕ���'L���OZ�B�.�	Tآ�0H~
U`Ȉ1��	ل���ع����w���ԥ��EV�S ��D�T腭 �(�;�(�*6��Z���6��䝰G�,`�!l�3��)ҧ�\䰑+��Xaf�2$��J����9�'ɘ�4��>�Fǎ�U3t(Z���>{pAj������6���̉��g~b"�5;t��ԡ�|X�Q��/\s�Q����N��V����O�a�64Z�k��D�@1���L��4�A$@��8�Z�_��,k1��>��a�#N���BԦ�f�B`b>���7 #�����W9Y��|��<�	�)xq�>d�Γ�4P�O�:��1�W'A�; �>O6)�3�ܒ~r�� #�8� L;�_>�Y���B���'ؖ4����#$2�Y��ÆN̺I�'f�pQϑh<|�O1��A�ፉ">`���)�iX�A��8y��K"�W�o��Z�FEq(��g�X�!8j���g�'âг	�,[�X��-[�j�4!	�>�Se[�Q�IrR���ɹ$/o��D��F���z�zR�-Q6�.E�pQD��7[�*��w��f� �b.@WX�P�e/��%j,A 4�B�T��b��^^���RC*�9@D�) RT���'o*I`�@C�^Ғ��5\Z���yo���'���Br*�(���7:�t�E&��T+ ٹ��)�W��Cϋ?~+����̒@U���3��ȓG��LR�!$eQc���E;���	bj�A;4M��c�T�QcE���aig�\)� �7R쑱�>�~���Z�o�"x�WŔ%W��qЋ�N^ՊР�}PH�ď��hHa$U��p<q���b��p��<o�Jq�G|yR�A�J^���gX�X� B �I���'(J�_�&x ���>�P����ŕ1:Xx���ٻb������_y���j�'kj�Y�ͥ2P�lI�lO,�(y��'n$�Ѳ�J9`|0h͓5uȸZ�fҙ��Og�`!! >i̪mj�+� �fpҍ�ē�0n�����5��O�I@��äe|J$�(X�n� �d�O$%�s"��CȔYk�e����-�����y��F�J��j�F��2F��M3�(߫EU@��E�(}��)�2�(
r Ѥ4���SiI
-D)���"MR�>Y6!ɖ!F4����L��$�ݲL҅��/ש�@�E�>q��D�y�Vu�Vj�>i�,ǒt#2ĻM����\;Jx�����A��mG�'j����#�6Y�Qd�I�H�,ac�'�.��ek�*P1A<���c׊B�N幔_��@�!]*�U�����͟A�\ �GJO%�?�0�#.��{Vaò�}#�C]U�'�DH0o�I�5�r�JL9:Ĩ�p4	�����	PL~�?P��c7璡�P�1W�S)
}���ɣ!�(��d�سq~6��; �n�Q���)��}bw*ѹ/%���!�!?�z�-:.�{�(��[�L� �P�W���&���{R��!W�a@J�x��+̋��D;3<x� ӯ��Oj�&ՌpR4�u����
��U"R��ȑg�![\Mz���шOR�b$j݃?��
Qu\���"q�u���yB�՟0��-&�tP
*=kb�� J~�x��U���$�&���C˃�G�R�����^<0��i��"§6b��'��Y�Vd�_��%�>���V���c$EɭD�Ȩ@J_hJd�{��߹C^��']c���⯕:+�E�v-�j6Xϓ/�^���g?�)��ȵ*��"-�j`�5f'U�� ��i��R���[&�%/�)�NX4/#4Q�O_qO��sS-K8*�贃"iâ��a� |��|���K"8��ɸ�ԥ閥�k�U�����J�P.��/S���Q6_�l}�1��H���:�ŉ�>*R��tb�^2)4��+3[����D�L-h]�-O�`i"O��<���%�IM���'����(C�3pd��T��LeT8	�'|:)��(�:���r4�1?!�p3�'�Fe�s�-EE6����56u*1��T8����$��<$��!W����fҚHU�aA� H��Y��I%Z��T��'[��`mƙoe����	K��'oXQ�r��&Jl�����;}���I%�?��=1� [8�ٲ�S�!�$K��T}��em����
 �d�%�9�t���ntAc!*��A�,Bw�9�Di����&�SԠN�v�虇�)�  ʐ�D
K��1W��"q�8i9C���	T��dO�p l%��'�����
I��q׀� u�4}SL���~�@����N�j�Bd)�l�<��j�2���""�4:��f쒌�MK6�_2vOZ<�&�U׈U�Q	�e"��Ųj'"d`m�$��K�I�,a�ˡ,�{R����E���=�wM�IV̔	��P��B!�`K�!�ݰVdW���� hԂ
�����'D�]i�/_��L9�@k�~�<	��
�Sp4Z��װ
��R�%^h��_ζ�[�\;��HJ���b9ʧuT䜢WO� �H<����-0����{�`)B��?O�����h�`xQl�	?��u!P�ؽ#�z��F&Ĝ��#k\B��;�Z>KV�O/v^!f_���k�?p�|����!�Bк�+0D�Ȋ%j[@[�c���6bD�092�˭Y��14O93�y���%����x2�	�!K�i�υA�4@2�Z�x�H`%��o��\��.�P(���/JR��Ժ��Ɔop�	�V�.�Bʉ,)�a⃍�â�� �<62�xR� ���'M p�)�]�SA]5}j,l&>%��R��@����&�nT2�"0D� ��?ph���Q�4���ңLJ�N���c'K��֬x�O˭=ʠ�}��x�I���oq���g�(�~��ȓZ�Ȉ�@�"G�X��g��E��4U����	(���X0�ڣ)�џĹ'٤�6�A�iə%�^b�$|O��q�"�ḎNYG�,�t,��6��С��9_.<`��2��qqǕ����&$��L`h�Ԃ4-�R�
�b��h�^Lzƀ2���0F�P�*9�5j�"OTH��ĥ-��Tj� �<J�=*IE�UJT�2���O4L) �F�>���E.֠d�8E "O�䱠kT1\��4ᇍ�'����W"O�Xi�BC%d�q�LN?��YA"O��s�J���)R,O�u)�dc#"O*`B1 	���TX��y*��"O �d��!u 2`W��@͛"O�[3C�;���#Mȝ,���s+ �4�40�=�M?�H�-�	�=�,mrr��9�Q��C�1�:B�	�,�5JX�qW4-X5��/`6���L+Ί&�����L���S�'wZ�h ���5`n��ѣ2u�`��I�Zrt����]��D_B  *  aH���˭[��-�uD@b��WY�$�?�' >���1^�%�Ǌ�x�5��{BEٽ��A�	�@�Or C'$��=\Ƥ�p#�8�걐�1pH6P����zX�d��p{��rD�й
q��҆�̄'��9��(}���X�d�T"��eس�v}��˞eŪ���i�=̲�C�(��y�Eǡ
�`��BB**0�X��,\p� ��+!*`���Ïc�(@��E'}b�iө(sn��͍�l���0�@�z[�zB��<�$|c�^�<�Ō6���h��6J����]�\�Is�>�c������ɗ�XУ+�o	T� 팊+���t�FD�{���퓋U���a� S>�d��,RAP�yE�M.,���'>s�l�%�j�Y�O�/UWL�[�ð�|dXJ��j�V>-��#�p��bZ�Ph��S�9VE�=J��B5D�2w�Q8xe��iM�yx�0�RgpӬ9*WL�2o�)��O�dV�2L>�|zEm$v��q����$��dy��k��$;��	�?^Ґ��:OB�`G-�	u��I�C�ԔTڈ�i�w�qOƁʌ�Y�4QT�^�a�^�0΃�'b���A1�I3dz�� ���?��"�,~2�y���0x�Ԙ�q.8D�\�e��N�bu�'	
mB�PqBYgWD��o6}Ds���DحJ��E�7/ٜm1Nx�w �!���th�cE(��(�W�ö������)7B��0>Q�L�8�!�e,�!�tI��MSm}"M�,b���=�1B�\L���¶O��I�\x�y�%��ev� �gI	L�!�Lhz�MBG�\�F=T�R�Gڅ$��n�r�B�*6CZ��A�|~Z�Y�O̶xaA]3�pp�E�4�B�w� �Z�%��tG�9؁���q��J\�&R�R'D\���0p_��X�]�������8� u�fM	o*�#�C��v��P:烝�kKʴ��)Q%W�"�$�;:��i2��%L����J�^l�,#�'�5̰=�a�[�� �Տʱ �P�x4i��<���0^�43pK5}*���%�ĠO���ش%�$��KqXH���-Rm'�L飭�,ay�"G2k�0��z*�0���	���DX12�L�ҧYB�B�͔F��2%�����lZ�:
*apHI��l9��H|�E���',*��iρO'b!�RiE�"/�	5��-IHı�Ub0(�N���?}D-dY&��!$�> ��Zʸ� �Lh�ȑv��}I�ڙz�`X���	�	*Ζ9-kq��l����,�@�RAJ!B�ʴ�ɼO6��(��,��Oh����+P.�ȕ���]%O1X=���5�(�B&5O�Aʴ�j1�e@K��'�2�	4	��+�H7M�s(p��b�H�!Dq)�F>rg�3L���H�����Ė	z�x����K7L'�٤��h#�ɗl�^�cIH��L�o^O�	��H�R���=)�𡄥��=?&y$���t1vQ��(�O���k��FV9i�ʞ5$6 �y6&�0/~0c��U��QSr��IU��ѡ�����	�x���鍭IS� ��fw�)��ɚh��̲t�KR�/�Ґ#���M�:��ы�>�A��1 @L�wI��]�ҧh���A��a�� ��M1=����]�7D@�m�qO�>*VKU�029�G�a[bL"}b��5����D�<9w-#\E���&:�-W$a���q2��,��u�"�2qO�� �`�ڕ�С-���$V%SVrPJ��& 	�!+�:�џ\�ai�+�����3���Y�����RC� ``"O��k�������#A�Y�t�J�@�"O���#�M���� �����[�"OJTH���%Z��V+d�8d1"O$� ik%|�@]�h��T��D�<���/�N�ɠL�'V�0k���^�<�B�9fXx�b�>��D��K_�<鲯��5f���^����qR�SW�<����m��Qр� a�����FUN�<aF���E��ؙFoC�1���[R�^�<�G�4`�l̠�o�c0��B1Js�<q)U�l�D�P�m
�pw��:�Øo�<���$c�z}�b�۾`)HXF��q�<��&U�n;d	Р�־a��0�w��[�<	f��o	Fqc��8e�;�$W�<A�#�@=9W"�z[��GN�<�Dˌ�Q� �xn��]�=b��D�<I��ݎ&����EB�lS*�+W~�<a6m�94V}Sg�N�~����y�<����W�� �0O��2��A��x�<	�
9�H�! � G�a�n�{�<�aj�%q�,Er��P�9�χv�<��ϖ�?�ja:��^�.�V�X�`�r�<	�aǑQ7*l�`
�!H�&En�<	Ь�Xr���t�B�Z��@Rg�<�������qz�'\���@z��
W�<�w�<�Nt#i�T:�xj�i�<)�
�X̐ɨŇ�bפU���e�<1���)"� i�a�*�v�H�ma�<�b>'�j����]~���T/�F�<1�oM7 �r�@I��|@�� �M�<I��� p"��.��H� j�	w�<�BC��|jV�2W�^�P 1���K�<�G�y�m�vh�?<_h�Dj�~�<'Gl��6 ��u>�x0l{�<���?a��R*�8#�T�e-�~�<�	��`4���'̵yɰ����Xx�<Y��'�v�+$i,s�hB���u�<a7�]�T���3D��*Zl��Yd�<1�K�l�(lʆJ�4{�"��`��i�<�bbÍ�Y+��S����h�A�<1 ��*Sr&E1�:\��ǝm�!��U�P�V�_�{G�m9�c�2+�!��7d�ȉ�u�1a�|��MR$!}!�d�zYx�`�L	"dA#�̒�d!��_I�V%J�M��4�C��[�}�!�$�<�ܪ�B2�T���k�!���X|YɆ�8!`*�j��!�V.~�0��63:���h�3H�!��1R���M4(�F��,�$"!�� ��)s�U�e�e:�&;̸�{6"O4����H�m���RA��8���P"O*�H#�`��8YA.�e*Hk�"O��#�`��f���N�4���@"O��%�O"j�1(�[�w�X���"OX���E�ub�Ae�ՆE�l���"ON����S|��У�M+j@*I"O�x+� D�;5�x�7��+rFl݈p"O ��eܮa�	� W�;JN�b�"OL�"�;h 	c�IB�Z�0�B"Ol�[/ֹ ��@*G �=f�c2"O(u�n��l�c�'˥ *�cC"O<�
�D��<��cE��8VXK�"OX�0��?.�ΐ3�E�'_2�Y@"Odm���]8I�y�ыF�
�l�`u"OHtJ�
��;�ة�B�*���S��,�si�gTqO>�Cl�0<eP�p!��+d5P�`0D��������iHd���XA2Ǌ;��E�RU�;OV첁*�+���&n��3�B]�dl�.��A���Z��H"�׌VGN�袡��@�i��+/��u9$D�/џd�݃��$���O��hR$߁%� �pB�O�H�@�X��ɓ ��@}�O�F�8 �R�T�ai�9ol$0�J>�A�F�lk*,�B�T	����1	�D�t�B�!0���R�IcdT���db���B��>E�Dc\��<ڲ���\"���D>�}ѐˢ��DW(�?�'�n�Q�G��YS�(	�&�YX��>AB`�*�4��՟��Oj��UC�H����݉h}�0�bfZ�6�>}2���-�ƭئǏCX�t�`�(r� �5 ���X2�mZ�N��I�s�Ƀ]"		%"ۢa�'O�"��KM8)���B$L�.��'2N�\������4i��Z
M���E~�E¦:Ax8x��{�#@r~x��
E�&-8*œD���ɇp]�h��2�@	4���Cwz�'I	Ɛb��ѻ��4�R.:,�x�ԏ2;���������������ƽ4�~ҧ�O���kN� b�@S5��9L����0��z���h��M6V����Ȼ������g�D�3�d!�)�@�ֺi��y"�+�r�pmQN���$fֲ"���Zw�i��+\�@�<��	;o��kX ^�P��$%M\:"m�q�	V�D���E�MU�l�2,OB��+�7�jh�����r-ZRöv�4C��&��=rѬ֡#?>x{�5�n1 R+ �z9r���t�6��b�xdAT��X�WLJ�(��?�Q�ЄSXp�"��h�4� 5k�ʔ)!�n9��Ғw�����3�T�j��>9A'H$"uD_/A-tb�>	��^�X��=��ʶ3��=O荚��]#��d3K�b?����M�" pt9%�\�fP MާL�B���@�Q��!x��U�t�TI8��K%�F��`Q!e��+FN��Y��<�eԐy�1�O ����/-���C����g�>W�f����׈t�℟�eHf��"�ˉ9�{�$V>-嶀���F&}�R�*�!Z���0Q�C�dp`�Tl ��T-i.�I�?�Z=yզPm�'x���%V.�ys�EԖ>ȉDzb΄�nn��r��W�'1���it�U2,��(�ê�����'��iQ���R�Ĥ�W%.񩏳��)�z�@��<:R���Vɶ�m���Q��@��S�O��\Y����48��#��<LL�	3@${ӣ`���*�ŏ����q	�	�NdڂO�>�Ǆ�M'Tp&b�>�CG�$ihd2I>���H0"MB1ȕ��sN,���U>��>I`�]�zf�11��\I⨲#*K:1�4�����^�l�,����`j*�)§y�V�#�/שN]�E��C�9~���Fz�%�I�֡��K�g�'M��!�#�Ϩn�~��6�C�	�t��/��[��+����2.N?`ɰ$n�1p��`��ԳZP�S��M{��0}iCǘ�O!�e�'i[u�<iաؐ+(tXX%!ؔ���'k�l}�CB+˲��wxx���gi_a
8!ÀE� 4H�qU�*�Oj�ڃJP]�&�#�/�ep�PP��ZА �Pj���yG�TXܥ�=E��*@!BϘ[b�\z�PM��	1�hOJ�* (�2dƔ"|b'�'?����������91�V~~��ɼr &	sc�'7��g�Y�TE"ա6��/_�ȕП'���Yud]�S�ӯw�F���?4��� ���Xк�,�{���POF��(Ē C�2�� m@�Y�퉶{�Z$I������Gl�1gl���ԥջs+�E�@"O.�ñ.,G�>y��ώ�f&Q�W�R<�(�"�m�	��𕧈�BB	lOԍ�բ��M`��yb-ٱ8�q�&�vL��%JŞ�y� �Od,� 7�:R�P��� &�ɴ�L�\�ݺQD�(����'D ]�*X�>ԙ������I7o��CN�i��ݒݴy��PU�@ǃ�;r�,�pm��4d�A�?�F�0M���!�%ss�b?�%*X�\ab��׍]�c?T=�p`$D�y�H?9!򤊃%�:Q��y�$�DA���+;^����O�}�V���$�$vƴ�(V�*˔T�ȓ��l���<�AIE�U5'�ژ�ٴ,�l�r'_�+�"����W5џtj�Q25�ʜ�fQ�����
 |O��(E�Z�I�`B��Q!Y����&�>y?�I�ƪ�D��	�ui�.�?�t�%}�%��5"лp� N�{�1����I���l2~o��N�S�V+��� A�rH�pr�'Y2��f��k[�-�7`E+%ž6d�6��P@%�˼`��8�X$R�>�I�Ic��`Tqm��"ckIs�B䉌$���AL3b��0s�X8_�v�x@��\�sfA�0���Ռ�Q��k�@�L��X�b�sj�i8|O�l��',\���Sr����6.ǤV�t���GS%���e,�8o�xD��	���`����L���b�m	��$JR���68�*�@�z���ď�/�h��.�/�i(�?�yfE�V��=��C�yf�Hatf�
dX��N]�J?�8���Detй���O���a��! b�9T�I��ih�"O�q�K�CpD���Ï̀`3� q�r�S�H
�i�1 Y�nB F�jޟ2�X=Y���M1@����O���=�4�\j���J^�3rVA����V�s�D^�4�H'���x2��� n��M!��!r���IjMEx"�B,+�F]*���-N���CD�+_	��ׇ�m�C��7Q�J�1&.�,� )>f��|���b�@�"~�	�1�>	Z׋�V�505�ɟw$RB�	> ��2��H����`B�ɢ0)��k���v�u!N@B��5[��p�U�Qz�P8����	�nB�I�L,)bDkA?�=��W���ye��;�ZI;�!5�Iz�"��yB�¼}����T�*s0� ��yV*����=�|��Ԯ+q4��O���M�/Ϙ$�wU32�T���"OH��"�C�6L�E��'@����5�i]�l��&��I1\P�DH��z��&�b>q˶�Ԡ@c��Qk�A.N�I�1\Opܲ��P
PgX}I�'�|x�(V7f21��O=]�!X��I�`�'��Qs���>IQJF)siɳ�$U7z�~�X`�	gܓe�~�Q�R�Q6N�}:�K�Kz�8���O�1Z=���O����hi���d͝�x4�rfڇm[�y����	���9�͆.e�T ˧2�0D�RN�FUT� x��� �� �4;j-`���K�4�0�R��L5if�Up��ű4m��_6u8�nTd�J�x���I�铧�O؂�ɗ�X!-�)��M~)��דAOX�� ����)dd�Kbf�<EH��B�+N��"��Q���	U�l���O^�"3�GKjN�Q�"�@Bv�p��P!"�NRw��h���r��`����O2B#Ȕ�3�8#_�1X�j�>ѢΒ���b$]�Zä����/.�"E�� ^���	O�!���"F�ܷ��$]�-���8`��|<h�OS��!�D�G[�8E��Q@*�vě9$��(˃�8�"
bՄlǄ�J�)�SUe| FD�xJxL�ECI(<���$��d�hr�O8�yb�M�&w�����=i��Zw��/��a�{K����A�N]��`T5De���"�ĉoiqO�D!�E�15�Z���ǩ(hP��C�e�P���˖�TB!�E�'	f�ZR;�l�3�K��L4R �)'��	ȣ|�'�)��b�8�m��"R�!��'&�8�'�lJ�I���O7��` � pJ}�$ޅ�0>)��e;��R��!>�~Z�#�o}������=�ӁA�젛�(�V��J&<��ͩf��ᔭT��!���'G� }���̶:G>8�C�?��mw�hH�ǖ�4t&�ȤhPd~��,-c�?F�I$
���8����3�8��d^t����P�K$��%��e[�\��r",�=d� ql��X���'��a��$)��<A�/V��xq�ŗ���|K2�Y�'j��ja�-j���}�v��	����� �u&�|�$aЦ�bv���J ���$lO�����0ݲ��S ZGlxZs1O�t p��.M�4�M�ʧ|��Z�CR|t7� ����5h9`c�,�9MH`F�|�l��8O
L��I@T��a%s͈	Q,R�y�4�'�9sR�Y�a�"Y����52��M��i�P�j�H��%+W�.���dVM�)Rd��y8�<)��"�t��e��$F���5��3D�#�S�H+�؛��I�5��x��$06�±�O�e�R�B�;�ft�vʗ7-��|�/^���ONM0�G�h�@���KY/
��!��n�.-�q!'j�?��)!<�Fɉ���2@~ĥ³%�u�ӯ. �\B��4x��m]�i\�I�"h��Æ
x��S���<k��Q���צ)�U�Zb��Y�	�4��\Ò5}��ҍlZ��^�T��$Ұ'v��3\���sqZ�>ņ\��Od��g���Uu��r���%t��O��Rc�3 z�q2���!XY��a�+Vf@k3cܦA�a|"C��8rFB��xꬨp�Q�K7�SB�E"!�t���N
��'r��3��D�&�hT�O�|�ge������C�Td�Qᐡ��O�Ha�/
�8�Hc?1�R	�,q��jQe�R�p������0$�Q�b0���>E�$*�70��:�"N�8::d"�lW���dU�s��ى{���z�3�K,!���W��5y��X@4mwNi�*��ݣ)[�AZ�[�*�,���B;aZ(�Sdŋ�+5i�"L�=��rD�C	Mے�B
On��T��:�fYZ�NA�7�J�p��	1s�\�u��.R}V�B鈿o�x�o���y���6s��#�a�La&g�9�y"C�*��H�dɆ_���K��2�y��FxZ�{ �ZA�0iY�dŚ�yRL��L<�̹�`�&r�|I���O�y�IL#}]Rd��cm�eȆ���yRET)/�̚�;/.h���K��y�B�'��A���	7����k �y�'�*MU�̠�$�D�H���y�Ɇ7_".��*ǁ ���`aҴ�y�fܰ!Z�#WZ+jV ���Ѱ�y�FI=t6�$"���%��͊�C8�ybQ�(q~���F�-I���PM��y�JX;ۀ��M�(��s��y"G��;nZ\Ӑ%� t)B���N��y�
�>@���YP�q����EoT��yR��7ʴ�p�ޫA���W��y�fO�ư ��Ύ":����±�y��5����v� �f��@���y�D����}�ӂ�H��IR���+�y��N�0HPP6��M
d� �.�y��P�����W+<&�hS��R9�yRd�Q��Q���,IX��5��yb*��JU�V�t;*��'��%N8vB�I)P��U3��~��D�R�_� B�I(Nz��Cu�3.re�C�1O�LB�ɪ0�p�J���>!�(iZ&EO9TB�Ʉ*����CE=iQ-"�J�ZB䉚pl
,��E��@�F��NWRB�	#7	��� sצ�S�Ʒl�VB�I�;�|1BkY� ����E
B䉢=C�[W��`��%v��d˸
 
Y8��g]�P�df����0�cĥ�!�DB�H�	��[�<���YE‒�!�dP	(�#��+v�fJ��
	!=!��2����Tʑ;,4��t�X�!�!�P%>��A�#MU�l Y�Ƥ�!��� �9��\/x^lp��Q�0b!��\�����ҹ5J����?LP!��%|E��+RF HZ�B�>��|BH%}�?w�d��Rh�s� ������J�{�m�?)�t�8�.���*�q	ç0��belN,���F�,X��,�C�V�dD�Ԣލm�"Ɋ��ºێ��޼F -�b�ϧ
6�X�ʉ�-��c�!�".g�x�`c�m�����~�)��2�9[CH��31��F��S�(9�'����wL[-O�L-���)g�|K4�OrM�')J8��ٔ8O�����x�0T��#�[}���M>y9:xB�
t��}H�C�"H����� 'E�Hר�G}
�g�? ��J��N��-��C{��l�"�/$���I�+�B}�E-�0|ʒ#�n�f�s�'@���2��p��g��i}"�YW�
��)d>]���I�3�$��7��+#K^C�o��(��poڤ>��O��G���u֒���GĐ����a��r�^5Qw9�S�O�R1�NT�Q��ÈU�
d��'gq`�d�	�l���i��P��OL��d�U����6#��t`U�Ԅ8�!�K6e.9U�.�ҹ�!CO�!���=�<����^�Za��1e!�dX�}[��'�]d�&�1�j2pH!������ш�	����
A�aI!�$�5[0�tU�(v6ě�鈅j3!�$͙n�H�瘉 jLc���R!�R']���(�W$}��]Kvi�T�!���pPl0I��_�= ��+�!��';&z�FGV"g��@X�%S	�'����ɢS��)�`E:��=9
�'z�}����3���0!��}oL�k�'�vc����ب����G�f��'�8E	��?��
ǋ��B��p
�'���9aAI�I��,�fϞ3���	�'`p���ŕ\�5
�Ǆ�%�Hr
�'\y�&υQں����^ L�Ƒ�	�'┑���
n-��k��\96�l�:�'iN`	DT0�%$� Ƅ�c�'*�u#���3G��d�\1Z9��I�'Y
��#h��nU���Mt���'��1�Y0�vQ�����&�Q�'�=��a��H%�4[a�T�*�
�'w�	��̙�R�A��DN"�v��'д��!ꖎ��) �0rܐH�'�|��T��d�+�&��S@ы�G&D��z�	��j��`��
	��mi�i)D���C���\�|1�Q*��u��)��(D��9��rp�50��� l����A�(D��h�*ީ��0�.
�{��ү&D�T�W�<!z0���Z��E[n)D���aH�,sx�m� ڷM�n��e:D�81Q�]\���-Y�,K"�eC#D���q��xc$�$�K�QJ&H#E?D����I�&vܔI����h�U+�, D���v���)7<(��M*I� ��2�?D�8c�Q��
�1͐�t��aj�l>D���-��d���#���6�p�p�0D����FܑOH�qڷ+L&P�#�.D��)��6=���Y�D��3�f0�k-D���vB�i��^$.o4���A+D� "�dI��Z�0�l����x`B3D�����޴89~�� �cC�I�(��:cQ�*�����&X�Zd*C�/:p��ۥM�6Q��P��T? ,RC�IHy4�B���r��{㥅�(XB�	FI~0���F�*'B���O���B�	�Q����0C��8:b��s��G��B������A>b�T���8�� �ȓPc�5��E�9)ހ��!C�;��q�ȓO�dpآ���P��䈱�:��H�ȓY0�FV`t�P4�X1g�nT������gǑ&wt��*A�)U�����6jr�Q�d�n	��t��	�����i����4Ç^�2��T�GR�p�ȓW�*��iL�kZ�����n!�ȓH�a@G�-XX���O�y�̩��?נ=q�I`yBK?@N����S�? X�A�!��LW��(�Ȍ� �,(#�"OF��/^)��06n����h1g"O>d��F������R 3�l
"O�`��1^�cw-G�5m�Y"Ojms6`F��UTB�d4"6"O �3���=FM�BH��	��"O 1)0�K/�%8�hX=#�4�{�"O	��KJ4�,��&��(��"O�xq�k�+- @U��D) )��"O2����FH[&][���*�4�
1"O�d��L ![ ��B�/K�$r "O6E���2�Z�Js���02"Dx"O�l1��N.�@��
C*���"O 8�����b,�'T
�1��'r
��m�	d�P���S�&\3�'{T�	`gV�L24�0��2!��	�'� ��W�f
����[b��h�
�'�2<�����t�ኦeD!X�T��	�'�85��M�1g8Y��"WܼQ	�'&~��I=B|�09c�y�j���'�4�*��R�e��� @,�	�'J,ip5Z{�y�`�n n�9	�'\"P��W6\S`�\��>��'��4�W�I9bld{�'B��.�X
�'
:���Ŝ:��k�n^�6� )�	�'l�-�@�8�I1�I!,R�[	�'�� 3G��=m6P�u���*�\���fFuqs"#ԖHbr�_�"�e��zK���b����8
$͓8 z��ȓCb�e0EB�$$t,�v'B�k�9��"��9��:�b]����*z����ȓ'_���EW_}��*�&O��m��?璉��B(�$J��C�Y�N��ll�ɘKV�̠��#��G56��ȓZ�F� ��ag���E���-��x��k�	kF��	"@�DJ�bef��ȓ@�P��1�W�_�l)�� 6-=���ȓ�^����K��u10`A���Q��&���aO��W0��MJ�H
���S�&����!B��b�V� ����^izE" I'�1[�߉b'����Xb��g�3�c��VZŅȓP�$pQU�B-ڈqVAƁiS>C�	��4�mD�M�  ��Ο5.B�ɡd�B@h�߿BH4��PI�4x�C�ɞPq�a��YF��L�%v�B��(J��DR��ґj�*���+�$"�B�I:��$E�4�$eP��B&L�tC�I�=��� d�4֌�'AV�.HC���に�^Ҫ<��P�9�C䉨"�j�'b�]�l�1���P�B�	}���3���0V �yҭЍ/�
B�(a��rkJ�}���
�(��B�+{8|(Zo��@i�fo�C�!g��#�ʇaF�H3e�:a4�C�	;gSj P���F�r�
T����C�ɿ~?t�ct��<(N�	�F}��C�z*
9��"��3ユ�C�	7\���G
�bB��"끡)�C�I�E����ȍ�l�R��J��`C�&h"� D�� �bɁR�E�)�lB�#e�eW��8J���g_)V�C�I�F!�-y���(k�4m[����O��C䉎f�Z@Z��p q�W;q��B�)� �E��A�� �¤艑&�9��"O04+5�P�P� $�bV&["��[�"O~��"�1��Q�f��:*��B"OxÇ�O/�6(�'A�fFh#�"O5*V��hT
�S1aX4Sy
�"O��`�M�/k�LMB��K���ʶ"O0���K")Rlr4�@�	��T�$"O@�[p`�.��@�� �pYj�"O.d�F�55���Tᑈ�hH9S"Otp�M�;!���rf�l��a�r"OLT�6�å]��ŤX8[����"O�H{bgJ�m��œ_jT�*b"On�w�U <S�8Qt��xD�(�"O����.[b�2ؠpkK+�]9�"O�,ӕ�k�	H�(�#twB�C"Oh)�OL>$�X0"�I9w�=�D"O�}�2皏�j	�A]�5kJ��%"O�A��I%�x�e��E[2h��"Od}x�*^�o$T	"�cR#(>���"O"��#����T+f�Z�5P]�"O(�Bc�	�o���lX?5U�ڑ�%D�����r��5�T�
]�݃u,?D�t�dK!��aZԯŘl��Ix��2D��P፟�zv�h"6�	������0D��i�H��z\ڙ��+�,jlX�d�/D���W��(��qHP�
�P�Pȁ�*1D�Ċ�A�~ ��b���?;l���;D�p�3-fhd���	p�UIԂ>D�Ĳ�I�Y���k ���~1s�;D�PҕIV��4+ת9��b��8D��yT�N�aM��	����j$f5D�lR�k�Ju<���ݵZ�l0ٕ#9D����.�x��l�;^��r�"$D���DN�]�H��i܌5�Ju�q�!D�\�^",z�5�AN��1��Ar��"D�|s��D��2ْe3)	B��C�ɩys��Ɏw&�I��I�1s^C�	vY�B�,.2L� R��A��C�I�5L����Y�?�*e�ܒ�N�XC��6Pz�lB�t�$-:�)�M�JC�I)=�����ߐz����	��(C�	�vPb)E�%ɂ B�#�]S@C�I n��
��V�)��2NM%7k�B�I�I�n1 ��F���ˣ����B��)c�nmS�'J��a�MSj�B�I.h�d-�D�ٿ����)�C��B�I!ܤ���M��Ҩٵ��n�VC�	.�X��bh?�fq�Uȟ��:C�	�� l;|��4�4 lC����GQ�sc�S�*L�q�C�I�/����b� .t-{D�	9��B��;E`�j��]�� �d��Y��B�	�E0�v��2V�Y��dE�YĊB�I2
}^��`J
 �t8�b�v�bB�ZS&x�&E��E�� *6ET�a�^B�ɽ�N����:͐,�cR�/8�B�� b�rf�4D�h(��-��%c�B��M<����M- 6���gMG�B�ɜu�@T��
:a�\-�s-͐��B�ɮc��)���I�N}[��πg;�C䉳�a�Ư޼
ц|�*̈2'�B�	�f@�HK�^�&hCG/Z#�B�I���`D^A���A��2N|bB�Ʉof����tQ���pF�bhC�)� (�q�Y$m���dj�g�R��*Oj!x4h��Fh��ԧ�.mi��#�'����Q�=дȪtA�S�^�2�'G``�a�د7�Y`w��K��I!�'2RՓ�D��t�Ì�%?\�xY�'���뚬�Je�#)Y�<eJ���'�1��D�W�ppÂ�'l\��'��H�'/�{�(�CWN�k��D��'�p�BAA.�s�K:^N�S
�'}��h��M9
��4)�M�[=�q�
�'��P�� )-����(O4Y�Ĩ	�'��=P�"C>�v����:e��'(��24�D�x�l�zGA��b�� ��'�T��RʛJ\�����fL��'`��AT��kp�
D��"ci"D��'� �  ��