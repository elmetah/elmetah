MPQ    ��	    h�  h                                                                                 1>K=�<�?Y�����v$|7k��Gz��!8���'/�x��o�2R󄠻T�:�s[����
�}�8V:�^�&;5�H���< S�+B��M�� ����3L�lsg	�:�+�8�ZW��e��)���0��^k���P�D�+D=�P���ȮT�!��j
�E�gV&����2}�-�V$Iuϖ2�*0�R敿�������� �M���`�+\2���D��wS�����I3�ߒqR����X�J��2{ԹG��L&?d�G�l11�
��</0`M�oξ�u�m	<��hXÆܟ%8%E�4�-�ֲ��D��yy;e�bV�n�+&*h��Y4 �Xʬ�o��l�$��ܠǔn��6&�m�ve�Y��?�Z_;I�g�gE! Fc�ϓ��%H�A��i�m��{p/Y�+Q�E�sͮAFc�L���1�w�o��tMi��u����x���g����FP)=Ĳ����2��In��tA��;��sjL+�r��<��n�2S�v1��)a�WK@��1\�q�	t�槎�G_"�A��}��PUD�?��؝'|}�Zg�|^�
�6-Fy9��hq!J�K�粭�������=��+�#9	�F��{
#����$�ȸ�Ѷ��7
��D�U��((�a���u�?���s���j�T����͘�K��#n����I�d�z���n� �����h�z�=pO�����Y���vW�"�ٚ�O�o�5�9 d�)��Mބ���Zg��3��V|��P���n��~����ݽ]5I�p�x1l�W�'\3���(��}t���}��
b<���w�/W�%tɜp\_E��e��g+�%�C���?e	� �O7d}*Л�_ӑh|5�&�H4 �D�)T��m�������[��~�Yo:�QiS9mZ��?T���^4��Г���%���Qu����j�Zæ��%UX��s���/�U�y� ��lɶ����Wi�Z�a0���=UV����	A�*ߠ��a7�yNϛ���%:w��c�rjM#��F<�B�j~���-�KG�Ք�?��#L�����c�t�A˰�9�#�[�J�.��!�N�M���{Bo�S�Q�p����`��OQ4��j(%Op��{��Vnw� n�#��q[�f罨�MЧ@�̾x�;_�r�pO��w3Dc��ԏ�����X��F-G�@) ��b8�ի'���-��wE��n��.3���_�j���D39��(�34�����A����2�?���޿'���BRɲ�g�(�����!*�]C�#���O]N�վ��wS��ʩ� e�����W���x_m�CȀǾ�|ԺT�*��!�~��̊�^��7�r�U���$?30�8�p�al4����5ׂ�=5w����O��C�����7Eǫ9��E��Xcx�T���L�Nl�� *�t���J�^�y�7U{Յς�z��ZPDT�0���>��+��V��N��'�ڶz�>g��>Fe��5໊�*�\�0�\,
=��?y�u�q�ϓ?9f�1"c�fQ��*��	���x�#�|s<�v�����k]����R� ���Uz=/�[��u�`�l�,�x��^11sa8Q�/�Io��k[>G���K�)��pB.�a�ۧ��[xpG�z_����!�5�nq�~�*ASf�ޮ��o33Z�k>�5���n�f�!�_�NK"�)�!O��C�3�}���<-��݈��<.W�509U�����Hz�7��u�j[�b"a�]��n�>xq��F��}�C$���f$�"}���#4x�R*P�6Ώ�@�c@�5�Cٱͨw�/L/�y�d�#� ��o tOm�����t��D�>ڼ�u�C��}��P����}�$�桐����ME٦���&Ia�� Z\�6�ޱ�l�O��lO#��|k��������Eb��A��_3r���=�y�~�t��(����U�LEh���d�8�o�6�͖�Ǫ˭V}�N5�Z?���R�'�\t��M:�[��T����B��c��u.X��V�7*��X(�ƆV)u&09�����L?-yx�@���<kď��Zm�hY���'����v��$2Pe�a?�bǫ�g_�f�,2ܨ��Y��q�ݠ-mA)�b2�����M�=�k9�'��V:Ҡb"������a���Y&,�{�\�N�
i~�9QT���;��%�qݏEs�̀�EVo��NQE��3�/(:i v��%��C��{�����E;`� �^[�9J�<16CS�U�&hu����Я�<ng�/pI�����I�XS�~G��8����a*O�>"��rGN��,�M����QS/����o{�1s�ć��3G���
�	N�`+����t	��2/�Б���w�?��!�Q�J�\0�V�K7}H̱���%�U:U���&
o��Y-�i'b+Mn፬㈠%bz��ɽ�\�K�g�m2��+ �K�����G��,_N�N�uc�[�K���1���U��͠��ot���Q��>�e���4�s�Fe��x!��tm������%���:��9��b�j���p˖7���h�p�@�dBL�������{-b_��L�JG����V�{W���O���۠��=v{P%űL��<3��mF���m˳1Ҳ�O!�B]nq�B��GB��ũ-O�<�=2�.q��hy�-0} Gp���r�4"���_]��C{�vH�֬�g�@(1i4$s����	�q
�i�c֋d�^݄��C�I0�8�Ғڟ�Fg�"��Zzؐ�����ݛ�KU�w�� hJ�@�(H5�22S�.�a��_/H E$#��~k�=I���A=�c��6s%�����!��7��]�w�n�Y���hL�gW�mL�D�c-���?k�"!��^b��u�u+���cZb��`Y5�`��Ԙ}^Cz9!\���;��Y�i�O ��3���@-O`�1$Gđ4=@���/�/���LL� ��[��B�w6��i�l����d;�H2�i	���?k�7S�����ͻ���o-���}	��W0ыV o�Ӵ'2��	1s7�9���LN���e�d#�T�Ճ��l4$��l%۝~"���uz׻������|�u���gj�,���̢�de�z5���G��&��6�E	�t�:��4� ߙ*=o)L���W,|���
@搁8�t�-���n�[$�M�[`�֦\��x���x��|��hb��%)��"R�Pw��jF�i������b��L��&��������8�s�ߔ$/��0��v!�uGm������IV%�-�8 �4D���E�_�y�h%�=3Lnأ�*B�Y/�����{�׌)����$aMD��ŏ��M���e˗��<�Z䥖��YE��oc���/�����d�r�{+c�Y4t�QdT�s��*F�*Q��m1�����k��2"i�7��(7�xe?�g�4)��{�=�QC�`5'2d��nZ7��;�ƅs��x�详*�ɟvS͡/1��)�K�*lY�s	o���`_Á�A�e���+`P0�\?�۝����Z0��]�
�!6F�{�����~NK#�X�Fh��z뼘�Q+w�r	�sO\Lx#����A�@��
X�g>��7�n&����ý(am/��u�{Y�JÏVN��"E)���u��&�.#��A��b�_�,�ok�)����S���Q��}Ҋ6D���&W?���z$�j�-���� ޏ��d�sM��o�ʹ�gݞ��q������K�,�Y+M�6�,]ТDp��lN�e����;s�sӣ�0�(b�K����I/vl��T�ɷ�\�<"���`ǢSd%�sx��?�?l�b��ݔ�j�'}�R��O�̛\5!�iH/�vD5�K��ƫ��F��{��6�Z~�:���iN����.��7F��4�M8��!9��_B��u�tS�;jMɈ��U��s��F�jZzU ��$寋n��iًMa�`9��!�V�d�1%�A���J���yi���ah���kw6Q�՞#;M�����B�ݞ~̹q-#��K",׃
����Q��e��c@�A��9SYP[t/�.�&P��&L���JVoFyfQ�M��n`�C'O�����\%JL�H�I��V�?r{9�#u[��L�C@fТQ��d;���#C��3I��u�ªV���4Ϗ�y?Gxi);����L8�f�'�B��K&�}*�������.N?���1����3t������.�֤ ���{������!����魚sLbɭ�g 7��Q�����P��[�Os�]�/չ�Zw��4�d�QU�B}��2��2Q�m-#��O|/�8��;�<�8�z��� z��rD�i����?g�b�����,�Gl���ș׽�5�>���NOm3�������!���'��է����E���X^�%TF[�����i�B��Oη�.��J�Qy�6tֳ��=�U��;�DϺ\��7�3;7CM��IO�'4��z�s���
�e*m�����ٶ7�0�X,eqa�Ѧty�,�q3�fT�"���Q�
}�L���J�>H��Xd���懱��{	]��c�M[RJ������=�A�[�"c�����,���/�� s��Qۧ�I���k�EI>�G��)�����"��=a�>r�&"�p"�j_7נ��iE5��,��F*���f�,L2ɶ3�kyV��`���a;ܺ��Kݵ�) 7!�UC�r�!���{�����R��WK�R9p�$�^��HU��7�P6��]���b���>��������FC_Y�D���Q��#��m$�����-����۪ЍP٬PGw��/��WJƤ��d �l�[�mV�K������ǫ�w���v)�YQ=�+(qM��}�[�ẓ�0:��.��U�ѡg��5�;��э��P9Ox�'�����|�oN�ҏ���jE��F�<�T_� d�A�ӝ��-��lg�B_�U[��h�ghdw�l�*��I���ơˈET����Z����'A�ߠ�o�v�T6�������d���f�7���#�ơ��u����i%@�@,-`�@�k<��c�T�ȉ��n���{��mv�x�2�8a�4��,V�"V�3��,�]ڨp2�L���x^Cm<����b�s잶rMQ��k�Y�F����{]^�MӃ��!a���Y��{�M�N=�
n9L[�lpJ����q�x��k����o$���O&EȦ*�+�:ϥ�vӂ_%	�4C�R[{T ݝ[z�@ؚ�{�[�{r9e�K1���S�G�&�B��$�M��#��g>��I�um�U7�X.EG��ܥb\]⿙���PsN������J��2SjA̵n��,qf��+3���	�@}+����T�MH���ZR��_'?صM!�~�Ÿ0�����h}�L��Bȗ�MJ�i&%ŁՐr��Dp+��?�Gϳ� ��QRLx�f0����ֆ +�~T���5_�;}z
_�v��=�����S�tUl��͛��oώ�¤q�Y�_�`�=�U��P�e(�x`�tȆj�h���'7��V��-���zj�vЙkV�7x���#-�[�Id��W���J�)��-�a^�G�dG�~��֖/��8+z��=I��S�={�P �SLG�ǻ�~���	 �@�;��'����B�F�q�.uO����vu�H��<E�2�	��%\�qj}���%i�r��.�ۏ�]��{��k�t�f(,�$�s�Y�wq%m ixkH�?��^W�A]7I+�-����=�=<o��+�������6O�U��]�[2�J��(�5 ЁS�{E�OI/��� @��\k�fJI�� A��xcz 6���Q�!����˟wQ��Y:��l�Vh'�'W�k �ߒ�-{H�Ϛ�"�|^}��v\+� uc�kO�����[�\��@�C5h�!w� �;�΁L���껝�
B:�/Oi�1?8��I@�/�Nƍ��G����t����6�|>�� �~��;�r8�{��䤬��8��0�+���Os��A��G�K45ц��o�Bc'��	L%?����e�
�&NeI����l0x�'�P?�e��e�xη9��u�䈫�J�9���0~���ɧF��Zǋ����z�R�
��G��w��ץ�`|�td��a��ԋ�=
����LUW��x�Y�`��i��݊�{Gp떐�M.O�`�=^\�˺¥�����õ!�Ua�R%����� �cר��}��L�U��t�����}~�ڑ�/�x���x� ��m� ۋ������ %Ob�8�64�{�L�x�z�!yo���0Bn<]*���Y*]���������i$��w�}�k��\��~e���MZ�Zլf��j3Eǅc�Uțjb�w[3_�s^b�{�vYO?�Q߂�s���F����1�β�%S����i��v���)x@�Vg��|��=�5߻�P2T@n"�A7hf;��s�ʚը�m�0��$i�S���1,�)W�EK��y���ڧ(}	jF�D�y_~�A���s�vPx>?<��]u��z��2}�
q,cF�ݿ�^����=K^�2��_��d��'F+2/�	��<�#q�s�|���8m���kko7�2�A.��K��(��j��uFIk�����a���tD�͎���)#䒆�"�ҘZ���6S������^Z���Q��Z�F������W����<r�y3�+�w �;e�M7۲�śHg8�պ,�b�������4���q"�]kp���l�-t۝�޹�
F���A�~��@eBbr0���G1/���盷���Vk\:�؛�	�ݛ"%0���ق2?ǉ����b΅a�}��o�!��5�{(H*�D����_?����.��D��?~.�:߻iI��?��;v�'^�4,x���t�#���0��u�^� jX�2|4UN�s� T���Q� �|}3$�)��i��a&�$��%9V$�2̋�A=�V|h��`�y�'x� R�yc�wq��9��M�<��dUB��~��-��K��;�K���u44�̏�ur�c��sA�v9ή�[O4�."ǲ���A��P o�DQ�JV����`t�O�j��Jo�%E��ǣ���V�'��$�#Po[��&�޽vН�#�t��;�0��>~3X3�N�(7��E?���0"����G3�j)V`B�tc8w�'%хc�|�x�J�R@!�S.i���U����t�3�c4�O�:�)8`�{`^�x�2;��5�����5̹�v�ɨ@g[pm����t���g!��`3]�)մ'�w	���t6��*��.YmI�m�"\����|�?]�9��W����X�g�K|r�
���o�?������G�nl*��{�����5�����O�۔��]�
8��-B��x3��2��EI. XY �T�.2Ò]��)����ǻ*�7�i�J���y�U�1�C��Q���<�DJ�����g�njJ�c!�D9�'�	z[������e��Ӄ�ٻ 7�?�0�B�,��ϛ���y��q��"���f�Y�"��pQ��k阮f�J�q�Y
"r^8��O;��R��\^]�8d�]�dR�؎̏�=%��[f����(��b������ps�BiQ�?Ie��k�P�>�r	���.)����&#����a��D���p�?�_rH�W�5���41*�`Nf����)3���k�Ҍ��Ԡ�\}��L�K��e);v�!E�3C�+ ���r�F�A	���WoY9�� ��u�H0T�7 �ꕠ��X)�S�q�e>���<��t!C��-���\��´Lk#����>f�,ih�:��0���k=٧�w<j/p��0O?�>� k$���Fm���0ه��x�2�l�f���D���{�E'}E����󒌋��������0g����p��v̍�l~>��T�OӘ����T0|a���H�3g�EJ�ʽ7|d_�m�����W�tV2����}>U���h�id�Y���p�9����cT���ZZuE����|'rE��[M����LT�?���Xu�ـ�G?���b7�/��=�Ƽ�u{n�D���{,�-�g�@|f�<!Yx��h�������^��v�2�*�a���`��N��N�T,	�ĨK�P���S�<Qm7��ʏb�/^��GM�Jik�O����pCoX�,x(��A@a�6Y�O{a^�Nx3
�Ł9G����v�g��q�Qi�V���'o=[ ̈́n�EØ}��\�:��v�v"%�]VC���{�G]�8��;�Q��_{[{c�9�~�1,�lSlY{&ޏ�⿮$����~+g���I�?���D�X	�G�K���v�W�1��f�tN�N@D�CK�]_dS��*�	���'���=�33����*�	D�+��K1��}���C��=h�?��?!����@��0t�h�	d}~�n��������e��&@;1��=��|+�VR����@ǜ�f�EX遑��cw�3����/���7�_ŋ5�>��Q����o�FX��,FUj�͖}o*C��_�T�t ����s��%e�^^x@�t#f��X3��J ���cۼBZ�?�wjR.c�f�7�����m-�v�Td8���aWM�dL�-���Bq[GQEC�a��ֱ'���&a����?=��P'�L�-.���ؙ����ڷ���,�ţ�B�?Iq�:V�>�ǐmɩc�p<�@_��{>�B�1��}�Ա�frk���H�]�p�{�._�L[�p�('�G$)U0� q@�i�&��r^SI�ܖ�I&{S爋L�JV�X˜P?�oLj(����>U��W��i�J}��C�x5{�}S{踋�Q�.� ;
���t�k~�I�O�A3��cU�6�+��,��!�Z��oX�w�gYUm��� �haWW�(�zx�-v�l����"�C�^�َkO+fn�cДcŖ�O�V6 �N$C��!�@H{��;��Y��kʅw��q��^=�O�BM1ZIoć}-@�Q�/�C�+�>B�X�<����~�6�x{�b��YXM;�2���z�Z����j�k�F{e��=O㢰�,���0�сV�oU�1'�v�	g��/�@��
��e������ء���Zr�bƺ�S>�tbu�\刦�e����������"���5���1VzO���jGT�H����{1t�(��& �
=�Zյ��W�ҕ�8%��]Õj�V�!���M�bp`��Q\C���u����.���aÐ=����R�-8���"[l
�cQ���)VL�e�ȝ;���`ng�ծh/A5��N�Ӿ;�GmzC'�a^��7��%�i8�u4�b ������y�#���LhnN�F*9�Y%ѕ�i�ٯM(H����$W�w�X�b�3 ��>�Fe�s[��CZ�����j�E�ʇct�
��0����Zq�ʋ{�*�Yj*�QZ�s^��F����1��zπ�`�?�i��3�J�x��gQݼ�3�=��b��:2��an=���L;���s���C�!��+�R�SC�M1G��)�_K�����Bj�	e�ѧ�Ӓ_9�'At��� P�A0?w���!X�������
,W�F�_6��a��H]K��@�|w���oռN�z+��	,.xRM�#L�;���������� �7;s$\�,��Z�(�����Tu�6u�lV���⅙(_�2�	�u�܎�#�_���јUt�%"��o�����K���r+Ε�n�l�@��!;W�)E�񠒁��� ����DM�	N���Ig����<����*�A�o�����t�]�Op�l���X㺹���i���Y�Ʀ{�yb5���ߴ/,{��V:d��0e\�W��vl��%�2?���_?"L֒Q�tΠ&}�ћJ{�Bb5WV�H%*D�[�ز�
����«쭔~it�:�$�iD�nk�пp_*�B��4~*İa�@�^R9��I�u����&fj� �M�U�T�s����$�l� �`ڡX���QiNa�i\��IcV_��g�Ah�߱g��%�y���v ��T2�w��j���DM�W)B=]~(v-1 K�����T������U��ac��uA�9I$k[*YI.]�I��q�b�� k?o�$gQh��uqG`O�,O6���z%@8	����t�V�/Bq0m#+�[4�t�y[И�?��i1;��C1�B���3�t�c)��GC�L��W�DG��)q>��}�8R�_'`�A���ş���H�P.��d�������f3�Z��c�$�E��Q�r�)�M���2��4�pι����ɣ�'g��(.�f���]9���m�]ҺկoOwd���FnQE.�8������a�mcB�����|���[���r��p���B0���A�rz�\��M�?���ih�b!~l�V�oN��3%5Hw���O#��t1��%�7����S�4�m5E�%XTt�T�!2�Mj[��_R�8�ػ h��	=JSa�y��f���ϳ;W��]�D�#��������1y��?C�'�Vz="�ae lf�ƛ��;n�m�0��,:>�G��y���q����;�fʾ�"4��Q*��&E�@$�t�%탸��$��'é��k]�� ����R�\��\�=�$[A.��(��Ѷ�fB� sI�Q��I�S�k�{�>��?�;6)���ǁC�_$a	e��p��_��!���5�r�׏|�*ref�(�(L�3�||k�nF͖���W"�p�[KS�)V�e!�3^C~W�.P>�y���ӟ��W�;D9�_E�T]�H+�7;���;�SIǯn*,C>�����!O��C�f�7�\��ϴ�b�#e���x�����ag-�k\���٢��w�6Y/+c�Kt���d F��э@m���徾��UB���C�v��OXA����#�}�G���L���
O�~p��+Mї-�KCGƱ������x�O.<����:|ܢ���!��n[�E�t��2k�_D}7��.���(y��J��|Tv�={U��\h���d-StӠ��T�婏%��>�Ҟ���Z��⁅'�i������K@T,���2���F����7;hh��xJ�׬�u�P��˶L�-J�~@w�%<|�̫�KL��p_��ᇣ9��vU��2!��aj��sW˷��p�i>�,���&�����r��9Wm2�x:�bcT���MGEk��n����zS6��#C����a&2�Y��K{<�?N�
:��9B�e�"���"��q.�C����yHox�<��\E��,�@�;:E�v	�M%���C}@�{ʩ��ӎ��6r��1�	[6k*9�}1��kSG�V&���ZÓ~7��ҡg��I�)a�Kr[X���G6������R#=�O9[/l�N.|����8��S�'ݵ����"�JĘ��3x0���	��z+ZKI���G���6��L����I?N��!�Rﴻ��0O�|���}�����a�f�� j�&[�Ն��a�+���}���ǜ����޿Tugf��^��a��\__nz����Ό3|{�%����U�k͑9�o�[����W�VR\��Hp$��e^ˤx@t~er���)���kۗwD�zs�j���a�S7.W��qё(d�]��<7�ϟ'�-3ǚ�=.G��h��P��?g�.B4��3F�Q G=G��P��L���mv�����6A@�� ��B.Xq�fS�I�K���~�k<;򷸿\��}�=�X�}�ˬ���r&���"]m+{s�"��b�8_�("O�$�V<��/�q[ջin�p���^�[�w�7I!�����szR��v�J.Hc 3�l�U����+J8�x�^��5�j%SVu\��y%�0^N 6-����k9�/I յA�Ϊc0P~6$_��f�!�H����w�`Yp���b�Mh�C�WQ�ĵ~�-q��P��"R'f^�4"��M+A��c��1K�Q��ԩ'�C�%�!��&��1;s ��7�� SY� �h��k
O�<�1uzS�җ@x5�/G픍�A�=�~����s	6� ��?4�;Y'!�:���u���H�%���a���E(���/�g} ��M�|�o�� 'ck	��F��"��E�e���e��ҝWuO1��F@�.����fuKO���A]����t�`�ɝ������Fz��� ��G�ߙ�</�tZ]����J��=@#>���<W=.S�������D��ɳ1I���&Md�y`�k�\�	��0FL��^��p�ky�˯/R[���`����.ﹳ�NL]��x"ڷXz	q�����/�܂	N3�V2�m����<�y�rQ�%�+�8�P4Uj\�½΁�!0ye�n�Ή�n��d*Ԁ�Y �����h������$�vC�3t��n����e�� ZK��ӊ�E�ucO[��������U�jS�{\��Y�5�Q�?Ds9�EFO��U��1�_�ۙˇ�.yi���x���g��Ų�:=����qp�2��GnX�/-Q;j"�sV�Z�ޟ-蠤���[�S�߲1b��)MQ�K�&������	`P���_�`gA:+��i�GP�+2?��\���{�4��1
�)F�U�TG��ݬK�肭�Y���d���+���	G�8�}�#'�S��P��n�F���!�D7��w�I�A�^(��0��-u|Dw�-��g�Y�@�`zPḧ́hW�$�#ZͅXl�P 씀-cZ��3]��T]������1K�����x�WP<  Z���!L� o��jjMmXAŻ��g�b������!
��L3��&���2]�o	p�ll_&�����(	���?�40���?�b�Yd�{��/�2���Q�+\	���QY��S�;%f�6��hI?}.��λ#}��i�%�$�}��5�P.H x�DF�s�Ր̑%W�|�-���Y~�m:Q�i?ݼ�0�+�b�]�04�H�<������f�u����kj~ձ�h��UD�=sh2�ٟK� ��~50M��?�i*�ia��b�]V�B��cA���E�M
:y�����i�/!�w�O��o�}M`w��B��S~��-�{;K��4��)���̷�+q�cq��A79�9Ĺ�[��.�g�}��=��[��ow��Q����Qf`*�'O=!����%;�I�YQ�z��V�W��[6#��[o6��ГDX�*�W;KH<L�Nt i3���/�{p	���K7G�[)�<8���8-٦'�g�����n�@�����G.��1�K�I�`�3%r���b����1cv-�'�hë�+�^c{�ޫ�D)cɞZ�gZ���g^��'�8+�� �g]���ժ׳w�x�ʕ��l�������G���m��Ѐ�ʵ|@Df��ɍ#���V�x����Rr@���K�?xh:�$���}�ul ���JA��ns�5�6��BO~��/%s�@�΍#���.OS㨎�EcXO�TW5�������D�����HH��m&J�L�y~�9��nE~���D@���e�ѯ�(���:m�'E��z��(�/:e�e��:��v��
0�4,vά��+y�*q�������fD{"���Qz��]�C��������h�䘈u�bS��Lk1]�.���8R{7#�J�=��[��L?����{�p���0s�*Q,�I[/]k~�|>3�����5)~���܃RY�a$(��5p��_�����[5�^���*-�f�����3��k*+��1<��R����X�K{�)q�i!;��CY��iVҨ'�%��c��W|(9�����dH�!g7vg0���N�����$>�m��23@*E�CD��q���x�z�# �:���"��<���D窡��ٝ��w�x�/���f���� !�J��m'N��l,���3ڨ�~�K�ʋ�㼰��!1}{ϐ�Ņ�A�5�9��G;����&�(����������O���XJ��A�|Wl�c��odE�|�-z8_�k��r����8�j_ �W����\�U,�h��~d�lH�[;�o}%�
���y�:�Z����&
'(�����(���T�tЮ,y�O˃�����V�7����D����^uFT���f��w-���@r�<�ma��1t����
"@��v��T2�o�a	p>����S���Ə,��]����+�IWUm-�:��bΞ�M��,k�{Q��I��4�N�9.?k��-�aA�GY�s{�kN��
ՌQ9=0h�}���ݬ.qI�}_��\u9o�)Mͺ|E��7��: &v$��%z��CX�{,��nX��1o3�x�[�9���1"��S"�A&T�R����y�ޯ4�Hgo:�I4��ƿ�X���Gq\�3��M���+꩏NI
|�9\���S��?���+���c33��3�'	:�[+5�F��m�I��uB���?	Q�!�4�6�0*� 7\}�����X��G���H&v�����
X+9���R����b��}�d鷳��Y�~P���7.��OR�+z_�7I�����Iu�����$\���U=�͌�3o��Ր����~�Ѭ=ˠ�|_�Ue�W�x`�tل&��(��D�깁��r�^��cj����\��7�N��Ty�ѬO�d.N�7C��"�-�)��8��G�����w��}�s��ی�=⃝P	#LXN{�("ʙ�����Գ�i�;��Bɐ�q��l`����]��ǎ<��<��]̧�=g�i}���6��r�{�,s]���{Nf����m�(1�$�w(��|qv�5i�A'��*�^ɍ�j�I�^�>����ف�I�F�n�%06�=����U�� �l8�J�N)�yPJ5qhyS1"0� �n�˭� 1p��m�k��Iz�A)vc��6_���b!j!�V��%Ӈw���Y�m���'�h�FW�&յ��-ls�ϫ�z"+�^ί�a�X+��cFGH�����L^��K^Cf�!��,q�;Ny��>ʻN��.Z��)OLV�1���}FN@S9/�l��a��8���.�6+�-�X����;���Տ�p�:��$�����|�/��2_�6��{����w�JoQ/'�S	��F�%x���a��zeCY� �A���X^@�LC�X��	~X꘢u�ao���0�J�<�a���9Hu��X��w�P~�z�k���DG
0k���᱕�t�T��`߅oG=������W����������`�����G�nM��`�2�\�����ũ�`�x��F�!��1R��Y���o����*0��1�L�tj�S)���\���o��H�/����Ֆ�q�hmp�c��jí>�% ��8��4����}Я�ˋ3y�^ߛ��Dn�Ķ*o��Y�;�&8��Cw��g�$Mo۠|@��5�t�_e�ϊ^r^Z����1E�1Pc*��-�H|P`o�X{r]Y�`�QP�{sDoF��,��1�j_�6mև�m�i �%�ݴxѢGg�!�Mj�=�s��nN2PQ�ns��uK;E�Cs����y��蛎��5�FS�4�1}w)���K��X?��xMl	[ۧU\�_�@�AU���UP�5D?��.�7��m�C��
��F ���Lyh�,K9������导ǣ+c�	bh�H�(#C��-��	UF���|�?7�Tk��O��q(o��c{urq�ڏ�����ӥ��NE��x#��΅��K���X�}+�N�$�ώ������ۊ��H���?W����A���$���ȏ J��P�dMǌŶ`gI�ٺ]v��1eQ�7c��FO�"yr]<I;p�yyl�ҟ��2�C8�_�������$bC���vo�/�	(�̟c�#EQ\��N�,f$ǎ4�%r���?�0J��Te��}w4Λ oӸ�&5�kuH��D��볐iJ�@G!������S�~��N:� i:!�s���x�y4t�������Ā�#u�ľoj9���n�U�G�sC뜫V�t�� ������Z�"iE�a��=�'V�!��VA|�g���y՛�l��
0�w":��
*/M
�N��B�\�~8�-��K�SɃ�.�F�k�
���lc,��AR�&9?o6[�~.�g�U�w�8M���}o2PxQ:��kRQ`�rOx,��g?%6�fǴִ5�$V���g��#�?�[��l���xЎ�l̅��;�g0c�3� ��:������Ï'�GdbI)�Z�s��8�'�3@�4Z��i��c�N�h.��F��# �;H�3`��� �@��%�����.
���K>�$��2��߲Sə�gl����=┃��=��;�]U��ե_�w ��P�����.�Ӟ��Fm�ក�P|��J��Ҏɨ���fG����
���;r�
���i�?�E���Y�٘AUl�}��%Tש�(5~�έ�k�Oٔ���8p�[yn���"�	��~E��XJ��T�h�ÇD��+_�. ���؎��J�X9yyrIBm�)oi� D��@Ǿ��|�g��5��'�I�z���8{{e�σ|�V���p���0�! ,т���py
Iq��:���f@�"j4tQu����b�{����&�.��c.Z�����"�]����n�R6�.�W�=�C�[�a9�����3����ܠs���QG�[I�*kY1n>ne	�R6-)y	��7�c��a?��|cp�!�_#\�(��5�j4�Es;*��~f
�RO�3zޟke��̟�M���&%K���)�A�!�̗C4��A�C�x��|��c�W75�9܇�J��H�857�Y��q;vIx�$��%
>��E���CKA$�m&�	�]�r#���L���A�!:��LS�<�٘�wM��/��-�[���� �
G�0m����:��=!�c�����E���s;9@�}���^y��[�����-�1э!�����'讂=��� �O�����-g|�U]�>3����E̨�(��_�y�-�O� +?��	�2���.��U��$h���d���kv��yͩ����@�uhZF�҉��
'��ߌ�n����T"?�ЉF�� a|����$7�f;��M}�1u�[ɓ�x~�,�-�>�@m�<2(6�@7����p���ģ�~�v�es2WB�a���)�����n	,zK��݌�8���Km(���b�"̞"�GM=� k�Aģ2ˆA��I���z3�rԇa\Y�3�{�PHN)x'
p�98����I���*qd] ��7��o��1�U��E�.�����:�ةv?�%��CC3�={@�-�	Ba�,�^��4'[���9���1��S�N=&�7��L:t�h���g*:I1^��A-vX��2G�w��U�Hi��>��NdD����V�SV�>�������N�3���N�T	��(+���;���i鷾��NAl?��.!	���2w0�Tr5�}O�?���k��_�G0&�]0�|!���+t�����}}��A$8����tK��h�+/��r6�������_!�f�6�����)��xC��?�sU��t͇Io; �0��e��L'��{����e��x�t4���S8�_p̹�Ք�MA���s�j#l�W��7���/��Ǽ&d�^���V6�>�-i�7�3�gGb�Ӛ�Z�п�$ٞ�N���,�=}q�P��L�b��툙�U0�,nu�xߜ�v�Bd�q����o�������<1��u~���U���}�W��r�]	�G4,]Ɨ{)2��Кn�n(3$:���E�pq��id�I����^�e�I��px�{����8V�V� R4ٚ�ݢ��U�/����NJ�����*�5�yS�3�;*��f� ,�#��[�k��%I6?kA�c�76�%�����!��P����w=*}Y���X��h�i�WǤY�K�-glO���"�N`^�Jaܰo+�w�c���g���G"�_�nC!c%!�r[�(;)�8@6�Vj������o(	O�h1�<����P@.]c/����.�3hߧMF��l�6F-������d3;�[ڝp���k�d�����5���`�;]�t�^���	���9�r�[of@^'٦`	�-�����g�e�
���N�ǟ��m�i�ӧ���M.%d2u�����-������b�TP<ɓ� ��򐾋T�z 	��5�Ge������̈etP���{8X��PD=vX����W�D��E�K����ۣ����V낁jM�]4`��\Tv/˦I�*������!Q(�A~R�i��l�>הGU���wL�I�.Pv��^%?�Z����/R*��}���P�m�jT��sk��K%�t8�4�4�8����y[,���c�n��<*
��Y���z�G�~u�ݎ$ȇ?��'��)��e�����Z�S�	+�E�c�r�V[	��q�K�Q��{�E]Y���Q�|�s��(F��D�1��{ϑ`��p��i;[��֐x�ˢgJ���5�=�LU�'�x2;_n��=#��; ��s�Gk��M薘����St�)1���)CP3Kb�����V	V�����_j@�Ap���_0IPw_f?(W����:C��:$
]��F���Jr�Cg�KJ���M~���P��_��+Ə	}5�>�#��t�h'Ⲥ7�5�׀�7l�$�N=�7-�(J�8V�<u��c���Qⶼ\�v��zU?�m��#�d���`�FxM�6���3M�iY}�J�b�_�8�FJ �=� ���W	7v�R���e� %+)3M�U0űcug����C��L� ����àh�]+�]�B�p��bl��ۉ�g�^����m����,��b���qg�/=燂��>C\�o�������$%�AN���P?3S䒂�C��5�}�����Fh��{�5(��Ht�D�ĳKb,�[WB�r�ǫ}�4~��:��1i5oM|����_����4����������bu���ʰVj����T3U:�s�j�����+ �xp�v�S1i`a�a�˃u�V!�8f�A6��¡���3Ry�W�^2��^uw]Dե{XMJ��h6eBn�~S��-�pKi-n�74n��f��LP���Pc��SAm=\9�D[��`.�F���Sɷz}o�gQU���r`��O�W����e%1�_�|���V���#��[���J�iЉ�}��z%;�߹��jM�3f�m|�±!��`��h"�G��)μ�v8�E'�ͅ�-�dA'����yZ�.�̣�Ap�$�3� Y�������������o�!��i��!�r�z\�ɔ�,g�2UY�57<l�����n��vU�]� ՠQwu����5��൩ ��y�Yj�m4a%����|��o��M�í��῅��g��7kyrK�����A?.C ��CٳlA�� ����o�5_��t|O4����l��v$������@���E�p&XE��T���~F/������Y��:�U�J$��yt�������8��D6����{�Zg�J�v�0!�'��.zG[�S�$e�ڦ�W���<�>�b0�V�,,W��xE�y%��qy�Z�ay4f{��"��Qp�>�ġ�6���R"^�A�>co���@���]������R�~�8�5=�[�A�������9��|*S2qsz�|Qb��IQF�k4��>�K����)tj�ǒd��P�aZ���piW�_^M��ä�5��|נ�*���f%��� �3U�9k���g#��H�?܁�)K��K)�I!1ɦC������9��[�eVW�a]9�K�����H�o�7�kF���D���DV]��>�f�(8!���C�^I���E���#�(E��s�+��u��;Yٓ�ew�]�/\l����� ^ �C��&m]c��(��f�n�@!g@��R2�rVt~}�����i��3������H�/��e�܌��b1�؀����O?����H�d|M_��l����E���#��_U��軟�\��`�>����i��Ub�h��d>������ݩ ����Ϙ��҇Z�Ky��Ї'ޖ�G̸�� LT�)��d���ŕR�.���H7LՊ��L�(#�u�ꓰ]��gm�-��@h�!<�K��\��
�%� ��/v��2�4�a�����L��Q��6k,������s8���9m#��K�b�^N�=TM�� k['ǣml�ܥ-Dj��՛�-��aw��Y�H{���Nd$F
�93^!�3�֏S0�q��U���͋o)x���(�E��b�Qb0:v�vZ�?%p{C�N{{�[ݤKG�'��B�[gB]9�:�1�S��H&�:�+�qo��g��IL��ܼ�Xu5�G���i5�C<ȿ`pI`�LNT��/�C�>KS�q�uO�G�ĩL3��i�i	0��+룑�7*��T���'χ��=?X1!!ִ,�m0���.}�
����w�u�Qf�&�S����o��+����NIԠ|2� y�+���UQ�Om���֭,���������_p*�!Ҧ������
(S� �z�Us0Z͂��o�T��K�f��<�����V�����e/�x �t�#��D���zV�w�R�(�#�+�sj�LߙR�7?C������IRd$�p�͖y�Py�-OJ�.��G�Z�M��HH��T6�)���s=PkDL�Ȼ��˙�Б�4"�Su↱(B�a�q������|����CM<��ʸP��.�W���}�p�8NrW_�bm-]"�{N�88L	�L(U�$��� v�q��ai�p؋�8`^?R<H��IoZ���1�6����G�<I�ۓBz�=�FU��Y�"�Jit���$�5g�%S��g�v����� 'VX�#>Zkj�IQ$�Aqc��6ոW��E!~���ͭw��Y��W�Ӯ*hn�wWCR��N$-b���a�r"���^Wϒ+�evc�y}�]��BGԺ�C�1�!��g�/;��s������l�ʶ�O���1�Ͱ�s��@	��/�ʁ���D.�������Q�6a���N�z�S`;
&���ðf�
�Y�aV����W񶧟OJ����Rc7�m�o�O�'���	�?���	��G�eP���������I�Ʀ��N��ۿ=T`Ou�Y���k� i��בo�ox����롍���J�z����G�0��m�����t�!E�V~���Q�==	��8kWN L� ��2���Ve�»�뽍M5��`� y\�\��a��4.�n�*�����|��R,hہ}v-��e�O�^���L���	�,�	���M���b�/�f��:Ej���mfы�e|�#yC%VI,8}�4f@ѣ�Uށ�2y�ś_ �n:�*���Y����*��9߶�)r$C�o���^�m!��e��*��Z|x�$�E~�c��u���j�~�9F�?%�&{�9�Y��QFKs�_rF b�&��1�r���ṡ+K�iV\��
�x��g=�UŃ!�=��s߂�b2�D�n� ���;��s��կCb����7oS/>;1��,)���K=���ڮ��	Q�ԧe�_%`?A����*PR��?cܒ�dx�������
BbF6���ŷ�\�K�9���C���z��{�+��a	�"+>��#�b}�����?:����z2�U7'�B�&��M(%B���ruM-N�0N�x���q!�99��{E�H�~#ɍ�)���Ad�����
����Q��:6�΁���0��=5Wa�f1�t�7���!�  w���_�M>,Ŭ��g�F=��/��gM�-�{q����]r\p���lp���DT�y�]�UW�ŵ��gw by�&�l�/���B���Y��\zn���&���%71n���n?����=Pf�{'}m����>�.o�5� �H"�DW���{r�v�K�����XyJ~U�n:"{;i0�י�\.$���#4jdm���J��7L�u�,%t<j����Z�U��gs���̵: ��CF����i{Ra��3��-VK@��lDA����"�~x�y4�b�8���Gw�n"�@��M �q��z)B)�-~n��-�KD'#�ri��|C�� ���<_Uc�O�A��995:�[�,s.Iȭ��]Ў�l�o���QpS�a��`�B�O��Q�d%,�4�jA@�wV+��]�#��[ "5��SЄW��;k�;|�>����#]3AL{Oݹ�L����f��=�G�O)��ռi�i8�k�'L��j!v�_�t�`��4l�.�Iݼ�P���3�w��V���u�BW+^H{��m�Ph���\C�&�ɏ�&g"ώ�R[~�y��������]���՛ωw�n=��Q�����$n��T����m� d��#�|Q���G.Q�ޢ �\XO���rr��c�{�?�`s�U�����l�$>�����5���ߝO��`��ޑ�ō��h����YZGEPQ�X@�Th/s�9%��x�$�ջq�	��ZJ��}yo���@ϟ"��S"�D�u���N	��6崨�+��'V��zP��ns6e��2װ�'٧B0�l,�K��3�y@�q�X�<#lf���"�-oQk�9�n� ��W����Yr�����0���]�k�$+WR���S�;=��[�A����g�i���2$���s5��Q}�Í7kg�>�Q����)o���K�!au1��ipD��_�^�^�J5������v*^2)f@�F��30��k�6��s�C������K?`�)�%!��C�F�-��y�R{k��t��W���90h�@;CHwơ7'����=?=�ڐ���>5{������C������O������#Q� ����J�Z�W�Ǫr��َmw �/Z��HV��h� ��x�qm��6����ٸ�2���;�Z�MYA�ܦ}L����T�R,��j��cX6у�;�:-Ɲ���sԱ�H;O�	.��)�c�|Ȉm����Zl�EQ���g9_��߲�ճ�6�%��\���U�zDU�zMh���d�xӌ�����U�{cJ˪~��\�Z|���Հ'9;%���(`T4:�?�w� +X�6畚f7�厊u�@�C5Lu�淓�b>ˢE-�m`@c-C<��������%���{�1����vA��2�G7a�A��,7��"W���,p.��s嗮�x�p m�h��bO�T�X'�M3-k6-Z��-�w��?f�?Q���a�jY��{��N��
�'.9.%�׎vf��oq���Ћd��(�odOw͋��E�2��3B:1�]vu%�SC�O{�r}�?u��"&)�E["��9��1�T�S��d&����UAjQ�E��g��Ig*�7hAXP�eG"���5#>/Ŀ���#N��,����FS�t��x�e���3d{�+g	���+�V��r8���i}魰�r�?:�!<?3��/p0�Gm�G�}�����Z��a+��l&�i��r���f��+��<���O��#�s���6�W��ʑ��v���[�� �6����_�S��&���ٌz�.�j���U���}M�o�k�е���f�B|*�1��eʽ�x�|t���]��ԇ������ήf�tjY�
�M8D7��T��,���Ed�����ϋԐ-�5�)�G0��<z�8ฅ����=��=��dPL�LiﯻY咙*<y�"۳.+��왒B���q�Vaq��7���<'�Ӹ+ J�i.s8�b}���G��r���}�v]��4{�)R�s���Y�(��$�-��"�q�%iZ8Ӌa�^z���I|�O���,���vz�[����`O�d��
�U��`�}^�J$7��>q5� ~S��ˋ�Z��\h "�H�~@_k%Y,Il)AA���c�o06l�3x!y@_�6��w��*Y����N�LhI�W=����(-]�}ϼ5�">�j^����+�s�c�BvŝM��=
��uoC� C!�0��;�C���Aʌr��;��%eO}cO1�~���c:@�~/3�#�2�")|���9�_VD6|E����s�b};Ed���_�ab-��������[�1*��S�c�����hRo'O��	��7��8�ni1H|e�������R\4҉��*�ɈOۚM��ZNu�Y����ӄ[�=���ъ��ɉ+�|H4�a�zV�թ�7oG���(^��[tF���1���6s�=��ҵؔ]W�ۉ��Y��M�ܕ�FX�������~MФ�`�G�\
c���ʩO������ר����/Rǆ �xh"#m�
�K��AL�zL���ҷD�uי��/�l��,ھ��m��ً�w��^Ɔ%�=�8��4�Ǎ���+��.yQ':�:��num�*@?�Y0��0�&���<�D'R$�l��S�ZЕ�E��e��Do�WZ7"�?KYE��gc����@���Ai)��M{HM�Y�Q�9ks�LF;ۤ�e71�&	�G������iq�=��)�xb}igx2~�-�=�*���)2�n�n�al��;ֱsBF��J���{�F��S��01���)9�2Kb	���I��	L��f_���A�G��UE{P-�?��"��`���·Tٗ
�hFQ�`�@_�p�K�锭�ͫ������B+�Qx	�/��#�"���}o��\V�� ��p7���Ѭ-�( ��Uu�0�q���PJ�,ti���p�W�#��#F�K�Ď8�<p��F}�զ�@����μ�Ŋs]y���W�UV�f[�'�A��T ����GMM��ŧ��gZ(���<y��񗥨*{�V+j����]��p�`�l˗����D���a�Б�Ӡwئ�t�b,B�g�l/�O����q�tS \���ؽL��?��%�@F���H?��ؒ����'�c}��ě�V��i��5^{[H�D��������<�h#�3<�~�ˬ:�`=i+��2R(��l����4���������B�Ҝ(uאv�W�jjP�Ԁ#U0�xs����+��" ��R������i�c�a0���gV�8n�?A�	�x�9��y&0��=���
wӸ2��~M������B��~~�kO-��!KA胭�*�@���KY���yc]ʜA���9�O�[q�.�(I�&\e������<ocQ�٪���`��4O)���~;%'����&f�VF8��I�#r0�[[�ǽ�O4�H�̖{�;7�G���`3�^��R�b�yCG���)�t���8�ܣ'�x�5�Z/��t�=���.6�7i���;�3d��_�D(���'
��S��(���7ޗ����Ɋ�g}���Tm���� �2���]&9}Ֆ�^w+V�ʁ$o��J��ۊ�/�oϺ�mj�Z��և|��y������3����� ����r�*�v�,?�F��T���dl(��L��Z��5O#h���O�m��4�ެ�}�9��o�3�E�QJX;�iT���#�&N���lûL����>�JZ;tyj��SH��Z�ñn�D,Z����f��%$��2�&U�'��z�d,���e����E�b?t�0� �,�_h��dYy[�qo�?��f�";��Qf*���"���վ��6TO��,*�N�T�	y]z�����RgN�n>
=7[�a��8�I���	=2s��^Q�p�IGݭk�1�>x�#��)j�]�HŘ��a�t���p#�_ԏ��5 5�Na�V�*�tf[����{3�}k\t͝�y�>��7�sK�A�)�,I!'"�C�GUt��"�vm-���dWh89-4�̻�0HR=@7b�,�B�T:
$�5�Ӭ�>Pj@��2�C��ϥ>�H��T6�n�#�*{k�:�'6�%Ъ��ىe0w^��/�g������V �(��m����d$��*ڔQTM��Ŷ�o�(|��Z�}�c����<��D��%���~�D����O��#� ���O�L�DEM�~�o|C�7��=)� 6E����_ej�^��Q�V�������U�fh�=�d�Z�GY���-6��B6˅Mx�&WZ/����'��>߽KY�3o�T�^_�TB�;�qM�7��Vd7�h�0~X�^g_u�[1�f������-Q5�@^� <C5�q��@���c����v|g�2(z�a����:r��?��&�,���m������m��b
6ߞs�M�qEkS}��b�:����L����a�HJY���{�c�N�ܟ
A��9)���<���3�q�X8Kx�Ȥo�F��&�jE����%4:�΍v��>%f��C��@{�t��ھ{�����)�[�q>9"Y�1כS�d�&@�q�a
�e_����$g[E�I��@ܲ5)X+GG]���TW9B|�5~��N�M�%��nS�G��D��	��_gE3\���L	&Y+�)���f��_��YL�_:a?���!W���"�~0��Q#�o} Q����M�-U����&⟘���A�O+%�������P��<ci߯�#x5�E��Js�#����2�����_&�E��3�3� ��		`���i6U�S��x"roL0�������V<��PKu�ee��x��tEB8㺓%���a�m����_���d�j��H��7����@���dP��v���O�-:���$�0Gs%Ś��>�S����)�����x_<=N�AP�LVL��ޙE�)��!��	�'+�B5�q�"��"����7�@�<�I	��)���B��%}�~��r�����?]u;�{�U&��f+?�(	�#$K=��v��q�.i�:�<��^���~�oI�F�u���������2�Ɛ�w��rc�so[U����U�J�T��x�5]��S�`��"��7,� ����b�k��I�NXAy�cwG�6K?#��K�!tΰ��HTwn�Y���ɵZh$��Wxߟ�z%-X��k"�y�^:�|Ml�+��4c2,�8^��8.�p`CR/H!4��]�
;���U�'}��*y��3(O8�h1�O�iX!@��C/n���͂X$6��^���{�6�t�D=�{��;��At�\�ˬ�?��#��%�ޝ控.�����cV7owΫ'
�_		�؜�b�vlh:e�!���o����D����\�D���u}�օ�uR줈������M�ѥ(����W#.�<��z񡱩���Gv����9"�"�t�n�j��q��=G�lW�g�v�7�h�&�LH�x���3�Mkx�`���\e���׾T�jEv�dLyò���#�RbŽ�sz[}tT��]�:�BLypȿ�i�%�퍷��/c?Q��4N���m\�n����Ù3�%�R8���4oj�i[��7t�y�T[��?n��*۾�Y�X��������_�_$9�4�z۽��S^��q�e�;ʧZ򩟖Z�Et�c�̛����8<r���{�uYM�Q<H�s���FvtJ\&�1��yϢ�B����i�h�� �-x=�g��ZŹX?=��d�8�w2<�An��o�GQ;��s}����P��v��jS��
1�g�)���K�@�Dh����	G����+_���A�����fP�-?�FƝ����l��؁
���Fl�����ԥK��ۭ����Q6�p��+O��	�\�4P�#n�Y4�u����o� �7����6w��3(�7�<:u�h�Ҳ�.ц���5 ���(v����#����_�Ș7���GF����wٻ�����v���&�����W,��B�@���. �n�<N�Mt�+ŢI�g�)!�Ii����#r[�1bS��]��p��l&��ۺQ9��4�K$��{Y�ݑlb����b�/N�D��ɏ�
\p�=ؘ���z
%mp֝���?Dz3���w�Beh}cZ�l�&Ӥ�25�H�:D�|+��G����~�	_:Xf7i&:	�*����9��;�4`����ڟ�)�m�u���Z�j%�Ȧ���U���s���B>�R�r {���U�F��i��;a��胩�rV�ޟ	ڒA�#���M���a%yALKX݉�v��w#7�v0�M����yc�B���~�rF-���K�z���3��\������cewA���9+��[L�(.�����$�d��"��o'�Q����W��`qB�Od����q�%"�r� ,L!��Va uS�#Mk�[�.ν��zY���;�2��<�0�3��F���R�z�y�VGP�k)]�_~�8tm['�$���h��U�ß�L���.&lݲ���w�3LƧ��;��6�����|��Ǣ�6��s��{��K�ɅK�g�g�����:�o3o�L�']�]���Ց��w�]A�<B�!|�i��
8
��m�	���| _�	$��.�R�F�d����*rux�q!l??�y�˼���l�KZ�ߚו��5����O6OE�y��Ǎ���=���߫uD^��,aE�r X6��TvTïBȡADZ�&ݻ'���CCJ�Ƣye���&��V����#D�^q��V��5��!�'�<zx�����ei���4˻�+lKk0ڵ�,=�כ�$�yveq�m���f,�["֦�Qa��$��g J���ؘ��χ���SA�]u�����R"$��ˠ=�E�[c��s'��������d�"s�GfQ��I�Xk��>Z�����)eM7ǣ����9a�������p��+_ᇽ��5���ױ�2*��cfv�
�#3�!(kQ�f�8n��9>zܒ(�K�C�)�e�!�~�C�����:үp�q� �*)�W#�{9HXj�6j�H-��7�b���a�5���������>ky�홯qNMC7v1���ٸ����d#ǰ�Eu���w����ͭ����ل�w��6/��E��q�vY� h�'3!m.��堲�w���O
�hw��1mp��%�9}���!�}8��&-ٙ�[�y��m� ��􂩒����OP�D��?1|�;.�����дlE�����f_f�i(�l�,�ѥ���&��!U3��h���dOˎ�>M���~�qB��`<ОaѬZ� >��?�'��X�x���N� T�����v��� ��f\7]�b��x��y�uy�V�A̾���-��@Yú<�Q
�,�9�[��qDϣ[~1v�R62���a�m����-��##�O,f9 �H���$���P��m��\ub��힎-�M)�ik�0�~���5������^�/a�F�Yyy�{^T�N��
�./9$��D#Ə���q�A�Ƅ��@ o�]���BE����b6:��v���%�!C�	"{,���u(��@��Sfc[�9�9=�1�y�SiV�&{,,��ި`ǩ��^lg�2I�F��-#�X�XG�5S�:�C4u�q�x��fNг5��6�Z��SB��F����ĺ$�3�ė�	�ܕ+|����%uq�"���"�?��Q!r�����0qc�^�w}�����bї�hwꂂ9&��`�h�d�7�+`t�����8��){�$���>���:��>��^��V����s_�uR0P�N�ό������+�UD��sxo����|�_�1U�8Q���#����e ��x��Yt���u>�˸��+�۹T����j����C.�7P����E��3��d���^$��-����+,G�:+�~�g�npR������۳�=�gP�m�LP���\��`��Hq����b�gBЋZq��'�<ǭ�� �<�j��A��߆�n!}�5}���r�$&����]��{��ʳ�-Yږ�({�$���1ܫq��iP'��+^�hx�|I���b_�g���5���z�l��Ov���U��B�3mJ��� ��5�;3Sxb$�'���� �^�4�)k�TCI��7A�adcR?j6�2��i�d!o|޿�7w)�hY��D�Th�4�W�����?-S���rF�"��^U�@��D+c�kcm5$�ӎ$�3r�����C^�!O˦؎�;��$������9���!O�F1A���lT@�,�/���h��򧹿��տ:6�݉応�V��;�D��܇ �W��j:���{�Mw�'G���}����#���^Ƹo�=['�Q�	$6!��=����,e!iK����q�����W����PͦѺu힎���7�Y������i�"��2��w�pz�����"Gѡ��5��8�rt<E����߬=�v��ά�W_��1Gy�P���i��SN?�nrcMlK`���\��C˒Т�����߸�Í�c�-��R�#��n����׀�ҹU��L���Ț+𷺧��J����/��5�k\ƾ��m״��^����I%'��8�tA4w6g�$3�R~yG�(��n�}^*v^%Y6����j8�z�5$�)ɠU����z�{|ce�e%�3Z�r��u�E�bicql�BTG�O��7��6%{�ԅY'�Q�vGs[��F�-��1����mn�\�vi���{��x��g���T��=��7ߓF�2�!�n���;�9�s��}Հ�� ���3=S`��1�i)/��K�?�BS���	Bn��E_V<A�F�K��P�F�?,~�5Z�����
��
I�F�n��6H���|K6�V������<.����+
]q	�&�@6#Ix�TTM����L�C��7X��o�#[�(��BB�u6��Sߏ�qC⢫�CS�f����G@#������p�2�a����N=���p�6f������2�;������"�Wr"vb�t�]�U ���wu�M�/ŝ+dgKc������ϥ�٧��,�I4�]Ci>p���l���u)2�����[�V[P��0bJ�A�]�a/��sM�ɪ��\�'�s�ǵ]i%���1?�Βn�f�]
5}�^��G���5�ЂH�Dh��7�����׉^*��!,~h�:�)i!@�"̿�ي���_4۟+�^�����S��Ou͸}6~�j�MS�
-�U&�s�g��}�*�� vt%W&ˋ�i��=a��4���MV�]��@>A�]��.����4y\�.ӜԈQZ_wI�/��M����wBZ-~���-v�]K�Ԣ�#�7�M�������Mm#c�vA���9��v['��.�H�\�����}��o�l�Q�����4�`L�O�D��"�q%b��{Q�܉V|�)� L#(�U[��H��*��u���L��;����BVg�3�� �y��񜐮��O
G��).�ܼ��K8O�'���;��P�ş*���ea&.A���-����*3����'�,�H��Sk�����
\��7?�ğ�^m��Bɀ��g3d<ED�x��iZv��bJ�]\BZՌ��w����)9�U������E�Em��p���Y|bR��x���/B����t�?Ǌ�#��r��ơl߇?�x�����BMl���l����j5��Q����O��v��{���6��P���
F�E!��X1 zTyI��j�C�\Z=���"����AgeJ�r	y`�	%@������D"�J��
��Fd���N�	\'g�Vz3�����e}�;�Ó@��e��̳0�j,��F�d	y�<�qe(U���sfg�"q�\Q\
��ߧ"���1��J
��v���T9���]p��5ʶR�e��x�=���[>Г��
�:���:��ssf��Q΀�I=�^k�'�>�$q�Yڌ)`.���<|�a�Z��y�}p�n,_JR��/G5̆��*���f�����3���k�4��q-�4����~�Kpes)�i!��C{
��bK�J߮l�o����W�T�9c��̱1PH�M7���x;�0���5�I��>��:��tL��Cr��t-���=�$��#�s`��կ^!$�V}�C:���w��/H���+��� Ccwn�Hm��� ɇ��f�
��gŬ`]��!�`�1}O␴;�c�����ٴ�z���HC�N�x�D������O�3@���|9�P���`��WE"VҽtW_�������`��Lz�yoF�U�NU�n�h�Qbd���ӽB��F/30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�&ڜ4�z^�27лXo��R�|n�?S4��{2�в��3�i��R����@��r����>x�<%Vֱ)#�׳��'Z[�Ϲ,@"����4����Z��mg�U�f��Go�����X"�q���D4�y���O|�:�G��oT.�t�U���8 N+[II��
U�v|#r!��HQ�I1���7 �dI -/�,.y��1#r�.$�����S�����ڮ 0����o}�#��o��O\u�s�4p����O�>Ԣp0ut�U`��D�i!C����k�z��( ����x��R�׈ӞX����jI�����q#;r���Y�t�����ه)�9IhnB�v��r/�#�6�ˉ�7vCl�Uɽ>^M����5���Ve�)[�����R��O�>Zp�#�؆P�(o�\����9T�͋�k��Gt�_ÜH�e���ʽ_�	��l�ګG�;Tx��ue6�G-z]L��^�nؗ~�!�w��t�}T*c�w�����Bŕ:������2!�,�f�)l󌄷r����b��<��}Փ��}�����څKrg������c|	��e1MI$�?#�>^a����Yq-�锚}C����vb��C����H��@�nf��a�DX02$ib�!�����t5�QJ����ݡ����~���9"�:@ȏ��SJ_�Ѽa;a�y�N��
-t�5Mw�P��"ߛ�v [�U�ڝߚc���d�t� 1���M(��G���pyuZ���c�)�ê��\�t��j=4>�~�a�p�!�x�:�o`a-A���B����=��Y���F&�n�ZkW�������N|/y������{��$�NwEN|i0}�6�LiU���h,n��	��3N$	"@�0�<��욕�Un~P4�B����6����;��Bl˝1��9�1~���c�=�g�����v��x,y������mP�`#y�U�!��g9氷n��$q���j��3��2���PH��}j��2w��Hv��,\l �> 2��3���D0t��J���z�j<��@���o�� -y�BY֩w�Au� �H15j^7���������G;�4Y��kt�+;(A��3�24�j���=���Z��T��Z�@��©	38Yj�Aݭ�ԫ/D���oz�N3%�@�Be���	��1�b1�+�3{� �ʇ���L�DƮ�Fc��]�h�����q��9,��sK�K�U(��������R!�9r x����c�������왩e�83�e�n
N�j.��"�2��*��i2cs�� z��"�N��R3Pr�`��d�/�IC-�	 @��'~��u���%JX���ͭ!&:�}���
6߂��;�u�&y:�b�Gl�(F[��O����Vb_��gB���j���#\et}��O|l�T	Yr������m)a���h3�\���h{��M���B��|��)n &����z/��Z�}���6Qy�՛�����!������_�K�����U۰'����i���ơ�5J@���o��A�j��K2�ݔ_�3���������S�8
fjj�SϺt�|p2:�T�����_q��u��/ w	�,HJ�8��� R�WE��i���V���5\�WFė�mx�"Rqcټa�k,k#��lsA/��BA#�0��bOɽ.x.����xk����ϲ����|Ĭ�E�k1�Z:gx��y�V�
�c�i���ҕ��2�hE�Ѯ
�b��sԜf�]��l$��z�7�4��e�񃈰�,��1M<?wߝ�$ƶ�q�s�G`��P?��1,ޛ�ѦtA��/6���q�i!��|���2�U>�5 ˘�J���\�Q��獆-Zvk��9�j�?�#�����3�t�����X�	?%�k��L�)�$d6�E�Sp��ׅr�����[:���qr��rh�2~8�臃y���:�X��ϟL��_뚃Ԕ3;�� ��������ٹ��[H�a�y�"��%N�9�o&���əb�$��O�zahF��wpo3ȥ#�43;��<���J���� �f"��H�\�x
�;�Ї��Cz�-݈LEW*f;VO��HS	�m�����9��n�<����ڲ��i���?,��F�pe�ۢ,w��O���Sn��XiE����^�B�1A�@2�5�ɶ�̊r�t��u>���τ}m'�VP~��=���Pʢa�g"\�CV�������V�X�;rҘhGy�(��t��Q�t����M(���(ܠ��52}�O�q�9��g����B�\��9c
���n�}j�TB�*�O��PNQ��W�e$�cy�
�o���^Y��dB83�q��W��!\)wR���g�+��1�xY�L�d��	�p)�p����H��P4F��1#��v�l9w$-���G�����g$��bK�s���Hl>�т	"Te�f5]������@&4I�+�=����K��	'�,rC��S�p�7X��7�@��i�oa��ue@ґr3C�פ��B#r	���]��yÿ�^���A�P�P򙁎Z��l̛�/q�^��y=4d#&�f���0���m޾mk�K�)�,s���t�[t&[M+�U�8�4�W�:���c!&��s��t-��o���$�M�䜎�A�����$��qR}����ę�MuI�"����*l�'�̨�iW��p?�Ok��m��D�~4i4U��'~b2,Fwyg���x��f�Q�J4�����I�P��Ǝr^t黎�5EFaF���83R*����if��sSs�H��]�ɿw�o��5����T�E`��-�i��uﵟL��x=F�c9�6^zN7�ك��B:̜#e�>�"4@z|?�g�熾,[�����|B�7<�E��TVC�������@��T}�|B �j�� -�;i�*|$.�+Aq��.�S��]�W�a�i!�s�<;E���RȼC��+Dpr���7M�ӆ���C'rQ*P�J���C\���;/�v��T����ݔ^[�8P��u�p����rAZ(?��Y��u�M@�7�F'�~����Pd�[��x��^��Fe>t�["�[9Bu���%� r� ���"�Iޯ)������[���$�E��V�&u��q^�!��ǵ����������"��.�6��$^�8C���ph皏ܨm����YÜ�G�0@���� �G���z8ƭ����|�y>J49�����]�����u�J��WC�V7xn_]��뭐���w��$Ѫ��[��l+����h_ꜱd9�ݱ��V�]�9Wc�� +�lY��.��'&dݍ�^Ƅ�' %�9<�~��T੊;�[�̩���ƈ���e�ؕ@���'� �DW��;H�-{�H�e=p�$PLL���.p�3 ���Ev?o��TW�=ztm�[�xA����+�����C����H��dz�(�~�6��|�+�����&�����C3̿�7�X$جb�9P� �y>��fi��E���.�����O��ӻ �J�0s#	��W�{y�|#�{.�s&5F�@33\_nX�hT<)\>�{��� M�*�H�P��J�Uʿ��i����U���y}]��g3�F��U8&F!�'ep�&pQ�/��а�����B�G����8����<>�*]薑/��4����a�N��	b��ʅ�a<X7��b���<�کD�k���չ	� N�"K�Z�^�&��X��?�({5�>�@_�ǻ��o�>�PD�{Eh�QS5ķ����p�
AW�D�G��k�[ǂ��x�J���+-m�G>�І��<���4C���{-�JG���\�|��b���}�Ŕ���FdלJ���(�	�qn�2��Ť���I���6<)ޢ����_IWvq��l�_�C��B�`�K�u�L �A�B$��	[�d�/��DX�����_Km��椝��\	�w%pAfW�iX]��}���־mIn���WߓW��%c*S��Ӱ��s��h�5����(��Xl�����cE #-O]-����>-�y�Q��B����,�{�������[��Ý}��fu$�At�ٓsUC����J*M�-3��(�f��LK�,�x��'��-����a��~�΢�8�Y2�C��*0�E���p��,����;R �z��E������ g�R5��_;��^Q�g��$�c���@t�,�"�˗L�t���=�g	l9���&M��gA�i8��Mt�19p�W�6��R���/��CA	��4W�!dM���ox=���ΙJ�����|����G(&)�ͪ%�{��L�m�^,
ה���6��(l7M�'��L>w�}��qc(��M�����bL��!��ϕw�P2�ւ�$��H8��� 3Z���AG�9�7ϒ�^��*!F,1`p�̩��3j��ܕ��TJn@�|M���6y��� �������{ bA�uv�pk(�c6>6�y0�8H�� g]���#r1�����E�_�h=��>`]@;>�. �}���}!"V���w�jK˸�]�l"Zg/�x�.�lN7�'�py?�ZO�O��Fn&��jD[��e�k�7�W�<���9����J�%�\ҩ��D����g�!���郞TH��ʯ�D 
VɅF�Oe�b����9���Y�*��沃��y���ov�$���uu뒡Op�0<=�u����ea����:� �f1��`$�H&RL��3�~��uj��������/_�(I ˌR�Q���~d<�/�K�Jʝ͂p_���x��S���`0���y�a:4o����]Qm�>sx�A[��Tg�z�y	Bu�;�K��^�SsV�T��-�0	�g�'��7J��`�(;�3S�.��Abs��ХdS��-��cnCm�`ʌc����DQ�u;�OU��)\�-vX*�>�m�xr�����|و=\�[hl̡_�kA(��V�5ψ������Yp�y��o-�O���.9�֞���q�4�v�/��n[��ϫ ��>�E&��>��2{X������xn���Sxf��[�����Tqi?N��E�Y@ ��d��K�� �.��&��|8�s@Z��p*"ÆB
���c�>Zٝg`�f�?�o{`k����"c����4w�{�Én|y���T�o]qt)]���( �bI�z
���|�T!FL�f���<�ֆ�z7D��I�I�p;v�����#6�=$�
�֚�����k�CO40k�ѳ�1#G]��.c�u_�4��e�u��>�3092�Ub֔���!��$����kZ����)V��Ϸ�Q����L��Xʼʊ.�M�������;��4���s���a%���)gA�h�B-�:��rs,���׉Ze�v7@U\�>"�0�L�L���2|��(b������6s>�#��Pi$0o����bk�9�4��>�r9���-�� be[X|����M3�.M�*b�������e�X�*^��7��6�ݒ?����8�d�i�)W�t[r0��Lh�dmT� ?��<Df$Α��X�B���k�ڽCiL�2����[�D����ܦ-5F�7��^e���l�9jpi��G���G��m�I������ ʆU����x�aDE�Ö��Ͱ�\��� hm%kw̒+�!���Z���;K`�����HW��f���ѧ?v�(� Zu?��t&l�3��z����\�`,��/֬,����8Cñ��Q�Bx�Ҵ��[Y�a�F��`%I���Y�o����t���D�S\���L+T["��\P|�u}��� ��)?���h���	�(�[뵃�Y���l��5v��v�#h'3ƍ���d��Yj_���rY��-�5yb����^	n�	�a`�eɰ�0m�'Lp��,��s-z9�>=�$�8�c��a!����T`�bA���kf
�7�O��R�gxFv����{i��R�.G����:� 7��9��V֜vHc[Z~��pT��DX���6q�ì�-HH^��M�Ե�(�����`�V>��3f�bS��@��*��#�&���}�bm��ouaWn�d�w���#�G*�Rr�D�<2�߰��ɲ�w��|	C�ɔ� ��QPJd=������)����������ʈ?΅�Q��&����#�Cy�U�+E��,��ދ�=�
_��fF�8���ى*�+�򍰦�D}�F�<N�Q��FTY8�.�]�jd�'�)��*��Y]s|�$�Yʧs�������x��Hg`R�X��Ŝ���-��5�C���Y&Ӛ� � ��.1x��p�9�����zG���OﱑP6�~�&�]���F�W�������T���ʗ�
�e@��;#���F?�!++�NX�V�w�/��J�A� ����uXM�s���VmfA���n��sż��2� ��=��*��l�m! �2Ra�?��a>��Ge�����5�"f_�����W��D�Te��u��GZ\�L�Dx���Fؤ͜!{����T$����{�b�f�����?!��\f�l��y1@r5��'��	AA�bٔ��b(�����'��_�;�":����,���M�
������I���@�-)�����d�c�mb6�C�VՎ��l�ʧ[��6
c�Fw�0���b��T�Ͱ�t���ᗼ�:j�.#+#�����d@�Lo��/J�!�N�ha)�zN���-A��9�w��ȉϚ��Q�[����*�Uc���dИ��)���ś(���G��pfmw.c�(�aP;���kt��Q=�^~�=pt��-g�a�J�ʁЦ��=�=lh���a3Xb�2#��_�}(_�I�o/��]ܧ��{	6�$t�E�(�]�K��i�*�uW��el.�V$���ɽ���`����~�·�O��d��6Ϊ�(��B�.���)S���~�7c,���@������y{W?��UP���q����F2���{��g!�Q�Fj���� ��2U_�oH���j�wz�Ov/߸Y� l�2�R����D��"����E%��V��̄٪Z�e,v���Y�d��Q��1��\d ��M��HQGH�}Yj7d����+(�����3D�4�V��l���nz�V����@�e��O{�3e\�F6�A.�D���L�N�,�@�3Se��6͸1wHH��}'{��w�<�[���1T�ӮN犯�h��X�0.��FQ"���2K>���BSc������Q9yK7x����>�����{�6��e�oe|��NDa
���^��3g�F�����u��-Z�����NP�3]��`_���f���I����6L� 0��XK�.,ua��r?���&�:��:��-�]�TL���6�u���:6UdGY"�F�A�O,��И�J��gO�%�ؠ� �1\R�?}�EO�4T�&Q��'<���6)����\�������E�������+�ѧ)�y�nmu�v#�z�f��d�JR��%�Ŀ�,n~�+��3ٱHx-5�{9�UH� �L��
hթq�[�5�*����Mjo��K?@�A�l������l8�=lb8�P�j����ǚ�|�32��ў1���m��
T����	�aKHWt-�{%�R�1����io�%V���5)�����7���%�o)�c�}���
DkP��l@�gV N�0j�9O��x�mm�5k)��Y%��s�|��oE<�>�� x��L��J�
��3izX#��d�?��EO��
;1��~�a2���7���4�RA�7��S����{i,�oM�[��$�`�qS��'���X�=�Z��,�m��3�a�	1X��&Ԇ�!/特��a�>���˅}�J�.Ӊ}�Ԧ�\��wk��@���pC����с-�JD�X�*�%�R�Y<������@M`��r���Ѱ|�:9�������re�oM<~��;����!:>́�ҳLx9���<�  �aׇ�����&nchGa��"U�ɔ�.9h� &������O���aD���#g3�����;3̓<}��=���:� 5��;�MH�i��Q;ܹ��fR,���|LRM���V�57H@`ImL�m�5��9W��yAm�������*Z�V�e晰���p2�c��& �V��MWnSj����g�cm�.UE�X�Aj���b_�c�!���c�ɣ�z.����m���V��J�J��ɺ�D"�T�0NlģL(��4VQ��;y�h���u�W�aQ!Qz�S�ݠ�(�G��r𴺙t}L�ݾ�=���lxը_~B{�m��
]G"���s}B
�)O�J(N�t�W�6l�0p�
e�o	�*��O�\��d/wP���gW�p�\��Щp��8H�1�u�򙄎d�	!����44�0�X[S#n1�^v��d���J��`z%j��Kڣo#п�f���Y.��^VHO�~�3 J]MT��S�1�&Q�����=u�x�L	�_r��S������z��B̷u�����$u�@�vlr��&ױR��Hϧ#����J��ѿ��L�A��P�Y��.�Z�;�̈/�q�}�^�X4=C5&dɳ��R5�U#��gk�r+궣s�@�t��*&�"���I8-KW:$���|!�s0Cg�AH�����dcM�&���U.	vR��ZR?����q�'�ֶ�;���L?C��k�׋O�F4|��U�V'�S,��yRW�ή:�^�\�=4\ ��:$�.�q�m�]
����I�CFl��P�R� ��6A����	���msތ!�O��������z��H�`~�-��H���ϵJ��������Z�C�zy���a�B%��#�*����z�N���E���ԙ�����gB�ϼ��)OT��������a�㏲���d��UR xJ	i��*�)���vA<�N. ���&�H��WJ-�i�Mm�~`;����AjC��D�I��| �m�V7�'}�P]�T����CA��ln��ab*T����S^fu�PK�vu�B�"=LA�I�ȘV��2�]��Qx��騸C���xH�7�p@[����C�[DxU��%N�7�+`��(YI�dD�X�FѤC��!�m0��Ԗ�#.uhh^��K�#�у���m�P�"�4��Y���qU^�c$C�8�py���o۸�Y�R�r�0�����μ��!�%E)ƸFZ����D��J<���+:;ܥx�@���x�xJ�	�WqaxVd�_�
�v��l>�w�h�$|���f1�lz�č�p]_�6d��������9���+^�lĚ�UP`�R�0����o�\'K4�9�4l~�*����|b#�X��s�\����@����� <O&����6����e(��$����:�.{�� �EA24�Š��
z_p2[1و�uvϲ6���hQ�������H�z�i���S�aay+�a�Y�]�v�nu,�J�� ��Xi����7b���ԋ�Hy	�\f�гE���.����� �~���U�isnTh��{<��|�5�.�bF�@ވ3_y���?)'8@{%�r ؕ��3w��2U��;��O��y�̭��\��yQ*�R�JÑ��U�h�Q�'�RY&;��/����#�bnG3���[���Q<�]]�a/84AS��������	��ʐF�<Ï��-���E�6�e���V���)�	��N(S�ۍ��Z�����@��t�E�*>({�`(�����H��ڇ��[�Zh�g5����]�����O�{�h( ���(
��#�J��G+b�G��tm��i���g��ח,ۏ���J��2��E�\|%��m���h�8�_a�qj���S���{(:�oq��B2�%��jZmI�6g���f�q��_�L�q9Vr�jz�C�*�+��K�q�L�
\�-���i~e/��XRD��+vK�gФ�A��=@\TŽ%�Lfb��X��	}֏A��9I��岉�p���%:�������3,����G��SK��<��0ıu�cP �0(-|�6�'6~g�Q�}&�Jl�����%��
�Ƈ^����}rZ f��ǌD�>����#�*[c�X䤴Q�If�ͮK�ހxV�b���4�9��aT�y��{�83Xd�����ۍ�!1��]���@�@SRKy��w&̀��R�C��X�R@ϱ_�ݱ^�fcgh����{�] �w$,W�yˢN!t7I!��Rg4��l��̹�'0���AeQ����t	�8;G����OD��i�/�:A�;��?f��t�'B8�h�A΄���!O��Y���dB(�eɘ,�6b�1m�m�9�,UF��57�6�z (�L;M�D��8��^cs���p����ͶZ��d'��(�P��7���V瓹(�l3e4>�F���-@ϽDq�z9�!1��`�I�b��j��� {M�8�nkbbM?�$6d2��������`�Ѽr{k}��@������66�R%�
�H���g��Xz�1M"���������Ŕ�O�]�u;�9����0�[<*".�7�X��꣹��KR]�"�"eң/eE�.q��7Һ��qQ�(�O���ᛗQ�Dƪ�eq`I7��<����$T;���vgҴ�^Dh�_�s�S�Lz��M�Ӟ?��-��F�Vԁ���fb}��d����ٞ�!C�����\��FU��Lԙq;f� Yp~�u=�k���1�~>����h�Ċ��#�R72�3�ţ����l)�e+ �S�� ��[R���~d��:F묵3*�My� hŤ7�j��0�By�_p:?���?qFQ8�>��q�+$��gΙ�y�J�F��Kz���)q[S���TK��������l��7U�`74�9Sߏ����q��(ud��-��hnNA�`5⢅����h�QUW�:h�t�G-!�l�Is������3�E�ƈȘ���(M��LT�kL� "�5����k�>H�Y[vҘ,���P�9�X�ܗ�lʋ�_>˅�ިnFܚ������w&)�I��=J2F��G�ּ!��nr�$S�B����
����N��i
Xʻp�@@�;SOӀ̖��j	� ?�44N��ZJ8v���"���U�s�Z�n3g�qgf��o���V+M"N��4"����5.|�˝V/6oC�'t��� �[�I��4
��|>��!���*�Q��q�7�E�I�n�{�jIs��Ұ�#a�t$hzօ>��Clv�
ZR�0���~��#r�C��-�uJ�4�Ho� �.>#�0�KNU-�3��!䌊���k�{��kgT����"����w��XU=�_l�M��g��;�p��#�:����w�ܚ�))R�*h�,���r~���e���%}Dv2H�U�"Y>�S���б���= ��X.M��h��X��v>	C{#4�PN"o��ͫ�9c����EX_�ݵp���[%e��������ș��5�*����aq��s�et�e9x�*i�47ꏖ6�a�?�����n��T��W��	��#LӍrm��?&��D�!�u��Ѝ)�������L�^/��C7M�%�i��~�Z*8�^p�!��j;���� �D�>���:�������A�� 5)������ĺ�xfp�E��� �m�[T�<4 �J�%6ɒVo��.Z�&O;�X<�v��S�G�!���7e�jU�(�_5Z ����lB�5��a��Qi�+훧�	E������x8����IB���`Y���Fŗ�%�dy�%|o�4	�K[��SǴ$�"1[M�+\�Q�`{�d�� _�?���h�	|�[���� ��C%lؓC5!5�v*6h�r���!T����Y�����oX�6�n5$Fs��g�Ƀ'Pэ�!����%l'�%�����s8�����=�h������ ao��$��⪭�H|V������	���v���PfV鄧N.%��&�`:d���&���͝v3�[��ۈ�?��	��Sd�q�K���8QHӰp��L� �`�V?V��&���"��m�Fs���|m_�qG�%�8��C�`��yJK�9Lyz�����>U�w#n/�f�X�d���] K��7�r�!�(�\�n�%)i�f0�XV��}$0��[�Is�������%;o��N�|����:����z�^-ٲGP*A�lĿ��ct&[�-�`�(-�L/mQ(?ِ��v��1,��˺�?�r.���}@�f�>���l|�L5��ݫ��\*f�g�fF4�p�f/�K�txd�ЗYyY���^a��@�|8���Py�j5��β���%����tjRY7����[�0���X��m�R��_4n5^&	Yg-TP�6cs��ِ�,e�6�p�tŇ;�VݴgB�{l�D��;�B�yAs���m�t������D��n��Ά��/C�(A��s������P�t6���o����&l�c�f(f����Ƞ���mO5,�N�C2�6���(eC�M=�դ�K���4c�����_��7K�[[x�:����(P��p����f��zi�33m���9c�R����rX�H)_!�x
`	eϩp,�jh�܎{�mJ�ny�eMb�6��՗e�����ї{�+X��Ӄ�����T6f�0�H�n�g����K1�σ��n[hՊ�9�K��]��z��Ӑo���J"<�c�&0T�1[��Q�]�_s"3��/���.���7�Α����x�OZ؇��	I�e�DT�e��7�'�<o} ��Q��i\6��҂h�D��Z��K��Z꠵
4��s��cJ�wV�*Q�H�<b�"G�r��M>�){3�`=�������`��R�������5pL��=6s.�c�r����!{�3�
��]������C�R���3R=/ű^B�푆������s�a� x R�uM�B��d�SK�+�C�v͛�T�.���j�(�0:��y�~:H�͙sQ�0�>�g��1n�
gKdy�%�;6K���w�S�n�T�A];�� �z��7#�`ŸBT.�S�oؚ�y�QDyd�-�&�nZ/`�F�2
��v�Q#'m��1����-/7��zZ�q�o�&�S���V������,]��+"��h� ��QĿ��g/�(_y���˴��}ֺ��r���:v���5B��7=n
g
�*��}��wB�!fO���N(�vWm�"��#~
onoS�)�(�&.�d9��H�XWr��\�ȇ�'G���1�+�c7�d��E	kW��'k�Ռ���b\0�ED1Zp�v���n���U`.�DW'�޶=�����IQ���cй�7�٣L��{�]"��7)�Y&&���(c=����י	��Jr�)rS뽿�n��N�9�m3�����S�@i&>r�j.�����=#�p��hH���]���E���K�WP�˙��Z��̒�#q��^9�=�Fq&nFp�q���
����4k�d�� �usY�tj��&�	s��8��&Wz����!���s�Ʉ�^��E��%�&M�׎�܀���������q�)j�}����>M��@9�J��dYt'`�ըG��Uh�?�?�����[�t4��U�'5��,�4�y��B��Ư��hA4�)���*ƺH�y����������N/Fx���{R�ˍ��m� �ӎ5Zos��R���x���
� >���
�A�`���-2�f�ݑ������ˆ觴����z���?B��#�3��Y"z��[�^C����y����	�Bq�8��~GT�x��^"��XD�m�׏>M��R~�� ��[iC��*�'����AH�.�?�	���b�WV�i:�î��7;<���)�*C�[D���Hy�*��⑵'���P�h���sCͩ�x@Õ�u�T�/-^rm�Pגtu�J��ɮA����Tx����ewPM�]���un����k�xT*���������[P��8�%Z�!��*���޿IU܁�d;3�0�p�-�������Bu&j�^0�����S'
�z"�׫岟�}l�^Ls�C�9~p���������gY��`����0׀���<��3���}�vVI�P�lJ��©7 �hMQ�LW���J�IW��1V��_+p���}��fw�M5$4��r��l�ȍ���_��d�z��8�"�6�9�3��7�lP�/a' ��9��$J�����'W��9US�~��K�Ԋ�����d����{���X��̞i��L �S����ψ�� �e�[�$����ơ�.�7� ���EM�̲Q�0�;�z��[[=:����Bvj��d����ǅ��H!�Zzc���ծP��,+�8�����b��)��V�9��8Xu}š[RKb����Ȩy(�f Q�E�I�.7�d��E�
}U�a{�s�s�J{��t|�.#���C@j;~_}��_F)3o2{�̫ �Ϳ⛌�UL&����Q��+kKɖy�����tÝ(Uo�']~'\p�&GP�/g��/ɨ�>f�G���B���b<5��]�|�/ċm4Ma�O�����u	��ʜzC<OE��9L����N�q���<��6k	0p�N4ӣ�`�Z�7��aU��^�����{����w���0�f��'�+�2;�h��25;�X���A:z�[����A1��Q���S�a@JB�"+n�L����Ϗ3�������SG�':J����ւ�\l�yYb�����k����j���邈�(Fm�qF<�2�!פ���I�3�6����&��$�_�!q��.�v� C�7��7<KkN�L�x������:x��E/��sX�Y�����K$�}а|-�&9�\`2�%��\fn��XT�W}�K�%�I����H����=%�����zǿ�?�.�yր����E��54�=�c\x$�?-�K=��3�QQ&�7�VV��cG����� ���~���+}~Df��ǘ���28)�6��4�*$����@�]Zf-��K��vx�����H��s>a`I����8?��H��(-��|�[��d��#z{��R׵�'EY�^x"�W��RL�4_2S�^�sg�p����1q���D�,���ˮ�-tÊ��@og���l�Nҹ9O���
�A��f�t���G����;�%΄]�/kA@B(�K�(���� Τ�t�����- ��?,����2(�Yɤ��Wo�=��mM�9,aC�����6��(c�M��b���μ��,c�����q�&���Y� ��S��L�5P������N��H�3q<�����h"�I�Ԇg�!�~�`�*h��Cj�D�܌P�+��n��uMK��6������%����\y{�k�L�D�'B����e6d�M�H(�g�r���1YA΃������ՈO��	s]wܫ�E�/�HT�g��"��P�d���/�p�\�]"UK"qV�/�J?.}}�7^SD����O���}����!�DR|ie}c�7CJ�<����?�'V�\A7���'D�xL����ت�Yڣ��K��!"�{ݶV���FL�b����� y��{��'q���J}�������}"��I�jp�o�=4���!B�Ŝ����1�6t��So��*.oR�+3���/��+k������q����� �WQR�ŧ� ՘ds�yF�"�A�T�Y�������C����>0�,�y9�B:K�����QD�>*�"�5�Qg�V|y@�2�R.�KL�5�ES*��TW�[������7a�`�1�ǫSk P�؊L�O�d�j�-2��nZ	�`��p���~�\�QaE#��b��m�-����U�Q�o�H��z���ֈ�Ҿ�~��Y�Q���IkX���T5�T��`�J�'Y��8OU�\բEJ�
޹x�����R�ư(n���G��u�O&5�;�57{2R�W��b,�-�n��S���+�+�ږ�i���(p@��m�~�̢.n�7)
��W���x��ډZ�\���l":s�a7s���Z�J�gWϠf��0o2��b-2"�P��!�4����]�|p?�b�o�M,t�d��*#A �\�ID 
���|ʲ%!i��'�$���u�7���I]܎�]`�42�ޣ�#�E�$t`���A�Ow��f^N0bQ�ъ�#�����_�u�~H4.���j>/(�00��U9�2¿�M!b~�� k��B������U3Ϯ;d��a�jhXa~��jj�Y����y;�`)䯠+��׈��ܦ�)�eh	���q�r��,��p��1�v���U�H>�I/��� �0�g�I�P��'ۈ��v���*v}>��W#@bFP���o�h�YV9o��o.dYy�A�j��6e�Kͦ�����$�G��i���c) ���2���| Dk6%�9�A��S�����j�'��sC�T�Yw�����1�q���*�����V�G��Y����T�+6���a6g3�($4����z��B,���z�*I@ӯD��3�ao�\�S�OϙD��I�hQN�چ@���e�~;�Āq1�m��L�{\>M� ҩ�(�?�ޡd��h�g�>+���"�GK���P'xRn�筯^�m-9�v�x�x���Q�Y������!E��g�e�:NR�/�~a/�mG)s ������
���5���N^��3+\�`�z��0�*@"Ib�r��e� [{7��ބu�Fk���ܨ�0����:~S2����Z��|{�u2b:��Gg��F�=RO�p���{�"!g�=&e��N�!\`�3}N��O7X�T$���
g����)������\���sO�d�h����nW�7)Sb_n�	D��g�z�,n�	��N���R����Ⱥ�yp��Y���[����UVXg�7�ݤN�#�W��r5��ʢ���Q�j}��K����ܴ���H��s)�:�ͷ��\8%j��ϕa�|�������ߚ��S��0BμJ�	��1H%)ޑ	tyRR���i=
�VFxg5wU��*-��ڑ��aֽ��c��+��dk�#l��ku�0�Z�Od�9x)�A;zk����u��Q�|�EE�Ά�u�x������
A��i�9F���_Eݐm
�	a�/VAMBB����`z7~#�䠹��#��,�,	M�#7�G$�!qa ������%Ӻ�?@,٫s��ᾗ*؝�QS�䶓�W��mr�>0#˓�LJs�_�%4��$���:k��0��������q����ؙX�1%�+�'O�_Zt�7�N�3.h�rJ�{���c:X�~�˭Znr�F*}C9~��ׇ>���{:L����L�5��.$P��]�sZ)��M�4�6�a4�Y"���  B96�~&Y��m$�P�O���a�h���3�B%��oC;���<�܀�K����� ÓB��
H�=��q�;j#"���^���L ��e��V���HN<Gm#'�ì�9�}��t��^b�H%��M+B�d�M�g�z�p� Ϣ�����#��3eS����� ������S�]=�Ax3���
��U;�q���	��ڡ����mBI�V˗�����H(�e�s�b������뗤ĝV_��;MƱhP����T=�o�QHވ�k�(�H�������}ڋ3�d���\��vQ)B����P�
k�$뮸�}�E�BXW�O�h�N�T�Wqw�~{a
sb�o�A!�(����d=�'�̇(Wv�d\Dd��+O�M�1g���Qd��	�5�+j�����f,v!D1^Q�v'�4rE����d�C�zʾ�JE�=��M���mйgʹ,��*����]za�!��)&�wj���=C�y�"r	B7,r�E�SoZ��r1��jM�����`0T��b�@��r�J������Z##+��e�he#����Ě%O��P��֙�k�Z2@̖�Tqs��^=�D=O�N&r����ٚ��!�Y]Jk�.\��Ws]8*t�y&�5��M�8�'�W��B�Ίw!�Aqs�����]Z��5l���hM�W���\��m���о�q8mgځ:+���M�R#�����/'dFۨ�oL�Y�?�H����ɋߕo4x8Uu�O'9v,a 2y�28��c�������4���gƾK#�����+�ث�_RF������3Ran%��`�܄�ݎ9�snB@����^[�F��ExN��H`W`-6_1�aӵڌ���諞�,��z	�ٞ��B��#@ ��]�z�N�b���!��[6)
Bu�z� ��T���!�윛�V��z8�BPs������R @iGg8*�M��.A� .�������Wڲ�i>�S���;@���C�
�D�����Lۮ�����'�EP����y2C�����o���RT�(`V^��*P��uHi��PAuG�X\�PD5{E	��Q*�y�:��B�x��Ъ �q#���W[����B7%��'���Q�=ڂIYH���'��4Kޒ���[ݩ�8��snu���^4޿������s��"jb���լ��O^PgyC_��p��:�w����kY��0[H��zv�"������H���zp5����J̝��+Gl���Sd�EJC[W͉V�A9_�7�:3���w��|$������l
��:�(_�pdTl�<���8��9�H�����lT&��MH��0ݨ!���|�'�y�9Y,�~��Oˇ��	��b�����e*��;=�Q�Z ����2���N+�)��e��$+�����.�, �Q�E��ѲU �r��z���[��b���;���1�v�ǉH�уzg})�Y�Q��H+�����"�����������S�X��H�_�1b6Hz���y��f$��E�T.;��
�����s����2�X{�PC|>ǵ.'&�H�@np�_�Rʈc��)��L{�� h����� ����UP��=�/�	XR�=��O�y����{S�!U�Uspa�ۇ'`~I&��/k���H��B֩G����F�B��3<9�G]C�I/��4�$}�S���)dZ	�}� `'<S�>ὢ�� -��G��4���.�	4y�N�����lZ?�y�e@���ږ�a[{���{ބ�V���j�<�����6�h�\5?w��3��E˵�ߐw��#� 2��)8�.5�JF�+���P�4�k�ȏ7W�������2?�J��m�Z�\���������>��<�7G��T�(ʹyqJ�2{�r���IR"+6��UD�}��_$��q�mM����C�)*»3�Ko�aL;\���Z[���%g/���X���i�K(�4�J�*Qe\�J�%��f�ߦXXU�}f]q�0cI5?�$��2%���e���~��É��}�� U��Ip[����A��c�I�(��-�������Q*A#��:�g���E���ޱV�����}|�f�"��=��k#�B����w*�h��h��}�f1�`Ka4ox��������a�W�����8Ù����Ĭ�N��� �tF �'�T�"n�R�Xr��H3]�r��lˍ[�dR���_6)P^h$�g���~*�u�}P,�F&�2�dt�$ڕ�'g��5lT��=K�Z�A��R��t��������0��Έ�/�+_ADp���j����W������+�C�Q�%��(!���(*�[����mQy,���.�6gd(gh�MO�ú�B�i��%ca����ݺ�f��]b�|���P��PM_؂��# ��)�3�=���"���o�M���
�c!��`K?s��N�j*��ܐF���u�n�QvM�e�6�EY�]a��)�a�:{��]��̎�+�>�~�6h�Ur HUwg��א�e�1�����W0�NՌ/锍��]{�����;����),"��w����3}�˓��]&
�"��e/�P�.D�7b������|cO�\�����'�DVF�en7G��<1�z��7�ȫ�`~	�D�AD���C����	��ٸ��;�����gVd\�J��b<����
�t�o�+%���'�NB�ϊ`�������M�!p�K=8�����&Š5��Fc�5����W�����R�U3�kD�3U���X����q����M1 :gcR������ldw�����E/���t���9���b�Z�0|q�y=�	:�K����Q���>.��\͜�g^ߨyDB����K
	�ʹ��S.� T��(_1p�B�n�(7�`����5�So_��\���S�d.{0-6n�J�`��t3p�`�<Q�K��떛�|-�y@��H�s��Yq��C�Xzĺ�<�)_�܋
k����}�5*�[���ιY����+��� ��WBȸ��'ʦ�MՅJ��n�gφgQ�yϩ&�ܳ9�%2ִR��u���vn�sSSx����������i�ձ�  @]�&��&ל�;�֐�����N�`%!Z����� ">���#����Zthg[��f.�o6����l�"ހT����4�TB�^�|t�0��\So�p�tD�0�. m�IH%}
4+*|��!��!�J��.`7KnI&c�G��N��b��#��$�kK�b��i�bOꋱ0f/��y�#�I�<uھ�4�n&��f�>��04G>U������!���!Тk51�����~�ϲ���r��aFX����2���������;QZ���O~Q׌���*<)��h�W�uzr&���^����9v�3Uw�>��^�'*:�4���	 ��i�_{*�zP��Z>���#���P���o�~3�]wy9󿰋s5��@s�E���g�Ge�4�E$i�$����*�\�(�e�t^�����e�?G*��'7z{�6'�e?I���Spu���NW��%�"���L�Lc	wm��`?�_�D��b�J�_�i��X�L�j~�9D��f�������������^ ��g�Dj��O�sk��6����$�и�׮� �TE�GJ��T
-x���E!c��;���H� cv%�//��N�� �Z8*�;&��
$�㧝����K�����|(2�Z�^���%l�g��6���-�ջ:K�O	ެG�����O8��� �DBߴ���Y.�~FU'%d�$��o�Z���"�Ƣ��SW�=ҧ�i[ݪq\kc��G����� �'�?9�]h�g�	�h[�0��t�	�llh��5�,nv�<h"��r�U���Y���k�Y�Ɲ�5��[�=��Y/P������q&« ''��gSsȷ+�x=8�YTJ~<�a������青��=C�"7����F�Q���v����A�ߪ.�����:�fBöke�q?vä�[5�{�<��3����Oq@�l�gH-Hc��(%kԐ�E���ޜ���Q[P��"Tbɚ��[��*��ט���*�b�:opI]n�K|w����>!b*7�я$<m��zp����$ŝw���|$X���Go��Q�;����t)g)��|y���j��?��Qꄾ�7�#��=���d+ N�,�j�?���|$��?z�88����.+��1���h}S�><)����~F�x`8��])���r`)���">OsW_?_�V�BJ'�����X�#߮]o`mpc�2��������/�C� u�:���Z߻N��:�E1��p����
z�;g�J/z��u�~yQ�]U�F6.�� ��/�i�)���Ţq
�����k�΅�F��n+�=X'r�wx�e�� �A����:���������1�m�g
���_� F��c�2l���XN)��?)�G�Ym\1�2�?�>=��G �X��|��WH_`�K�چ�/�T`4�uM�G>�L�]-�F<����!��e�\C,T&��_E��L�}�D�qy���!��f��t�{ry�q���{�$0�ݫ����"��=9����ZI��}�W�Kx}���$M�ކ����&��/���|-�p	�e���~h(b��C�·�����H�V)������0m�by�Ǩ�cto�2'���3�݉��N^��� 
��@�b��{JG���I��a�8�Nlo4-\18�w�C��
/��^m�[�?Sڅ1c|�'d�	0q�\����(�BPG}q�pa�rr�c͕��|���ubt���=^�~�~�po���`���C�a����|�x�$=���/�.H�V"NS�蘘Z��$�/a��⌀{��$o��E6C�!���i=단P'�7:����$��������ޙ~8ګ�*~/�J6�k��#�B��˅�N�!�+~t��c�w�O!5��O��:	y��8˾ĂP���a��S������D���NE����j�a��k�2�����J����j�uGwuM�v���L �g�2�ϭ��`D�)�+ڌ����Rs��T���I����a_�Y�qPlg�Ks1	�S<�h�<���G#T0Y�Of�S�(+#���
�3���4��h�续��]�<y�Bu@�C`�q3 ���)�����D��oWz9N"q@���ei����41��>�,�{i�����B��,Ȧ�.���E�h�3���'��!zy���nK�P��=���6��ډ��:"x9�Bx�b
�K�,������:��&�� e�ײN��㯋ej���v�,����K���YF���N��38�`���L���NI�!'���6 (
�}���u���������͕h�:��7�x���@�㉶]u��?:�78GTXFC7&O�E�г_4G��g*�]�^޳� \M��}�-�Od`�T�ɒ�w.����m)I2��P��\�Y�v������5cO�*�dRX) �n3I�q�5z�bB��e�1������d�g��Ɩaߕj����3�����~U�v�#��Q�p���752� ���R<j�ҜK�?�|�\������/8��N8�jR`�Ϣ�|X�����a�G��]x���u	k*�H2Ls����Rkl��p�i���Vs��5D�$����4�U���
��c����S�QkXl[�b��)�{0���O�� x�^wk䮎�t�\�n�|��9Ew�C�B��x��_�>U
ng�i�)�}���/�E��f
�0�8��+�z�1��Us�̀	7��1�M7�p͎,��>M$6�q�$�Tq�#��ru������G=,ƽю�A��kB�¸�Q���d>���m>}"ˀ��J })�DC/�� ��Lk��טR��ֵཽF�\�&��,XÒ�%�p�4�$����;���nrwl?��Ϣ:����<9�E�r Cj�{~ �j�kU��_�:��ğ�WL����$�G|�p����錴�١��C�a�qA"�
x��9�>9&�='��?�O�}caP���_��3���j�;��x<�����<��l� p.(�УH���`�~;�L��<a��NL-*���V7��H;�m�����'9r哢���kU��y�ښD�Q������̒�pMI'��;������Sk;���~-�e��B�*�A�Ҁ�?�ɞd��ZU���w��g�
���*m��V84\�%����y�o��O�����fS�ރ�V�v;Z��h�~Ǉ3-�\��QՃ飘uE(����bC��x%}����Y?	���\�4�B��ա�

؁���}RȥB�/WO�JN9t�W�!�K��
�r�o�+<�·��|�d*B��Y�mW��U\��@4�(21�PM�4��d�$$	|��X5��ݴg��v4.��1�lvt�_����S����(Y�O���JY�����ﺜTTZ����
���N�]|��n���l�&�@�Ւ=���3�h	��r+�S|)��ж�1��p{u���ߡ�@�:�r	�׌�����#Z�:���m��/1�̥��g���o�P�;��i֮Z �̃��q զ^j�G=ݰ&ߦ�������K'ަ	kޕ��&�s��t�<�&CK��U8hL�Wխ܀��H!�bs���\v��WhǄ�G*M�dI��Y~��u�G�N�q����$.M]1
���!:+�'��O���N��LJ?�B�쨽ڋ,G�4�R�Uz'ff�,.��yO�$��2w�K�9��4�?�����r�ʤb�Zd��LB�U�FIc����R� ���d��Q`0���gs{s\�E	��_H����g�<��`�]�-�?��nⵇ<��|H��iD|>6YX�׹�i����w���F�Fh|>��/�R���۲ݥ���i�%��sڧ<��ɗ�~��Ķ��������`z�-"�o��+���?��A�H����z����
TB�̪#���I��z��ŇN�=���l�q\��GGBa�[����T}0��+���c�]��.}Ȕ���Ѧ� tU�i3*�*��?��dA8��.�_@�'���>�WFt�i*tg�zVN;,Lߺ�>C���D��#�����%��'y(cP�]���urC����h>z��1�T�A��b^b�P���u���➹�A���D$Z��	�g���M"#�e�Mu�KxDT�� ��	��Y[@^�L�%J:��������KIEh��TE�� 	�74��,���Ӝu(�^ Q(��:�����Gʣ�m�"�}��b�mh^<ߖC�#kp�Õ��	ĸ�lY�[���C�0���Ӽ�����KƴK�f*��@�J��ة'�^X�
�<!f���UJ�W�V���_�N�rh,���w�{$�+��b]l��㍦-^_�YOd��2�('V���9~��'��l@d�QI��Ι+�����'GK�9E+�~���;59�����aTF�������ؼfI��� ��D����똕^Ee�W�$� �Y�.w�E v/E=�	�A��i�z���[-�$���2q���Z��)�u7H#zS�������G_+����<W�r4G��9Y�F�x|�YXe���K��b����.y��fQ�E�G�.'^ʏ�����Q�Ps�A5�SS{��|�.��|�3@Z�s_�]�Oj�)#{��� ԝaͯ~[�)AU<q<���҈�!]����;��y�`��[IÍ2}U_�NM�&'Lt�&7��/W?���J�.��G���2Mғ�Ǒ<%�]���/�;�4=Ё?����	��ʌ��<?)��)�������a�c�Ҙ���	 ��N$���	4�Z����Q��p쬖��u{|�,�g���\�V���!q�"��h�|�5+3���l�12�K��������&��ϴJ2�$+^lʽ<oC�׳��#U����旨����uJz�Q���\��I�i/���B7�[�'���R��9��r��(6�`q6V2����['I�56�8�d��� �_���q���fx�C����'�K[~|L��������k�h�/�Y�Xν��{�JK��Р��>\P�v%�<f^,�XD/�}�t��}52I�������&%��0�ъ<�j��/M��iˀ��6�5�6�o �-��cL���P-x�t��#@z�<Q���F�H�S�.����Cױ� ��t_�}n"Dfy��ǈ�yٺ��?���H5*0T��X��M��fQiK�ыx�1̗�@���w�aP�}�u�b8/��rĉ�'8�l0�����n�厍�R�e~���I|��Nbm�G#ER<��_"7�^��g����a��,�A˞��t�^��xg�I�l��w�)�9����A��l�t���7pv8���t��/�$�A0:C�;ݢ�Ēp����d	�� ������/���n{(g�ɔ��G�t�-m=�,Q�!���36���(SRM�����W}�����7co^8�t�o�o\�Ix���U5�<9�P������h��~�� 3a�S��d�� Z��9��v�!�j�`��
��Q3j���|����]n���M;K6�Ʉ��b&�3����{�rA�<��Rp���6T��͙H���g�E��+�1IZ������z�x���N�]gT��5>a�|��WY<"����TԸ�������]�^"a�./�n�.m�7N3�������CO��m����wnDB�em��73x<��s�����`ZL�|ҰD�|�ovk��j��I�#���l�k�V���6@bby �����)8��h��|�:���� )�f#�m���9��pz^=$���Ō���2�!��dL>�C����R�eQ3 y����q���ϖa�<�Ϟ� ���R������dc�#6��1�\�I�����3�����0��,y)ڝ:;|a��z�Q4/D><�ȓ3�g��dy0�.�B�K����%��S��TGQK��w+�`7Q��`����ZS[`����å?d���-"��nJ��`�̅�rH�L�QQs1��6�p��-�<�E-��_���\��H���S�n��I���z)kH����y5�&�vp�:�3Y׉u�(���v��5��NP�hkR���e����n«�����e�&%@ܳ%k*2B���Rx��n�S�= �Οq�ʺ�iqK���@��~�̒H.�'�����Ȱ�q��l�Z�,����"*�QA敊��Z��gGӦf��o"J��R�"����4�KZ�ʓ|`3"�R�po���t�4��| �F�I4H�
��T|��!��S��� ���7�l
Iu��ws������U#���$d�M�27�?��ݕVd�0R��z�#�"���� uƺ4������>0 Y�U)�_¯E!!п���k�V��硭��;ZϞ�g�ާ�����XQe����~�I�G��;�6�4�%[�xL�ܖ8M)�q�h�~�a�$rz�����"�!�yv��}U�®>�E]��S� =�9>���+��z��f���z>���#0�FP�x�o _+�Iem9_k"�_N�Tw��1�r��b9e��;������=��ZB*	�S���E�`���a�,e��*e��7f��6�¸?5;�������M�W�d��)7�1�LO{�mB�?��yD���ѵЉ����x��x�LyO�t(޿/��!��������^l@��Stj7���_`��@Ƀ�xh(���-������ �J�����@+	xb�&E#�Y��ע&�Z O(�%2�גқ����Z$b�;�����̒O�b����� ���=u(�W%Z|���
oll�v��"E�n���'�;�����T��O�8�Ձ�MB���q0Y��6FA��%����o��]���;��SC���T[ɧ�\����/G�`�% ۺ�?��h�e�	xsr[�Y����o�X+3l�j5��v&��h���j�sY�L�W��2�.5��5��)�E�PL�r���D��'�t�S-/s4���X�=�ՉE���a������&��Ҫ��5����+Ю2қ���v����L-�� N�.!k�����:`~�âp����v���[��H�(�������U�q�l��SyH� kA���7/��]��u��=�����b��\���q*�A�Cސ���bt2�o\� nPg�w�w�����*#4����<Y����l���/	���7w��T|�����"��VuQwX�D�Ʉ��-)Ӝ��]x�|���V�?B�Q��ۖ��S#rn���+�Zp,T���62�Qrq���e
�8��p�P��+�*Ͱ-�j}?�<�`�x��F[%@8�Gp]��q���k)�\���sì�K�"ʮ�r�����Ϧߚ�V`�=�q����V�C	�l����ߧ��l1߸�p+����fzN�M�6�6��~e:q]{[F"�Mr��3���󮋱�S
I�:��p�:8yF���+r�:X^w䓗��6`Aeio�&���������Bm�>i�m����Ń�;2XY~��X�����۳�mH4D2Y�?ۋ�>���GwE�w����۾_̩��	����TL�]u��GJL-���2���F4!�J����T��������E���[�]U��]�!ѓZf�j��`�r�Ь�����Ǯɳ�������.�
Fg<����7�2�:E�M��Dj��P�l�-����Q3��zb��qC,�յ%+�s9��B�U��*}���0�+be(��"t	�D�;O�����寯�ش#���\@Й����J���5`Oa��3NXhr-�G5	g�w�I��������[�9���=�ch"�dW�b]�����(���G�4pM���!c�����a��t�>�=E~�Bcp[��̀����a��v��b"��w=�0���Dƞ�]�?<o�!_ʰ�n/�+>����{y$[�rE�*��[��i)������񌢙�Q�$���Ʉ�A�y�7����edF���ߠ���;Tt`r�dC4�>֒���������ZB���! �	�i*ae*Z���ŁA�ٲ.:��P�����W]Oi!���QS�;�����4SC�DNn��/���1�}�^'P�P���|��C4�<ȿ5ǕtTkl���^9��P~��uK���)OA8 ��{Mċ�YV^M�$����� 7��yAjx�ͺ�#�?�Y7�y��[�t> �%�d2�x�� ��I|�k���w?���6�9���R�t�xum�	^WO�%�	���gԮ^����"mzƫL�k���^s$`C�]p�2ŏ�W�Gu�Y!{9�eV�0��?�ͼ�������ƋQ���ך�J/O�~v��l��S[C��<�J_7W�I'V�R�_{�&�ɗGwi $���9��l�淚=Bl_ d�_���h59u������l����%�Eȋ�k�z�"y�'^�\9<�'~��� ֊������&w���س����ʁ oC��5�L/��)eۍ�$���].N�% -�EԏL����5��zI�[D����G��	����	��y���f�Hh�0z�Ep��Sq���a+̄ԌD��	3n�a`̝�Y��ZX|9"�B�?by�9Ծڟy���f���Eڮ�.^�b�����(,�s�׉�5�:{/�d|�.JG���@Qf_�(���)��{ +ӆ��^'�&�U3;�������E��@X}���y[15���ä@�UV�]$�'_�&��/γf�v�E�eP"G%�d�)%Ξ|<ܞ�]F��/+7I4�yh�v�=���m	���c^e<��<��=��8���w�	�����	n�N�����sZB�������$��4�{�-T�^�Ǚ���������K�h�5b�4�>B�(&`�"Hm��A�r�>����hJi�Y+ud��3j���龎���R'��J�ȃ��;�\��b�@p4������δ�d$z�����^(M=�q-�2���~�IU��6Z�����$��_�fq��R�=��CP�¾Kұ�L�HT����9��/�OPX�n0��FK��E����MI�\gG�%�Z�f5	�X���}i����v�I�)>�<�ٓ��%����N��!J���b���Ề�z@�lN{y��$�Rc#� ��	-�N�sQ�1xQM�D�]�L�J⸚������Y����5K}��'f���ǟ�ٱĊ�۫O�*�:��K�Ǵ���fT��K�O�x�r��^���l�aa�|���_8�J��Q�/���cxKη���ʏJ�%�R>���n�g��7�e.4�>r�R�_��^k��g��A������,�k`�u��tj1��8[g'��l���`N5���TA����h�t<��\�����JΫ�r/f�A'����Q��O���5���o�74��&��h8o(�k,�+A���5����mti�,hl1��56�q�(
;MR<����DU`X�3�:   8   Ĵ���	��Z�tI�*�� 3��H��R�
O�ظ2�>���& �H�O�QS�� y��]1��S�x%�D+QlW���K�4;B�^�?�vR���'�V7O�`����4y��Y�t�B.3	*���ņ�S�B���4A�qO����D���M�`��DO�꧇�=rF8��ʋ^y�?l��pS��(��$֊wo(Q�&č5o��I�	*��e�Sg|� 4l����	��'�'Y����O�牚!̀��t萧��ʓ%ӎ9��J]�f.v�h�џl���O	��07��hy�E�{)"�ҵ)u~2�ݠ0�T ��ݺ��
��rE���NHb2`SQ�j� H��(��|�(���5A��<�`ԑ��Q��y�.Zu�'�ֹDx�U�Y��''7�̀�f�W�+ђ"<�q�%�!2P�o������?�����ݶlD�x�O��Ӊ��ْ��'e^����$M��(B�Ӝ`D Rݴ��#<�Ҁ'�MP��h�)@=H�h��U�}�iɥk�\�;Z�"<yc�4?��.Pᢁ���_=�x��aSoy�JT�'.>��?9�KL%�����>������)L�:#<ɂ�(�|Y�����+����∕g �����?�1O��r��$���w�|0����]�v量[E�'ƐMEx���M�'A)²
�A��m��/�sUÏ��W]�'|�i�;c���ˆƳ}�{�JJ#.�qOp������I�8���F	x��Hf�ݿB��JJ#<yP�6�V ��l� &I�4	5$�Rq�ȓ	Ĵ   @�?�_]H��O�#�(�ñ�3D��u�   �                                                                                                                                                                                                                                                                                                                                                                                                                                                      T   �
  �  !  �   �(  �1  �8  �>  )E  K  �Q  X  Y^  �d  �j  %q  hw  �}  s�  ;�   `� u�	����Zv)C�'ll\�0"Ez+�'J�Dlӎ���4Om���'Ԙ�5`EK� yw�:u_R����՗��HH�h��$�^�ׅD��\�DHc�!aӇ��?q��d��?��Jپ	N��$oǶmEqq�D�����`H�2�B"�e�d����u�$@�d�']�|a�^�8~�:�jZ�S�"� b�ݥf��8ë�O�X���T�]&���ƏΦ	����ٟ���֟��Iҟ��rT?��Qc�/a�J�GDF㟘��K�^��4���O>L������$s����L��N�T���/��:&��Op������I՟���R��x�����?���:��iѸf4�p�Eؚ�HO�">��4!t|ı�
]Nհ�
�3���wZ��F|B��K�b�'�L*��#N:d5�$Y
"@<ܑ���Ov���O��d�O��OV��|b�w)"�"�#m{9Y�)7gN����.��Im�Vn��Mk�H:��h�^Mn��M[��J}��1D�?|Vл�Tg�ƹI���ȟ���o��d �4c�KM�X�y��.Z�k�A��M�V���mq�NHo�1�M���Rk���t����g�E#
��!`�$5�(�MƵrn�n�K3���Q�]q�) 7oΏB��9T��Ź�4y�vEq��z1�R)1$<�e�N�&�yJ�ʏ�r*e���ԬP�Hnں�M���i}�����u�1�;d,뎁κ��X�V�x�*��<#�@��~ٌ���Ψ�ٴI�6���׋ڃgf4Q�Q �>��=Qf,��~$����O��:I�ud8+��n�4=��^!%���b�GE��
h��c�g�����X�Z(�T�&a�h����1j�Zh� �i�$6M�Od�����j7���e���p��O���%�M"c�C�R�j�*TH�O��$m>&���O�ӗxf�P��g�R��%Kǎ�]�1�S���	�2� �!��V8yBm�8��O��	V�	/h6���^�iՏ�	~�P%2r@�`҅�6��;�F �U�'�����?��OİsS��06҂q���:i�y`�'�b�'��OQ>�zׄ�Qt|�I#怑�)Vl��8Y���.RvtN�P��K�w�`��m�3��E��9��|.��F����U�
T�}�s"Oҩ�6�7�0��wǇ9X���ٱ"O�9q�X!J�ԚW��?	� |��"OrDS�M`� ��s�T���d`4"O`��!j��R�&.�C��{�"O�H���ڔ[�+��:�}��	ğJ�
)�S�Oy���>n\"���·)�<�(�v�<AG
A�u���Pe��U,��RjPv�<1��\ % ��lF*E�f)�/�i�<��]�0)�U �̣3�Ƥ�գe�<!୞�HOm�E� 56bؗ�_y�<��.ȁ��)���B5�X�ӢMP~yR��8�p>�c�4��\CQ%�"��K��x�<�.ԗ�X%�%@�,À s�Ϗp�<�J�8dN��`FK%J��0�X�<��a	�.�`wmӝUp\��(�U�<��Dh)X%H&8��T3��Ox��b��M���?��M�O�v;�j].Um�@f��?y��:����?��O᦬����f2��F\�>��ĳ�e��!�b��(v���6,�6�"?aR�T
Ŗ���ȑ�X�����@�|�����2+�Ԁ��!C�*�L�$�N�\ˑ��R�n�O0�$�O"��.M��h@��˼�{� T�m����?1����U���+ 	�+ ����h7X{�BH�O"��v��U|t�
[nX����'5�	�c���Aٴ��'�����?1�j!O|j��qC-G]�
S�.�?��u�\+c��0����"��Y�AR!�%f24P��H�P�G���gi��g[H+!nF�����
�n�U�Є[�lQccF��uw�J#fL�O�LZ��%>HY�@� ����O~����'=2����Ȟh������9���V ãf@�'�R�'��� �&z_���V'��@����|�OR~�M�1m�e	G�K�e"H�g�i���'���Q6P�%3��'��'?��1��g�6�JnS:"uVس��/ 4�9�_�N�p�+`ؘ�1��1&��	
��}FȰ����D��G܏y�>��A�Im�\p�+ֳ`�c>���ڳ����=j�e�E�Z 6`Y)�&�9Z;L7��|y2�J��?������?���$�,ɡF�z�Z�"� !��'JDXv��D8t+7�1<���H)O�Gz�O�2T��3� �)�n	JB�^�i���pw�� M�24�����\��ğL�I��u��'�"7��y��d��u�6A��������s�Q}!��O�C��D���C2�����i�uZ�|�RO�T���>�(���_:r�9�j��AY�O�L�"�чR��� �N��"O�%�a��7+0̽@�@Ÿ) ��q�|"�z�B�OQR�^����������"�6 ���`g�%zmd��KP�,�ɄR�f�I���ϧ)���I
�9Bm�mݢ/Z�� X]�*�&{���kĈQ,z΀�agXn�'���gc��v�b�Zj��r��/��8q�pG偒C�v	�6�J��.8�'"ғ:�����0�'��`*�\
�� yӈd\������?�����(��,�Qm߻t�,ь�X��a��'�n���5,Z)�2W�R��ιh��Q�0��٭�M#��?)�"8�m�Ox�CĊ3/3Z���֘?��"��Ol��׵<.�=�2�B4R�ZMs�K*/G����Ot�ӯ�R�/!d��!E3u2�OnL�SŇ�)��6�ۚeG$�B�b�� ^��$>q����>#�И$�4���3?�I�ܟ��I`�Ķ$G Uq�h
)]^�`�sl�
&�%�0�	d��ȉ���8D��D��T4Ш/����>�3ĩ�Y��cPm�:vʺ�j5��y}r�'""#֖jӲ��D�''2�'"27��TP��Ήd{RL�fǓ�kj0rW��w�� U��QD�"�!�^b1��i'��i��ʉ)I�B��O�g]�c�Ą~�T��9d(D+�@�8�b>�Z���8���v���	�_x6���
�HA��'��G�]���Y�����E�=r,�'�~��4�7�܄�H��hतk��l9W�R;(�t5�'�R"=Q�'�?�,O����a��A#��v��<�����`_�Bάo�ԟ��	���O���k� �<��A��Fj4$1'�םy��!h�-�I	>HՅsհM����(O�X�O�&��-��ϝ�J�� $�4�����MԺD�6d��j�'�ݢPmB��(O(8i��l����*� ����*�y�R�'���d9�'6�4RG�-�����X�??�Ȇ�2��=؇��U�։�Lݠ��%�tY�O0ʓ'�Ph���i���2A�AV�
>�c�
U;����<q��?љO@i ��/N$@�bO���d�yH��P� ^CQ�u�7�Lj-N|���PcQ�H����S>n��$n �[-�����j� rcID�6Ɏb��U�>"���C�9�Q�� ��O��D�M��E]V����:0��*�/,|zɗ'b�4�zc�ȹɖ.4���R�$|:����:�OP�m���v���dK!c�Zu��p��Dc�4��D޷_d�o���ȗ'\����KfݵQ�֙�cώN��|���������2`@w
=D�c����b��E� �
����n@�r��+�N��"�ғ_�<B���б� �7��L����yYT�H6��	#p@���~b��<k[�4S3"B�gS%�z~�FD�?��-�&�'��O��	�-�<a��]�a9�i᧤4b��'5��T~�-@.møMQ�����p7N���OJXo��MS��T�S����%�#5*��U��?q�n�1������䄦d�	�h�,0��hE�,=�!�D)u+|�3��a+0,!�����!�R1BP����C0'��"��]�r�!�P��@�z�>���a�Q�!�dB����[+�N�@����!�d�z̮p���&٘��$`�d��ɰ;?d�����P>i�(
�EϜH:�D�]�!��I�2�Ȣ�我l��,aE����!��]�q!s*�&W��9Yca��;�!�$���$����G�� 		���3n�!�W�G��X�E�Φ*�i��E)x��}R���~BÉ�VAl����ش<]U(�i�8�y�(,��v�`��ΗIp�(5�,D�<J&HFahH �s�+T\�Z��*D�PI%��a��e���FF1)�M'D������2�T��D�f��\x''D��s�Ɖ���\��Oߩ?��st.%�k�\F�4B�Dx,1J��ְq��L�����y��>a�4�0Ȁ<A �l�'�B��y�сM�f���5?M���rfQ�y����4B��G����iW��y��N !�P,� =�����!�yB`
,�Z�kT��,>hI 7eȑ�?9uE�E�����LZ�lE:T���&	� e�Qsvl8D����a (]xO^�o`�8R�1D��z��Z�1<���k\*"��Q�c�$D���u�#~=�Iy3BV�K��Ч�"D���w	Oc�2N��N�i��+<D�`��[�N2��JU�Őiu,,�t��<ATĊB8��Z��D�_��bB��+zF
����7D�� ,��G$(�v]��I�_ �%�"O�])�hҤfĹ"槔�F���u"O�yaQ.R�*shi�RL�,l<$��"OZ��mԤIT8�Rk(\+�	v�'�,���'��9�C��9�*��ò��
�'`��A'.gN���KE�2�#	�'=�"v!RzZ���B��
H��Փ�'������d$ �AJ��T�;�'XV���� P*���"�8z�vD��'�F�H��َG ����ŝ td"�����]n�Q?%y�c~G��� 醤[<���n*D��CBl�2WA<4����0\�zu�F<D�d�n�$51RA��*���S��4D�$c�D��m!��ӥ���3h>D����� w�iyf	�9|�`9q�(D��8�@�/7[h)�C��t�7��O*�D�)�'5M,UX����Wxf �DC��`�a	�'��:���'>mjm[h�����8�yOA24�켫��)�����W��y2*�E�vǍ �$��Ǌ��y�N�
)H��r%�yL�CB�;�y���D�:,x2OF�p1�����f��|�a
/Dۖ�Q� ��	���y/
�M�2\���D)��B�nS5�y�֫4nL����� DX�ٰ��yR��1���o��N��Ę�I��y�)G7&x�<�&C-J|�s O;��>9�ϐD?	D�Ց/�d�U���u< U[@H�|�<�2͊� ���3��S���Fi~�<����DNޕ��dK�>�iDz�<1s�7.{�Ա�ǝ�GvV=@�m�<	��.s��}�ՋAuNAp�aj�<	��ÓA�fI�4�ƥkV��;���A�'�����ąq�ƈ�u툄c2�:.�@�!��s`4H�aJmҦܚ� �Y;!�Bb��Pp��q�:i����{-!�8m�p9d�'���%�J�m!�Ö���c7�^�DfE[!ʅ�  !���̖�Y�r�(�/R8%
���Of�D�)�'f��3�R�gB0c�NC���a�'�� cN�8��-p���3q�̫�'�l1�:A� p�d�&eO6�+�'��p�c�R��(�IZ�Q��!R�'���4L��`�N�`�HXC��8+�'�ޱaT�ǂD_`��%A4S�y�.O�z��'/�Q�׮Yu�4�c�^2(�x���'�T���E%��℘��Ek�'����MI�7(&0�&f�)~A��p�'D�a��Our�s�*G�61�'�8��e�l0���ŭ�j���n�9���<%�M�~�	(T+?���>��HR
�N�"(أ����%g=D�����B���E�,,��č9D���R�ثS:�A�)ː�����F�<��❗5Ը@QS�K�{o5�z�<)wl�<�����D=ws�U�˞z�'4�`���U�3��R1�������EN]&�!��X�!/�Բ�'�@Վ=�$�1�!��
a*�a��*t��`��,ߌI�!�Ċ�F�1�g�ք�N�i2C��!��@L���WOP�Z��]X�i�3�!��ͦ:��p�#-����p�� �Re�8�O?�"�	�/}��	�	E"�ry��^�<�gB��$�LZФ��,���Y�<� DD`��ۙG��k��;c[� �"O��#���CCd�A&��`]Ԍ��"O��zPE=����C,px"O�����D�x���0Z.qڗ\�-(�O����m��rT��p4��5K��"Ov��ԁǌk̠��H�6Jς��"O�q�B��c��
bH��L�����"OȽ�� \A�q���v�.�hQ"O� ATQ�<4^�:q�L��ഓg�'Ih�'����1m�{���؂̒2p)�eR�'[�y�q�M2w��鱂)WZHL��'묌d�[pL �b����|mh�'�^��fG=o���a�o}9���'�葠w!0�����J�vc*���'��p���d��CEmZ�n>�uی��L�;�Q?�Qi��� i�͇D���pF.,D��c�Т:�0�h«)e�Z%���)D�|���õY�H�����IZ�H&5D�\iD�6x%niS�A�N�t}y�-D��s�'K� 
�apaý_���Rn1D��;�n��-��e��� �f��i��E�O��#5�)�]$��@�0�d}�7�L w��|q
�'@bd2���~�2���t�h�p
�'�f�G
��oJ�p4�+kE0}a
�'�� �6@[s����$M���1�'�`��%�½vEة���]+(�T9
�'�BYW(	�Ycf�C  I� ��)X*O�pbB�'}�- �����cԄ9��+
�'�R@p�"�2r�)*t#,b��P�	�'�>%�3���g'�Ty@���Uh�1B�'�R !�6-c�Уh�Q����'�
L�ơǡXU*eo�2GxN|��8�����Zq�11�E�&�iƥ�s�$���%{QbV�(6p�ҩ�3����xU���*�5[\=!�P&�d��.�Tr"B_/Xs����B�I9"x��Y���A%�+)�P5ң*��58xq��'`N��JD�^�(���
�$J���E{�(�'�����`���R\�a�-���@�"OXq�B	�D`�(� �R;�l�"Ov ӄ�6c�h�XH�I4&�"O^�;���m�hY�f�>O+�@)"O������F�T飇I�%$ƈ��"O�`#PH�"kxЗ��#8�)��'z
�э��S�1��۱�ǌ $����És7���ȓx�	���=i�, ���-%T<��S�(�
e�]�[vܐ@�K-K0��;�*8��26����oҨd���ȓ/4��V# n��Y8�cOlɆ�F������&k�T� ��Y�F�'gRL�
�[���!}_��!A�<���ȓD+6 ���7*i��s��ԮH��L�ȓ>�:%Ӈ`F�?b4,���܅wla��c��娄��SĞ�y��R�2)�ȓL02U�v
[$'r�G��;n�����	�Ad�I0�]���� �ȱ���v> C�Ʉ+���XG"�@'��q�/�8$�C�I(���Z��ZRK( ��m%p��B�I8|p^a�0H�$k25�W���Z�C��$XI�`s��,ʶ�8V@O<OW@B�I �nx�q�\n���N��P�ʣ=��/ZI�O&�����B	�9c )��ۘ=��'���A-�!j��@I@�آ`w<!Y�'Z#��_\] ���LlA3��� ��s� qU�80o��1���4"O�E#qG�AĤ���Я)�Th��"O>�qq텑:��,ݗ�N�[d�'(��R���ӵx���A!c��A7���B��`"���6�$�z'�O�~9�`Eҽ�:Ɇ�s�y�"�S	zh��R:
��ȓe5c��C�&Q�L��e�b� M��G���X6�'2}֬���[�%�\���^�J`bI�v�l�[�AH��1�'�&�H�7���JԿ >&m�X<�A��*�Fu u��7@� 0ఇ]�p�d���*�����Ht�P���S�F�؄�lczm�R��$�4���NI.Ѳ���vζ�x�*���@T�1%�%[\`��I�Z�����:lDd�d�P��s��	^B�ɤi��"�A,�����uvC��4p�0��F�V!�A{KN�L�,B���}u��5o�ȝ�uI�+��C䉤"����-�P
�M*�h޺:
�C�	�;,St�\� �B�*�L�b?ў ��1�j����9X��ڣ� 2Vw�a�ȓPE @�sf%I����� �����me���mED��/B @��=�ȓS$��;�T=!��л�NA;sN �ȓ~~����H���ik�Dؼ[�Xфȓg�bHj&��M1�}��	D:c[v��I�f"<E�$ɟs��-iE�X�rX��mW!�ʒsLAg��#e���F��K!�kf|��ׯ��6}��C#B�!��
�(x��d�e6&A�b�+�!�צ^���y�	�:+�(�gbO,u!��[ݛ����]��*��Ŭ'Zџ|��h���M��j�.�?��O"�����(�`��� ^�tM"�Qt�2��?��q<Ph��� 4� 8�)�Y��O�$�k�D��8sHX�bP��BQ0���[<@NX������D�|�Aՠ�R��7!���c�+�A�'�6���?)����Ώ�X{0a��I�ظ��N��D�O��$I���+�ǉ�h[�Ʉn�� �'�I�J�9���(q~Ԑ�fgO��e��a��B��	�.O��'���v��hկЪ[l�I`�)+!d����^��}�6@���R�����p��S�E��2���ڸ"�
w$�'"�\�Q`�X��y"ğ7D(�Z�ρ�5HNU(���"(�)���z�'^��ug�M�~���8��	�l��Γs5���I���'���Ԇ�d�	U���j�P6쑸�!�[-J�q���ׂj��x�*X�$�ўH��i��g������>�z4�TΒ�q�4����O��� p��� �����O(���P��ث_��kp([�i-q�JBW̶�O2��D}8
��?#<)�oV�tҺݛȈ(I�������� w2���sm�Gp��g�'ڄpB-_<Fm�{�t��O�x��'6b�	�<�'ظ(̅��	1��	y���Q�<1���eĴh�-�b
8)�o�ПT
��4�X�$�<�s��5N�s���8vɠ=�Ł����R�˸p�@p0��?�������?Q�O�NhA�&�0Om�h��Ԁ �|��B3u�d�`��΅AÌ���S#E�l���ft=�we?;J�C�-ԯY�Q4��[؞��5��O�������p����BĻ%S��"C��Ob�=���$�N��Ki�'*d�x��ֺZ�!�D���"@�$=�T���LT-~��I��M����'c�H*M?��8K'�,��
�HG�0CG�?D���bZ�G��!�c�:]v��%�<D�\JAcD<�ꁺ�Mݿ{�Hܡ�C?D��k`�\��d\۲nF��8���0D�ر4�V1!@0�A��<B���� $D��ZUMM4}��)
8Z]Pa#��t��#<��Z 1�+���@a��AS-Fˈ��F"OD� �W	p�J��ʗ 	�L��"OZ�pae�%\E��V�v�+"O� $�a�D&'���	��S�
�Ip"Or�z'	$x1:؇�ќ`ɶ� "O^)@wK�M4>q92j�9(&}��J��O,�}��#G"K.I��t� �Y��Շȓ>��B�dR*���k��M,����E��C0d�����۪���}T�M 6�O>I���¢j��dx�ȓ	��$��N�YĤ�8v!����m���[�$3{�t�I�3\����	J�,��d�R�l�yS�
�Ob�d� 3#:!�� 5�dp��)��Yn  ��<2!���\o�����Y�;�)����X!�$�r��mZ'�/����0J��.-!��w,��[��Y� �4�p5*>dџ\(sd��M����?��O���+ �\�2�IR/�Cv�@����"�"��?1��1�|
������!��8��׾}��U��ۈO�X�x�Ord@�c��>(��?P�P���΂�ᓯ�
X��'H���qt��=h�6C��18��p�4�	)_�Y�BM̵p�"���Jy��X�GD�a)��){ ����eH�����O��D%��?��'��3ŋjW��H����yZÓ�hO�\s�j�1"����a��%�&��`�BO��҈��"J���鰔��#ތ�Q�*ـ��I{?�
�T>�ɢP$��%(S�"��x�ۿM[��K��Ia~&>}�H� ��	���'�	W��"X�ҝ�C>$�ء��/}r*���E��'�EP��U�s�Me��(�6��57� ԥO�P�O�ꃑ>)�V?y�ȗ���g'R�0��+C��dS�[�pE�t 	VS�	���1@&�)�� .�B�ܰ��Ƀ��ɻ3���'	�7M��>�S!߭u�r�$��o�ɇy�(ҧE��1g��`�Ā��+��k�	�t��4�'�Z\	H���<9���r~�'��J����"�⡱��]�dTj��$[��㗦ǟ ��-��>%��U�~�
{��\'2�p�"���OX-��'�&�A�O�s�܊Ub�����ED��ə7a�80��Q0��OT��aoJ\�����^?\��r�<S������.�)���<}0��G�N;�R�lZ埀$��@���I_�ܴ1����Hw6���"ϡF���'E�'�ў��;��:�W�u�:\(4�@���y'�xD{���a޶w�X��q'Z�Qr8�����yrE�p\.m�bD�N��8@���yb�T�e/�p�2�W���"7�y"-��d��`���m�2�yRl��It�KR �Q�lRv��y�߀keFBG�4��-��D��y��_���&A�WC0� G٫�y��)�T!҅-	�P�����yr�Bm�Ěd����P��ʢ�yrL�f�A@��$�%l8�Ox9��O�{�'O<k(h�@` I@��	�'��Mh�l@6A>l]��`��'�aӉ}�HE�z�~�2��H1���u  �|�lD(m�\�$LO�W��H�j%*n�34�¾_����������g#u��<Z�JB�c���m;k�`��Ϥk�Ę#'_�iJe
*�R̌���M�/f�u�Q'W����0���)�:�i!Ӻ<��3�V�ga4��Hݛ�M��遰;~���Y)>	$���
�=�r�'����%�i�An��+:�H��HU0.K�)r�Z?�"����Pu���d#��g�}3ҥ.�D�fX���bG�uq�Q����u�DQ�V�'肉�U�9���x�e���le%�@3��O����O��?��L��TR�HK/Yb*�ؤiR4v�,�	mX��DJ��\��T�U�S5n��?O��Gy�gۯ@���`��SA��i��'h��n����ȟxC�Ϻ&��\������ğ�N��Q�v���N\&%�x1v�܄[�0|+v��7M��Q[�Kp�l��6��w̧B�,ٹ�I�O���t@��a� p��ѕA��A�{'�}{5/H�'%�]v�R+�$�>�Dk@��y��&]����0-ø�^�!�?xj��d:?9c*�ٟ�>�D�O�6��(g�~�S3˗0yL�s���;6�*��ē6���P�Ե$�,p�R�W�i�O��Gz�O�V�sˆ�R^r�;��4VK�P��۱)V��۷�	��?���?��QZ�.�O&��w>U(�!����x�lD�\o�ǉWJ����ꂐ7����X�P�&G�?�Q�H�� R� egE�tʚ	R㒂 ���#�Pt��z�n�=]nC�cӪd���B�'�4�Q��G�$I�)����$���u�C�?1�����h�r���-3���Ջ�7bY��*Z��y�:/6�����!q&P ����)и'��6��O�˓'��I��W?�n��qe�޿B�j�av$�5�(!���?頭��?1����T�R#9�BMq"����yAMϰX*��L�1M館�Q�S�;X�"C���@����ˤ^��0v�Ɩs��CM�I�H�%dߒT]��1���f�'w �����?�OR�F@V���m��	�!�r��1���O���$�`>�)�w.ضF𴬁`DE-�����LT,���1M�����C*o^����d�O*�5��QR�i!B�';����l�m���ё�9 ��QiÉd������?����?I�y*��I�ʩ#%ϦC��U��i�O�����)�ӧ[����T�����|�j;s�Ov%�P�'1O��R�p7���]�S���?Cp�)�3"O�}#��(M��Q���*"B�HRG�'\ʢ<��K;�`r�,�.5� �o�@?�	�(�t� �O�4�XPB��A�Z��%�ȓ�Y0�ks�i	f�$3ZP4�ȓ"F�ɡ���	����"&*R�9�ȓA ���ɒR�R�E�B����h�b��ўQ=��Pǩ
 Z4��2�e҆���{��03��)C� �ȓ/ �}��,ڮR�^uH���Fڍ�ȓ?ځ����-B<h�M���T%��5������l<�P˓�(�����\��1
���'�4l읽I�C�ɧZ"\2��7x�z��ޅGbDC�44�HL@3��.i��Y`a[��B�ɓj_��#�ř)��8�Χ#�B�ɪ�k�ز#/
�e�Q�Z��B�	=SG`p�򌊲Q�M��j�X}�B�3V����,`T�}ɒ��a��B�	qK~e:��)��h��M�jB��"\��lA��@,&Ѽ���H��	"B�	,\�5����k3�X�OV�4�B䉴
Ȝzb�_i&��R#�� �B䉙`�sc��U!T)�`ՕGo�B�I�=�L�2��xP�8��O%z!vB�ɱ42�0�"��7@8-0RL� �,B�I�L!�tI+�9���y��!v��B�I�[/\H�3k�j�ʑ���@+	6&B�ɑ2�~���W�&ݴ���J�>��B�IFY��ha擿}���I8X�B��x{�Ih�.?\e�葻~jhB�I�5͞���!81�>��`�ӣbp�B�7ɮ%s���MCV�ɔ.ͅ�fB䉸`{>�+���bA��D��ئC��U)S��͸\&���b�ίd�PB䉄J��|��d�6h&��S�ha<B�I�AE�1�0�Z)r;\��'Ə�2YB�ɩP���@ ����<� �#�M�B�I.�@�f�&h��͝5q�B�ɨL.4�(NL8� :�$K	w�hB�	
J� |K��y:f��GFA %�!���J�4��!��S��	ʔ���!�DH*"�-�6ŖT̓3�I�3�!�d�Ǣ�0�5F�}J�җ�!�ė"��4Z� �K��2g�}�!�D�|򖘣���=�ցJb#�}G!�%
�4���#a�T�W��)E!�>Y�H������1d�F�y2!�ę��Jy�OO�I����85&!��A�WJq;k�:X+zT:5 ��!��c0�@�g%f��S$!�� 6QK�,ݖ`��!��M�n%ѣ"O���C[eĎ �E�#3�F%!�"Oΰ�A��&�Zt�tdXa���˂"ODu�dE��3�h\��c�61VY�"ObtX0L�m����3���%#�4�T"Or���G�I��X��w��	�"O��h���>��^$#Ԏ�q7"Ovq�!�N�,��K��X�A&\u��"O�Z��J�"�.T:5K�z
�@"O��@�:X�v|�͙2���"O(�p���_QZa:���e���HV"O�Pb��ʶ?���(V2D^,F"O<�9�Bˣd�����`2�:'"O� �t
Ә�|�PB��0����R"O�q뤩]^`Da�2o��QsFYC�"O�-h�mƀ! �$k1�#/{�}�g"OAʥ��	T߾mZ'M@�l����"O�E�.E>����ʠ+���"�"O��@�*B%sK|(��AN,(��,i�"O��5fڲN�L��сW�=�5��"OxaH���@z��`��,0P<{G"O�"qb��gК�(��O�"��"O��P�#H_�0�"�R'n�֝h�"O�$hP�D�w=��*TMW2<�Tl�"Oa�f�1JE"��Uj#C���"O�����ǫe|:J�cכ]�B�["O��!�#��XTi�%��B���a�"O�P  dS�Sx�ݡU�B;}*YI�"OD=�5)L�����n�x�M�""OȈ�)O�y��ȩUk�;A��{w"O
�(!#<�Dȧ녘Wr9��"O��*�'���V�P���
8`&"O<q���Gn<MU%��y���j&"O���V�L4E�]ƤV8$-["O I+ ����h1�ƌ�m+���"O~�C#�D+.
�!Z��\�a"O�Y��D�n��UΔf��0"O"d��(
��4΀�)���P"OZ9a��C��E��j	S��y�"O2mZ���0B��<�t�,��5"Or�8��E>bV��PWH��V(�!�r"O@E0��L�4�����>4�A@�"Oz�cA�xl��bE
C!�� "OL��T��r�,	��n���7"O�)�F�,H����P�Q>\�a"O٪�`�uD(���BH9��T"O&�b����0��Ƶ(��,�"O.i�ECؚ����p̘(l��q"Ol ��g"���� ߂,;�՘�"O��0�l�P��]�����-!�$��M~FMa�˙	%�Î�n!��V2�ar"\�&��8����1T!�D�*2�}�5�U7hx�M�̐,Y1!���5tc�ٻ�,�TYp�)p��<"!�����
 IL�xޞ�� O�82N"B�I?&p��R��1U2(�>[B�	5o�\�i�����'Zz��C䉎SGz���ҏV/2��4oٲ%�C�I*RX|5�F-'7}a"�)גt�C��o$�M)C�]�O�"Z����p�C䉪48���gmE�)�ȵ w�G�K�>B䉙3hTqe��'���c��УB� B�I6$��uk���+��pd.�`�B�	7b��|�D%ZM,�EabB��;�B�)� �2��:��i���	S64��B"O����P�RA�@ a�,x�5a�"O�l*D�e��%"����"O|T���S-Ud�q�*D�B���"OЉ1S�͢�*���A�e@�"O1P���j	�D��)sl�i�"O��S2,�@���^�-��iX7"O2�K&D
��Uj&眱2���@�"O TXp@�#i}2h���s+��Z	�'A�ST�ܡq��C�A��(��	�'��`c!F�1E,�x��̦6'���'��dď�!�zg�� 4KR�1�'6u��K��z��V�2
F���'ԡ{R���=�FF��$��1��'�0|s�c�)sdMn�W�yq�'���>V�b�2GjJ~�8
�'��	��H;qs�[�W]ƼP	�'�R�*�N����%a�>:H���'��,��=:� �����u"���'��t�<_���P�!���r�'���ړ-�-g�ҝ: !��%o�QP�'�jрw����:P�ґl��'�z��ˈjB|����lM
%��'��8�"JC�T9��LM�k��A��'E�s©ڦu��EzpC�l�DmZ�':���(['t��O�*Y�l��'G`��QhQ�G���ϘP���q�'>��֮�P���0'@ў�ȹ��'��xkb��9D��iF�\����s
�'�ȣ��C�0��� �6K�'��]q�-ߍ���T�ђ{&I��'��x+��k����T�])H5�8��'�,<�j�=z�	$�߸/�μY�'� \�ցͪ�.�:�!��c�'�\��3
JX�=�Ao
<o���'|���#/�0�t�p���L3��B�'�u�Ռ�1j��X8!�H!W��I�'q<��_0�쵐gL
�O��i�'%�P�p��:\����=:0�
�'�葘ԏ��\e����OV�l,H�	�'&��@�$�,Z�χ�2$͐
�',��b$9L��lPf��%,�����'Ʉ��0��FQ�͋u��\�N��
�'"�}U�V��H�4D��B8���'�\Uj1`	܂"�k;|?:ec�'���[�f�%��鹓��kf:���'���y�!��#I��hCd �h��5��'��)���J$��cf�N�Z����'�>�ICfW!f�VL�E �W�*�'�(d9G�ޡG�	"E��I� ���'�$�17섁�$��O��IW,}�'[,����|�H�*��8:`$A�'1>�	�'w�tp���(L��'��M�'a�l���2���w���	�'��Pv�ܬlu�-#R�Z
!�����'\��#�JN�<�Ȱ����'��u���[�/��$
��P>�
T��'yΩ��@p� 9A�Ū
l(�Q�'��b�)�*}�	V%�8��'{������5���{"�9OB���'>:��dϙ�JE����@�ص��'O,�����V�1�1-��Q��'�Hd#��U�B�$0��)ό#�.m3�'�1S�I�,��Ѣ�+$:��	��� �4+*t�|���7D� t�"O��	�bH5q]�u�2�X�U���i"Ona$^�J�Qw ��>�x骤"O`X���5
.U�F Y<���f"O����7.&="�	�C�X��"OX�s�L�l����d.Q�N�����"O ����˧b��80��$4���"Oxd�fV.�n��B��3|x�I�"Oz���ԧv��y�Dj�+b�֭�"O��)Pǂ�\3T��	�"z��<��"O�œ��
�6N��ͽ}�V�"O���"�	��܉K_;"�ʑ�"OΨ!ӣ��R=����=)XP�e"Od�P�P_���f�h�$	�c"O�%"w�P	������6vvycb"OFM�n�"<P�b�e��fp���"O6��&D��*\a���Pcv�"OTY �"A�"-�I)6F,!i�X�"O4�`b���b�8[&cƧz�^��S"O����� )��haA׽G�x��"O���a�,�N��O{�PXSs"O��B�����MY�g~M)%��E��!qE�AC��{�߄r��y�_�KB)�!�͝�`Q4����y��#c���b#�U9đQRhS
�y�C�zQ��[3Aޟ!�ʔ�E���y")��<|��1�1B�źG*ƍ�yR���L?�Y�7�#m йإ� �y�O�Wi����[�E@š=�yr��Mv���mU�Q@L�k�
�y"�F7�=�S�(�`a$E�#�y���!�$5�w�̠6�D<j#�0�y�ŉΥxb�:-�L�gT`�<� �:K�H1bg�YwHTZ���P�<��!��#�QR��KP�#RCAd�<���	�Қy�s"��(��C��a�<	��N����R D���h��a�<1#�ITX*�@�ep�N�}�<�h/[(�p�i{��sw�Rv�<��'��\�<|�DkU���8�&�y�<y��J�zs�T�c �"pg@[�<�׎>S�9��섍.��*ӏ�W�<1�	أb���o֮ɸ
T�P�<�4��,pB�E�1��mt��[�͙S�<i�E��ѣ@��B�9*U�l�<Y��f�� hy���b�D_g�<ِ���x��	�n��B�*Ca�<!4 ��k`��Qg[�0-��+��@z�<�DA^kβ�+S�Ȏz�X�p'̓y�<�`8P����Uo�\4j\�C'�_�<���~����t��~�LI#��\�<1��Z!y�>a���J�M�(Xh�%�Z�<��c�.5ZH(j�D�~C����m�<�vς�Z(|���R�fX���i�<�# \�2.p�a��	J< ��I	l�<1�GD�=����@�C Yt��[�p�<�'��x�BD*�	В8C.A�ŀf�<��Fߏ~��PBb�U�|�����Ox�<�eɂD�@���^�_�T�Cd�v�<��&�q��!�C�
�j��#.�n�<��
e�D��pB_y�l����A�<��G� z��cAA� ��Kw
g�<Y0͎,O��ꓢ�
) Re�k�<ᑄI)-�����a߹8��� e�<ـ��ق���D�XC������<� 襡ǧ,�1b�Ú`��f"O�q�Rb��Na���-E	X�����"O*��͟U�"�M��FL��C"OBl� r�>�@�#�"u�I��"O4Pa��%!O mѡ�K"����"O���mH!H���ن~mx<�@"O Ej5D *���*K'R|8i�"O��:AD]�I:5IU��	u"O��CR	�{Xd�V�$̦�hV"O�襂��B0A� �۵g6�-c�"O��JTN���$�� /Hk�"O  a (���.IH��,"�X�s"O��*p�]F�Q���^ls�"O�ɓ��9=B�9��F�,`0��f"O��HՅy�(��D��!;V"O���c_�%5�[��e�� #"O�a4c�\�z0
�O�flΈ+b"O(|�7��G�椺�A�Hɒt�"O�uJ�"�nXgkʋS���聬)D�t9$��(I	+�!^	�R��u�:D�\�œ4��MP�䉼2
T����8D��q�%Z,D1x�fLȄ2PTq�%D��u�ܷY�0Q�&�K~�|0��5D�i��%Zӊ�����a�0�&4D��b6aT��B��hé��(�vO'D��JU��7����"�-9�L�E)T�T���ul�E�	S��(�"OP���ڱj��#���W>����"Or��m�tH�����"2~@�"O�I���#N�6����ӶuZe��"O"�B�i�&O�PDpQe��j���"OZ�	􄎝Wi.d�����~�[W"Oν�c�� ���Ά�`X[�"O���S�
0/����k�4v�b"O�p�ޞ^x�D�C �|�kS"O��%�_���pg��^��J$"Oz�p�FS�@�$�G��6c��2a"O"�3B��9�\���D;Q"O����[hs�,�V���7�H�""O*�Ï�%�aj_�DPȂ"OV�(f�U,9z�; N4>�^m�"OJő&*@�9�����ԓu��$�p"O��fo�!q��%@�dV�4�X�ȧ"O��ؔk�Au���a�%&w�Y�"O���F
?%���4s1L�>!���ŅۆX��$*WH�>8D���"O*q
A(�'�Q)��5���"O9`�LV(&D�h�Ȝ�w��"O�1�(�L�����AQ�X�"OH���y��U�7G۬`VF{�"O�q��`��x�E���@�T�1�"O�īF�-|<�Q4�څH�����"O�!sc�Ք |�q��
`���"OԬ� U2$���k�@�]԰P*!"OHi�E�^�i��[^�p���"O��#Go�u�ؚ��j=�Eا"Oʈ�F�;Ĭi�a�M(���"O���ŘqyLh�"+՛0���"ORDɕj�K*�d3wC�Ll �"O���.Z;�LI�emH��KD.�y�$��q�|���'�gU�A��Ą�yR@���{���"���ɟ	�yTjv	" )�R��F���yF	)R�	s ħTZ�!	]��y
� dȢPnD���J!��#3�<9"OD�P\ �ā(§��x=��҄"OvaYu�?[j �A蚙N5��"O�ٻ�M̮Gx���Y�	\��"O``���<���%cm$���"O�����+8Rt����>lo��9�"O��0�J�_�mq�/�KkFh��"O
U���"|?���bɶb��w"O ]���Di�m Ќ�P�±y"O
D"�C*�t��S���i��"Op5�4� uJ1��,÷&4�f"O��b�C�'XߢYj�閪/3$�@�"O�=���%���c�WT�D���"O�,k�bH6�qs&B΁�(�"O����K��.Z�����E�Y�:Q��"O����OH9�P4�`�+4�\�s�"O�-H��)=Q�K��?*g�u10"O�y���ߺ{w�p�3���5����w"OT�
��K�
��1�)@�ٙ1"Ofy�6 �(aCv��3x�L1"O���iL�lƤ� Æ�klA1�"O�]��@RWR����5;���"Oh�A$��)�<�s���
uqT"OĻ6�U#m)j����ܘXXHȩ�"O걩�eAbx`�5��Xu�eB�"O$��5�D5���a��@�%�h K"OD`�Z- ��I�v$�3e�xS"O68+��*$�,`A$�<?�4Pq�"O�%�G�9�*MM	Mۢ�3�"OԐ(�܍|��0��n^0.�
���"O�|����,R�E���єg�<�3"O0���V?T�PM��)"Is��X�"O6p@VA$Y0��2)�Rj���"OJ��Q�é?.I�)wNt�Q�"O��#��,�"�@�2O$���"O:q��0W��A��Ym�rd��"O�}9A����T��+��F���V"Oj�ѕ#t�6YxqA_(��|�&"O��ؓl�x�^��� �����"O x��ϋ�7�:�ص&àM�F�I�"O�ii���.3�z,���V�� ��U"O�q6$�0. X�W����`:r"O��Ag �4F㦉J�n%jQg"O����ϑK��0�7�8f2�qr"O���1  4@(L���6n�r"O�� �d�=+ѲmÐ�R?3����"O��[l��� g�!b�j� "O�QS�ŉW7T��tF��[R��h�"O���'D�+"�1v�<#L��[B"O��Hb�H�huz��E)H$\dHq"O�x�V�_�'��#"�U|:�3�"O���	51$�s��7wJ��1v"ORaӱ*�K]�!�	�2v�l�'"Ox	��K�8)�� �(Ͻ�<H�"O�98�Ra��Pqf�"W���
�"O�I��N��{�f�+e{ldj�"OU"��E�4z���+�lk�"O��ɰI���j���
^
6k�7�%D�|��7|��� �V'n����F)D��qaH��>�R�j�?=jJ�bU+)D�xsl��1�V��gG8_J@��D*D���a�;Sd�㖋��r�(t���%D�Hf�\�-���W�8:JI��h D�\����oj�5��JٻRBF�!3D�� \���h��E�X	ѷ�/(h��{c"OX���A%v^(���`�M��4"O���q��B��`P��O�%��ٚ�"O���2�L8N�|d��V,�ƅ�7"O�<����f�]�í�X�h���"O��[��0x�D�W�j��"O�Q�ÐF��B⍝B�T�S�"O8$A5�Z��D� w���T���A"O���bȑ=vî�3�L\���IS"O�x�rKO	\c�	R7n0jdP�"O�����e�	�6-<Z��$��"O���2���z%/,� HgB"�y����-Tv�8����D�*� �y�L��H�Pm�9cZ�2o���y���5(��Ug¥0蝲g�6�y�ܦ��@y� [�r���W��y��B>$�t��#a\�DN,
f�(�y2�˸H�,��� ߺ}朽ł��y2��>hA���RB��c@L!1!��y�.��S5�}A������jG�-�y"��{��p��S�*}�̔��yb�׏�Zmb2n�5aK8ԩV����ybkO�>rK��G�N���hűnW̄ȓ���g�K;'�^%qXX@��"D� ��-��V�N1�R� zT ��F>D�4����^D ���_oV��`oR#;n�����M2Ϟ��b�hx�4*�AG�6DbU��ʅ/5��� UF#D����+� tl�vbB76H�(�F6D�T���Ɔ�Ը�U/$D�lhG�?D��!�艁k#�e�4 Ųw0;�F9D�|)���	v����V3��Ebg�*D�hPm�Ns`a�5+��b��{RE>D���[y�{����2)�UWO:D�H�E���@��ɢ��C�Jnɢ7�5D����Ǆl���P�OBT�PqPL.D��k�(E�e�e��!T&�F�P��-D��y�iZ;����$��z����ӧ+D��a��U4h�{��A*n@�Sm'D�I�bN�T�< "B�:��A&D�,x�j��]hؠ�]#K�]0��7D�yE�Όb@��D�(��0D�px�� Z�<��d�Ox�(2'/D��C5�Z�;BV�A��I%]ν �D:D�Hc�N�b�ȸA���,ƑY�$D�\�5A��nd"��(��y�#e"D�Q�w#~���.�7Q@ف��!D���.�2��"cO�0����<D���!�?77H��@$]8��%�:D��@w3�:;���=F*ఢ $D�������a��)�B����'D��X�4�\z��#o1a��I2D�\���.��!����ek2@b>D�LI�D
`<lQ�c�,�J�(��<D�h�1Ə,�8�طf	>��J` %D�|��˨@�j:Ae���p��%D�v��u@cdN�P91f��$* 0B�	#0iy��/K'p0	�j�	L6&B�I"0����f��Wm��H���C�I�v8�
W��.� ]1F)w��C�	�M|h�7��0f��H�u� �nPTB�	+��$kG-�ia�*�M�7BB�I3%��A&dN���ʳ�_.0�\C�	<L�`��Q^K��y�i]�[WC䉣`0q���7#���Y%��2��B�)� ��x�Ʉ5m�xm dj��Z"O��ؤ�Kkt��W#�&<K��;p"Oh�J�	�A��3�C^�/"ly"O} u��:Ů	Dl�+%*L�1�"OҔZ������k �^�#PXX'"O\x�e��-~I< 0퓜d\���"O�8@�DK
���LN!?�b��7"O�ȕ(WIΑ�Q���"����"O��񬓑�H�v���}���"O詪 F)�L��D��n|.���"Ol�� ؈{��z%�C�V��6"O��[��(6@�:����!}��!"O�;0J+S:�k�.��RH� � "O��R`"��Ⱥ�
@F�s�"O
5z�׻i�0횳NZ*�赠�"O � �- 4��s��9�J8k�"O���.[�Q X�:3%�{c(�H�"O�58d��*�R%�"�	Q���sE"O�$2Q�Y�(�X��`͢UYx�"OZ��r��`v4x�NSD��ze"O���r7(M �#7�L�}	�)��"O,�Ie�-�F�j���s�E"O2��#JÞ#��H�6	C�Mˁ"OD�!�&؎~�zݩ��߃7E�jf"O�$0�K<K���j"�i�V�
!"OZ#d�;Q>0hS��*�2�� "O|��)��z��`G� �$�;�"O�d�С[)�^�� )�<C"O�c�0��w�>P����"O���$��	%"�q��ߴ���"O��x��Eªy���g� IY�"Ov���MX�v����Q ��<p"On�+q��F�&��0�Ag�8�8u"O��x��Ԑ{�d��v�9"O��sgR��ݹ��gr0ԸW"Oll����^���8�#��g���"OB�1-����kS�^�^ �"O40`�.s�.1�de�=
�A�"Oh�a'
�a���a�$\��"O�u �'��@R�eBǆ� �^x"O����
��X\s&��~~��3"O�,r�R�%�MA3�3/y�ԱV"OH�9.].6f�F�M(99���"O��AV�]�;�u��+0���"Ot�F���Ub@u�.	%C�Sw"O\i���-'�h���Cy?�
�"O|��@#�x,)�QM�)2"Of�ᅠB0j�"�)I�IA�"O�D[F��'p:���A���P�"O���p��;] ��� ��F0����"O�ԩAI�-U��5��·@��p��"O�}3�O�-�r}���R5���u"O��M� 4vF}� 3sn�q�"O��S���*�|�FdGQZ00"O.i�@��A��x�a>)E�9��"O�q�0���.�D��uoF_?��y�"O
@�$샨L�L��6Y+tF"O�U2���mҨ�Z���-#tL c"O��K" Du���FH�1���&"O���� C X�����.p�9�"O�0�Gܫ� ����5S����"O ��e_8��תS+Q��w"Ol@A� /2, �n�'1��M3�7D�d"A�����A���9g���D�4D�� 2� �)��00Q�Ŕ�`(��"Ol��e RW�1���jd*"O��S��U$�T�R
�xs�a�Q"O6M@Ҏ�+�� q�NQ��D"O��ҋ��D��6nS:e6����"O ���9��s��Yh3HQ�a"O�|Y����>���
(d+jT�3"OH�F�ȇ6d�1a�~#ܙQ�"Oz ��ɨh���1���7��Dp "O<[FF�)�|}T��#I�����"OʵRb�לK$��!@�Ĥc'�5p�"O��֊�t���0���.\� ,;"OJ�%��_�~`�hW�f��"O" �'HB<g�0Y��	a:X��"O��`"Z diɲ�B�s[^�R�"OP�ssCP
i��yq�%�@I Lȶ"OPU ���G��0�dM�R����"O`��w��R��B�U�h��0"O�t��*Hl�x��+^!}OйВ"OB�Pҏ�� at��엂3���"O�УsDڐ5�0����	*f0�O����N���Ճ{gู�����!���^`�𠫇L�U���}�!���C�J���.�8@�\R��ЎY�!�$�8#�jI�֏@���!��<H�!�d8H(���e��[ՆH���^�9'!�$��#����f�7�� 3�@�,�!��L 3I�P�T�O�OF* ���_��!�D�3j���wm�5 5����G�s�!��M�F{�%����9NfI;v��%F!�D�� ���õ��2(1�Ń��P"7�!�$E�L��ْ��T~�a�
�*�!�G�<h��SB��Z�hq���G�!��R)�T��-�:S�|	y@�:�!�d�T(|���Y�*i�'�Ϳ^�!�@47h�驦�T!\�
Q��ԙ+!�dg� ��ퟛA���3NIE!��!&� �)��B�y�\��@k�w�!�d�<S���@�A��l˪�.�20J3"O���	�P�]y�D$��	�"O${5L�\��)d셕c��1P"O~"��^�1���9��a�Da�"Ov����Gd�$���D�8����"O��8U��t���;ր^�+д���"O*�b��Y�d\0pi2�|��"Od�x�A�%� }�WȆ'K��	"O
aB���tm,�J�%)7M ��!"O�8�#,Y�*z�2&�,6���"O �P �h�vl����� �F"O�d[�.���e�4ԑ=�BIC"O���ˮ%��<H� R=A���0�"O֔����E���+&��5;m2��"O�A���Kso��RG�->�,qps"O�x��jA=w7�!��#.�j�b�"OBlP����d�ݺ�nR�|NH��"O0,IQ��^�<�C�	O��,�"O�UJC$@/a.�mc��ѣ{h��"O��p�ڵq�nLف�S�_��:�"O^ ��}�^�K�b![���"O`��D+�D�&t[� �)2��i1�"O�Ű�H[�^ڴ`��Ӯt0���t"O�TR��͘rI^(R]a7"OB�W�ߠ,��y�)��i�"OeT��g���h$H��a��"O� �P���.=@ ,��_D����"O�Y�2Lõ5>�y�p�O�`��UZ"OZ��`E0F7M[��X�C�$պ*O�=!��ϢAL�#cAƪd��l`�'=�s#�_�l߸��i�L�J!�'��  �O,b����]�I���'�4@��G9@tL���&��0��'yr���O��ȄBc�A�!oR���'*~<A��V� Ύ���M��!�'�!j��!���J4�P��'�]�eiQ(H������H�|�)�'"��"f9;�<��G��>x-z��'xr����\�g��g���oh�P3	�'�5)�N�#�E{Q�CV��D	�'�du3Ez.\�Q@��F�,L��'{ (V�ffi��i
<p��'t pSN�.u�:�iQ��/!21"�'2 ��]�0����$>���'9��"�˗L��8����	g�����'���H�����+�.�7N���'��}#&@�_1�%��C�4AU���'���j ��J�RY36�G4=�h�'P)�G��-R����e��J@]s�':�(��LT�th��� $u����'7污Di�[&0Rr�]�:1�m��'��Y*��7*L1���#1�,���'u`$��z����)�1����'��`��Á;F	L8y���s"J��
�'Ū����x�����.@�Y8���'�2P�
�$`�ܴ�/ֻW?��`�'� Y9C�
���*4n�K�:��'��+D�
-]Y@���"=zv|��'��{S�͸e���)큁F�!��'%� ��?���j��	5D护��'�ޜ���D+׀Xb�H9*����
�'�0\*#�
�rOf�����53.��'�����̉���+c�DaH(ph�'Ѣ �G� cɦ��É�7���'��+ G�0�ޱ2S�Չy��AY�'Y"}Df] Q���{bΒ�j@�8�'G �"�H�+�U�1�Y>y�(Ũ	�'�V�8M��Y� "&5al�8�'mTqq�]�D��pV/`��L��'���pcF�90A��\��yA�'�"y*4���mh���SM)Ðq��'sp<Ȧ��T���b&GJ#ɸ���'6f���`P3n�¡� �ѕپ=B	�'Q$9T`��͈��s�m��'�H�h��.Cv"DX� �0a����'HJ�w*Ͷu��j�J(}+<	�';B-[P���1�*K(�*([�'Z�i�H�܄���I�s���'V��:��{B�<"G�7g�*`��'t5�����͎թ�O��\Q����'i,�rD������A\��,p�'WL�1�O��9�����#[{��{�'��1���0�b)a�ٹD'�h�	�'G��`�
;\���"4h�5@E��'1�uY�G�3Ach�cn�%+��@;�'~��8���4�}����L���`
�'C�M���~�������2K����'X������(b|��!�I�Js�'�V9링3)<���4�ȿ3�R��'���p/?`5*��Í��+@��+��� �080��2#���x��?:N-0b"O��
���&{��(���˩"����"O�����Ƅm��"%W�pc"O�]�qI)V9@Ļ��U�����"OT��`aB�sI��@D �%��(�"O� G�6� ȁQc��YЀ�a�"O�����2~�<��GѩE���J�"OF5�421
��1	�Z��؛�"O �B�%�JA�r͙6v���R"OB�R�ʤ9�0@b������}3�"OTyr�#@�����e�B��"O�,�4F�-��Cu.�8{�p}Y�"Odp%�R=��m޿}W��"O�̂.�9S�:0:%Z�Z@���2"Ol�E��,*�P�k�&��"O��r���3��|AG��Ao��#�"Om�n��������(dJ	�a"Oܰ�dJ_!>�S�JR�:�"On5+a�&qEiI$��# �����"Oh��q�ٵ,'*��� .Q�č��"O���@�,R�P1'@��}�0��"O~�h�,B��0(�ŅP�	��9"O~\`�	�3.APJ20����"O�����>Е�fķM���+�"O�iy�N}�H�5⃶c�&5˲"O|!��f�fi�%� $դi 0"O���pe��o�rI�u�U=wL�"O�ct#�r�XX�BX�+�R�)"Ov��Q`��'7>$a��A8Y��Q�"O.�N�C��d�qoXl�V��"O
59�bNJ�`e�G@�_�t���"OV��L�,1��A��4��L�"O�$	K�\s�cD��-w谙�"O�	�m��-D�i` �tmN9�"OT�	�F̱v�XtB��; AW"O��֌A#O�ʅ+�(�+`x�"O"����p��|��!Qb�}�"OV�(���XXD�.�V �"OB!��o=���(U�{�8�`"O���-�6˂�SwMW�[�J(��"Ot��r�Y�u�6�ر@z��G"O�ī���T��2��17f�@h�"O0`#�S�3���ڧ�W�[R~izr"Oxs��Z�<U����]��sw"On���(�%M�IP���wR�"O̙�¬ѽT:� "ʎ�!��{�"OXıU/� ��p�r���{
p`e"O�����Q�S�rpr��#��"O^�!QGU�6c(�#"�����:r"O��zaE\�Є�`���8ό!�"OvD��<e��5
"�d��	V"O2��'�*k��y��Gۺy�|�1"O�����s�prRF�
c���:!*OҁɁO�k�(̪wm"L�\��'�6�3�NɻR�0(�c�KY6�j�'��l���0@�x��;��z�'�
	���C��I��:�(
�'n�A���NI��Lƥkb��	�'ؠ��B�8���F!.�`�A	�';t�Ҧ�P�
�Iy�JҹV<�,b	�'����S��6�p��c_�I=�1Q	�'0�Y�U	1 �񗥊T�<a��'��H���4��})w��P	�y��'c���[��\Lᶋ�t~����� $�i%��)l(�{Fb�&��A�"O\��C&�2����L�A�Ł�"OTp�bO�y��]��I�/kU�Q"O`���^A!�4�ՠ2��E�"O���E&�9h�@�g�g�P �"Oܐ(AC�Wh:�RU�Q;?\,A�"O���!iF�q�~����'Q��˖"OFqpF�7dH
}���::/$�"O� ���25�̓6툉8���"O�  �j��m��ۃF���	�"O��R��7'�ɋ#K��W�0y�4"O$������O��\g�:*\�;�"O��CH�#r�1���8b����"O�Xx��I U��`�j�VK�<�$"O�H�נ	xc�iPi�
*D<]�D�d���<�2��*�hu�2�Ԟp������[�<)��:x�|zm#0I��(3�]���x�K�	hgDM�r�L�,!Roޘ�y��ǂ)>"���Ϛ+m��)��R��y2�S|,�-��ca4xt	v�y@� R���T(��O!DA��C�y���$?:��!&\E���ٖ	\>�yrE�11���N�D`�y F	"�y�BQ�S��9�.A::=�Id�ߣ�yr#ӏt�L�yP�I�8� t���)�PxR�iC(j4�j<S&g�3���r�'�8�;�lB
m����u*H!h\Q���HO��#j�		�N4�w���z)ܡ�s"O�hS!,��U)Y���!?kJ�A�"O�5Y�ċ�.d������4�( "O`��%qT�ɒ�p|b�	�"O�=��S�"1�%!���t�4h�&"O��iŒ2���Ս˭/a$H�t"O� �w���`�P���}�Ԍ3"O�E�GM�!�P�9�@æt���g"O�b B;y���bg��xj�-YT"O$�3B$tbրX�b�2�"Oڔ�ԈD7z�t����BO ��r"O|<�ŗ�,(l�q�iζI
�s"Ov���ץ0�hd���@�0^�W"Ol-�$�Á,t�#����>�S"OJʑbVt/� j��ݫG�b��"O���@��
K�Y�2��@��y�"OB��#�ʛ0�"H槂l����"O�-:`GQ�s|��˳��j%,iK�"O޼A"K��ha�S�C�F�"O��P�bԿC������z@�#G"O���Õ���!�գ;?.��"O����܏x�Lٙ�ǉ�SXx11"O���v�̜jdI�QS�=�.���"O$1��
:_T � S�;�"O4���׏}�$���kY�D�&"O,�ᄎ�p�F�h��5R����"OE��-$2��0��`� $��"O<��C�\�Z41rLSP�>Q�`"O2���ȵc���P3��5����V"O���'I���Z��\~���"O��6ǀ�Ls�����al��`"O�Xc7
V�j]�L#pB�3\�1Y2"OD��dgJ�I�Ľ�UJ�0/�p�V"O깰+^&<똅B�+�:�)��']�Xʓ���u����g6*�	H
�'\D)��O �o�� �m�S��
�'�A���d�6�z#hF�Lu���� �U�!�Y�O[t���ڕiq�8
"O$�Q F �fw�9H�Ɩ^j@@�U"O�� �@z�FmR1��lV6p�"O��a_�s�2���N�%T0I��"O\�S&A�2��r�>)��"O���aާ=�Ƭ���/|P1�"Od0��/ :EAH\: IZc��B"O�)�$�7F�г��B2B"O
���k�8*��e�Ӫ2���"OV �*�"�
%:���t"O����Û]��Ze%?�z4:$"O���P��e�PT�E�K�o���R�"O���mL�Lp	�R�h)+�"Oy 7�R=4��PÒ��*����"O��؄Q�I�jDcM�t�X� p"OTQ'P@&E���@2HnyF"O�y�Y�sr�jLV�FUh�c"O��i��X2\��=�� ^����y2�_�3�8H+��"~vR����ɣ�y2#�kRHR���,``�%2 %I'�ybN�S��c�,תW�d�Q��P!�y�*%#�`����P��q�K̥�yhR�m8v�;F F�I������y�f[�pI����C�:�FS!C[��y" I�}4z�Q&��,�B1O\�y�(Z�N�������)$j��yrꌽH�5�P�
zV5aD�?�y�'
�y�bQ#��H9tB��B����y���<�*��U�*�0�#�V�y"�W�L�A(�#��$k}����y2�P-LГ2�G�P+���b���yb��-�N�1w�_�B������y��S�:�4��e�#5 �0AT@���y�[ڜ䒠Á�0x�����u�͘�|$Hn�}��9O������"��R�L##���-��R���b�D�0
4bш��w�
Y����'eJ2S�ݣW��6"�pd9W���MS�L��k�&=SC�����ɇ�^��H���Ƣ���*�P���c��&5��F�i�BQh��?��i�R�sӒ��"����h�$��1XC�9H��O���9|OX7X)�����i�����ae��dZQ�P�ߴ�?�M>��'�M�] ^9��A�
�6��A��O�ɀig<X�۴�<Y�[%4F�WXbo>�e�Ջ~Eb����Û@��}! �	uC�iY�O5�DxBk��B�fX�M@�L+��&eھh 7M˚5^<��j���~���Ȁ��{̓ ���	ھw��[U`�B����'��s��?�$�x��'V�X��9���p�Dpz*��gA�Y��K���G{��ɍ�:���'!T����i��^���S�4LZ�f�|�O%��[�Ȫ�˽>>�D���T˓9`D�XP��Y]�>�����\86�ׇi��3E
 Y�%�RiG�_��h�3��)%'fh �b��������9f��ARE"K�7Ȁ�/��G��3m\�Y�4D�����-K��&鉜	m"�D�4DTte{����*�z5��V�3y�GŐ��1��my�'��O���pӔ���,�6��6B��jNt�KbLYϟ���	xب�`w��]�x-i�Mڊ>��I�M�v�i�I^��X �4�?�����!��P4h]�q����DM����ȟ��	����VB��F0.Y)�Q�D����-ѓs#�)���9H�N� [���`H��L�a��Ph��F�C�R��u�0Y�1 ��KT�{�#�V�(K�@��HO�w�'r�~Ӹ���~���&���Va�>$��Y��+\zp���O��2b� ff�8FZ� I�����A���OzN6n:#�<w��S���<7R����VP?��D�\כF�'m�i>���T��"0a�aE��Od�� 7m�n[p,*A$ڦ�1O��3�r�1��F�M���}���ߝ�6b�O5�|8�9V,�� &f��D�/�.��!�#e�f~�@���I3�j��~��)�=+��J*i?��e��)�p�mZ�f"��O`H��Z��i��ɆC\�/���Q4�İ~6�!����O���+�$>�u`M;&]�SB<��S��?"���Gy��gӀ8n�]���u���K�`��|^f�S���=�~b�'QLT"CA
�_���'�'���]�xoZ�o6���&Aҧ>�J�����<mf�M؅E�&_>&�k��Z�"��Ū�Y���?�S�? ̸I)!r�bT���O�D����  �<ZFn�&n�� y��	o��S+b^��r�B�D/Pp��vAX��vt��	�f�T���j���I�M���~�'h�_��{���<b�d�5y�PF"\���O^"=�g��/��RViT�.Ɔ�������Emڱ�M��ƛ��'_���'��'�5E_�` |  �   8   Ĵ���	��Z�tI�*�� 3��H��R�
O�ظ2�>���& �H�O�QS�� y��]1��S�x%�D+QlW���K�4;B�^�?�vR���'�V7O�`����4y��Y�t�B.3	*���ņ�S�B���4A�qO����D���M�`��DO�꧇�=rF8��ʋ^y�?l��pS��(��$֊wo(Q�&č5o��I�	*��e�Sg|� 4l����	��'�'Y����O�牚!̀��t萧��ʓ%ӎ9��J]�f.v�h�џl���O	��07��hy�E�{)"�ҵ)u~2�ݠ0�T ��ݺ��
��rE���NHb2`SQ�j� H��(��|�(���5A��<�`ԑ��Q��y�.Zu�'�ֹDx�U�Y��''7�̀�f�W�+ђ"<�q�%�!2P�o������?�����ݶlD�x�O��Ӊ��ْ��'e^����$M��(B�Ӝ`D Rݴ��#<�Ҁ'�MP��h�)@=H�h��U�}�iɥk�\�;Z�"<yc�4?��.Pᢁ���_=�x��aSoy�JT�'.>��?9�KL%�����>������)L�:#<ɂ�(�|Y�����+����∕g �����?�1O��r��$���w�|0����]�v量[E�'ƐMEx���M�'A)²
�A��m��/�sUÏ��W]�'|�i�;c���ˆƳ}�{�JJ#.�qOp������I�8���F	x��Hf�ݿB��JJ#<yP�6�V ��l� &I�4	5$�Rq�ȓ	Ĵ   @�?��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �   Z   Ĵ���	��Z�JvI�*�� 3��H��R�
O�ظ2�>���& �ث�4�?y�f6TU��*�S}�!æ�Y`���k�d�DDٟ��+O��M#�'�u��J�3����
\��D%�!^-�r�o���'SrDx�o��y(ED�Y�,�;�+�u0Du�f�<�ݔ@�"�Q7����u���NH _��ɥx����e,�&}L��D��)������қ]@�a���'��ݮi����ql[%wL��'a�q�
�5�Aq�#Pad�cBCқ6g�<q5dK')�}�F)(?i�A�#wQ
���-p����'18dM�%�6����o.�'��Fx��I�Is����͟=4�!h���.�I7L#���v�	<-��S&q�j!�`�	��:� ���L��O���Oi�aN�$��dj�ՠx	��b�>1��"�Xf��x�?:T2K4��}�!IGm����𤏛�O��V"$�h�CQ V��D���I��O��ي��7��d�&8v��[�G�.�N��DG�_��	!!��� ���	�lː�#g@��\�x��P��Uxf�2���Ь�O�b������N��^�*��
P�t�<хC0�/��OJcf��;6}9��@^`���O ����$��(O�K�m�_Ʊ��(�%�1�"���	tj4�"�"�S��)��=���4��>e�b0���4}zJA�Z����Lt�ēO��8�g��_Ӊ'�48@�V9H}a��(�P���O4@�O<a��ԕ{K>�'\���j\����-_�J�ȓ.�b�   @�?��|��:��'���D �L��I�#L@#z]��� ,��	e2]�5\�unZX�W���'� II��%l��+���~�HTk��'���"6z�KH=`I��Hvn%.@e*�ၣ��S+(��0�&�3C��,QgV�(,�F�̕8w���q�����5_Hx&�rN�Oyx�e�O����1i	�(j,��O�=YS�'Ob��D��=>���B�-�J�*h��\Bt�'���'�l=��H 7hܐlBfC�.s��Í�D�\�O�h���*f��L{E%�Mv�1�$�i�X�(٠{>I���<��Vy��5hqJ����� ��LR$�)}���aY3|12Q����5bL5���	�, ���'�P��� ��u{uf<b�6��rmE&)�(��-f$L�WH�	��O$�
���T?�,Ӎ,P   v
  �  k  �  �(  	1  L7  �=  �C  -J  oP  �V  ]  Sc  �i  �o  v  \|  ̂   `� u�	����Zv)C�'ll\�0"Ez+⟈mZ�@�	�1��D�{ H��P�N����G#�r�֕Yʁ�8#(��B%���h��偟��ٮ�;�P�i�'E-(�0�'��Ii�
bA�ŀA�JbĄ9&`��{d�rƆ��a�H��5��q���ӳ�=Ī��&�$C?=;��$��Q��/��:�$��7�,�I�*q��U�|�<p�4�0�z���?Q���?��aj�-0�#ДUr ��Ƨ�dL-z��?g�i�)�TU�<��$�Rl��ԟl��#B�p��B��N��py���@�$��I���Iן��'�RL���M�a7O��d����L��E��!�d���	�
"=A���`�rY4���K��B �O�q;�,S�D}b?O����{B
�>>�%��&��h���#�\�o� u���O�$�O����O
���O��Ŀ|Z�w0؈�O�^�����N������[X���i�nmZ�M#��?	C�i�2�~�
�Ă�H��fl 
EH=J�ϗ�a�>�=�4 2�=�4�'Di�U�L�!,j�i!gJ�0���=Ŷx��4%A�ƃy� �Iк���S��h���U�E#H)�El��f 3s5����E��\�c��<��k�N��V@Yj78�N6M\զjش1�(��b��S�-� �960B��.,�Nx��g��*��g�@�m�w"<(paII,}��Ǻk��`�)��y�т�H�8.��)���[$A*���*K/8�v6�R��U��4�6�[�'T�p�u��%�"l	� �;��Y3`�5d��(q'��&# ����<�(��ǖ%������7������>�8��fm�ݶpB5	S1E�"��b��
~�v�lڎ�M������'t�구��O�^-��eR�y�n�|�F�9��L ��I���D�O0�$�O�BѬR�5����ST@�޴ �jh�`�ÛW�\�C�FP6r�P���ɓ��0Im.�k3�W#C�����%�5���7Ak!𯜏S�F|0G2O�� �'�������ĜJf(hh،oJH��OF���O�㟢|��dL*oc�Ԛ�b-+M�X�0�AY��hr�V�~QH��Ϩmd����DڃB�p��II�kS� E��2�Z5JELոZs�� v����H��r"O �Se���%' 3�&�s��F�y�Q&�伪ЬP�3I�AB��<�y�hʅ�|�	�[�*t�m@�{W!�d�)@�M�CN8�eb����:w!��Q�UT&dJ[�F����(/�%+��U��XFx���ʉO�*A����?%|!9#e b\C�I�OZ0��*B�`�5�����FdHC�5K��1D$�#�2%�o�(VhC�Ɇь�y4�Ӡb���R�Ą"�B��6���G�k{`��!�.Ld�C�ɒHqthi��ϭoh6[ I�-UӢ˓AH@\��I���� �g¦nA�%�^�FlFB�<lj��#�B[
�, ���?OXB�	�PZ�쪑�07��$!V�u0vB�	��*d��m�4JW܍04��1Y�:B�c���3V# c?�=c���j+.��ĝY�-oZk~R��٢�І��j�,�a̟�?9(O��D�O��䂢\�d���*<o��i�@Ә�M{#�H�<����
P0S���Z3�Fq��8�n�F�l%�DB� X5P9��B9�ڹde��t�����\):���� +s"�'���'���aU�:���Awʃ3���gS�t��o�S�O"&!*s�S���B.���@�	�b���k<2ػ���,)80ڠ�Ŀ�?!-O��d�Ϧ-&?a�S�?��5����I��
5y��˦Ww���Iן��s̜�1,XlV`��$�`��3���D��BJ�	8��`#[�F�:s4���h�HK-*�&ɻ�n�eY�	re+�')�0����5�b̂�OfE���'7`� ��?�O~���T��N!xj��
b@�����?�
ӓ�\��PaB\ +�HJ��~�E�,ڧ
��8h'��Oĸ:�(�{Z8��ش�?�-O�i95�����O��d�<ype�!�@�q K�"5�"=�vؕ?�h�Ă3�67�=w���*���DN��89ª�~B�)c�,�~f�S�gӂQ)ħWmpeh��+�3�ɣ<�Zy�3&���Zsb�Y��8nZ���DSA���'K��'�<H�qm�4Q�g�D+76�t��"O^LX���� �@�O�_��ɓ�^�����4���D�<��$V�q�7ղm�Z��@ľ()B	�k78��������֟�Zw��'��I�>X0���j�(	xV�{­�3�20�O���,�%_�`�q�h�j�x�D:;6!�Ď$_���S6�]�F���ʊ�!Jx���'f!�D#rx���=k��Uo� )F!���5Tx*@RLA20� Q�&���r��'-�6m:�$�	We��m���x��
`"�	+�a��j��t@1D�$tD�����aOğ��	�3��@�'��� ��j�Z�o�l�@R"U�'�\�;��'���f�����8�l�t�b��GZzd��� ��P!V�ʚ�0<��#�P�	��M���D�*�����m�><���ٶjS`8/O��$(�)��OvQkU�ɕa����eŸ_�:,���'X7��T��`@�-`�L ����>�ʑmZ[y��ŭN�r7�O���|b�eѪ�?9׃]6rA��Т.���Av�ߎ�?!��%���������>qƧ�&�  ���@k�`�R��l~2���D�ʉc�[S�Ӯ��D/X��#�Y	/L�^�,��������4�?���I�Ղ��х>ԩ��۝3u�'��'vў��v���PL26�6����W�ʢ?�1�iڔ7-3�S4"��Յ�o��' ]�nfT�'��Ɂ���SX�'n͠�K�!�����!�p�>����U�$I�Y����!���UQ�&�YD-E�|��\��o\*T��0N�����ѥD��c>c�����O�; $���W�0��M#���O
�D�OtqJ�Olc>��?)\�c�8T�ei��R�(�de@�yrH=Y���9��P�"�
�CvNM���|�'U�ny���r��T��"aBh��*�9Y�R�)tha����O���<�|�g�=t6��C����!�ވc�nLMK�(���Ӷ�*�91,��"�4��$A�Th���v�Te��eA��ڲ�,����%}h��T��N�bɆ�	(J�ҠA���(r�K
�	񤨀���O���Oz�tG�$��9~cp�	#��-�n�#wM.�yr%\�
�D3���+{��PH�3���I`y���:o 6m<�o�N����N��5�8����[쟬�'�B�'�󩏉[O�4K�H0}t�B�R�U{P���cۼ�0D�Z:i�4���'���FC:�0Tp ��jɦ��r� ��wdJ��@m�@8�܆ቄy�*�$�O1oZ���ܤX
�XK�A�=kT���my��'��O�8�I�PRH|��`�$�f}T���:��D��J៲P[Z�I3�(3����NM-�M�*O�ٕ+����	ry2Z>��I2aGT�+�GG�tR�x��g�����I�@ѥ�;4_`�RLC�S)��A@GT�Oڼq ��6C	b�xq+܃<����O�Ò$Z00F ��oV/i��U��c\L�	 eN�nI�8���{���Qܒ������
�4�?�K~Z�OKd9H�A�?��%au��Q��D2K>���hOv�1��DЇ��$l΀DJ��΁a2|�E��}�do�d�'r6�}���S�_�9�gP\
��	�S����?�g�'-�)��aXWY�\�M��zx�
�'�̡���B�3�<
�F�$��	�'qڽ�a�ܤ;u��q/ϹN2�@	�'���{4 ���zT��?�ФZ�'y���0�[/�]3��E�4 |�
�'4q�mȥDAH�б膯#���)O�����'�qɂcO�4�渘�e׊h�j��	�';x��n�&L��i!��[-$�8	�'$��R��x����/$+lpb�'q"�K�ףc͠Y+�f����a�'!4�y�E/�pA����h���{V���r��{&��fD����=/��`�ȓCw�#Ŧ�'������j����ȓ{�6ջ�ؑ6���l�87m&M�� R���<n,P|0�N2)��=��.�:��%�\Dp��ҔR��I�ȓ�(���X��u�V �''΍D{������ja� IL�/3l-r�28���`�"O��Z2��&&���<m؄��"O�)��V��`$/k���"O���'�7*�)���H(Q/�D�E"OؐI��ȇ}�x�	6k��joj�k�*O<�EJ��4su%�}����>�Z�Gx��i�i��Ղ��;C���B�J &��B�I!T��la��>w����,I�F�B�	ALh�4 K�+<z�SO�#W�B䉒0�r�x��_��t�u�D�G�~B�&k�Z�
6	B�%X��d�~B�I�[B����������7���%u�����f	��9d�
{��E����O�C�)� ��I�ڶ|�����φh�t��"O����7cf��"ǹ]K�"Ot�r5��:���b�+024�"O�h�'G�+zҬ0KP���W���Ñ�'[Ra8�'�
�Q�mԲ>�d�ݯH �Q�'�>q+�ݺx������>_�4 	�'��䭙12Z�xc&L>4M�H��'�`Q�!��3��S�-�\5��'DH�����\��@���ğN�t!�'��p0��Q�U�:q�F�}?�|Ѝ��HK�Q?%)P��I��$���e=�`w��<�y"�3p��D�l�~�MI��&�y���<�TlS���P\۳A�3�y�=\Y���/F7Iڔ�cs)���ybjE-}h(��ͯ9#f��!���yb�2�ԸI�C5�^�z�*,�?�V�Rd����T��׉ϴm�ܺ���N����F6D��7��I�@�0dGƼ9l���3D��I�$V�p� �-Y�H��N2D��3�,�/J� ��+�g�(p�"�/D����h�L��$��bʣ..�}�B�1D��yv��P�����e��rk�IibG�<с�i8� ք���Y镊ڄ}ne���.D�x�ǫ� ��I)�H�+ @R6�'D�dP7@�4E�<
G��y�:�$D�Ƀf <2rh�1cF8�h L$D���r+�&AFX�J�{�>�A�a-�O��a�O����%	��tE�,�3}.�9�"O��NȬ|�6x1ŭ��Vs�e��"Odu�u$�5e2E{b��8E�Z%	�"O��"��C�1D�m �V�,�j%��"O�IJǊՔ3��-��j=1�ܩ�"Ob���N	-�B��	A�|��t� ��g��~
���d�Ը�j�p���ec�C�<��_�d��80@@�G��[EgW�<�����?R�p�)p�+6�y�<񧠐S��50g� +!U�#��x�<q E��` +`�R��Hq�<��e4z���VC�<���"!ğ�X0�3�S�O�ɘ�D�9Bu��2���5��0�"O��3�e�0`�&���K7<����"O�]��"��HM�`b�ˈ?k�(��"Obl��Mh��e�K'h�8��"O�����V�ai��j#*ݓt �t��"O*�����9�Ji{�H�ʀP�V�H�R6�O.h��ц.A ��+%�� �"O�@�w-+h9#��)E��"OК�cR.�t����6��E�p"O��p@EY�F�@��0G]A�*ѣ�"O\����xJ42�-�����'8r�'������Lź��R�I�ohj���'�&Q�7K�5w<dRs��)Z�<��'��b�)6o���'eȁ�'��0�@�h�&8%���V��ʓL��y����eH	�b�R�ĵ�ȓvvu*£�*A�t8�'�ޗ7�>MF{�]"����yr�
F�.Cx(s3G¯z��"O���	�mJ>eH���G"e �"O��F�(W�\X���jIRY�3"O�  ��̳>n�H�����b"O��@RF�`$����B�x�8'"O�����1��G�qx�Y7�'s������R�Wi�%&^y�BF�<�d��<8
�+sA��Oe*]�f��dr���S�? �,��⑃"�ț�k�~R�pg"O��ǋ_�d�Y�S뙃6FB9Q "O�P�͑m���92K��I0*= "O�,�&פ��%˗b6�L�Q�h���+�OFL�2�rx�$�s*K�&ayS"O>��gFB�$��jٝ".���"O�<r��̔)�����	K�< f�C1"Oмb�8s�L�V	X&�!1"O�̒��1�����.Tx5�'�Щ��'�tIg�[��H�b��%�� +�'C�8�H4�ޘ��
�w^�0��'��u �iƭ�>@E�Q
?y}��'u&���IY5a���{��S�e+\��' �eE�"v�)Q�%�9N �\�'AFY��S�T�
�CDn�G����ĕ/.�Q?FL8S�R���dT<A���*D��3W�_�S|l�Aq(�0*8�!�3D��J���c�
��g�G���u�1D���&��W� x`1fp��p�:D��y$EW��� ����T�d@8D��C��Ad�b*���YߠЩ#c�O�I�1�)�'�2%�`MNun��!KM�Z܉��'��t�F��25��8w%�*R�:�'"��BjÞ��B5A*V���'�<Y)�E��{ފr�jK5-���y�'��	Gj�S�d����(8-"�H	�'-@�s���b|�$K2�4�L��(Ot�e�'&,�Aٱ��<[�A�!���q�'��]�7˔?��8#������	�'@��XwU��8��Eǡn#Dl�	�'�����dR�)�K�׏a�Dh*	�'.�5����44%�:w�,/��	�P�	�� �)��ǎF��+N0EΥ�ȓ/��آ2cED؜���7WJ�X��`{>=��Ê�r>�:�)�6sv�ąȓ<	�<�f�W�p"a
@��6R����/$��b�(m4����Z3�x�ȓE2�2d��O��4�ň�b��D{�M�.�ȍ����6D�l��H��L�1�#"O
T�S�Z�0����35c�x:U"O0 �QN�y}�{��Ά1>�[r"O8��d�0|�ּ�6�րeŢ�X�"O騁.o�ؽ2�ѮX8�j�"O^Ԡ��"_�Q9&aH�qP���0�' @�Y����7	[�0��C��Df��S�`Z(:pU�ȓ���h�� �h���{�m��<ir�zB�K��sr��q�N��ȓϘ�
�MW+̨l�w��6Y��ЅȓY��doL2?L�xa@Ƀ�{s��ȓK�,�7@Ȥ�	���' Sȼ�'l�50	� _��j��&�Ԡm��ȓ`ئ�q"m�O��1F�m�x�ȓhAFڄ��%�*@�R��
yW�ąȓ4���j��Ƶ0�\8I��%:rL��+ޢli� ��.�Yq6��-9�<m��	�F>���_�����9 �<�4���"OB��bcһ���9&��~����&"O��;���$Ԉ"D����"O~|iԨ�!`ʙ��X�t� �;D"O��(���!]\L�Ə)��x�"OP��6�;w��t�4��b�I�k�L�~:��M( �
�2"+�7�^[w�Ky�<��ӕ/�:�E̯Ys&U�`�l�<���_�@q�Go�~I��0F�Q�<� �(�J̛H"Ƚ�vEKD�ΤrW"O�C�Q�B�����#�h�.U�1"O���g͈o���c�,W6%�0=�')r�
���5R�F`H ��*�^�`c��.ڵ�ȓ5@�Bh�G�&�`"�]en0�ȓK�䱂�B=*��Pf�*�`�ȓ��M�׈ÕquΝY����0}&��ȓ.�D}rw�N�T�0���,T2d$�ȓIx����$_�$hz�˩i��'l�4h�n�6�!B�^-f`F��ԨY'4� ��E
,���!~�IHDě��x�ȓ�"���c�S�UAA*ɥ�⬅ȓ)��Ě�Ǭ�J�(�+�c�ਅ�P|�bB�A<��X�f'B7⭄���`���f�:���QF8�`.)�hB�ɱ[>`ևY�iT2��t�[�l�4B�	��:L	Wl�;?����9K<C�	�\�pP�mȮ@d�u��51�@B��kVDE�!g�o��%�È?M%>B�>���B:�4 ���F�=�R`X{�OM<T�bĪV�����I�c��	��'^�!d+���}xBk̚dL�L	�'��J����=�
��rAVZ��`�'OF��@�4[���!.��}�H�'�R�ȧ�[1Z�Q{�D�L�X��
�'f�l�J(|�)з��'>O\;��V*|Ex��	&h㬝jCfY�Y7tI��[1D(B�	�V�T��S�_l��Õ�9|�DB�	�,8� ��kD�C�呲H�4�nB䉸����y\�I�%+̣,qC�� j�h�H���/a��`zG�K�, �B�I�$���;��Q)}�"��F�>��UE~�,ؖJ�H��?��Oh9�%��~��) �@�-�v,���8�ia���?��#M���P(�A�Vɀ�*��O~��x�MR�ae����m�f�\;��ą(d���j ��x=�6ʳ|�6k�%A%���ŀN���I�'�`m����?����N�-��@�$��$+�|&)ް��d%�O��[v��-����#�,N���C0�'Cd˓u��E�E%��+0Vp��H6{�z��'p��a��'���',�2�� �	؟ġ�П[��M���!;M���5ڟ�9w���Mn(���6h����4���a̧I: ���9zچ�Q���� �̓"C04�Dk6ٚ�ؓ+M!I��cݥ��Lg�S�B ,�z%*�WX<�bȒ"@��I+V���D�O��S��P~�@��|�D�³hD�@&$��y��ǈ'��e�[� ��B�,�L�����y�ON(�iV�� AXZ�g��DS�l��'�R�'�$�U�^;* ��'8��'U��'�������m@�-��F��+�P!3��2\��6mF52��bv�3t�R�'��'�
�`'�(U�b���m�*QL��0/A�(CL�;|����E\(��ɕ��Mk�f���$G6�����Id	����Bt�ɣ-�����O��=1�'�VL��(�9¦e�`[ �N�
�'dK�a�6t�qʐM�?~hM3�k⑞�۟�'�V���H������̙<��$#��M�EN���'���'�2�O�B�'��里���匈j^܁��꘴�t���Nu1�ӎG̺ ݴE�џ�#w�\��0��:I��B7%_�@b�b�*F����[����d��Ŧ!S�D�h��T��ɳZU����4n��,r��|���	r�'��p@U�88�I�%��
1�Q6�"D�D��GP�rؒg�O���	����<ᗴi�_�t ��F?����O�S;(��u����|��I˭\B�,�I���A����\��_3�iHZD|<�G�y3ry�i>����tpH@�J&�Ĭ�â6�zt� ���[=)����&��ͩqf։+d��?a�ЪG��#|��!5��O��d*�/h�T���&|ps�B��U�˓�?�	�U:zHh�;a���R� +ȅ�ɿ�򄒍e@���I�"	fui�n
���I�k�j<�	V���	V��
��F����'N�g�^,2B�@�:骉C�'�H`���:����������6�Pd�T�	 �$#��Ǐ�*>�r��c-�@���K�����[���@7�A|�\w��P�֐���e���Ç)[܆x��y�.�?!�����4��� @4��_"K�\�0����#��$��"O���z50�S�V�l}x�%�I�ȟ���)^�yL��I�_�H��в�D�/g��|�3�kYƉ;���;]Ivث�fħʈq�ȓ
!x��D��M֔�2��*37�|��]��(Ф\,Z�}Rf�mEĆ�_=�$��J̩F�Uu��(9���ȓ'4@�"�
@Y�b���'F�rd��I�"t�0��X*-�s%k�,0���!�		������������Xw�r�'��	N,.��t2g��k�bDr�&Ǭ1���K5蜥ZצP���
=n���V�c�~��(�:-dJ�����2l�Q%�.�n(��`�pR���Э.���RQ
Z��PN0�~k�䒌v���'��Oܢ}r��ݪ=��|��IY?zH�X�Qi���yL�5c�IAuK_�m�rU ̊�����֦i�	Wyr�F�6Q�ꧧ?��Ot��#�7�n钶��I�j�Y�RR,����?���]$&Tj���.�;��Nޛ�,���PA�M
,��`�?K��%��I
(^ Qc@Ę����oV�d��Y�⅌	��� �H�&`��V���V'��Tq�O��I��'R�I�9]���I�ӊ_���t��4'��`���kT���5�4 ��Ǔ�}u��3$$�O@e�'��@!'�U4L\��dH�'0��(O4�D�O��d!�SX~�$�	#�m�%��^��j�BQ��0<Ɉ���}���+�n	���3F�Ew�O�(�R�x��IT�Q6�M+F�� ��"��ݼt��%�~2��<���|�8��q�A ݙ6fFh�����/�������D_c��Ёt��̉O[	��R�}}<(�#%��L���Q��
z?���9O�l�Iߖ%9�����F�0�ׂ��=n�P��|]��O� �O9�1Q��M{�8�A�
9���G���O�+���"u����T G�%5�@�q�T�	r�ɸI��'��'���(L���ڴAߞ����T�h�nG�[<2`�'dDY�O�$:��Iѵa�%9R��*1P��q�Ma���DTE�O�s�� �N'?Sɏ�\�~��B��C�&�����	S���-O
!����O���W=���0擊}3��j�LɜZJ� �!��Q�8�$
*�~�����?�ɣX�(�	�V4̀�AX ��d��N��������?	��P"W�^	� ��	S�ɑV��X�<Q � �&���t�ʂT��:'$�Ѧ=��W�	������M�7/S�k58hZq��w�PK}r�'�Id����ج�@�:N�`O�������Z�'�ўb?��o؈9��a�*��)`R��eE!D����B.N������/�1%	!D�@���-�`E�k��sh��!=D��9�k�x�r1��`�8o�-�w�;D�t���N�X"��\�x%�l[@�7D�������i�� Z��5>�H9�`o6D��S"�?|�~��$ɰ=jD'G D��QЭ��y|x��7���h�[�a=D�2�� ���Rs���	A!D�tR J�!!��)r� A�`, B2I$D��P�]� �7 ��f��)8D�\	Q�[ �5A']�qA���T�5�I1p�b��b(C�%�X�rN@�I�D��E�&�T2��t�b��vC� {�LY�f��u��a��E�b+<Y�N��Z�P��d�@��D��E�G�k"�?Z+i��B%GH�h�GH�)y�T7,�6,%t���ŏr�9�ƌ�G��BA�2w)���ގ0�O��R�T!��A���1�d]�"O0����I2eW2��R��O���"�"O&�!EbA9M���� \�E+fUD�<)eG��/�ݠB�R�H�2%p���|�<i M����J�@����/ZC�<���=�t��	�|�L�hg��|�<Y"+Ң�p(	�/6<� f x�<	�O�q�x����]��@d�H�<��R+`]��$^�mH�&�k�<As@�'wÂ4$۽l8H���j�<	�͖H�0;�K?@(����d�j�<4��Z�e�DDQ�:*�q�j�<!�HWF�����9#��|��ba�<� ��딫	�K�VE�mۮ~��8�"O��*�g>V�|�R� Avt�ۖ"O�-��.V�����C�no\%��"OBU��	!c�֌��c�_v݁�"O �0vc�>W�እ�M�D0q�g"O�аuBW�z�h@���\7xL�""O8�z���WZ���Ђ(�S�"O̔��j�n�j1�d�3n`�0Q4"O�D�;9[ =�ŏ%]V����"Oj�!AƊ����.)!���"O\�k���	Q
�%�"1
��p@"O��8���� ���#M�
���)�"O�z�͸=|씱P�>|�z!�"O��@EG�-5�r�#�����1S�"O��3�.ӌ��*�h�f��g"O�����#,� hQ�(��x��"Ob�����[��$v��@����$"OV|�6脵KR��R�)_)|��I"O����mt9}�G�����|@"O�-���@0^!s���0�"O"}�K�~}�`jw�мW�x�1"O��b�.�bDz�'
y��t"O�l-0�4�H��B�q�fP�w*O���m@:a��� �g��A��
�'�~�C��S���f�Y�v��	�'��|[�i�U��1+�i��w�2��'8�ᑍ��	��ܐT�r;bY��'�����΀O��:4&��S�LP�	�'�L|���[6��u���	 R��'�t��I�1����Bb�7x!�eY�'���yQ�I�n�{U���8��'��U�a�6hZ.T7)G��2�''���q���,]�V�4s�'�|A��L��_�(��F�H��tx�'�Thr�n�V/��SU�K�F�.��')�����R
�r��37�v-S�'����c��";r8�3I�+2��
�'͘h���t�<9B�BG,Uqh�'���!sG�7%��`���W�TQ�'I�4�D��:j��Ⱥ&c������'hŘ�F�)H�a�B��y�01�'@�d2����=�Hl�Fę�rL�@�
�'�H�e
���eD�`���	�'a���I�17��i���f_�Q�	�'��X�ŎA�L����U ~|��'*�R�0��ͰŁ�U��щ
�'E
��pk��|��=#� _Lx���'����ш׵�L��l=Z��'�.���EC�
M����}��I�'��0y1H$�%&ڢI.�];�'�:����V�� p�W�@R,��'L2͹BJ�,�L���. D`|b�'����0�J5d�L� ��4@����'6����I>i8�GBX8:b�$��'U(}�a'T'vt��K��ߵ.s�Ey�'�A�`f�Eg�T��'ƗY���'�Q3��SR@֐���Yݨ�`�'戂�I��jO�8zD� PM�a��'z*dB6f�W^��0愯@���r�'�Z��$n�/K�vm�W㊢6�H�x�'n�� u�$r���"�%�)��A�'���b��\����O�IV�Q�'���(�>!.�r��RI�ޤ�	�'FRd���@�~�xY*U��9����� Ba��	�w"hS�)+�V]+�"OTcR/� 8M$�&�V�"���'_�죡˻������@ՆY@�'�,0�r�0�\�d��)C�9�
�'3����0V��9;`J��
�'T8b�)�A:��G���H�
�'[XX���Q�H�0͚Vn] ��,0	�'՜q�1���N�kAfz�1�'=l�ª�$)�I��Javݛ�'��i�ri��9��G�>�m��'��5rCg��_�8����0
�i��'�2eӄD�>c~�P�,��A��'�	���S��V䕱'�B��'�b�36�^��*�c\�M�5��'�����6�>�`���� 3�'��R ��2��S�I	^\���	�'6]â�Y�x�ShX��P"O��	��5
����r���-U`8�"OtQ+���CR��BA�iT��`�"O�� RD��7���ơ�*Eh��Ӂ"O$��B�Eg���F ɌjYx)!�"O����#H�D#��#�^�3"Od@�r/Ƴm�l@A��ٴ��"OҤ
�/�� A���-��eC"O�	0��Ҧ/8
T�әU� �9�"O~(Q����Q��
�������"O�E#����	<x�� B���"O4�0f^�:�tu��#�=-f(��6"O���l�%@��x���d�]��"OA�ʲB�.���
JԀ�"O��
���)N�%7���"Oԉ$��[�@���b܆'{H���"O��1凷f`a�!�<\r�`"�"OX��(ѸH�Lq�OM�v�,�"O~}�����~d����@��r�B�"O`hc$�����P!��~�� "O��YwM�,��jV��p��p�"O�hSR�ֶqC�̩t�I�H(a0"O|����E��]J��_w�hpQ!"O"�j��/7>�꣥V��Xi9p"O�p�C�Xލ1d
�&,�J�"O�%�1�:� 0��CP�EAp�s"O�t�,D����0(d�"O8�Rqc�� �<ʵA��;<�qu"O�\��8g����.ū8�~�1�"O~y3d5�Y��A��5Q@"O������S~)EMU�d�Йz�"O�xJP�Ȃ
��M�V�R�P���"Od�*�NA(� <2�;5����"O�|@wA��mY�jQ�Pe��8"O\�%L��Vm��NX�5�7"O�T;V�&NZ���/�80�q"OR5�TkG,_�x�S4@='���"OH��gŝ7(��H�n�u����p"O��x9��p�nM�h���"O�(�Ūۼ#��8cbN!8�@�"OZ�b��ހFy����C�
�~h�"Oh�e��zZe�_�@K��d"O\,�eK�87�Ұ����G?ɱ�"O�M{wLDX�8�j�<�̩�"O�5���	}eI�����Iâ"O� �%�P ���ѕh�p߮�&"OЄ(��cmt�s퐅L��P��"Obi!��n��i`�� {��Ū�"O� �J!���r����We �$q��"O�1"����pA;��ͰH���%"Oz(�0CU ~�d3���zp��P5"O ��Q��W�t�B%Ԅ-tB A"O ���e�D0eϕ�.^b�R"O~Հq��'4��ie�G�D$�"A"O �.�(:O��4�ܸT-���"O�uOA�Z_T�F�Z:b��	�q"O�ٺp�I�#}PEp�T�:�|aq&"O���1��)$���fC�(f���"ON=��m�0�H��u-�3S�"d"O��9�LD�a�ĉ����8.KvE�V"O��� c�7�`  u�1YM>�1"O��+�\l�X2Cʎ8L�Q"O:b3�B4�.��d�"D/L	4"O��ҕOK��D��SA���"OP)�������P��\S�"O|�I �Go���:s �0#��Y'"O�8ŏ^!\m�$	�J�{�"On�bpF	�R�6���\�>�|�Y�"OT�Qף��0;$�p&�/W�ZA1"O�e%��xPӇ�
%[�̀F"OHEq��2�����S�{�`@`"O]��.@�0�2!f�уq�F�y�"O��d �$[2�$�B雽V�$��"O��k��Z�V*���*T��Ir"OX�"�IN��	2g�'�`�
7"O�����3��0�'��H�p7"Oi��蒱`�B`J��֙K����"O�����
)��E�jyՐ�"O�aҤ�NlX�IL<m�x3�"O diB
ǻh����n��H�zH�"O�=A��%2 �Bv�Q=�(P�"O �2uhWҔy',F���a0f"O���3`�&q�őD
͉E���"O��I=?F��I �Cj���W"O��ѢP15nT%QR�
lJT"O����L�H���� Y�$�|���"Ox�z��,�x��D�\�MP�h�q"Oi� �Gdz�t'I�eE��J�"O��E*�����a޵w,��Q`"O��Af��&N!d�xv ��K,�ᑦ"O,�)����^LTR����s�"O �A@�N$I�D�`�$�� �zQ{"O�|ч����D8�Q�R"O̕v&��7C��z�!�~X�@�"OJe�I�z�k [�\WpXAw"Ol��!�b�za�u��=��i�"O�`���qp�5��`[�.=9�"O�)���%��͊P˷>����"O4�;Ň�@� �q��JlL�%"O�y(s�T7r������U�
�p�"Op�6l��Xh"�$��d_"m�p"O�囧O�.L]fX Gc�L:�`$"O��!%h�n[$�  !�()P6"O\h㓩B����i�D�*@�*e"O� �aJ-	1�6��q6Z�����(;m����C�I9���9T�'�Dt��.Z�x09��7u��*
�'���&$*NF��P��\�4S6���'��!3�H40*zQ��B-A����'2�2l�����üPԤ�a�'Ȯ�)�N]\6�;?d,��'*��[D�\&F&-U��X`�{�'�Yӆ,�98�t�t���4zxi�
��� 2�R�ض\���5�O
Fw,�R"O���MJ��K�-	�q@��"O"�K�n_!s��hf��'FX��c�"O)� �Kh�h�0L�A�x%(e"O���9$ז�X���3G"Ov���׏a��p�!l���w"Ox�+�@�t�䭑$O�i��H"O�ƮٱT=h�Q��d���r"O.E��GeiI6�H��<���'[�ȢT�!T�s��2oR�Ő�'`"��t�T7-�c#L^�%2]�'S���2�$�BTȲ, �Z�4�q�'�N�1��9�,�GV�Q���'rhC���13X�m��.M����'����#cn�BR.C�CN����'�r��ْ�N-�
ؾu�j�'� 	M�b�^��Gd���
�'��NV�i���.ߧj����
�'NvX�D̈́6&/�u�d��L\:�'#��*���L��I�蟞& �	�'�F���D�6$���C�2�n�R�'}nYБ��wG��
��0�DAQ�'�$�K��>�� C"D$���;�'� `�����nD���ՋF�XT��a�'Ŕ��5��8fx�!
E-M�|��aQ�'5����!�gQ&����_�'骔��'є9�� ��Z}��X���kf��1�'0�Ze�8ZH؂w���l���'q(y!����I����(�T���'�Τ*w�
a�����/��
����',8y� �==�ș7oZ�.�b=��'��š �X#a�(�2' í+:����' F$(E�S�u
��$�Ĺ0 8�!	�'��!���Q#2Ȍ\s�'Y:���2�'�d��4V?f�zР�$��$<z�'����£U�j�+bm܆c����	�'��(�eˋq�=�%-�Z��'��sի��f`��aEAǅ�Z�H�'�``j��V�C\���T��P�8<��'Vtk��:k�$�$@�I*lp2�'.JX�Ԏ���Z���޸�'N�-ڒm��pA�g�O"x��'�\M &��
A8P2�mλؐ5�'��[�� �����u�Xi�'Oj�����+t֌!'�\<�%��'+��u��%T(�m��.!J��u��'
�8cѯ|����$+��h��'�U�0G->nL�Pҥ�Ȱh
�'0*U9e<zQLS��Ѳm�)
�'���3�ޗF06� ���
�( ��'���GD�+~���`Ra��'�N��&��&8��c�-@�E�$�'����%C�k�]�*1�Re��'�b9j��}�*E g�"�@c�'���	F;���%�Ʀ!m�x��'�b�ps��K������m��'~|L@�D�8\��u9���,�ʨa�'İm��( T��=�g��)9�(P�
�'��p{Q!�
m�h��g
C1��
�'��1��#Q"��<"7c˲0����'@�y!�W:8��!��3��Q�' bɢ�ۘ[t��a��B�цy"�'-�$*Q�d��AR�B]���{
�'*@�CĦU:0�h�h�N��F24���� �9X�H�0yR4cDB�/X�j٘�"O*x(P��"��ȫ�@2Bm~��!"O��跋Y.]]�t� '�}�,��"OR��H�)WZ����Tw�� "O�=���#z'���g#�#b<jF"O��S��RUXpc�Ȁ+o`dS"O��`�Iq{a�����+��Y�"O�ٵ��"VL`�Wȅ�]>H��f"O�кG��6l�`�C�o��4:���1"O��Bs,Y�eUN��ׄC�Q3|�$"O�q qn@�"u"xSW$˄}fQ�v"O��h��6?r	SB�;��+�"O��
�� g�2\���M�E��J"O�A�w�Uv.X��7��/��\��"O
�(��N�v5�#�؈#�8ԓR"O1��%6nHB��I��`�9@"O��SF)�>�Tq�5r0ܡR6"O��5���Z��X2
*G}�D�Q"OZ\��"D�x)� �)S *��"OpxP�Ө}�Hd�S��/mȁi�"O�HiA�ڈ�� ���]Sd]3'"O��K�# ��� �`Y�'�N(p�"O�@�g�G�@ʃ	M� ��"Op�@$˟=O��ap��r�"0��"O��	�9k�(I!�
�@�0*R"O*�Tl�4��e�U��Z1���"O��z G��O�X�RAM_ �0C�"O �X�E��J2��B'��xh�M��"O9c�o_	8��m�!ٌ;-�%��"OT��a	Y�O���+���(�Y�B"O��*�ڮ�
�A�.
,��"O��S��*j�4@cԑx����"O�@�r����#�A߃9��q#�"Ot��A�58����ռ!��:#"O>��@-o���V!��w��З"OX�{w
A�ne��Z��C�2���)3"O@d!v��(X�ZQ;�W�ۮ q"Ot��3�K\3����)e��H;e"Ox�S+�!L�dI4��*k��4K�"Ob�h5F�K(��h�N��ce4�"O����X���*B-PY虐�"O��&UGp�J׌\n�̳A"O����>s)X�IwӔ0;H�:�"O�i�`+Q$y)�!���vC
Qp�"Olq��!��٨�mD 5�F�v"Ot�§���y?�0���ʁ]��	×"O�r�F�j?�$X�6��$ �"OP�ᣏV� Ԣ� ʖ�p�\�zT"O��qb'^�(�J����'w�5k�"O�!H��/-����)�.k}4r�"O�i��k��=��M�E.�zq�4�v"O�PQ�/�#)�rxÓ+�)W,9I�"O|XS`��>#�1�,Y���XJu"O*TA0-�7N*�bl�2/����t"O�P�,����5 �C� /�.� c"Or$*���8��h �m9
�'���  �)~�5jh��q�t�'~!�kD��0���\#U9�	�'��\�$Â�J I�P�L	B���'FV�a�'V�xh�V�I�I�.�	�'bҝ;O4E��#T|`���4��I���A��Aз��Bm$��;,���(�:��=H���4H8�ȓo��B�3Q��R�j�p�����S�? ��a���=K ����g����"O|)�`���LJ��,yL�e��"O���=�� D�S�CN@�U"O��A��2��D��P�J��|��"O�Ȉ�g�u�x�ۆʔ-N�ġ�d"O|��˝ y������K�_�����"O80�.P�d���
���p"Ofq�䟶A�6	sb��~ ���"O`�q��_����0CI޽Qf�)J�"OP���l�#��5I0.��PP^��"O�]ٓO�6��a���@�v,c�"OVP4�^-�&LC0�E ƼL�"O�q�G4LP���*�6>l<��"O� �Ҏ�).�.��jJ��Bt��"Ob�1�fZ�k��c䗞����d"O������?9��0�1��-y	ĩ��"O`0�mЖ$
���ώ)��A��"O�11�`1T�j���oޞDa�Y�u"O�]
ãűT��!S�NT�erH�ڷ"O���H	%��4QQ���`Y�Y�"Oz�di
�0Ӡa����}�Z-�s"O�8�r�C;z6U���ř�����"O@Ȅ@� q�x��E�V�`)��"OB8S��Pj��Dڰw�8�u"O6�y�풅+���RTi�n@�"O���5�ٚ.{2��Zh@8"k�-�!�d�A�4s��b��;�$�ai!�L
Z\,鱨BQ3��J��QX!��vi-PV��/�X��m��!�$Wc:nٛ��N������A�!�
�k2� j5�֢��cs'	�!�d�&2��jvn��;�@�5�!�$C�v�N����J_M����]�e%!��^�P43��^Cbs`�
h!�F]�Tl;[x��ӗA�0B���J����d���S�ԏ`�B�8s��ЊV��CN������d�B䉄2�R�H�JR�h�o����C��6Z3� !#�5k�<�)�B�z��C�	�|���� �/yt)���*�C�	.'�ȵ�1˂;'�b�DK!F5~B�	�>ۨi0I�#��]��H�m�2B�ɵz�މJ���!�n����t��C��\x�#�cبZ\n$#���s��C䉮Pm����X�,�@@`��7'�`B�	�Y�d�(ViM�!l��Q�	a�C�I�f���X���hL�@�V#ϴB�	�W���ѵ[D|��JU�H�NB�ɝB�|�"1��
h� �X=��B䉟����&cދe[� ��	��B�#-�ʩid��� ��ρ�>�~B䉧_�f=��T�e���c��A�G,B䉺 �&pZ�
�bvdK1	@0�B�I�i��`�6�5�JD8��̊,1FC�I�h��h���|\�$�Ǧ4C����+���MH�<S&D 3�T�y�-��IՄ֕1X�i��)�y�N,o�j��6�H�8w6��fOד�y�lɜ]��
f��,�p!z�H��yb%�y�^9�EK��R���1�(��yRcM�FN���!%%<>���C���'���D��:+�5s��O	9���K>��	�x��D*�,n�x����r�<�GHJ4��	&��i	��s�!�o�<�΋�����D���V�<� �Ъ���E�â�)� ��"O^xxP�[-�Nh[�,?@��X@"O���H>�(�CT�B�Xq.�"O�E!2DZ�p'5Buj��"[���T"O��z�N��%l���g��HNp�"O�*�aH�	p.(�E��g0�$8"O( ��b�.w��s�G�&��"O2����0[]8%��H&.��8ze"O�U{2�{���fgI.FJV"O@�#e�ٺ"��ۗϜ6H�p"O��1���-��b��5o)��b"O��؂����,c6��+輚U"O`��@�תS�(TS ��i:Nh��"O"|�6'��|�!�r��x(�a�"O",bc��:���C`��$$�R"OF��f��56
 �ŊY�.�0}A�"Od0�+?f�da0$��u�X7"O���"Y�)	����۫\�E@�"OV�x'N#Ut����S�z
����"O�8��� �,���	aQ$A��"O�,C��L�37L�ѭ!���"O
Tq�)'+W���`���� 2�"Ob�ѵ�s�И
�k�s���"O21��"�O>X�"�H�8Jh��k�"O�Dy�MZ�:����u�U'KfVHq6"O,���Ȅ@��#6�T�|Z\M��"O��(WC�_Z�ФIM0�bI8�"O���u�B�4h$j�*#u�8��"O���]4dhy��]���U�"OҬ V��2�����$�p3"O��� �k�hu!����N���"OHq�'�ݞ`ɎԊ��33wl;A"Oբ�Ɉ:?�&����V�"1ip"O*9X$��5��&�%Ji|�SP"O�(-�TL�L�UEHc��3"O�����%������:�&U��"O�ܡ��L�QDh��\�"�k�"O�,86h',ި@��ݜJ����"OJq���݈n�D�+s`��x0� !�"O6(8�`��@�0���D<|�6@��"Oht�P��]a�©Oq�ĨQ"O@��JX��тuß�4Vh-��"O��������&�=%`n�F"OnI���>QZų�ʉN���P�"O()���h�DAj'�ʈ�"O��qKB�Q��(���H
��� "O�y2�A=oOzt�2b�39����`"OĘ�&�F46�l��C�Yˠ��1"O�	��O�.�id`X't�^�PR"O�<�Ǎ*��j5-
�q��pC�"O� Q'���jT��7�H�(�"O����r[#l��O�4�	�"O,eB2�U�v3|t9&A�]ɖ)"V"Of�+!D�_� ����h���"O����6k�¤cT'�y℩!�"ORu:'�$R�`h�e�7����"O��n�2�U��dYl����F"OPZ��ς%9԰#ƛ�%�����"O0h せ-�A励?�R�d"O��5�V4U��mY��E+4	�]��"O�ɰ�k��6$`���"F��eC�"OL`*��DdgM� c�hi�ݘ"Oԕ�&�L>"֪T�rg�0Zl��q"O�,��'�Yjv]��.Pm� ��"O� Ԁ:�D̀0w�$Cp�� ҄�"O��aՉ�1a�����6E &=p"O�t�6�)�dWm��︍�@"O&Dr������U���h�x1��"OBx)aM�a�b���a�;�\�7"O�X9@�}�t���@ـ#^�8A"Oj�P��,/ߨ�� @]R׆�
�"O�ԊA-�=g|�"��Ԫd��@�"O!Q&!š0.��-R4M��z�"O�ɪCE�2r%jd����2R����"O��k!� 	�uFmQ7�����"O�%��N�;I{^�k��Ĳ,�R�"O<xbEfI�Y��q+ @�$8@�"O�<��+ܺ%�p�D��^0��"O�p�G�H��:�Ӳ*�i؂�"O�$��Ėz�P�y�o��X�`h�$"Ot� %lP';2D�V�_� ��"O����^*t۔��LX ��X�S"Oh ��j�F��J�d�9v��\�`"O8�ʀ	�<R����F��XU.�i "O����a91K<ԑ �gH��"OX3Ŏ�<(��`�6�4d��"O����LX9���a�iY�o�b��"Ou;G�J.�4����D\�R"O�\��IT�/�P�qGы>�4� "Ob�Ul�?n�V��EX�g��CU"OR��eH�U}:�;v���~v�{�"O���kU�[�N�� �ϣc��@{�"O�3%" R�v�I��Ц1���j�"OLP«K�:�.<��(X����"O��R���^�0h��b�K��}C�"O�0�!��_x� ��9,ค�T"O@-�PJ�"D!�(a7�d���a"O.$�!�=T���E��.SN� F"Oj�9q
��F�`�9Cȏ�A��"O<��@ʑ6MҲ�IE��5�*-3�"Or��򩃾2T��H�*�K�D���"OZ�j� ������ 
p�dXU"O�j�C��?*���2T�8A2�"O�Z�`�>H���ҕ];$M��"O�4�T�N+W`[5��k1�e�0"O`��cA��N�đ�Pj΢O��"O��[ǬW7;���:)T�"��V"Op {W�X>H���͍�耛@"O��3���(|�'NŉX���"O�4(��1�i��?Wj�(A�"O��FCe���7%D�\�h���"Ox� PB�2Izh�#οd�\ɪ�"O pJ�㜖}�RaJCEȞk]����"O���eb���F�9G��'H0�S�"O%�bI�@À�@�.�:4mX�"O&�څj�Z��o��[�֩��"O�|�`�<(X`
eL�zWN�Cs"O�����8�r�r��L� �a"Ot�(�½.VV��%�F�@7��6"O��[�f�9/Z*P���C!`)���B"O�����LBpc`W�F�����D7|O����	��j��A��)rK���P"O،cCCʂy�q�׮ĦD��5"O�=��	3�x�u�"&�Y��"O\H
1lM���e[� P�G�n���"O���gD��Yq#O�=n�~\�V"O~;安�F��P�3�N�Tl��g"Op��E�Z9����.��T{���"O� ��WMP�a8C�ǅ�`dbp#Q"Oษb(K 7"n8XU������"O��p&&� [�)q.�7l�����"O����0yG�q��U
k�M��"O�u 3ϊ84�.t����B20�ە"OD��ό�>�D���U-?��"O*�Rt��_k��X�/J5L6�S"O�٢���G�\e�R/�9 �\��"O�p��Η��[uN�J��=#�"O�ݓC �-9*�L��,�o�<3R"O���M8X0lz���R�n4�u"O.!@�ΝJʹ�S�P7�`�x "Ox��%	�^��t��#\����u"OL��3�ؗ�ɳs�� c����"O�2�A�(0�j�;NF�A���c"O��#%�+f�5;���[���)"Ov�c��
�k���T����b"O��ЪA8T����Y�7���*O�1��_$�>�ؓe�hC ��	�'� ��d�V�Oz`�ڢ��q~rQ(�'�<I���<LL�(��
\9d�h���'1hI� � B������sЖ`��'�R�i�Hܴ�q*5'W.",��'E
�� �	 ΍X$�$����'oP�q�cK=�Z��A\�8R�j�'���"k� Av�X#S�E�g����'B����#Y��X�Ց�@
�' �h��(e�-�kR���@A�'E�� 5EB -����`(r�ޔr
�'�~�"�L��S�mP��gzn��	�'��8����ir��0���Zj����'T��T�	9132�JG���$2�e��'�aq`�@*�ʵ!׆W&!`0h�
�'`�X�G�� C߂-A'��%<=Y
�'�f��!%��W��� PDP�P6ra��'K�)�� 4�-�4`�;6k4�
�' �1�O�#�&�K$�]*�M�
�'.��s�İN�j���YB��q�'yJ�#l�n��R�!m 
�'�I��o՟	���9�W���	�'>^��uBT6��L�eg�"v1	�'���U�E;<�ʀ	J��C�b�'�&����K�v���eN(~_Dx�'�@�[ �b6��)H+zH2�'(uH���=0�;S�Qp�Vtb	�'���!B�]�* �5��P�Ȩ!�'�8���n�j����Z>08	�'��hi���:���BB�S�{�M�
�'����-�$s��8��M7}2�P��'a��ʖ�%Wvր"Rgޢu�����'�rY��@�MX�Y�ES%o�lQ��'d`���S�^�01�c�-b4����'	��R@��4z�BŇ d�� �'7�I�C&ȱo2�����T�Ej
�'gt����)%n�Be�KFuJX��'�h���)�Q�Ul�;��T;	�'ꖁ�5c�0Q�>i�lɒ3]��'��@���^Ǣ�"ԀЁ-v�A�
�'k*���B5�-a�)ʙo��TK	�'6��NR�9�P�� ��7~���x�'�ԙ��Cnr}2Т��F��L(�'gĉ���J�X۔��-�?�غ�'qrx�G`�j��#.�0�0ݘ�'�X�4kػϖ��o""��� 8�21��
c�a#���<>ʹh�"O~9�#��O1仑�����d��"O2dÑ��9.q�JA wN�]"O�M���P!ZX�NW;�d�"Ofл��P�!�d\��*��QZ=I�"Oh�����0a0aU*ͦv�4e��"OVs��1jF]K�����>� "O���@��-yǎ2P(A7cլ�B2"O�8i��S�w �0
D�I�C�n���"Oh�:�`Q$��y"h�
nT\��"O<)�,S����"{b>�"O�y��A�3T+��J�-ףabBuٰ"O���PV�5~]C��l]�D��"O2!��`K��`��4\�KI��
"O���,Ζ����J[tE*�RF"OH�E��/�`Șt�˨t<��"O"H;CD�ޘM�ԃ�l�tA�u"O0�3�i�S��8C�L��9u"O)8�
���2Ph���ZQr�"O���3� R:l� �	�$"O��cѩ9x"}0�/�`�P$�"Ol:`�M��d�
�P'~�u3�"O�����Fv4��@�՘�
�"OP��ǭ� s��m��>�ҁ"O�QAJߨ.�xi+�
�?e�as%"O�`Y;S��h	�����"O���ңˏh�����H��>D �pC"OB�j"l��.}��ǜ�:����"Oމ2G�"$�iB�L�xA��"O���'��F�l�@ w��!4"O��q4		�WH܉FW~f���""O:EBD�?�0��dk��x�x��p"OB��Ri�MU�P�ϗ�B�C"O,�IM	�ah��1��y�L��"Ol��鋿P��)Ҷ1f���q"OB��ȍ�a�М���uLehF"O\����0(�(	@ n�2��"O��aj�|���ƈ]���$"OLc4��py��``H�5],8'"O�4�ɾ%��!�
n�!1u"O\�A�̱!�B`��c] :�	�a"O�Y3��^�K$��h�+?�`� �"O���
��PCR皕h���2�"O�u�A��a
� :�4����(�ybb�9U����j�M!t$���y"*�%�*�`�]�50��$K���yb�_*Z��$�r���?~Xp�S��"�y���-��8($�H�#���sb��y2͋.yM�Y��""j�)�a^�y��ș �@�A
���[�GJ�yB葟�,8vmT� r ���@��yR ]�B
�����Se�TÖA��y2#ڪ[�0�Q��I����J��y҄�`��f[�=���WkV��y��0��Ipw-E."4�'ʄ%�Py��Ǭ\����@ ��w���+�BX�<A��#���Ȑ�6�&�C�̓l�<	����B8JY�+P!9�4A�v��l�<9G!J
W��Wѩt�������#�!�>U�J2�n�J���vF�:T�!�ā�,'�xYR��d��We�;z!��	q#�ja)D&A+����� v!�d'�!��@�91�t���P�3`!�^�L�\��T�?��X��K	p3!�� �`B�8o	�}�Pɠk�ZM�S"Oj��L�;o8Le��b(�]i3"OR�i�-->D�hU�*l!($�"OZq�S��]g�X�'�x�N��"OyI$�S_� Hq|�i�4"Or�W�,OO0���hՕ~D��q"O����")*�l�šWvŢ�"O��ǃJlc,m�6��9j�x`W"O�J�i��1(�	i% ̣DzB��a"O�A�쀴%ǬHЅӨYi(��"OP�z��%6.Υ�eݯb`%)�"OpE۵+�?|̮1���B\Ty�"OTAR������k�2u"O�Ţ�n�fy&�Q�R�Py�}�T"O��$Oٌ6)p�!�b�9B݉�"O��	^ ����b�h1St"O�s�e�kw�G��Ή#S"O��BH1#�RY9�eƬT����%"O|��mS�rz��膎,b���"O�9$-޾r��!2'�ǆ �^Ib""O�u �BX�0"����Z7,���+�"O��z�e.%��y�tF�-%��02�"O$�Bb�n�&m p ��j�Ʊ��"O������m��a���?��xS"Ot1h�,Ň��Г�`�+y�x T"O(-���A�<� �+N�I "O\H��E�����]�l϶-#r"O��3g��o	�P�U�V�o��`��"O<D�3�0 \	��|�1"OY%aE�mޠk7�׹H	�9�"O��I��p�bR
Q�V ^i�"O���[�sr�M#D��9{��K�"O�I vk�s|v �FK�P���HT"O�ɣ���:�
!!�J�)�E��"O!j�\�3�ejƊ��f:���"O���t��E�V5 ����"O�\�  Z�apNM���S) n��"OJ��4@
�2i���'tMn8i�"O�yx�薭慉�=��l"�ę6]!�F6x�������R��;^L!��Y�z�TB���*L���""#�,�!�d�^��U��fP
`tF=���
�!�$�f��83�]?V|���F�	�!��s���d��%z��� �d�p[!�$ތX�x8:�#A�'�:$'D�B�!�d��d��-�^T\Rՠ��L~!��
w��zC��#{4,��O!�$փ8v�-�B�ܳa�� L��!�$M�FzE#toV�AIXQ(� xE�C䉖E��*�C@�Z�v�B�f�*��C�I:lEE
u�9A�"�Y'haV$C��v��Nֶs���0��1x�B䉪X�v�P%bL�$>�K��"*�B��,,U.I˃$G)H���ЧM�p�C�	�?NŪ��ϒ����.�,9�B�	9f�q�uD�*l�~�ybF�{��B�ɛU��K���V�F�j5�ڽʘB��$$�y)��b��$)Bτ>g�BC�	�0P
��������Fk��4��B�m��i"�߻��x��o�"O:��BF���4â#B��y�2"O4	��GߧM��)1eBM�h�x
�"O"�x�M��g^2ѯ�`ܤYD"O���a�T;s�Ȼ� \33!��(�"O� $��P$�h�>YC�@M�P96u�7"O|`� _�
�c�@I�F)|��"O��P�&�6jfQ9��"c%"�"O�5��P1.\>�P�-_�{�|���"OT�d�L�Or�|�Rj�!b�N��"O���r��8K�f�{v�q���1s"Oh��r�Hu��J�J336Z���'y��+�� �o���Ć��R���'Z��񳣎�\a��4�X%�J���'^��8�`�y#l)���3f�b�"�'�y���M�t�䩭�mh���&6D���GFi�>�0�� �f�`�#5D��R�m"N���	�`	'#���� D�dr��Q\>�+v��w`�0YǇ=D�$c #
�X&ȩ�%l�i�D ��<D�l
SJ�v\��f��*��h��;D��
��NiS�*uF�u��Ř�8D���A>*�v��ƃ�"O�\=���8D�Th�MP6PEu����z�8!��9D����lz%0�p��~ l`��S��y�ʊz���왏C�*	�ᒖ�yb/˖TB��8�(W�3�j��.[��y�D��B�X��� /�HY�TH�y�ʃ9�Zu�r�]	2�RY�rOU/�yr�� !�t�H���'"�����#Q�y����`\��v�G�؈b�U��yRiČ��؊ ��,�����H5�y)@6RL���=t��S��y"J52�l��횳p�h�9�ɗ-�y��\=b��U�ҠIm�J袲(���yb�+A��@�j���XRAM�y2�����@*V�c4 Ya'ƫ�yr�F!{@�9$�Y�Mj��Є���y�mA>W+��c�
ƀ?7de��c���yB��3RHB�]50���s 
��y2O�E��Kao�.T(�P�B>�yR��t ����3&P@P�R�y�%&R� ����O>��-�>�y ��6$+��	l������!�yrI��$���	�P��ЁW��y�4��}�㋛�6\�
���y��=fa��!��Ŝ/�L��vkG��y�Czƞ��',A����[6�N�y��2}�E�Ǳ�01�Q��y��,DT�$�p�	��k���y��T8)A&��I��Z����yr�B(Z�$����(*7,Y��y"R�j�ZD�&��\�$�@`V��y���qub$3�H޽F|2�z��\1�y�瑋�\@C�=9u��{5�͇�y���68(��⣬H08�u�O��yҬ�&hF�y1Bԝx��ՑS�Z/�y2Q5x�|��B�&�2I�@X��y­�;r�\�r.���%*���yr��<�<1�n�{
ձ����y�kP%����e56?�,`T���y2C�X,9�b��+:YD@��y��U&v�R� j��+��uid����y�k�!7���kf�0}�q���/�y+:7N��C�S�~�!Bڅ�y�%S�a�P0N\�O�X���Ă��yb&�6���wd�5F�:i��y�G�0|,:eڔJN?#ML������y�7+�Q�jR� ��y���y
� 2���D��s��  b��x�^�3"O� rՀ�c|�y[���%{-d��"O��(��`��f��q;x x�"O��� ٝ'�y҆��$�����"O���ㄓ~N6������0��R"�Iן��2�%��F��ǖA�x��|߾�/$ƵxF���OXpJ��Ɠ0ʢ(�qd�$U)0�t�(���d�����K�N�fz� �����HO�mA1��J4
!�!-=�uzeP�|�pi\W���G��`�dj��A�'�D8���?w�i��Y?Qpt�O<i�RU BZ(�:����?Q����'� H�ǬI�]H��@��40����{��	��M��M+��ǔ8en}�UGū6GB�AP��L?��&�8"�	Byʟ�O�=K��!vL�"L�^FQ�7O��e���9`?��̀��<L�<�2w���g�V0M\�P�#I"�>��@��Md���8���"�W66��&K7W��>ט���@�/Ф���GzQP6��#w:�#z��9m����D��4*�옡`�ƔH�{աR�Q]���?�
�	 z0�q
ءX�6�"�/W�������.'���'�Ӯ 9��L?YU�(�B&�9$�ʀQ& �9��,�'��d�SFx�,��F}�&�j�텟RZBp.����CHJ��Q�`�H`>|���TIh��S/?��ۢĻ?d��HJ�?iR�'F�-�����4n�z��R��>C��',�����])8�G��:M�=)��ّ�?Q��C�?������gy�';��:2��k�&��v4R�Qa-�+
L����-�s��5X���I�<��rJA2U��3����D:����Ī<)� ��@�YQ�IU��t��C��}�.���<�����z�!�؜sk	�&aN����M�PG��ɁT-�|B���[6"?�0ʃ$Ϧ�pUeT"[���R!�P��A!Wm�28���A��tzUrF�ɹk��n���Se�9�.���Q��ԩi"M����?a�����i]�;���q��`E��#ǰ�ֽ�ēy�<��A�k-�t[5���(6����w���i��˓4v�HQ�@'>9�5�,�#,��j4�2����0:w/E4+���6��T�����9f��Ē{ڬA�Ug	�ZtA�M}��|� ��$T��A��J^|♳���<
U��O�7s��  ��!^S&pZ���HOd���'K��p�$���~zp��!d>"`�_d��@��Ɯ����O^]��IףVʪ���B��?	����')�6-�O�6M��S��-�Ǜ�����o>^���[�N���lZϟ$����'��B��rW�]�a�^�)u$�
�.�A�W�EU^U3���g2^���n�5`q�:�9�¹	e匛s��$�5	�ٴ�f	HZ�B���GЭUT�!
��s��k�̔���ѥE��ՙ0�`Ӹ����'T�6��ǦU�IW��Mˀ��7:db ���T<�f��Mf?a����>�S�$��<��ᎃ _��a�_?�L>y״i�4c?9�O@�<�FiӔ@�H�b%�:�͉�$�d'lORm`�  �   Z   Ĵ���	��Z�JvI�*�� 3��H��R�
O�ظ2�>���& �ث�4�?y�f6TU��*�S}�!æ�Y`���k�d�DDٟ��+O��M#�'�u��J�3����
\��D%�!^-�r�o���'SrDx�o��y(ED�Y�,�;�+�u0Du�f�<�ݔ@�"�Q7����u���NH _��ɥx����e,�&}L��D��)������қ]@�a���'��ݮi����ql[%wL��'a�q�
�5�Aq�#Pad�cBCқ6g�<q5dK')�}�F)(?i�A�#wQ
���-p����'18dM�%�6����o.�'��Fx��I�Is����͟=4�!h���.�I7L#���v�	<-��S&q�j!�`�	��:� ���L��O���Oi�aN�$��dj�ՠx	��b�>1��"�Xf��x�?:T2K4��}�!IGm����𤏛�O��V"$�h�CQ V��D���I��O��ي��7��d�&8v��[�G�.�N��DG�_��	!!��� ���	�lː�#g@��\�x��P��Uxf�2���Ь�O�b������N��^�*��
P�t�<хC0�/��OJcf��;6}9��@^`���O ����$��(O�K�m�_Ʊ��(�%�1�"���	tj4�"�"�S��)��=���4��>e�b0���4}zJA�Z����Lt�ēO��8�g��_Ӊ'�48@�V9H}a��(�P���O4@�O<a��ԕ{K>�'\���j\����-_�J�ȓ.�b�   @�?*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕP   x
  �  k  �  �(  	1  L7  �=  �C  %J  }Q  X  p^  �d  �j  7q  {w  �}  ��   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dlӂ(p2O�=�!�'�AbE j�80�eˆ["����.�4&N���ρE��J�l��d	�V���u��H�y��_�S �DB��a�,y3fV#2ԐGL��>�P��FT0Ji<��̉�]��E-�H�.��~�&����@뵢Q%4� }
���q�@h�`a�_�e�����?���[�t鈀�c�	p-���F�iW��'
b�'��E[?Z2��"�a�v����'�7H�S#���?�e�D�����?)��DrP�S̋�nt\x��O�?����?�����O6���i>*��J���7oH��ї/5E
i�U�	b�'O�,nڗo�D��Nʩp;l�koE!>�h܁�OF��x#qO���a�G$��,��&�B#Z�Z�������������x������Iܟ��O��Цb�v�n�p�nɈ�D=��Lv�T	l�"�Mk��i���'��6��O��n���,IR��MB���d���f��Ax�*�L�'3��F�įY�6��"�̒�m*����ώ�M	��Fc�)V=>���-� ��6ma�
�l�?��S�:yd, ��X'|P>8�rb��z�h�A�Б�z`��4/"B(q��^5ֲ�tmS�|pTK���]�����4,�fd�5�N�x���3&��� �Cدdu^+ j	x}k��h� oZ�MS�(�0ִ5�%ae�Q�]wy��]!K����%<�ZL�F	F���-�t�W<h��d�ӫ���a`ߴd
����h�x��U��J����K2uP��-��A ��$j�I��r�4�8���=4	�PمD���.8��J�O���u�I3&��`ɐ�w�) �T�ur�4� �!�M�i���O-�TŇ�oXp��ր�P���({؊hP�"'���ñ��37��\����֟P�I6Kk𤑄��$�h�JC/dٛ�n�������j�0t�
����˕�0<aU(�a� %"U�!?��j�灟W7<\BC��~��c�
�wƆ���	��O���.?	cbتCf����C4H����������͟�?E�$���S6v�,��0Y�������?9��'�Pla�dM�1�((�r�	��|x����'1�\#���y�I�7�ߠ&��P��Ɲ!#��B�
7D�D�fłd���7V����_b!�P3t�\��!. � G,\�V�!�zF��+v/�/(�ʐ
E�i�!�z����F3H����u�SI�!�dʯ[
�e��C�b@lq��a}R/���O?)(d ֝��h�B��_+�-�C]�<��nX5[�$�5�G�X�栉Q��Z�<	�l��Z�n��Re��>�ⵯMa�<���J�?LP��P+I�3��B�Z�<ɣ �z�X���=�dY�A�W�<�s�\,iX>�Z�k��L���DMUyB�
�p>���;D.��cZ�q�ֱ 6�Vy�<!���
 qd�91`�<� 4_�<i��#0�8x��Ŀ<�yh�-K\�<Pd3�P@"4KF�t�Mh*@W�<�l^q��顥ϹQ�^�ӌ�kx�`��jC��M��O���j͹+�(�vm�&��Ј��'����0��ߟ����J�� ��! �Z�X8��i�����ị�45�@T�p��@�g�����S1Ъ���D9k��u ��	�l�~݉���2��K�`�`����On���O �D�1A\d!#�e� ��Y.��ʓ�?ي���T�m�0H81)�0S%�-зEߛU ��/�O���L�Y�aL�'�t���'�	f��̈۴��'�����?q#�(m~�@�g�	d�0jB�9�?��9�<�� ��&���wa �i�6�Ӑv�@�F���8��;!E(7R��:Z�t�$��gl�S�蒙���D��N��Z���a/��]���xք�;����K��'�O�1�f��U#�B��C7F�`l8�|B�'�az�Ӌ��dx�Q�u�)
婓���O�	E������Q�Ȇu��`W���o?���'��I�|�:d�Sɟ�����'(�M���. $-Ae.P�Yk���GP8Le�ࢁ��̦5#�(s��b>c��0%�F;^��@Aͣ� ���Ȃ2>,xn��r�$�%%���|�<���Y�$􋑐b�|@ Ҍ�$��LmZ��d��fi���'c��'j���&��B�0��W�Q�W_�� �"O�]��� w���(��O�d�SZ�$؍�4� ���<!���
 ��{5f�\U���UnR@����_8�?I��?�����O�}>ɲ5��F82�4m��E��h�2b͎�B��qT�t�FU�!�:t �)�U�l��� �h:��չ;�hUy��I.�:B������$2�0{G	��W���w#��}T�Yѯ;D�䠃�!$���*ş]	�%#�+:����'��Y��M����?q���<.�!ȇD]�a���� ��8�?A��H�8�{��?��<m^�����Dx�� ��rp��:	�āYtQ"��̀%�',��&�A�s��ii�(H6S��, �&�d�CF�c�TtbW�H��0<�4+��L�	��Ms��%d��ڶm��a�	C�X=-�0/O���;�)��OT)WD�7}F���K�* i.)��'Qz7�C�T��ĺҎ�#
�=���2Q�$�o�vy�g�4r�7��O���|�
/�?�BF٥D^�����[��T��ާ�?I�F�������>!��Ȫ,~Š!e�0�\�I�Hr~rǇ+A8!A��^������>�"�i'��2H�nhhE�]�Y���e�������D��4�?Q���Υ��x�a�	6)+n 9��WF��'%��'�ў���6�<�"��;!�l�k���_�n�?	�i��7�&擆O5����Q<Z�j��A��Jy�'
剸A�4���t�'��H��CBxPd��V��D��ςm���)0�<b���K�iҨ����6�*��Gط�`��M��4��b*c>c��8`n��
��`5F���a�O����O��	Vc�Ofb>˓�?ф�`�Bh�m��7h���Ǎ��y�̙72���lK�2�<I�DjF��LL�'��{yRf�4M����3O��q�v�� 1ڤ��Ln���d�O.��<�|��CY�Q$y����l5J�e��}�P2�Ɵhθ��eɲd���dG'�n���냡x��аE��*�@��k�|���eL�a����	���N�rq���ۑF�*� P띸t����OX�"�In�O}��1U���.C6�+��(ovR5��'�dZ=ȩ��	�U��m�CG�$��*I��ry"	�,V�6/Zț�a)����E�%�B�!�ş��'���'u�	R������L�#z��ԡ>o�r21ɉ�L�;E�iJ Y��'��K�j�sp�j��ƨ��=�G���|�X�GS?6�4iQb��9�0<��R������MS���x��.��e&Ry2Ai��T��.O��%�i>��<	X���	�N�E@T�N�0.���Ŧ-�qD���dI t/:ԡ�(�M3/O\�[��N妡�	]yP>��IN�^����р$7�`�G�|���	��H���:tP�����|϶��C��D�O��h�҉ܥ?�EHDES�l��<��O*��N�.[���p�Üm2�������X@�T�	kS(͘	|��/�d���ݟ|��4�?QO~"�O�]����V�J�ȳ �$J�3J>����hO��V��ف�V.W��UAR��m�h�D��e�R�n�U�'1B`d��凚"�"�k�-�.
v��������?�g�'������P;OX�2&��.���'�~����	�`�Eꗻ%� Ik
�'@I�� �S!��8]p��0���y�Bܫ%Y�kF��Eg�Qp��8�y��I�x��X�v��Q��(�'�υ�yR�8&�Ԩy�:EɌ<�G N1���|R�̽�D?^�r5�I��{���	�'��r4EU�d?�Q�@
a�� 	�'�4�I�iBn�xSAL�$^���'��)q�"��n������4���'nJ{��P-\7\���ƅ
��}�	�uA��?���)Qb�>�`�퀿"����)`�i��ލ0��a���7V��y��X`���]�[����.�G(���a�Q"�"݃SJ���@�?뒅��Q�B��i��J�,Psk����SQtAc �H�]ѕdل|F�G{2 ������E��N�^,���FC�=GX �K�"O�!I�A]!�9�"��>p;�"O�p�v	�7�d�Є!G:J2LT`�"O���땹.�6ЃA�M.��"O���0�c�.���)�(�ฑ"Op0�bk��+�:�h��^���9��'I��B���-|'~Ӡ��3XP8
���7�\T�ȓkbdH���{�����:��a�ȓk���;��������?Gfy��g�M��m]�|�@�A=q�Ʉȓ�T��&��?̕Z��X8K�,�ȓO�����ꄑ=Ȑ�t3� h�'����3���"%�\ +���gHKm�����S�? ������X���D��4hQ"O����M�N���'�4t�P�S�"O�$��������{c��{����{�<��G��Eڞ�:�)^�:�9"��Sx�h��L���1���T	�1#.�/|g���#$=D�,�F� ;6��Cܜj����O?D���SJE�F\��j_%\��g�1D��:�ΚL]��c��	��)C��<D��bB��5�\q�G!��j!�i:D��u�E=��H����>Bm�f/$�o���D�$�,$o��b"*F�q�<PY碋	�yR�E�S|B]�5b#Ψ�V���yBo,E�H��J��[�"�q%�V�y���x�	��}��a��!���y����P��� ��t�~�Ѧ�ē�y���?VKx�q2MW
7\츁����?�BkHa����Xec.� {R����p�j@c��&D�,+w�Y)f>d)�HL
�t�C!/D� F��/0�ڼ���W3b��	�CN-D��x5%�{��{��T@�xz(6D�����ȝ�ƨ��#ޕjP�4D��JRB8�l�AG�*k�ƕ��K�<�Dn�b8�̳�oǷ��<�2�*s�ɓG�/D��A���QP�lbC�g�x��-+D�X@�O��b6���a��6��y�G�)D�0���Cp�0(A$��X����Fg(D�0��̕8,?|	��m��'"0�G�$�O�u���Of5�F$\)|i|�BV�<Sj�x�W*Olt�`�P��J��X	�yA�%>�y2��<[��j&�F�q��2�yBOѰ'ܚܺ*�����c���y�K�s���d�	��5����y2$�'��� ��@	��� �읐�hO������,z:Q�Q�2u��A�I�T�<C�I���� �L�I��mU��8']`C�?D�@���%$�Y�Վ	y�@C�	-0;�8���8=��"�X�:C�I�~
�5��҉X��T+��X��C�	�z�|�Zp-�p-�PIv�=P���$�z(�"~�Q���=�V�9�c�YzT�aQ��yR��o������1Q�4�P�m�9�yW1,(}c ƛK_��6���y2��x����a�&vsb�����y� �,���ô(X�a>(T84f��y2ˁ�;P�Ң����aҰ.����T���|���H;@�"�f)-�q�`J
5�yRm�.?$�P�b3��!7B��y"��>��4��aY*$��$�F�5�yb���:�kW��l|�zŚ�yR�J:b)�#Ӵ ���Ν<��>y!BC?�QE��TILsF	;Ff �a�v�<�M�Np[�@�c���D�l�<AEa�d*2�"5	�ln�$�ӏf�<���&(O�9ӂ,S�K��T�%J�I�<i���w����W`�R��u��TB�<I�F˫��(@��lN���!I~�',\*���ؿ2�L��ȃ?�:�b"g�O�!�䌅wD<�Tȍ�cǊXyp�D3:�!�$��`I8���%#�x�%��k����
!(B����ʇS��e)w���y���/O�x���C�|�(�Q��y�	�=�J`r��9:5�����?!�G�Y�����<��R9!�|�CV�L0\9�Iр#!D����2�$�����f�#%�=D�� �E!F��*Հ�C�n��B
 �"OP1f�y֜M��Mжe��9�"OZ頋�6X��	1�a5�f1B�"Oh,�׋��T�6X���}u�&X� �
=�O�y�u�H*�� H �?i{�4R"OB�j�^P�н�� k���,җ�y8A[���
Gs��-����y���\@!�'h����X��y"קl^�l�S�[�`���a^.��>���Q?�e#
P���ؕ��/0-zl���y�<�Gɛ/&k0�k��d��d�y�<� ��(`��=#E�$T$"�YS��t�<���N�TjQO������p�<�s�ӿe�"��E��,�F9Ä]k�<��e9,F髥�.A<}���c�'q��b��i��*hi6 ҆X�X��J]��!�Q�D�����y��IS�+ɑw�!�$��~
nAhV�/X���Ig(S!!�?�����T
8�"����-�!�D�	'%�U�� �	�8����_�!�d��s5�!2�_%x-�EE 4V�lΥ�O?��RnֻR�Π�T��0kZ��u�VR�<�3A�+n$�@ �M����3E�Q�<�s�^�&3Bm����y�
���OM�<�1�IM�t��ЋT�Zԅ\�<yB��;{�n�BcfP)BV(�CRV�<	f��
�x՘�$S
ii�W�iy��-�p>A��N�bQ#���T�8��c�a�<�ׁ3}U*�B��V����I_�<q�`�#>�\��ƶ���]�<QF�&���")�A����ACHW�<�qǟtC\�Y �K-GF�(� ��yx��;�h����&WT��1)jəvfFt9��=D�h`�%�=*�xQ�t#�)fb��<D�Ⱥ#AI��$��F�
�H�hQ�tL:D�t��j�F�5��B�Ly@q� l8D��j��)jZ��`i���j�1�N6D�
�K�� �R�a�E�X>�
�C5ړ*x�E�Tg�,��q�iG�=c�Q�-�yR��(~���e��$t,���Ć�y�΄�0z���'V�!d y�q�H�y���ΩzD�CD(�)��M��y"�ގ6��Ł"��6r6��̅��yr�6o5��pϕ�{�V���B�:�?	�l_�������1(�	K��RAi�/�D{�,2D���dY�/X�!sM�	Ͳ�@�2D���5�Œ$	��K�#_�6p�5�=D�@�Ӏ$!��Q�gI�A�����<D�4e��	IDĲ��EbE���
<D�K�c�+�ԩS@¨x)Xu�P�<�P��^8�H���	�ٱ��A�2�$�n4D�@�D������	9d���@�0D���F�F�*��T�]�#ъH��0D��z�LW��yꙔZ���B$.D�\3���lT��� �{`�	a-�O�h��OT�b����tp��A�5�~\�"O�l���T!d�mJ� ���\�"O:i)�H�=/�̑�֐_|f	�"O�(��C�/`��&C�0֤�"O,�qR�Ԍ����шG�Q�� �"O�0i�ٲ~�����I'��ۡ�I�H���~z�e^�lHJ��4+F&�������f�<�p*iEP��E�m�F�K�c�V�<�rG��fdj����Q!�v)�"	�J�<� �����B�Ђ
�%��7���:#"O���vK�L�[�td߿E���"O6��RA�5�j��%C�z�Tt U�'�̡���S�CL:�Q�2T�@h0�-��D����ȓ:�҅S�'Z�jx~HX �,�N���CR��L�i)F�
�!�Ǡ�ȓF��$Z2&�$p>͠ "Ьvp��ȓh���e�"@` L��Ɠs9�p@�AT�ɷ)*�9v�u:R�' XU;��~��.@=n-��o�?�D��{��P�� ����ɜ�.j8���Q����']> z��&j����ȓ
��3�	զ����-eslمȓP�̃���S7z}I��¯q��l��	�Iբ@�Ł�	-�,���׈<6VB䉵>�4 ����|u���T�ԁ �TB�ɚ���sE��9P��ǨvB�g8�b�C6eN�lB �zC�I.k�,i$��j�t0���_� B�	������d��PB�Kڠ%Q��=���J�O���5 .�)�����d踈B�'r* :�(sM���i���@Ћ
�'V�+��5U���Q���=�
\#
�'%��,ڙ-;e
E�J����':r��3	ش1궼�t��d�h
�' L�Y�<Y���4��z�j<Dx��i�.^ò�2&���p	C#��	9�C��lO�dbi(XШܚpє9�B�ɋ �8�V)�nhI��'k�B�I�0���f��(b��p7dɩ�C䉻Ķ��*�B@ G�d�B�D�TP&M �n|⏉�0ܣ?a��δ����O���n߮�E\�{2��B���L���<?K"�'4"�ȖTu�R�P�_G2�ȡe�O�i�wd�� ^�O)�ÈW��LȠ��8,8�XJvM�̜�OL.-�`�ܹ�6 I�� pP�Pl�'K(-���?����J��,T�0Ún`�yhf�N��d"�O@ة%A�1sY�D,.� �L�8!��}B��<ђOa�����2)I��ҡ�uy���$I���'��V>�I����p�II�^�IϘ�(���4��+yv���I�<�d]�߶|C.)��!ӷ�M�T?��|ZEJ��0�Af\� �LMJ��O�<AmB�)
�;�ȝ=40*�`F�Ɩ+�&�݅q��,'>�2VÓ9ʾa��oN�^�-IE�g������O��:?%?��'	�1Z�`L�y��X
C�j��52	�'�ҥ@�	;�,�:��R�U�F9����_�O�B�8c>vn�������n�s��'A2�'+�=�p�7y��'��'����'�UP���T���rեԮV�L���V�!��6�T�k�h(��H�����'��'Q~9��Ƕ
���u'�� ��c�)Y|����� h�YX��Y����Т�M�d����҉k�"1�EKCA�0���<1^�I'����Oޢ=a�'�@	�._7��!�I�d�'�teY1�u���4*]5!3���)�HO�)�O������ү����ٕA�%&����`�F��0��?���?����?������͉j���"�_�`,d����	� P�bN�ED�e"��0��/��=j�[!+ײ��:�Yݼ93d�O������	0�N��m�t�6M�E}~c��Ȇ`�O���-Օ A�u��� t�����O0�=ٌ�D�{!�Al�]|�m)�N3R!�߭p�½S�О|D�y`n�QQ剛�M����y.���O��4�^���@�,r'�`����i���2"�'�`-!��'���'��l���	bEP��b���]�T�4��Y���7�TId�J_"<S�ɠZ��%��DM�:��#�/�]�TeW;�F�;�D�-���
%m=ӈO��j�'���Z�[b^̻a��BL�!�D(��q~����8��	�=�V�
t�a�ꋟ;����T`y2j��l਄صO�cB�H���A��7#�����3��'��ә|��$����r��V��4tX0
�+�i���˟�B�2�`3b�	&!�I�4n��k�'v��b)H�T�8x�*�	ڔ�	�5���"L�D��ȱ5�Ţ����W��9X3�9��t�&u�c���
�]����'�<�1���?Q�O�O�)� 0L�g��{:~%`v�� E3���"O�TõE�1i:��$e^5N��q�퉏�ȟ�t"��!J>��L�+]Z%yQ��������3�y`Q	Юؽ���9��!3e�P�ȓ[ �4�	N  zP��Fe��ȓQ��u��R%P1%��w�<��ȓc,�T�s�^�T�lQ�""5�l�ȓxC�1�A/O
f$��	E|q��	�})r5�%��<�^��U��j_��u��^**T�Iޟ���ϟ�]w�B�'��I%B���qO�+Yz�5�@�߁kf�x�F���Aq8<�G�3Z ���P�x��۶gz���Z�:"08���ƫ+�VP���V�dq:��.<OX\���'�d]�w	�#'�������`�0a�'���d>ڧy��ś'�W�t rq��㟐eg���'�@�p��#®����3i�q�-Or�l�ğ�'��"��g�2��O����2H"G1���˴��-��$��9p���O����6,���1�i>��i�d��K�� Q�����$�7L�G�D�M�\�������>��@p6�Т��O�i��'2>�z���h���S���2�X�ã�?D�ԙ�hQ5+�BhAEj�Z�Iq'A<�O�'�¹yo�~g���E�K�¡;-O����O�O��e~��
�@T���AŖ�X��j\HrÓ�hO�t�u�ؓ b���f��)���
��d[��'��ʸ0�m���|
�g�=���{������'����N���<�r�E�oy�|��
.��]���:��}��O�ɥO����>�����h�,c�z�@��?M�td��߇R��4�O�����h��$Y!_�:��A�%\dD��"{�� ���>�r�>�D�Gy��Qr�$���Ĳ�M��	�E9���"�?A���S���EV�?1x F�<ָب���\̱��ԟl�sm4}�*}2�O���M��%á&6�袄�Áb\������Yy�S6��	�ȟ���A�
����KlV,\�Bk�s?�F�W�T>��>(9��R���P�+Cw��6g�1#�%jd			��䛟\���d�O���6O�c>����p%�!7�O� �x����Ol�Y�'z�p�O�s�(� +�������N|r�2�+ϖ$�\lSCF�OtR��n5�1�<`�)��Y�U�i�ȓN�#IF�<ǮM	�*ҝH||o����$�������f�ܴ�x�	a
Ф\� R&��X�E�'��P�(G{��ڀ�J�7]�V@I�:4E�����x��)�S(N�����az�J�/	�>B�ɯ j�h0��?{�8X����,��C�	�l��0������aW�X�C�I�7T��̀�1�Yy��:EU�C�I{�=P���;�|�2�-��vB�I�~�c!oƈ5q>�ag]4[tB�I�6��@+�&�Hp%�aܤB�	>9�4Y� C��h{��!|FjB��8آ�r%��f���#��ZB���a�nч!H����`W�
�RB�	6R�z��l���R%�:B��7�<)��,����
�3��c�T�셧q=�P�R��,�j��"ޯz�v���#�^��Ǡ��%�JGAʺ�
Go@�q�ٸ�l¥~e\Aqg*��J��$�D�����싔@}�J8K�iM�E�n�K�M�\�	GH
d��XfiC�^��d�pAV�z���@V��]��DB�nH(0m@�.�Ra(kBN�O��@��]<i^�ASզO�9���O�䗎��d �|�'���e
�2�Y��K�H6HjL<��i�i���O��)�SB�x_� ��0@O܁"L<B@\��,�<�~B��Ǩ9��L�V̖�R&j�"�K`�<�]�X��q�R�	>.��Q�d8����Ԝ���3#ȣ"+��`����D���8�OF�X�Ə�J�MІ
-nn�,�"O�]R�N�G�p��o�X�n��"O�2�J��wvn�P��N��܊�"O|$��A2�.P��(f�"
�{�!��A��x�bE̼Vy���F�J�!�ć�a5���b'�Z@��D�1P#!�]}z�b2"\�3��j�\�3.!�� �!�㩗(d���CD5�"A�"Ox�#(]�-�R�S����E+�XYG"O��6��k�e���P�#W"OZ� ?�8ySvL�$>a�M`�"OT�"C@���A��6�8�O�0L!�d�.�,����4�^|�j�wC!�I�	�6ax��\�� ���#�0�!�K�C�4Q��Z�D�b`��ʛp5!��
 Y[�C�&����'%!�	�F��4)R¹7|�\scJA"!��,aWFtBr��2n\���&S�\!�$�E֔���F
R�y{G�5r!��F��剦d�:?V����Ju!�ă�W� ��CƸ[>����-!�ė@��Џa* d�$I�0p�!�$��|l�v$=� ��H	3z�!����}T�0
�J 6;� B(ZC�!��єj:�{�`©3$�	�q�#�!�J	|�ҩJ��O �8�C��4�!�W"I 0�Ӊί)�lybGA&1!򤛧S�����&p)ٶ�N{���Y	�'�ε��	NA�i���_�4�a�'�B}�֧�]~"}���&	�N� �'��2��ج��D�6|O��
�'���RO��	���\h`���
�'�R��F&I���#`��	��E��'��MCqb .,\(Q��h�03f����'�� d��(�%��C°d�t��'�Nq�FM	t�t<1F  �(A��'K0R��Ѣhjޥ�ud*xD �'��娌-2� ˔IZ����'�fd�E�.{���7Ɇy,��'�%��F��{t0a��%%^�
�'�@I���1I�ֱ����z��'�����u:f�ҠOٙ���Z�'��M)�-��=/¹���1!N�h�'���qH.'��`�'��1� ��
�'�8��eF�Uh��z�k��
FPq�
�'Լl��2��G���8]��'�b���PGR�)�� ו�.q"�'���Z�*ԗ;�RV R�J0'+e�<��W�CYD�3bP�O���ǁ�u�<��JJ.(�1 ӗRC~��%�L�<�KH�!�<��R�F�tEưC kF�<���I%�c��vd�0��B~�<ID������
G�s���@D%Hb�<ѷk�(�F ��%f�VP�6��a�<�m�'uՎ5���g8.lHL�`�<����<�
2�L�7�"�D��T�<�b��,`\ڽ���<P�X@�6�Mg�<a���K|��R�7�p�S��I�<1U @�S���F�c\��"H�E�<	D�M~�<��^�]lЄ�0��x�<@6_�\�*`�Ӝ�|��$O�<!  J�h[N�Z�MU�)*�	r�<Y�C� $�((��e�H�q��j�<9�ǉ,Yn[�h	�g�����̝�<�ү��GPI$�^��B	G��@�<!�u�"I��K�*6�	���w�<��iO\��+�LW�OH@8ӧ�t�<!�f�PK\�Zq�
 �>�$�Z�<Yp���K�H1Q�9�6q���R\�<���̖���2�)
�o��LJ��a�<ң�2�����OH� dk�k�`�<� ,9�$Ɇ�w��!vl�-iRg"O���!!Ɨz����,��V��A�6"O��1��&I�&e	@+�	�v��"Ok&F?h X���H�1h�@�p"O~�9����y?v����[X�C�"OB�腄\�F����0-ƖeA"�t"O��I�l��AxL�I3׹4��1�#"O�4�4I�1#p��7�ԺG��cw"Or!����}�P��Ƣ�9bGr]h�"O�	��oh|�� 4E�@��"O^m̍0;x�I�U"K�n}�3"O0��D��G�<tC�%��G"O��$�F7Z��%Z���4�Z�a3"O��Z��#M��e�G�-��bd"O���ģ�M�eф�M�OCK���y�'	R񐁸"h�3b��H�N��y� ֻqj�2�[/%�tT��*I;�ybO+j8!�]�������ƫ�yb�۔>ADx�FQ�l����
��yBD�x��P{�͟.4&�d��y�dB�UeЍ�Պǂ��9CQ�N�y���~��q�(�l�*�e� �y��z ��G!ףd�0y�S���y2���8Y-�0L��R8�y2��fς\s�o˶s�li+i�7�yb!ѵ\(��A�4F���� ��yB�K:O�b���n��ݱ�ǡ�yBf0e��d�P"	�r��`cI��y��E;;�$j�؈q����!�'�yB�Gx�6�{�H�=�m��"��y��Z��dB��7=�rE#���y�b�:�<�/?��Y��ѡ�y�hS.n[�4[�n��/�bة�����yE�"c���$��']���&��y�J��$q�pE�R3v�� �I0�y���J�L���' ���ٰ�Œ�yBc>V*	�%��(w�M�p�ϝ�y2�Ţc�\��ʘY�0%�gJ��y�`��#�n����<�2I���y��O��5�	�&f)8����y���Q�5���9"�ak��y���Z���z�eؠ[�`hFa��yB��(eP$��#�1m�Y�� ԡ�y"ӯL���3���g�8� 	��y��"����,ρoR�C����y���~�́0��k�����L�;�y�ʖ�$
l�)�Y�hSh�W*5�yr&\@Dfɪ4�ȋ��tӦ�G��yre�^��`��<bm:4�T+���yb��4��cG�S@�<K����y"�Q����J!�F�2ux�k��y�M�B�B�kw��5=/�t"��yb��pך�� '=��Ńw���y��W�{�P�ÆX<q�I���yR�I�S~N�P��A*�^���ߕ�y����?��̠ n�= AVY�@��y��%q'Dൠ�����L�y��N�~ɑ�@'*�q�ǧ>�y��P7q̱��J�;e�l�b%�yR�8&� �?�v	R��	8�yr���z�6H2E��jd���荺�y��	�=6J�9b��jmࠚAj�	�yBB�d���cK $o�Pi31d �y2��F���de��nBTɕ��>�y
� ��	.V����&9D�E)6"O���Ӏ��E�JI�����$
���1"O��Y�x�B��UF��TW^���"O��	Q�>/5@ݪ��I�(Dn��"O"��5�^2w��p��S�l��\i"O�u)�(�UeV(�1ʀ�|��`"Ol��d�GL�4ٳɎ$q��aP"O�Aj���*��Yp�G�*JREs�"O-�Td��QL8�yW�
�<b�m"O����L�ಐ� 'H�6�>;"O��V�3%�=;S�g���"OT��3�E�	�~Ӏ��l{�"OHAbv�ͨQQ��HA�2��r�"O�%Ҧ+�̍�C��B�����"O�Uh��@�aq�Db�_�,2F"O�"aQ,F��r�+V~N<�R"O�,�FD*$[(I��To=��S"O�XbB/a�N ���5`��a9""O
���$Patd���M����C�"O ��蕈np���L�l�
iPb"OfP����2l;d����1a�옷"O������.*pJu��:Ʀpv"O�9tj]*M�������]���"Ol٨�nŻvt<�K�Ң%���y�"O�җ!�
s:��b�Ӿv���xA"O��b]/#Bt$���$B�
L��"O@q�P(�1&���n�9�Tq��"Oh���(\T`8zqN�%�r"OF5�.�G8�@ы� z���"O6̀4�N;$yNd�d�	:��@�"O��A��9Y(F�P�B��F}�}�"O&���HI6V�M���Xv�����"O�q�5�E�<H3B��;�$��"O��2�E֬Q�t#�O9��4�g"Oz�i3"��] @�@-,��l�d"O�t�pG���A���)X�"O�5H�JY�5a�EѢؒ&�"O�X˵�Tws�(��L�5hF"O�\�SCP�W��-r���;��5*C"O�T�Lč_CP�h��وW��"O@)Bv��9>�K�*���F"O�����I�4��^F�rs"O�բ�ְt��|ZƯ�8"ա1"O��s3�ԅ\�f�w�Ie����"O��q���I��i0y��d"OJ�C��&G�Ƹ���ma!�"Ox�j�͑�N0RE��H0Z}��"O�x�)˽lKz�v���P��D"O�+�ˠ�+�@��e"1"O��)��J{�����G�l\y��"O6�&	�/L~|X���%&�y�"O���aI�u�t�Ń��Z���"O����A��Xx@dH���?�ܙ["O�̰&�D4:�����@�	xx&8A�"O���fύ,B�h�c*shR��0"O�hI�D�>+�(h�G!S`X�"O�)PƜ�k�4�"�+3Y��[�"O�E�`h�+Em�����
�;>��`"O}a�쏈/:U(7ă*%�*��"O��j�h֝cZJ��G�
9
t�a"O���r�G�spHz���"�I�a"Ot�	���$F`5�ю:ph�Hg"O��3���VR�@�D99Y�t fD@.3� h'DT������%<O���#�ĕE��Q e�")�z 2�"O� J��%�@�j%ʩs�@$ʪ�#�"Oj a�$}r�˅�P@2,5�v"O�ls%�S;y�lx b�~% \:7"O��f��A�z�� #S-]���r"O`��7E ��bY�V����5��"O��y�b.~Y0�`�Eҋiᔈ)u"O��0c�8|Tj��d�I5���"OP��F�ߤ}t�� �X�> ��"O���v�H��Q�@�^&d���"ObE9��H��ɓ��T�e3�"O"�v��$G���)���H�M!"O qR�NF��0S�B�}NT�R�"O"\�Bc
(x@�(J���/�e�5"O �k�"�j��t�$ F���)�"Oi�f�C/;�(S� iCT|�.$D�H�$ʙ<7��!���_.�Q�$.D��x�^>*����t�Ǩ �$�ceK-D�`h����ܨ��ٶoƲ���+D�Ha%�j��1T��� yǧ(D� ��n�.u��kQ�['"���J5�*D��(ܾs=���r�̢�v�ᇋ,D��T�j�~c6 �Ij�%VD>D��Ua�?z��pF�w�}:�*O���3�&����i��k���5"O��;�lL qc��K��t.d��"O�0#d�� O�̐�ε"�`[7"Ojը���^�t���+ ��;�"O<!:�+?�hM l�0SktA+�"OX�y���*c-�=3���tL>��"O�E��ol����ރs��<��"O�;�	 SR��̗-47�0�g"Or�ӑiïT��Љ#�	�\x�"O��b�B�`����U��O����"Ol�I
_l
);��^6yE"O��s�/9Ў-hش_6>�ɡO<D�x#�L�����A0z�8���L?D���1d�8A�p����D �T�7D��4��5�5B�ˈB.�b��:D�0��@�!4��QÂ�*f���)>D�,!t#�DX�p�*�`�MJ��=D�$���(l�*�@�a���0�/T�Dq�}kB�I�%�Lu9�mʷ f!�C�x��̅$FZ0H㌷>V!��oy�}�r�$ZΌ�7�8&0!�$�l��c�ctJJ��F*!�<!-2<j5fN�
��rDɗ�)!�D�zh��g�ä.�*�r�Q2!��	�C���3H�*t�T�kR$�J�!�ě�i��"�A;Q(@"��Т���䕫HI|�
f��0�^���K�9�y�T2 ����`�� ��DB��y2`U�0�4�$�1�=�
��y�%ϝ)6�a���LBH� ����y򉞺s[�5s�lX�El����/Z��y��%`�z	1���Mfh����y��C�	�2x�a������2�)�y��Y�V`<\�peZ�u�$�Q3�ݜ�yR̉�x���#h�=|H����y�O��^0@Q�6a�$q�"�:�L��y�I1	=�U���B����]��yR��+n����>L�����S��y2�Z>`������K4X��.��y㐭�0�t��GA8��ӊ-�yB��6t�dTS4�
{��8i�
�
�y
� B��Pf�-�H���Rl@n}�"O����|�̛�I��v��5�&"O��d��?����邖Q�����"O��; )&C�P���\X~@9 "OLȻ�*3,P)�`���x��"O�9Dɉ�1�(�D��1z�64;w"O���'��].��Vl�`�ܑ�R"O�̂3G�8Dp���5fD���"O� ����$N�jg��	H�HK�"O^DQ���� Sl�9���S�!�Ė��r8���DZ�p�`�V)L�!�D�zT��PB��:��A2�˂�Em!�d�-A~D�DG�12�<Q����
g!�dN;ވ��Kɮ�R���^!��իI����6@��H�4,�'��"mH!���qT٥����c�`Ұ"�!���(�Խ��F�@$�)�*'2!�D�-�!����s~|J��Ry'!�
�<�X �C�;D-�w+�!�DB�C� y�h��������D$Y�!�$A);��g(ßw�
���! �!�Z'-<�v���)�T��0g%!����(���+�|xɵG�M�!��F�D����h����HހS�!�$Q.i�$`5�ѦW��}��o��4!��¡h��(2eO��d�:0n4e4!���>A��@�V=6\�ʤ̊.;�!��R�W10��$ƙ=�Xh��$"O�Ჷ`B�H�NI3��T6LU�A�G"O��Z�f��9�6�������p�"O~U�a,�xf�}��{��PW"O�QS��.�Ȥ� �3���c�"O�Hu�%s�ԙI0��4o�Y�B"O�e����9�n�Ƅذ;u�5��"On�0'�����ȡmlH) ""O��HoV=S[\a��$�?)���"Op��B���L����� FДA��"O�	y#�WL��dSu�^�P�2�*�"O���K�]�yS5ƕ0;:P�)4"O�{$��,YE��5��W�c�"Op�G
A�-��d��hP���a�X�l�8�"}B��6��H�I�4`��Y{�B�ɯ9�0��^w�6U!�S�#Ll�Jn�l�JJ���<)6	�vt9քD W��u�NpX����& E&��gL��ffh� �U�80NQ����GF4��O�DCT��Euе���U�9&~IFz�C���� �E矂zhq�8�W�&.���t��krh��"O򼸦��_֐8HR]�1�P*߫+
��a��dl($��-�O?�	v"<��tLܽ� J&pO6C�Iik*���c��z�+�
j��E��@�3I�W>b��FMD�'/P���E�#����S�P�ߓ{/*�2E�P���E�E^Ȫ�fėE���I7�8~1XUZ@�5�Op��E�.��-ڇ���EXD������%����<Y�IM��$e+��6�]�Q)PE�P��HB�S���A#�S�I+8�
�D`�<I2A�O=t�:䙰�S�0ͤ���#ҧ�~"À$�4!������H	0���	�y2ƕ�<c��|.9K3�Z
�\h0tÃ6�����j��t#���[w�Q���&$(������$u�H�S#(lO�A1���0	�j��!\I���jP�H8u����D*VGZՒ �X�F����Dƒg_lڇ
�8��sc0=��O���D�Y˞|{�a
�@�?��RL�����kT�� �˰�y"�#����'�g�89�g�R� 3��غ>���sbh��C�����I��(`�*��a5�%�"��޴�5�8D���#I?4䑄f�Q�� ֩>1��t�Ѝ��eĸD0���� �P3AfZ4Y����G4`�U`��'P�b�܈1Z����V~���%͊�^�N���Z�?�AΗNQ�� &M�������o�'��}�-J�O�ҥzM~�g�ՒF���B⡛�ˢY1GN�n�<aQ.�	��$�V���an��<1���j������"E�Ś�*v�:%�؆H4C�ɛO�á�K3�AhP�ہ��|fŁԨ �C���F!6���
H�t�Z��:	L�}�
I�jUfk�D���  �� S��
FK (e�I�'�dp)ܽ�h���[�93���X&��)��	H<���r�L�#Z�9U�׌_�!�$F�6	�LP���'%x��H3
��/���2t�<(�?E��F�YY��ӏK$.Z��'�yRH8f@.L�6�� ��@�Gۆ�y�+�
�l���Ӷ'd�1�1Ԭ�y"�7��s"��X8Yz֎߼�ym�W;6�QޅV��C�)^��y�?1R 3�N�z�J*^��y�%E�PH��
�V��7j9�y�#����tbW�!m���'M���y�I.���i"f�)[^|i����y�j�&T�24�gΈ��f%ҡ�y�靃M�ԅ�	��`@�Iz��A��y�"W�9�TSG
A�bTv�ʅ�y�,��MLh9k��A)n�^�r����yR�@$���{&\X����y��ر��W�6m^p�!�'Z��yB�֦2���P��	1��ˑ�/�y�O�5��<��X
� I���y�O�1F8�+�gG�N�y��	(�yb)?\CN��Δ��L�%Î��y�Cʒ=�OӤ�D�ҡ��yb���f/V@�⌑�6���b�N�yR�ЫZd̡S�^/1��yIčИ�y�"��g���r�ݵ���g�P��y�G۪uH�Q"rN\4T"�j@��y��v5�1�^8�\T(�%Y�y�c������vK;t� �Po��y�`Q����O�Ȝ݋5�^HK�B�	�N�,� ��AM����1��.֎C�	�^�mX�`A�jDd�@
Q��C��%�B�z���e)F�ٕÆ�C`�B䉃2[z4c�'�2+A�����ߑC(fC�ɂ/�HS��e � �UtC䉙�@�a�+�w��M�S�5�"B��(A;j�p5��yS���,�j�C�ɤ���P���w|f��+�$)|�C䉖~"�$�� ��n���C䉧V�Y�v�AN�4!�EFM�T�C�I�7� I�E�2f���%F�
.N B�I0��C'�HR��C�O�rG^B�;^b�)cb���9܌l�B��WE(B�qF���� 
*X�hB��|`BB�I�
f�с����")�F<�tB�I'~�4tq�<ee A[V�Y)C�4�<X0C��Vԁ�phҔ..NC�Ʌy�%�#��v�^}�%kP�>Y�C�	:NN<�@ 17S��M��Ik�<i%M�'O��]��BS�!�(���g�<�3�'\�ȵ{��ɀy��ғf�c�<���� [~	xg)��@����#z�<1��?:+j�J�mK�i�ोr�L�<�҇D� u�� 3+����SV�RS�<�!eFQ�@�u�0@e�n�<� ����H�,\��Q��@�?j�<�3"O�9���)Q&��gC8*�B@*"O�Y��4D�Ga͖��[B�D�%�~HB&�QTVl�!<O�@Q��+�<���u/*�K0"O�qh� =i���"퀔B'X(A�"O.xC��/X�L�B֪@.ԡ��"O�`�ج2�<�@�(�0.tq"O�	��Ͳ^�
�"��P/����"O�e�2lJ���Y��܍�d"O6��W�
�gb	����{�ĉ1�"OpQ���$i�Q�V���<&�"Otl�p$2W�$	�ul�@%0�0"Op���	��S�L0�ƫ�$��"OxI
�J<pn��*��9�.h�"OT!��LVGˤtB��Z���	�"O�ݨ���/:B�h#��&▅S""Op���˛�'�y�4�R�y��t�P"OL��v�"S���R�K#��s"O"�H��Y�R�����p��iB*O��5��f$�q�DZ:\t�Ȼ�'|4 ��e�G�(�t�#Y���'�v\�$2	g�t!"��*�5h�'�0m9��Y1Ik���!G�>Z�l�1�'��`�bP>w$�0:����m��'ܢŉ`/!|�м���A�,�x�'L����YFDP���8b;� ��'|p`+n�n��P�F�,�@���'QD���ӭ��pS�T�|9$
�'N�+e�_]��-�e/ ��ٸ�'���v�U�)�8,�$oMR�D��'�6���`�����ƹt�p!I�'�l��Q ܇݅�fe(�K�D� �y�EG(<�P�Ї��e崹�(9�y�!	��92�V��	r�*��yR��*Z���*P��NPvI{��H��yR)�t􉊤��D��T	���4�y���,,�P��b�>:�X��NS��y���2d�(�Z�&۞i���IRF�1�y�ڳBjxK���a����*�yB��qs��2�b��_��!i�D\�y��Ƀs�tY��V�>��!��%�y+Ƚ��P�D*�I7�8�T�\�y��C�VR�2~���SB���y�O;2�^���A۔'4�3���yZZ��4o�H�$��\���ȓl�A���ݭ}�~�X��U�F�����s��M�����V��/�y��j]��Vk�Z��m@�&Q�l���ȓL���Ba��*qMpa�1ζz��Єȓ�3øm�t�O�|��¤̑�y%�B�������r.����O��y"��l�-���՘?�&�{p���yR�L�3{,�`�TM��M0g8�y�̊j{l1b M�|#��Y�n���ybHQ	z� ��SaB�p^X�@i��y&�}9ڥ*uBޏO��Q𫕈�y2��"l���"�H��Jx�7��yr΅���೷�Y&h�=:GV�y�/R�0�Q �0A�t��V��yRĖ�`��P�Ѻ9=`���.�y򀇧T;���R�0��1�R!]��y�N�I�ƀx�KV"@�S�C/�y�>��Q�wD�5j�r�a�b4�yR�V�|�h���9'-`$Oȕ�y
� "����M*m�$�F��?�l���"O��r  MX�
Px%lW�<A��"O�q���^$f���A����>���"O>����I�`��1{��J��Ux�"OA:�#5�T	J�'�Z��� "O0���z ִ0�В|�\\i�"O�l�� �n�%�@��DX���"O>�ᷮ��+�J�q�N>N(���"OL�'�޴o4"����Eh<��"O�D˖ʃ�2R�9���G����"O�������|+w擉t�5�A"O"��GJ�	U~4ڧ�$7�&m��"OnB��@mҨ+��C�&��=�"O@��ǖ�1p���ц;��'"Ol�"ļZh"��EM��/(��"O�����<Z�r��FB�[+�+�"OPYj"�Ŵ �.���Ҷ
�B���"O����ϟcZ�ᆦ�����"O��9�FG5d4ʤ9B��n����3"Of��է�F�t����M�
$���P"O��	��#SJ��Q�)nC,��"O�"�K2.-�y��ډC>��"O�	w��q���9���]�"O���FMR�];���VLZ�x
�ᨷ"O���unQ�
���H��<�Dp!T"O��P4됐��{W*	�LjJ˶"O�9+1�Z�D_�y��	��, B"O^٘��ɜS�����J�I�Q��"OU�5@�#4by�o�X�>	)�"O(�c���O�ぎ��	#"O�a��ɩ[J�谬�E�0��"O�3l�Z3�{�N-V"O�V�7 �@Y�#�2 6.���BG�<qt�6`�&%��n�B��E�F�~�<�5BG8{7��6��x�̓��{�<9Wd�.4���	A�o9|e#F�J{�<�S���$X8�p�D�B�8�x��MP�<�E�M�L� O�Sux�	5��Q�<��l���ph�l�:�I��i�7�yRG������e�M���ᆧ��yr�!��G���rܭ�����y�·�sc"�3��cx��5ǟ��y(o�Q��[&G�b��7 W��y$P�}�$d���F��`#���ybD�>`$�y�[Bk0�w �6�y�ǂ�p��$G�����f�9�y���[Z���"oK�8����L�3�y�늀ʚP&f��*�qC�iW0�y"G�FT���V~��a��y���4j|��ä�4�B�V��yBA�+�j�Tҷm��y"���J�d�2f��Q�^Y�h�1�y�G��\�� �}�@�Rs*�yRɞA��tʈ�B\�I3����y"�!L���K��ѣd@�R��yr!GkvE�eg[��	��H�y�"G"1� `���N�A@�ȇ"��y�
-u:�!�a��vV������y�lG�3�޼q�lՍr� {B�X�y��:����� ;�V��-���y��I�"�d��Bэ7>�XF����y��Q�a�)���7?zFng�x��'�*�!&��$M��$�/?4�H�'ŚF���lH�yP��\>(h�ia��� ���jC5KC�Z�ʑ�i��	�"O2�)P ��+0c�|\�@�""Oj<;�̾6��K�C�#&bA�"O���F�ܱPY�0r�АB����P"OnE3!̛#NgBq!�!�s�x�H�"O�m�J��.3���!�"(����3"O�Qh��P4�s�I�(���"OH)	(��1��#�`��e)�"OH=te�<+����F@�PV�J�'�*��jZJ�����ЅS�'�&�@E'D(m�r�RB)ר{�<��'��*d�?8�<R� 7|d
 ��'�L��,�[(��f�4�j
�'��c��K�t����<�Q�	�'(�t���%sgM2~��Y	�' P��f���\�n�G�#(u��'��	8�,R�{��@gjY%
�LB�'�x,�1`ϟF�,IY�,�3�*y�'��\���$MW�̈vO,}�J���'sp(�'��;r�0.EH�,�$N�S�<�#��=I��0�p�S�ntA�f�Gw�<yWk�s���qE
 �*4��x�<y�LE,?��!ڦ'#�v}��e�J�<����8��Âo�I����� �H�<��"=h�g�Y�@�r�D�o�<Ad/\9_���q�R"v � �
l�<I��F�7\X���+Âb�(AT�R�<�rC�+ZPԴ�� ɼz\`��MJ�<9�˦e#�p�:�.�@�g]�<����u���Eؐ��p�<q�����I8�BL*w�� ��Yj�<ْa�r���.E�[np���l�<���W.E�$��Ɓ;%^��ƌJt�<�UC�8���J ���(�Yaf��n�<�5�Ԑzj��r��t���h��j�<1Ǣ�[��%�'�/@�`Ѐ�^�<���,��9�7fL�N�,�8�Zu�<��;�:`�6�)2j|ڧ�Ms�<!�Kڄy����Ɉ!��9��r�<iQ�<z������0n0ѹ�NS�<Yrˁ5Z�Ne��-�:��y�6n�L�<Qcc� n	<�لfK,@j��5��N�<o�Lf�@�D��W�ry��ʏe�<	%�7+���yu�!&�8�/Cg�<�P�^	ŀ��u��O�T�0��`�<I ���*������Z���yc�W�<�CQ� �<���|
�!9vAX�<����P��Q��-,TX���W�<�5O�4��-��,TU��7�:T��v޷KnP��	�G(��8��/D�����[.�,0S�BP
�E# �-D�0i�b�!mk�[�H;M(n�Q�B-D��ƍ7��A�! ��9�)D�`H'�I�	 �)�C�+l�<���'D���p��Sٌi���
��}b��&D�����`s$��$�A��u�v`)D���%@�O�p���׸2����:D��B�̙1{*�r@� �{նD��*#D���ek
�~<}R��:B���B�,D�:BN�FWt�׀��P���5�7D��y�'И'De�ߚ9@̲�i��6D�\�7@�]Qb��d�.;��T� �4D����MǠU���3"v���A2D�("�����j�%Q:-)|��ul0D�� �hH�͊�i�l��R��s����"OR +1�*^�r�pN�N���s"O��Pb�D�Y��6l�4H|�pz�"O,���&N�2���K�a�z�D"Of�*�������]H�L�"O������1� F5x�.9"O�����L L�,���P�M�$��"O<�Yg��#]��#�3A$��S"O��a�2"��dD��G;Z���"On�����!��m"���LZ�v"O�x��$_����3�
�#��s�"Ony��D��]�欆�%��Y�"O�x�"KOg�t���M����"O���+�����8э�7?Z|b"O0�`��2��T,����AR7�!��H[ 0c4$T�	�P	a�ϖ"u!����^(QS�%�6����;Y!��Ǚ#2��V���1�r�\�;!�:`�H�	�
M�g�4�@�K�X1!�N�d~��3�i�6�jE�����+8!���`
���@�!j�,�'�*3!�@���}S�� &s��c6�C'e�!�d��a���$ŴRTF�Y�	�f�!�d��>��!k��uP��w��N�!�D�<��D�� �P��;�Z6<!�$�?U^���mB�B��L�z�!�Dt���A��.MT��!���;A!�$�4���&�X:i(� PU��!��L%���(�fD�'&_"�!�$
3�ܸ���^��R���eA8}�!��9fA�K�1��Ya�$�+,�!�V�{���)��!�.�V���!򄊲\YlX 0� 	�WA�!򄏆n���g�H�����i�pD!��f��;ɇk��9�hƫ-V!�$�6=�8���e�%H��1B��Py�k��.�����e�*�|�A�K��y���~�XQI��Z�yt<}�'/D3�yroХ+���7/\+c�B=�q ��y	V�1���&�d�� [9�yb�۱e	phr�`ޞ��g�O��yb�ɤw_(馉Q~>�)Tc�
�y�[=}��+��a�3 �'�y�S�H�4tC �ܗ	49��o1�yF/ւ%Qk�v����6�y���(c6��j�/g^�S�ύ��y�o��C&�x����Y�|� #"�y"�R�*�T� ��Q�v8�gJU�y�13��]x��XO�(qq'JX��y�ʜ�T����e�}[�����y��M�PQ�Fq:!C����y�N#1ZP���p4I�TO���y2���_y��,ݎZ�������y"N�����E��|<�\�"oD��y�۞3NT4�I��y�v�)����yr"F�o`Tݒp@Dr<h�@B���y�$��a6�}2��U$Y5<��JT��y��χM[��EfJ;a�*`���y��C�SFe�S�W�S[f��AE���y�N(�E9����Q�@�+q�
7�y�o�P����
�B�x(ቐ�y���jF� �E��f@ �"G_��yY	i�t���
�YѐA��	��y��K�b�Z\
A)H����r%�y
� ��3Ўu�n|krJ��oF�$rU"O���jE�@���f/y7����"Ol�J�"q d� �K!QxM��"O�1*����؛R�J��kR"O�e��&����"���B�V�*""O��ڣXjL��ԫ�^�|�j"O���u�JK��C�J���\q�"O�[�gY7�8 Z�*D�z��<&"O�x�wѷ&Z�L:����.�t�Ѱ"O.e�US���D]P��9"OL@�C��94�`�
Â6R���u"O��{B�'^�mA�A�$j�>s7"OJ5�A�;[v b&��u���Ӱ"O��6'KO��O�
}�SS"OB���h#0��� -��- �"O<y�����(��i�-� +�<Q�@"O��CF�M*,�����+��"O^M�6GؼMf^�
兴b$ "O����,�s ,,�%
f�T#p"O��:�B�>H���gĊ=�&��t"O�X�q���cɒX[Q��?����"O�9�"R�f/���ebH�R����"OP�ׁ�sĆ:�`̿+���"O��"(M�h
N)��A��V��QZ�"O"�
��:��!��� ��uk6"O~ly��,t؆e��Z�Lzt"O:BF�R�S�i�N�=xkT#"O<ɲ6H��XU�-��bA�b9�a"OP�Bō�??��[���"c<�}0�"O]Ѡ�O�-�b�a�h6�`�"O>Q�� !h� ��4 ��"OzY��+�#�����%W A��z�"O�
�9x��s��$ ��:�"O~Y��R��}�%��3T<�F"Ob�C��ZǠ�X $�	m$|tcB"Ob;Fh��Z�|�Ô2(����"O�T�",ނq��h�"�T"O ��V(�_r�ђ��ر$�C�"O��ғ�%r��8z��_�'\(��5"O��  �*��JТտ7Zh)�"O���DEJ�#�P8+ua�r(�X��"O\X8P%�V<���J.xz���"On�ȥ�#g2��%�֎Y^�[�"O�9"c]�ZiX����M�7MB$�"O��iŠj�q�]�i1�l��"O�t[�N՟BY��r���Fe��"O.z�LJ/G�: ��L�Z�,"O�A��	ϖ�<L��Ă������"O��S��A�(<��v�R���8y�"OTUٰ�F���BJ2:�Fm��"O4�K7��61�2͛����d���rc"O�p2���6����
�Ht"O!�a�d��󬔋dTXD"OjE��!�$��ՌXy^��"Oȑ!D��1P�,l����3q"OАc.�x�,A(��	 �`!"O��	�O��^��P��N�*�[q"O�Ae�*p܌5閇"^�ꭣU"O��8e2:n(xB���/\���"O��Y�̗6RT\"����"O�<�1h�%7�ȴ; ��.]���x"O@UCfe�X�0<A��8>x:mJ�"O �+瀁�<�����D�%lX���"O0$�R�7[ͼ�/Q�B�\��y
� ^�ۦE�]� ����O9�9�"O���##LD�2�;�,L��{�"O65j�jD�W��e���0iF��"O�� ud�{��9c��*H˥�'���,#BB��&��� �}�����-D��a��C�"}�D�w��cW�D* G+D��[Ł��J���C() ��yGK=D���a
-s'v �B�TC.؃�;D�d��HLl�)r��D:N��N>D�@���5���s&(�����0D�(��7w���2@�R�(�
D��H0D�t;� _/���&kK�d�Թ3�"D�$1i�}w��H�ɏl�z�2�� D��J�J�0�v����-�d\�҅ D� ` )�,50(�6���:k����0D��l¤g�6�zbA�.8v�Y#�,D�,��/~@�l*�ɉ�	q6�B��5D�a�Ê��ᛆCIy��m D�P�/�q.�@��?R^ m:�3D��S3��2P���S��9fҶ%"!D=D��x�%K�z�xР�Z���'n;D��k0Ĉ�"R���处Lk����>D��X� ��_���3� [.���M;D���!'A"9�>|�m�82`����#D���G�D�LYx�"p��z�A,D�,aU��:�JQKV�)D-+)D��Fi+3
!�ď�J�R�:��)D�L���ѐ!�J��թ�8�1��4D�ܩE^ &^���&ҷL����(D�Г�&H 6;n|�u�>f:���P`1D�d��&�=>v�p6�g|�H���.D��c`�O!M��4l�$L֔d�#'D�Ы$/������iQ#c�<]k��?D����/�f�,![v��I��5p6!D��r�b��K.�|��
�[��a8�
3D���6䝩K�&�Q�F2<�^�{wO-D�d+����
���J%>�+T�Q~!�dL�s�H�c��ƨ>=���"Q�j!��ɯe��p��9���R��W�C��B��4\����@� Y�0	�CT��B�
?�rB�� �io����i�K�B� ��2�ԶK�⭂��O�4�B�	�_�Ve@g$�y3��pDc̚k�FC�ɑx���#g$\#���xdL�	OBC�It�4��B�\*i��1�C��A�C�IK����n�h��!�Ʋ�B�I�|D�B���]��|2M=5��B�<j���X�"���B �� ��B䉫T޴�bsƅ�@�6<
A�>ch�B�I�\B���Q��4Йpf�M+��C��jxA��؋l����С
��C��&f���	&3��y��Ƅ6�C�I�8�n,
`i�S��Uk�"�C�I�f�� �@@�1�}��/����C�	h�pȉTG\�_��1��
��\��C�^�����&6���%�Y��xC�	(@熅��fF=t��+֖P�:C�	)$��d�Ī��
����'H)�C� $RHmX�gR�8��E[F}�B�� ލ��)|�8�N�p�Lń�~9h��'�DC��s��D>󮅄ȓ .%itc�^�Y[��/U�u�ȓG�@U��	E) .� ��D��E�]�ȓO�	�ݤ	x"Q�ܑ/������ B��d���+(`j�'S*~��"Ov��N[�4b�R �Q�=<*�"O��x��ڎ+ �`{TƗ�y.��0"O��i"FR8z�<�F�*`�l��"O�	'�ͷR��uc_bn}�"OL��GI5*��+��Y���4S�"O���B��1��g��%r��YQc"O`�A�ψu��iV��7�� [@"O|5��������p���"O�<R�ލ	��i���;�Zi�u"OB�bE�H��B���b�������O�hq�����M��O?�ɷY�X���] n����q��i8�|�U.ؒ(��!�l��/�*q�e�*mل�>I���"����ճnY�0 ��|Ҟ�2��i��-{'뇔>�"(
�hՓi���@O:��C��F-(ךa��ʊjd|��h�ԦѠ��O|��Ϧ	�	x��M�歗�V�n���H�>u���L?�����=��4P��Qh<������0q���Fy�y�0��0�SԦa� EA�zVaz��]20#(*#����$��ȬlYX������� PQa���dLb³J\IV��0�O@'S�y0�"´�.������"<q g�
9��R��N@�H�����-10oϡe�&d�b���O}|��O�#<AP�8j�f��h"6yk`���L�:`�2@s�p좩��Iǟ��'�HB�f�V�4̡A#I�l���z瓥ē|H��F�C2�"�`��L5_�R-k1H`Ӵql�e�I;�i�<�W��<,J�Zv�]-3z�HI#�BhҺM�a�ת��<A��h�Z��2&�"F�2��r	 �mF��J�HH��:�(S�-��8�EG�{�X"?Y��Z�W�N�a��#��H,�Re`�j׮��F�인reN�J���	;v�x��x��1҆kɘ	2�A������ƞ�M����O$�ʧ����HkUy$�Ae=^�z��>���	�
K~ 1���
٘؁�'��6��Oʓ3n�mV�i�r�����|�d
X �� f��*l\��{��'7��zV�%���QM��������|�D�]�,���+�i|�((@�r�'�R���L܏i��}�V M�6��i��t>��H.ڄ�FbI�b��}*��5�F� t�I֟�I|�شZVZI��PP�B����N<��`��'�O�Si�0���补�F����g�6~;����I��M[��i�����nF��7,��h�X�`��;�~��O�����?-$�0�cN��GVu����N�4%��`?����""[XypA�'�ݟM`tᰐ�9��?��Q�%�<�2�I�q+z���U�3�����T9"�QSh��d�l�� �8#�D�\c��=�dGS�V����a� 'Bn2��4'���I����4�?Q���i�9`�m�$�U�Y!U��_?����>�B�M�`�lyQfE؏B�H��)Df�'o6��Ov�?�n�v@H�]>Q�xXX2`�R�
��,O�(�&��¦���I%����vƟ�5�&���@�:_ڌss���YD�aPi�;Rj���PC��Ҷ�3G84@��?:B�8�6c��1'�N�|�� ��~_����FB��0�!�`!�� dFѻ#�?{b���'�����'\�6-V.��Y���If}r'�"� �Y�cĤ�<ܹ�C� �p>�H<ig �3Xظ*0bʇ �|�p�Țv��6��ۦ�$�`�O\�'4�Ɓ�t |  �   W   Ĵ���	��Z�JvI�*�� 3��H��R�
O�ظ2�>���& �ث�O�=�p@O�rh���EL�G��-`1��Ѧ��ߴ�?1��'\ʓ���iӞ�I�6��I���F�p��Ŏ�b��9��1���	:�ɺ1H�l[ǹi���نU��}���	\Q�(O�r3Jˌ_�&l0�\�l;Ю�;,�Y��¶>y%���S��p�J�:o B�2Qlɾۈ8�u��a���`�\�D"y!�xs�K�<!/K�ϲH%,�o��Sc�_��l���kuӴ�'S�$bW�1p���'I�Y��Ɋ+�Nq�;+ӄh�����;�|+���#���$��(w�=�'�Z|�A�K<{�8�
Q��>M�'��8Dx�l�h�'`��A�<�&9���T$F�/�{��"<�f��>��I�u��P�-[74�����\�$D6�O*�0�{R���fLC PD��g ��M�Ԍ?|�d"<Q�o��	�$�����l�Pyv':e&��>1�a1�D��n�,�g��K�N�BV��8p��'�.]Dx��Z�-X��eޯ7�D-:u�[�c�nY+�a:��#<A�B�O�%�L�@TA�F�i��i ��䒋�O6]�N<���Լ6�`1��)�l� 	�J?iC�,�Im��<1���L[����?vT���)R@��F}��?�	�`2`��1�p=z'h	P,�t��S4P(��)GX�@�L�p�O~4��Bٗgщ'��E�׋P�I�*Q���d� Y�OTL�O<����{��UcK>��,��=��O"J�K��A�8��PB-D����(   �Z,���'����4!�:D��ڰ
�';��[	�'T0��;&����2�	�"/��	�'�����+Ne���������'�.58�&0�2싥�U�;i֌P�'t�#P��2q�9���)7�����'�5����8hd���sҞ2-��Z�'���y���NN\�
@Μ�0!�e��'XVI�f蓀2W���t3����'�vA���	*?�-Su����|M�	�'8�5SŤN�*�r��GJ� :����	�'~D]�7�źxajQ G���*��l��']<	+��R�H)��[�,3��;�'�T�����<d��{�#��zf�c�'Uje�̛���`�ūQ�z/<��'�Qy檉�,R�%�
@�$[��'.�	#�@@5	;�I�&D�"�Q��'��epF�B�?u���խ $��c�'��eᔂNP   u
  �  m  �  �(  1  V7  �=  �C  1J  �Q  *X  �^  �d  k  Iq  �w  �}  Ǆ   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dlӂ(p2O�=�!�'�AbE j�80�eˆ["����.�4&N���ρE��J�l��d	�V���u��H�y��_�S �DB��a�,y3fV#2ԐGL��>�P��FT0Ji<��̉�]��E-�H�.��~�&����@뵢Q%4� }
���q�@h�`a�_�e�����?���[�t鈀�c�	p-���F�iW��'
b�'��E[?Z2��"�a�v����'�7H�S#���?�e�D�����?��-�G��ɣ5ˇ�t�l��8�?����?a������O�0	�iy2�	៸CQ$Ț���c>Je���EzR�	ڦ�Ya�*[�@�!�XH�8D��g����o�H�G��.��	f�,�	?`��0ԋ�kn��?;B�'�2�'Tb�'oB�'w�μ�]X��XTɌ$J�H�!@Wӟ��ݴ5��&�s�$�lǟ��I��M��bt���'�u�kǅk4Za�tȄ7�R]*Q�	�C��?]���8�^�#�O�7���&�(*QN��C��R��l1L7-��#ݴ����,�	�bK�3Mb����/O�hp�e�ew��Ĵi/F��嫔�N�8(�!��"Q�L���V�_�z䬻�MS'�i�R7�Ɨ=D���1��r�4x	��ČZS$��ѫ�LF֦��JD7-F����L�u��g��s[wv΍3U�*P�إbJ8|p����8z,�2�M�Q+�ơo���o����}�Ls��g+�Y�o�/H'��[ ���6���T�P9�z��4��4��o�Ot*�/tP������'.�yA�l�%^2��G�
Z����U,֞t>Y��s� Tn�֟���?��U琥bj�kpW��0�T퉠r�8�0�jY�1�b%�CK�L�'���'�2��tE�9Bm�k�&h��h릭y��;5�9zu�G*]���+9O~0�N��&���c�	�H)@"��,EN�_1w ����^/1범�Óp�Q�I����'c��9��6�"l+p"ʠ/��)����?������(�>L��ǐ�tB8��l,Y�TŘ��'���� ���E�!CY���˓�I;a���S�7�>�ͻ"�� Dɩ"d����PU����p�J)s��/�bY��a�Dx\p��BW|A2�
N}S�K��c�^)�ȓc�����P����� Mx�(�ȓ�Z���.n��8� �@����a���@�$E20 Pe�@	H���	w��"<E�4,D!s����ԩa����P�0P!�d��D���bH�:�Dz��P;!�L6N�T�ơ�v�@�R�H<!�D�:Js��Cr�Pʲ4EjR�
 !�dʙ�,)���,e=�F����!�Ĝ!?����WmۖMU�0�S���
����F*#���"��EGT5�aC��b�!�D	�6�p����&&1x� �~�!�@�_+��`��K�5Eaʌ]�!��J;���QG'�5X|J����#b�!�$����y �
.lbΑZcl�5�yBD�_d�7�8?I�IԬeՈ�j�*��,�t�z!@����'Or�'�"S�U�2-��"/������Q��)'�I�-�jeX��,j:�X$�5O���v��)���ө	:	�N����,*dIQ��"YO�2hήc�ax2CH��?����?���r��`E���&�z��O�9D��+O~��*�)�'W���$B����pŊ �t�1��ɜ�?q��ϗb�ؤ83)��cd�� �-�ݟ��'7Р۰�l�䒟>�������h��6��/L"4�n�7H�v���O�0X�BO�-�&�WiW�_��y�t�O�V����]֜xS��O�6��H��O(��ƚ�mB-�E�~\Ԅ:�ᓊ�����d�P7���)6�R��n���ӟ�&?��|�!c3���ZTHJ�*��qCo�e�Iޟ0��3��-�6(=t���*,G6o7P�?�A��0r|i0 �gt������A38�mZ���'7��a��O���'+bR���B�*�1TF�3޸`qի VL�g,p���bWư����yB�Y�@iӮ� W����`�(�F�i �R�LXL6l`�������\h�	BJ�>�;RH%>?J7��Xy�!��?�����?��l��tpU���O�
0�֎��P`l��'3h	P�Z	y�$��V�Gn>d.O�Dz�O�R[�<��kŚ)�`�bs"J�� ekDKO+��$����t������I�uW�'��8����Р�y@���n�5oǞ��3hQ��!�DXOk�X���[ �fLI�\Lq)�O�H����a�y�7�B��N�P��qO���)[�PK��A�ܪ[*)�"O�=K�擌8����iβWK�	cF�|2�qӔ�O����%D�=��џ��bF,����K\�%�G�Y�p��O��2".�O`�$�O2l��C�O`��y� �q���Y,}App��c�M��P�'��=�aN.��#�(��@� �k8hz��Gh�ڸ���0<��@S��ɠ�M���h�\p��IR�6Xʰ�ɋ|!�u�+O��D5�)��O�u��gD�zȜrs+;{�p��'��7턲x�.�b���)Z�e��X�D o�dy��^���6m�O���|r���?���,HߚŪv!��qb�$:���?��bT�<�����>�:@x��R�a�7Y`2e��K{~���^�����D�Lߦ���Ӛ=׬$�4��/P�M�uM�iv��/_���ߟ|I۴�?Q��)��T����F�<��H���9b��'�R�'�ў�S(��� bEf�9²����r�?�d�ip�6�>�9Zt���f�x�c�W5�J��'�	�o�����A�'�:��Gh%j�V	!��K,�����R�$J�:�a���L�-� ��E@T����6�9�O��ao =	J�b>c���/��r�(�'۳7�V����O����O�9s�h�Oc>˓�?Id&I�n�Bؙ�o�)��5YrGI�y�l����K #�h��$#����^s�'�{yf[5s���W�5g�X���u���:��a�p���O�$�<�|��Y=x@�<���bn��$Ó�+��=���ś領`s �xT�����V��i�C�k`)���Z�XGM�@�V0�$��	4�f���	 �b�Cc,\m�`��d��_�T��H�O
�$�OR�PG���99�P=B��D�YBΩÓ�ދ�ybOݶf4�A&�V-'�f�B�	��X|��@yr�b��6�*rƬƗ{f�(���H`�a�Mɟ8�'2b�'E󉔃�l��g�+vR�r�U�^b)��G%L'��^� �ȩ�'o��R�Լ,� 89�#B�~��%B��]�����d�C-�Q�$J�4�0<�$Fğd�	��Mc�_�D�m܃2�k2�;ky�+O��d(�i>a�<�Љ�=���h2F����\��<
�4M�����w[���B8^����ic�I-VR�!ش�?�/O6�'�?�G�R% ��@"�ވ��i��?Q�Rԝ�s�I�f�z@_�!҉i���
�z}"A���B3q���*�*aB�ɑ\��t�X,c�J�8R�U�#|*B�_�AƊ�����Pİ3�aGG~�'���?���hD���'t�O
�	L�%����咴X�3o��ne�'��Iz~c�NI�%��}Wt��'�����O�pm�#�MÏ��E�@~��g��3ua�� �	�?�������Ճ0�uo	�D�\dkG�Q��!�0@��MZ�<��3�$;�!�Dlv���"�V:P��<k��O�!�DP:~0���e*sX���"��!��	@w+MmTtU��F�9q�!�$>UJt�B�c�O$�|���tY��0����DD�BN0��TK��AER�{�!�D|�ƈ ��҆zd��Hԃ�j�!���;��H�2��H�4tjc"�!���Z��N�ˠ"�

K�!�d@ҔI�Dꏡ0��u�#'��}�G��~b��x�4��T)]�3ՌX�� .�yb�Нɴ��'L�>0���啳�y�i$s�	ӆ�##�T��,�y�,B&P>�J3#h���4,�*�y˛6AR�P�mD��Y���y��*(����WS�Α����6�hO��K@�Ӗ�p��#��(y��y*��l�~B�$K\`HJ� T/f3$԰��ں[�lB�I5 ��p�J����THw"�
O%HB䉯���I�m�̬!7�q�B�	� �s��*���Q �ͳj�2C�	�J���"�A�;̨ S)Ao̴��Д=��"~�S��7���ӌR(D�tqg*��y��ԉ-�j`��: q�`*�
F��y��ފ8u����$:y���j����y�Q\��q-�G�lys�g$�y� �=�V����'\j�"Ն�3�y�$��$Bd���π��0�bTf���$��|�|B*Ψ`:��F�\
�PM2�ʌ3�y
� j ش��
&��A=O��3"O"l���K12f����E���k��,D� @�AA�e�ƴ�w@��q���d0D�����2<�� #
�^�@�S�-�O�5��O�Ha���40��Y`Ù�o�$�	r"OtH	Q�߁��H9�������"O��̭.��l�� �h Ճv"O�0� �3Vf�#��Z D�Lc�"O�!�C�0s�X{�J����"OL��ƭO�C�j��sϏcP�y���I�l�V�~
�$C�Oۘ1����A^�}rT�KP�<A��в���p�PhE�aB���Q�<� �Gr�hj���*��L���Ed�<y�kռR4�u��Ȓ'!�U��!d�<	�)�*Nr�H��[�:���QF��i�<c
N�1��rcїhX�9wLU�x ��4�S�OἍ�7��1nk�M#pe�r=
���"O��*��K�O�x����-i=BRc"Of1!$N����lr��ח^��� �"O��s(�!��Q���0�Z� "O����%��-�@�T܌M��"OP ��OS�OX��P��?��-1_���a�*�Of�P�ѤY�(��ց��!��0��"O��r��:2-nmJF��B/LtBr"Oҍ��^�O�J�4eҜ�a%"O̸���,X���!j9^ȴxB"Ov ��ʃ�l|���0�L�S�ؽf�'$&@��'４��	ɠA.�u8a	�f^I��'�,Ѵ�ȿ\t�-�p
Q`��b�'8y��@�=c|1��[�\�U�	�'Ƚ��ş�jd|#�M�WR �S�'�L�b�H�D���RV��"OzVY�
�'C�1B��%��nL�x���d/�Q?�XPE�s�r���O��q�Z��F�*D�hA����j�w��3��U8L5D�0xub� )|�8�
�H����+3D�X��_��B���㇠Ij�囧!3D�@JCɿ|=
l�G�E�s��|�׊0D� 9�G��v�"�}��X	�n�O��b��)�'U#<����E�|��]�p,c�J���'�P�#���nmڴJCn��k��,��'�2i��W�&�,Z5�k;�E��'�b)��F�V v0P���]j����'q�|0��[�$���A�B�M"h#�'�2I���^�$�!wH�
M�,O�(iW�'N�妜7�N�C��(S��h�'���櫓�"tk��X�DK�yX�'�T��R�CS����",��=!2Q*�'W<U&LX\�@"�H13�x� �';�a�!��o�ĥ���
�_�h!� �H���' qP�Ҹ6�p�0��L�h��i�ԍ��qFƽzvm�ZD����J�e	��)�u�0�
�Y�ȓH(	�1��:4xrPz"\�7Tȥ�ȓyL���s�����2D�' �����'j9CK�+eD��� B���E{�+6娟�l�0b�2e�lX���֥e����"O�Y�e�ǘ�&,
�C9oY�P"O�<�6��<�
bb>9T��zg"Ol�G��f>�D�/W��4c5"O8yNF�,̀qx �� Fdz�"OZ$0*W�9n���*�r�:��'^�8a���S�:�ę�L@ [�h��a�I;%�ȓ#l�=CcA�a�ʄ�A�n5��S�? �B�Ā��0y`�G�F�"!3"O P 6�̆Vɴ�!#g��+�� �"OLDs�j�G�lr�F��yȾ�F"O�:�o�<����p�S� !�):�Y�@��<�OpT�0�V�B����т7-�e҄"OV%�adR��F��`�÷E\��"O��+`2gJuڷe�k�tÆ"O��Q6;Z�̠s�L�h��"O$t;�+ԶI�ڬ��鈃:�v�$��>YC,�i?�Ҡau�%��'N�G�"@j��Er�<��̕\]��1ĊȰi��� �e�p�<�!��	�6�a��/����@�t�<a��i�L} ���0�,$Av�Yr�<�1D�x7��0�i����0*5dVn�<��ƥES*�{D@
/o���9��l�'O��Z��iW=A2�QЄ�
��%���[O!�$G�a.m�d�3��a�&�N4H!�$
� b)[�'��qM�5�bîAD!�W�6ں4�H[�m7T0�G\�!��0g&�ԨT)�}���P#'��g�!��q~���E�S�U�gDu�(@��O?��Р��4{�a9��*�D�a4�~�<�ՆH�d���"m[%U���8G�|�<���86�]aE��&�����g�u�<c�e����b/��\$B���n�<)�A�����қ}�
��jCb�<1�H^� ��	)D
���= ���_y�Kϖ�p>١��~@��Ŕ�c�ѷeG�<�r�R>]����@��#D�<y@&�
tL�}������aZd��<��
~�~=H�)׌��N~�<	d�Rd�)�EB�g�
-s2ȊEx�Ј�'��\P3@S�H�x%�OKZX�'�?D���C���"�����Q30	��*D�h�`��\�hM5�6!��Q��)D�,i�-��F3b���A8×+&D���(=,jhH�Em\l����$D���vȓ%Jx,LݓCbX!�D�=��!^�Oyp'9c
~$�fۢI����'L�c���Ih`��G���'�d�����
�X����0���'�(�����"m�Rea��4x�X���'Ǆ�Z�BN�`��UK4�� jTF���'	��P��W) R@��� ?ײa:��j�hFx��I�,X�@�'���`�.mY��HP�B�I�c�H��b,X#7 ���
خ1�B�Is(z��4ǋ����ivΔ./ְB�ɖ"���cG�ܢoT	�сE�
ǶB�5'jp,�$��t�JU�@��(w�B䉀A��)j4�	*_L(]��A>zz�YW�̆�I*'�Ƒj�G�<7H&���xs8C䉴��8b�6m�F��n�\C�	� �̘�T��*+@ #.���B�	��]��BY��B��{�C䉄X�� Gٷ��pLD�������}G��).&@��!	�3�d)�1w!�D
�Kd����hK*'�	J��� �!�6V���q#g6x35g��Z!��,��D((	��;T���>!�GPX�X�e�;]�,����"P'!��2(&�xڴv~@D��lۍ8xўR@�5�r
�yg���i6H�$�.ad\%�ȓ9)�$�BÎD4p���N*gǚY�ȓQ�$��ҋ;F<���EO���S�? ��G�:����GILTv�E"O�|�*��96^-X��LW���s"O��#�*5t&��$&7�>!J�'�\����
ڕ a���lp`d@T�1�m����9��Ky��P�`0'䶤�ȓP
�Pc�٢$>����&nq� ��;�ܬ�*˹@�~��g@�,��m��3d[���"`�\#Tn��)i���H�V�6/�N��{s��9f�H8�'��4�B~	J��U���|KW
5W؍������ך9T�a���_p\�ȓ|np�f�X1&���3y�2}�ȓdȫ���Yl��2�(a�x���\����Ҩ} �=���
B��Ą�ɯ=NX��$wP�pB�	t�D�S H:P+ B�	#֒�+�E��c�p�cA
�o��C��<%� -�u��x��³C1�C�ɣw�X��5�")[֝2�.�1m��C�	�>�zHj�I5�\��-[TlC�I8Ca|9rF�2��u���o:�=�!�g�O4. K���xј�Jc�רn˔���'��|J��c �2��h����'��pqk��r� A	q�«]h�Ų�'F
�S���_Ș�� �ND"��	�'�s�G�ⶠ���Ѩ\T���	�'K��P�Cr>�;4�D�����u:��Fx����AFfL���1;�p�$p:�C�	Z�d�햨>��[�b¥VGfC�	�+8:L����qz�ۢ��v�C��4�;F�ˊ�Vh�%�%9C�I�K�1UF��XF�� ´`,�B�	;g�b���d���*��$jK��?��ӳ���O���*U�F�B�H�b��u�%V��d��f�$�O��ھb�Ԁ�ª����f��4�F�ہ(OXB`�#�!����ɼAO�YX��5l슝@��Y��O��\�0��g(܃Tv����=��O�����'���)�L��-��z�^�X�$�� ��G���㢎E-xC��Z���&RF�!S�4�O:�'BD8��^PM��2��\W@Zd�.O��9%�O^���O��'C"����?9�̛<��d#
�A��4B��?IcK�uY~pXsbۂ{"��[c�i�'��O'�H�%˃��W�"sd����<��I��1E߸OL
t��V�nr��ݾ&�R\$>(��pڰ"�ə"t�H��b�g�\2 ��O���2?%?��'������`&j��țs�����'� ��KƓI�� B+�i2�<H���^^�OS0m ҠȮ�Tau��Q2ʁ�'Z��'�f5�qO��HR�'���'W���'�%(e�:��@�VN�ZR��S�UfX�7M�����S�G:C>���'|V��t�$77��QDΧwZ�1��H7x�^�c����A/��*ȋ����*�M����X8*X�
��_P��6�F�E��Ʌ,��$�O �=��'��4y0���4	vT2�⅂6� ) �'�N,96(Q+
c��\����|����՟�'��5�L�	SC�<j����+҆\�E3��'Nr�'���O��'W�)�5�*$1D�U!���C��)�R���͒xX�EP���*06�s�'?H�QꏊK	X@��P�ٶI9fN�=`����5 ������kۍR��nZ���0�>	� ����Pg,h<��)%���Yx,<�2���E{"�	�-A&i�Kę@���r�[;RC�ɶRM���w��܂�+X&A�ʓ웖�'��Ij�
�h���db>y�6
ڛ�9aa4UX�2PK�O���F��O|���O�5��D�\$0�`�eK,cyD8�i>	iHB�)������	0F�xȁթ>����I�#ܭqn�n����	�7bD<�{e,�;�vi���_����F��O���=擱?k�1M��BN��ɕ��H��˓�?���&��W�"e�jębG�E���+��$Q�Yv�`#��T�)3�m�'��	DC2H�I	Ra�M��R�D�#����'�|�E	�x���ȡIU9�Px���'d0l+d양��c�*�<93n6�BK���	M2[0�ҳ���R��i��ߪt�Y0"��+��b�8��A�i�	sXw�J감��m�t�����a
6�b�ЪȻ�yr
X-�?������4��� ( Q$�%�)��5S�R�#"O����TY
��uğ�yju)F��:�ȟ཰U*F�!E�K>S�Gg�$ZR��3�Q��3�
$$����#�6J���'��EȎ�gR���I�&\���ȓA�D��/�f�`��$W����_kb䰴d�jʜ�v� [~�)�� �Y�&Y�<�8L�0�UR������*%a	ѓ���1z�K�57ź�q�D�8a����l�Iޟ��[w���'��C&)�.�{����u<��"�`N�1�"Ŝ69Ti%%����VV����	;����/xyj灏�d.Ya�@�*+4���'c(Y
��X)��"mT0C����CIJYS��?q�����hq#���8��N�$.�0 �ȓ[". ���<���m_�B����'�*7��OZ˓ /z�:v�i���'t�)*9r�"��xi��EV�e"%
B�2�'DR��16��4��x���ZU���䮈7%�2w�x�Z#~2$W�JR�◯T3�	:U��\�'�,������^�u��;�]X7�ڊE�8t �"Orq��	2:��@W(�pjr1T�'���p��Is"eB/�����w��`�'_��'^ɧ��)?awУ)���:�JP�&)�"͙[�HE{b��S8� �G�?����-֯��'��J<a���Jҍ}�깨!����9g��2��di?qw�UM�T>�V���s �@!9ޢI���	3Y&��A~23} ���I���'/	e[+�+'V���6��07;f\Ӓ�.}rM��dG��'��B7&�,��M�` *���QM@��􉝌�I�wJN�'���'���k0mA�q<��Tȩ<���I?���'~B���)�-�<y;p!m�Q*]&0"9둈�O2Y3��>1�>a�ΏV�D��5;�էEqF��f읗hö�C-�<IZN���g�O������0�2w � U�ع�H�� ��	(}*��܂D�	W9>��Ex)����B�B���ay�l���'���q�'�1�z0[�����J���|\�y
��'�����^�����9O�l��O�́�������"%� �*	ʀ�',D݆�I�BV�@��Wt�Bcwᔜ:&B�I�M6rSc�~Ʃ�a8b�X6��O4�O�������|n��HK��F]�Y��c�Ȏ�A�nꓟ?�*O�=�O�2; �O�+��@�bֲ-� (�H<a����S$��1�̋u��uŃA��!���$��5����;q}n KR�3�!�!��� `�Y>`m򍳶� B�!�*T8F��G-�6.����w��83!���P������)����ȍ+C$!�d�Q�f<��$�:����ȕC?!�ΌQtfٓ���x��I8��̢7=!�Ũ�t�č���S��AF�!�ı�PyW�� j�̅:���Z�!�dea����o������!a<!�D��Uը)�G/A \�(�m�"[;!�v�j� �5�`�bBO��f1�Od��-ug���cC�LM��%K8Jɪ���*$7�����V�*�V���5s�� �M� �T�H��G;p
��:�Do($��[���bd�	xda0@�]����wd��D����V! k�y��I��uS+�ES,���c�׻r�]��Ϯ/d�1�RM:$z`('�i���Q3�ǝl4�d�E�@sO�}X�O���h����9�|�'�Э�R펪3X�# 0cQ2�PN<	w�JY���O,��Rf��87	*X��ƕW�*O<)��̟��<�~����k�>�(��W�x�|��s�<�QN@(vݴT�Q�-Nϸ�;��i8��(��d�*MȨ�A"%|\���[�E��d=�Oȭ �E���@d�"~l<�*�"O\�I�����S����0k�H"Oİ��"S\�J���7,BNl�&"O�%�D��,e��P��"9���F"OP��S�A/z��Y�e�:H&@�Z""Oޝ3taL-F�Q���ˊW���8�"O���.V)79� �B�E1)�L��"O� �����'tzIڄ��&�H%�"OR8�d/�e�����,�.F�\|�Q"O���e+�rpB�����	��"OŪU���y�>,�GIٯp�Bqc�"O)����1��z�e�;_�*�	W"O�H�[�E�@�YVeR��5�7"O�8�҈N��Ԙ����_���	�"O愈%!��	APd-��	JT"O>����'��h$�� k�L��"O�}�7�U)�T0E�/�X�d"O��	�흈5Y�3V"��S����"OJ��d\P�	Z�J	sDD�yR�]
)������n�KE�B��y�j�+v��h�K:gD������y�*��/���5�a�j��%�U+�yR�'��+E�Ȧ� ��@wo!�$�!:��1pmG�z�DM�p�ױ,f!��U5jJ2���%��d�����w!��[�b����B�#l���Ӳ�WB!�d��ec�!S,W ]�!��'#��k�(GY���!L��X��\��'�j� ��6cP�F�۾�@�'YF�2A�/Dڥ�u旿rȣ�'t����9L�J�A�*\�_R)��'��u0�o]���AcB�Iz�1�'�V�p�-�' Z�}�d�����!�'�	���D�h<���)�F�
�'~�#af�*h�3�W.dƘ�
�'w�uR�L�X���R�:0��'O<��N�+�ڽ��ʫB6T`�'�"H�햸p/��AУ�<�.���'LBqK/a7T�e��:KX��'儉0d�8S�5!Gm�%B%y�'��Q���~R�Xc��ZE�'\��������QD)�zM��'�.��D�	g�����"�Ti�'Gd͉���oK�Y�sL�/� `��'�PL�B�: ���S��̩m�u��'��-�qK�5E6��a�+o&�5��'�=p�hX�(�Z܁�Õo��I
�'���sbX�x��� �n�\Q�	�'�|9@�+͑//�M�BGZQ���'���`t'߰e2c�9O͆!3�'��)y���2v`z�avA�Gu�� �'��(��#=D��x9���A�@
�'�]�Q	_�Q��,�Q�Z�

�'�����@V����*��xD(�'����O:8RR/߮w0��'d ���ϩ �e�qaP8%��
�'F�#���l\�сJ($��a��'���VC�:g���@��p���'�f���G�[�0U ���g� h
�'nU�@�5&�{��=e�S
�'[� �뛼V��]Am�,%�H�	�'d�[ЄĤo�ޭS��_/L�NI	�'_�p�_�p
� Wi�G/���'�ҐJc�� rH�k�EBm�Q��'�(��g�^�ndh#4��R~���'�ąjWѺN+^�[�Bz���1�'�\�1�LQ�1���M�m��Hz�'��p�VG�>���kBu���)�'�ڹ�1�o��}U-�"<��ŋ�'ۖ��֡�3n`5�٩;簉I�'2���� XXVB�'谜�)-D�� 0��lB�&{@I�13#����"OdA�Ā�5�Π*��]�1&��"O�j�$S�����r��C@"O")�'�U��T���k^`x��"O��RQ�?	o����W�n�R�"O�y@�̍�rwn�y�&�mݺ���"Ov��ơӡJ�͐r��I���s7"O� @Q��K�P�T�#-���	�"O*(c��AM�,��a�.0����#"O�4Qc�d-�@����k��q�v"O� �&d\0G{H���~��""O���E�f��Bs�N�q^<�"Oz��]!.��P E�#*��P�"O�qw ��g��0��/7kBl!��"O`��P��*��T�3/���"O��BZ A��чFQ�C�	ʦ"O�Ea���$%P�}8 +'	&4��"O`�����:$3�Ģ0*Ǟ/��H��"O��Cf�a|��!+ Q�(�S"O��S��̋P�lm1īH�  ���"O����g� �|�J��H�t�~�!�"O�l�i�y&�����U����"O՘�՝�^�9�T�H�����"O�m�F)H�e�4�wjP���,ʱ"O$�H��k�6h2Q*����"O �ku�4�b�#t'�t���"O�h��,0��1��ϝ�@�r*O��	� 6MDX�oǷ��A��'|<����jn�|I7D�$�l���'@-;�b�:.@}�
���
�'���80�X22Դi V�T4(U�A	�'T8A��Ú�r8h�MK%�`���'�D��D
���Pj��8�{
�'���H##h4A���	�i�	�'d1	bI�&^�P�Dn��v�@��'���ac�M'�Q���J��'�쫒�Y#Q>�l���I2
��:�'��M�§d��Z��6vyTm8�'l���d �*^�U��H�@y<��'x$�Ck	�x8��ܖ/=�͊�'��0ŧ�(y$t�eF�0m<� 	�'	>`��ba��1+gBE&
����' �{�iE�UC6�1)H�a�=��']HZ��Y�~,����\� �
�'Z��XeV(�~(���[��ԩ�'nV��c�B�t��r#VoB��'�����Z4Gؠ��f��~vP�
�' � K�l+轚&�ތ��Y�'YN1��=Q(Ic�J ��!�'���j���[����cڙ�[�'��89��wl�%�1Q�D�Y
�'Q�m0 ݀`����d#�J��X��'X�SP�Tq�*�0d�Tx"=�'���RE�5ؖ�Pcg�$����'�d�1 B�3�<�����V�:�C�'�l킳)�!vT�X��@�F[� ;�'ld��7�HN>ʤ�ဋ/E�J5�
�'�Z|{b�W*q�t(�AI�18�f��
�'�m��bز
I���E���w��0
�'��aC��T�?�����K�,rr��'O�PI!ώ<]�f=k���P���'�:����(o%$0��G��J��y"N.7��y0GĊJ_�*�!��y�ѷ�ʱ�F I�ڔ��^�y
� ���t��tꪍ�Ǫ�e�ڭC�"O$\b��΄2��is�'OY:�Qg"O2�ATC�H��E)WC``�"O�P��cGAa8x�Y&c�*��e"O[%KQ77���8�Q*$r�тR"O�5ӧ��6���
Ѕ_�0<<R"Op�0@��Y�v$��D�;%2�"O>�Y2"#a�Dr��>���@"O�IⲌ4q*�1��Ĥ"fY�"Or1k"�\��I��%S�\���"O�d���H� ~i֤�3�y�"O��s���`�P��X���C�"OԸ	��M�5�z������A��<��"O:I�oI��@��`W�E�V�"O��g�V��X�O�brB�1f"O@� �X�G�РPL�-��xq�"OX)S��EO�����$��9� "O��#C`�cdN,0��7�z�2"O,8;� Y&~l�,�傶�����"Of�R���bZ�D�2ą�=p�	��"OʹS���Bά�#L�S�Vd��"O\��������b��"jhX9I@"O��ӇB8c���[�db�s"O$T�"e	9Gvٔl&h# �(c"O�u��k\F記#��ID��@"O�4ȧܗv����ߠt����1"O���#��-�­2���5�����"O�����A��q�	�:��L �"OZ�s��-&Z���p�#;z�� �"On}��M�`���I�#$l�}�a"O��lD�w՚�[!#N�/1�剀"O��1" �x���@耥Z&�Qs�"O��3s ��7ܡ��f�+ ����"O��Af�5������N��	��"O�P�m�/j�ؘh� 0C?�i�"O��8���^�z @��;0�UG"O�<kè��K�0�"kZ U>���r"O4��e�)V��JF�8�X�"O��R
���M�$�OW���K�"O��Яހ}�$M�U.��Gu����"ON�,tx��@��uآ��0ZF!��tw )��lD�)#N0*��K-!��@q�9& �)3*��bR� i!�؞q����] �9�	�p�!�%[d���,
� y�S-s!���?��+BW$d�&�C��)!��,>>�S�HX���(]���e"O� B�C~Tav.:)t�٩t"O�5��2��(RpN�f���6"Oh�8���)>��a���<N@Ѓ�"O:u�5��U�"�����7tY��"Otx#� ���@-C��i�4}��"O�4���O��B����	�z���"O�]�W ��x��9z¡�d� (��"O((p�@�.�Ԉ N0t��H�"O�PUa��F
�0j�n��>U�"OИ�$N�$9e����͍���"�"OF��V�.��r'�>z�x�"Ou����02�(g�ٖwWv��P"OT`�!x��	�q���+vH��"O����	=	",��?qʭ0"O���堞�QQ�t
�C��UZ���"OJ�8��pnڵ�ϖ?�X�T�ܚ#!��
u�^�}�|l8�#<O�)� ���I��W�bg�i �"O� ��֤\�2�J a�� =^��0�"O0`��["ȁ�� Р=�-��"O���g$��-���ֆX ��yk�"O<DI��^1F�^`I��Mf�L���"O��+ݾRS�����>��m9w"Op�Eiлb�0�A0�H�
�"O�SSe�o\P�!��4IRP�Yu"O��4�_>8��X
v(ֽ-&�t�"OL4��U����Sҭ��z�"O����A-�@��+q�ir�"ON�A1�Q�H�4��l��x~�`�t"OZ,�"Ô 5��D�T�Ǌ�8B�"O2��U�]�6tAiC���h�@"Oh!��
$�a�Pϊ1�0��""O �T�l�iCF���_�B�1"Oܙt�x��!�Ȫ�����"O��cp'���#��8H4�!"OFH� �-`��#��|�(��"O�����_68�,�!%U!Kr���"O� `�G�Gux��DDgN@ۣ"O��q�F :��3�B!n���"OmZd*�F����ӧȪ)]��c�"O����-H��{2�݇*��C"O��I@��M��9�����/��к1"O����-C�S����6�;LV�PЦ"O���m��R�$�k��B�p)�"O
�IFl�2|�u1�I!�(u+T"O�i�T,���$�_��M �"Op����g�<"B9<z���"OT��� �B�rd�"MUx=/�yR��"��J��V�*0X"F�*�yB��Ҍq���$q���� �y�<>� �$o"l���� @�y"���{˰�+��$n�sG�Q��yr�@=x���F'�
T��-�7J���yBo�Z�m�WOu�����[��y�C?q}=����Bi˓���y�MA"A���.~6 S�8�ybKL ,(��*C���I�XQ�(��y�C��&��msQ��{|�l���A�y�:>tTl�%��m|���0N_��y��T;}�x�v��N\� ����yr�ۅ8�p�g�L�\�S�� ��yR�ڬcʜ��.�<�ޑ�-D��y҅X�MD�꒘$�ΉB!����yb�D5=��q�dP.W�5A�
͂�y2bRD%��s�L�9���V�ջ�y���9P�콐e���7�l�a�D8�y��Ha&N�����;)5|���E8�yB��9�d�ãT0(��y֯�8�y���Cd�)��I�R�jfN]�ybCƽ���)��H�l|h����yr)���(���@���1���Pyb�ʒUG�]���|
�}�B)�L�<Q��\�r͞Ib�>s����`_�<����	;s�5q�*J:���[-�E�<A��<r��B�c��&�܋�K^�<��!�6B%<��$jyv<M��i�o�<��L�$Tv�)'��n���h��v�<���]�N���@�
� >�04�0��V�<�6㖯/�BP�gK�\�9�1�o�<�6�S5��,؄�=sZJ� l�<���:j�2E aIL9T�����%�n�<9%Ζ=�4R��K�uk�5�p�]m�<� Ȭ���P�W�n=yq�؃E����"Ol$��P�!M���6������"O��(OS�6%@�I�T��=s"Oz���C��=�F��t (���E"O������Z�~�"���g�"�� "O��X�I��7^�p�R	Δ5q�Xj�"Oh� 7+��VB���E��,ft��v"Oz�EA;3Jm�F�D�,S���"O��0�P�b,�Q���L�H�"O.��'ʏ���C'`f&��b"O
)��ʑ�T�Ve��'2t)�"Oj����  c�����
�9Iޜ��"O�1��N '�K�A�Vm��"O*lc��$K���x��$E)n`�"O7MN:��!l��8k�lR5�:D�t3��P)�Dh�mL�8Y���,,D�Hk��)^B }c$��&kņ���/-D�A���=�Ε;��G�b�t���*D�4#kU�l�EXwaǿ3,��B�D.D��d�.-���{g�	jy����
:D���C�wZU2ч>NH>m{e�'D����#U�n��!J�ɛ�ʔ��B"D��S �R9t�2c��;� [�j4D����-l�4��,~�V��R�.D��C�fM(Y���
"�H50�[�)D���G�tE`�Rf#�[��;�5D��K�h�!i��#��5!�
��3D��pB��M�a��.ʚ ��U��#0D��z�dǤL�p���������?D���g��H��bn����2�,#D����/�� I��a���� 2?D��� Mŋ�F�r���]�����;D����M�1o�\,� P�xQq7#%D�����N�>RY���_���U�K0D���hՂup
d*V���iP~�ce�<D����B�UD �W��J�ZT�UB:D��sL��R�����t!"%9D��QM�'��]a�n�u�L��� -D�d�@L�|�F���@nq��+D���3�fNZxr��4 IK֩;D� 8qƜ	P켤��gS�M������>a�-/���H��ͺp�fNv��5�H�u[��0�"O�a�"��^B-�W��:F�$б���Xv�޵5� ��I"G X�{�/
�J��0Y��ʴx����d�)q��K� �P����'�&A�	w��/�f�!h(�PK�e�:.��8+A+�o�^��1� ���6`7Ӝ����Dc��s5RY[���L	�	�d`X��y��c���t�P;GQ� �g��8A!(�;"���q ?6��9O��s�&��h�{��˃4�(�"OT��E�ӻ
��\�6NV  P`��F�O8���ۅ(cd ��!�T�?�  � :�VMj�fE�i~�Q�q��{��d��^'꽑$(� +t�R�Œ!���(%V�T[�U�Jea�g��`�h�p��!�<Z�`����'�z�dߢAR���
܃��'>�PA
:�P�b���Xpè8D����Fy�(��hC6��đL�DQ�#蝂_���2l���G��O���ac��?Q�x��L�uH�r"O����<Et�8�T+x�Լ���
M.�Q@��s�@���E�+p�2�\*E����u�N�����	c�����)Tr3�h�5w9T��b�@��Q�0��,|-�;�OI�+���pfu��TҲ�X8e�xѲ�=4�,��=�I�@�x{SAۮ"a�(�A�^�?t�%���gRd�d�Y�n�8MK�'L��!�A�v2�7��E?����Rub�k�)�1<�J�[�KK;?�.�S'�Z?�w��q��\sR�e6lɢ���t�<!�W�,���S��X�$
��xU�-Nx��'GJ$Sdo׋z�n��)� t,�g��&3J
 ȕ�����]c�'�l�Zdǎ&D�R�yEV�)/m��noh@� U���?�jڔEVV�S�dX5�@AO�B�'!�L[`m�̆T�L~���^����Eϲ'��}�%%�w�<�c��-z�Ģ�G�Q&N�0���<Ѧo]J�p�aꔑ����9&.R������ �Pp��$�<@	�B�I�6�Z����]�.� 4`Q�$0��$݊ jĪ�;���Fg@�q)cm�>qDI��	�}��+I�`�s�?Js8y�@��4.�,{t�@ o| ���'4Z�H�oԎ$��#�O � ً��E�txF�J����:N��}kA��,aja��C�;h!���S�&\c��̣tj��J� τh��	^���?E�$":Fu����%�v�>Yr3`E��yR�׀*���&m�$��ō�y���Y�ޑ�1$�Xh���<�y"�27ͨ��Gl�
W�$	 䒶�y�:��XЀN�q$��y���4G4�t���V
.�BH�&��y҄�# �lqi� E�J��W�Z1�yreʀi��5��־3`T��%U��yB�Q8D[29��Ezr�x�����y¨Ж"; � �Z��W �%�ybjB���de�-H�A����y�덨J���!@��4��525�+�y���)	�.d��C�^�ڀ%J�-�y�bѯ;����ƪ��h��A�Z%�y��H�4I�EH�f� w���H^��yg�1h�H+���A4<����yBcB	�*񠱅K�x����'�.�y��2>�����-Hr��1�)���y�#L6v�ͩo*|�y��@ �yr�C&���B�+M�"Ѽ�4]��y"�M68c�M��`G�
w���&��yJ�*@qP1�����a��K
�y�
'uR���f+D�6�niꁏ� �y�'�18�r �&)�r��юD��y�\���m�t��^z�D�5�yBM�8zY�e[�\Bp���y"��j't���];vE����y�
�o���ѐ	������1�ycI�90�`����1�:�D��?�y��Ėp�衈��#H�J�+�y�E�+���"k
qS���ҏ#�y2�G�U*zAY�D��dg��⎅��yBOͩO�����iV�\�����y�i�3Ͷ��v�ީL�N�@�V��y��/e���2�'J4g��3�D�8�y�� ����1<V<�T�yb�� ^�(H��|>U��Ά�y���m�ڔ*&u�� �	9�y2/�q*D�`J�A���S�׭�yB��k���
AΈ' �s�F��yB�6L4Z�
�vT�]��E�'�y��:
mP�r��#T�U�'��y�gVA{T�{�� _����rh�"�yDǹ ����`�L��ec��"�y2�W�T2����@[0D ��С[��y�Ԕ�,�DL,)���0�l�yr�� K4`���$�ʥ���^�y�%\�PNV�RC��Y��XS ��"�yB�Ʀ�0vĂ�W�D�h�Ȏ��yZd�Q*�b����1Ȋ
~��T��''���g��8H�8�פ#1|T��'&�0�㌖�B�8ғÞ�_J������ Nu���_qH��eԽ@���E"Ot��@��-��E�tE�(r���[V"O��+�^�Z��ͦC����`H!)�r(�w���{�Zl;�6<O�q��
�8?J��z�i͋U$`h��"O��)`��;���?%���w"O���DK��ξ4��&�a����"OD%��b��ڂ�CkF�U�$h "O�#'�I�&�9�.Yvxf"Ox��猞�_߶TYЎ��x@nE0s"O���޹��x�r���x9F���"O�A�Kh|�&ʍ;iJ�1:�"O�����s�h��"'E*z"4��'"O�T�Cѹ/�4YQ���2 �xq�"O����8P��h�Ş3��ى�"O`����� V�֠���]1Zi|��@"O�)1�E7FG�=!0#�{GnȊR"O���ӯ�JĦ�K�!��Dt��S"O�ajs�ج$��y�A�Ѡ	rҀ"O���g2����V��=��"O��6@X;�	k������"Oa�S&@8m�`4d.r
��h"Odx�'�ˇD`�T8&N-1�P���"O*�� \4L(�2�͝�b�6�[@"OP5x5cK[m`<!u.K�צ�(G"O���M�.s0N��!CϨ�����"OzPp���!uH`S㒽U�hd��"O�HS� .u2�vA:|̋""O.Mr@E��N ��-�yx��kC"O:p��
�b	mK�iz"O��b��7t,BD*<�>��"OX�h��r��X�R���kU"O> ��k�"@�ë��r	�A�"O\�MV�@R����'g��q�"O���u�-(��b��A���z�"O�� ��#�ܙb��üt���w"O�٢�' /V��fh�0= �Ya"O:Lw('H�d�m�J��� �"O�%��0rJ��b�N4�2��`"O����D#{��9�ȋ><�h���"O*���fq��y��!-�=��"O~���Ά�m��i��õ��!��"ObUKp`�vF�!fi�5i��t5"O"�����$y@\��U	W�.Ұ��c"Op<��`��s�8�c6o\/��� �"O��q��98����g�!�^�c#O$D�|�F�H�t�J��q��d�@�9�-!D���IH�1rP�vl�>-�BC$D�`��g�5:Q��U��%l0���&�&D� �G��.8gP��!ܯg�Ɣa�!*D�D{��$�t0R��5DU�L� �;D�����8 ˤ��1b�TQ��2=D��j���=U�[AD��ŋM�3�!�$�;P����,$|��,a!�D��̀P#]� �q˷g� uf!�1���{��j�xr��N!��32.����l��U
��]�Y6!��05��H��F�c�b�ꃋ�0!�$A�\�L���	��]��J�W!��]"�P��O�&w�E�q��=rb!�DN�B����,\*�R$h͔sG!򄁝"{��I�`�j����p�ε)!�$<`V�
a�U�P�D�5�4s!��X��"�&���p��$	!� g�8��"Ԋ4�PIREMf!�� ��@��*�"T@�Hܥ@`���"O�%�e-F�Gբ8����f���pv"O"(�ټ.*i#�T�b�L%�d"O�iY�f«@���"��6Y��۵"Ov�kS�W-�HC[i�e�T"OP�ৡņ	E��	� �#\�x�Q"O\Y�G��)�9{����=�L�a"O���%E�.�A�ԨB**E��"OV5�}�z��J
z>6i��"O��hX��+�k�����"O.����
7RvU����<F��`��"O@��S�
�W�J�&�U:E�})�"O.LjƂ��BPЀ�v	E�܌p�"OBxф�W�z���Q#R�8ۦ��"O���%M�Y|.e��U�b�&�"O �Q�Z*;���c�!��Kפ8�U"O�	��đ!s��5�!P+��7"O��c)&]5�i1%�5��(rs"OsD'^2Kֲ�z�����M��h5D�� �$�36y��J�f�2ў� C9D�(K�AA!LטAcƃW9r|= ��;D���Ş��434.�; ޜ�/D� �f�	�9fɓ.s�|��R�.D�h9��o<��� R�l�l3�k,D�41#�O�rL`Z� n\(��`?D��e̪�|5+Sfא���@�i>D��Q�
ĬXJ��&E��<D��Ap%�C1���`�R�� ec c<D�̳SG�n��3��<�ִPBo'D�S��K>$�����z�1Z��!D�Ġ@%��B"5�!�қ�1�� D��Ӵ�I�r��<٥CP�+	���?D���G�I��*�fN�1��}�ED<D��3�	�,ZI����O�&i�eB�!7D��;E">�1���X�Z���F!+D����N�3��y� �:eh��(D��&)� ��9{�O@.�j];�&D����j��w�H��OR��N��2�1D���a�O.GZ��ר�{�~ s��$D�|@�q����'
�7�Ȗ��K�<Y(S�/F�|��ŅG�&�	��@�<����$X��|a&cԫg��|)���}�<1� ӻP��hRh� y�J���Z{�<	�GҘo�P���>ghpY���KS�<ifK!Iy�9RqD[�p�h�b��V�<9' I9q-� s_���Bկ�R�<�D�]'$Z���V5N�>a�VR�<Y��WᖼA�@.$| �@�\J�<!u�ChE��{�g�LZq����H�<qf?�z����u�<HPj�j�<���۝k0�0����H`@l�%CFA�<��R"D��S��1s8r*y�<��	3yS"�K&ǌ"��Up�<�@'?CM���Q噃S���ä�Pj�<"�>т� �
+J�>����i�<!E�q<-{�@E�yz"�Z(g�<������(����̤?��MȠ+Cx�<�&��N	�y�D�۟L �(��s�<AT��\ڎ�b4�	j���jWdn�<ɑL�%����a��w@6���o�S�<)e�5�00c*�!�5Z�b�R�<����]����nU�����BM<���V�����<4L0�ː�VBՅ�i�����m�'Z��Y��¿ ���S�? �����e0T�%Ǟ���`s"O��X�O�����-P&:����"O�1ˣ�_� ��M�M�L!Diч"O@9s�hF/tZXx��ƴ*���"OL5�f,�3 <["���x�L��"O���Ơǡ\�Ĺ�� �>U�Lr�"O���2Fל�"�y�=���F"O������=�FA��T-Y��a�"Op�+B �+	�Q$�Z6ᖥ
q"O��l ,���F��a���{g"O����jK>B4/\�|]2���"O8��1���e �[0�O>HP$��""OR��F�)�>1��.�"B�!��"Oj�A�(I;n���"B�%�5� "Oԩ��'�;5B��dE�"XHK "OΘ���Wp�l� 61ܜ3T"O8�#��Y�z��L*sf�
?ۂ�J�"Odp�у�&b�^�6EG8,�`�H�"OTQ ��@8G��D	Ǵd0S��̴�yrI�1'm��H�W/ E�Jf �"�y�ԍc�킓h!!������y'ۙj��Y���؏OT�q����yB� "2�����B��E��YpL�7�y�!��=�ER3)�R��P�(�y��I�8	yq��I `��T �y�.�<) cb��	%z��jM��yR�B�B�x�RB�U�[(�Ib�T��y"�D!Q��*���;Q��bD�y�x~܊�/N�yD��0��J2�y�O�a�ibGe�}�vH��G���y�䃄4A�}��)�m� "1-��y"-��93: Bq�Q�b���ĬN:�y�M�_`��(�	��X� �BI���y��\���l���ʰR=�@f
�y"�=wr���̀�OZ�<0f�yʌ7Px�8�.�=@u�m����9�y�i�YI��#$d�@�ƌ!�意�yr��k"Π:�"�1[�H��Ĵ�y"�הA	J�0�ą�<����7�J��yr�	��x,��䅬}D�Y�6�	��y�$,w,:Di��w��@,�5�y�"�$	/�L�h\lژ����1�y"d�]�d=	�+U�5.��͏(�Py�%Րf��IP��_~��a�n	]�<���<c~�J��D�J��S�PY�<�1��L [�eDf<X�*Z�<Q�OL>i�45s7gY&V8H �m�<�`�?_38�f�ʖ�.�Sէ@�<��˄O�X������d+�Ļ��~�<9� Ɓ;��$�AU�M�2��#�_�<�i�3!�����3%����^�<Q�Я_�,��KN0H�>�!$�V�<I�bѧ�p=���2c����J�<1��ٕ. ��է���h(̅C�<Y[8`�O=gz`Xӎ\e����ȓ�"��@�^ ��D(�(�<�t��( �'"��p�a�:h���ȓF�0�cm��W+�!ᦂ�r��A�ȓ"`�q#�4)
���@��.Tў���\ºp��� �f�dEB� ��`�Z��ȓ0�V�{C��]�������:(pM��@2���CK�� D�e��K�<��:2�%9T,���+$�J�4�$��%)
�*aٙ!��P3g� �܄�S�? �;b��x��� �MM.:R4���"O8H���?OM��"�K�AFy��"O��(�,˙u��6�T_H1�"OL�B��R�{3��Yr�е~�b	:`"O��1Ď�.O?����g�/7$y�$"O :B(��T��l�#N��3S"O�U�u�^X�:A1�J��zD"O�:��ğH&��iE���H�L�b�"O�A(�,+-�esO�-W2���"OB��ukԫN�u�&L<8����w"O��@W�@?~��]1�)ݴp<��*OP)���;=p�K�������'�����k����1b׷.?N���'��P����U����#'����J�'����7g�xTt�:B.��
�'6NU@�䚋u����M̪P��	�'w�qrGKߵ;o�
�yY4}��'�diY#��2i:\5�	Ȭi���
�'{4�J���e�A���� ^2�`�
�'it=hg�B�A�`UT:���	�'��%s���(�@ C`Cε6q20��'�Ը� ��K��wJΰ/�� *�'�`,��	�H��1y㛫"YXb�'���0%Ͱ���(�a��'J� T� 7,��'�V"����'
�q�����]1�
J�
:�	k�'jT9�"^&UD �����K�'�NpQn[�1�����[�T�Y�' ����� �hzf��
|^���
�'�(� ��0c�<�C�ձ?�l�'\D��)S�ڽ�E�b�XXY
�'1t@��O�,�u��Y�*	�m�	�'����(\2Z �i��̆%�zI	�'P�y##i4A��3���!X��h�'&*��#DD�n�H�I�FW3�=S�'���#�B�<����=W��:�'� `K!#�	Q�Ĩ�W��.J=��'����׬4���c
�#�N�3�'KD��B�L�	o��k'�O�j��2�'q��9��$��m��fWs����'��$�ЍR�i�z4�u'N3z��
�'vΨ�foX6Jf��u��-b�ui	�'�*T��B�
bB�Y��aȌi۾��'>�a*�O�(�HG�G	w�hi�'��9y�b��~c���V!��!���i�'�|!��$B\<��&\x�
�''*�Q6��>`�	&-��t#�'�J��U�.�L��
�5bG�,��'�0�q	�?^��1D�;^~$���'�ڌ���Y-,�"�A4N�D�
�'�S��7Pe.dc�b��BX�)	�'a�
�H��B����>?Z6A��'��!��X������� !��a�'JD�����]�F`"�Ghn2��
�'Śu��3Z��XЅɣ@\�	�'%�E�	,��S犒�qg����'`1�F ,�j�(�mC�lj�I��'�,�Z�� Oڌ��g�*r����'�` �D�(R��d�3;I 	�'F���W�^�jiТK]fL0��'H|��A;*���rEP+4�Y	�'�vq��#��&^b$IR���"�H-��'������`5�J6�I��Е�'�½X4�۳t�j���L)������� �X��CY�`I,A��쇈x���"O���톔o��0����2��"�"O�k��˰ސr�+$�D�9Q"O�dY���+P�K��G#bL�� W"O��j�JM�$�>)Sʐ7E�}��"ON��Ō� �����qTf�"O�}�%ŇIK����63P��
F"O���6�Й|��L0Т"OL���j�(�2�%Y�R	�"O��k�&?r-�!��?�h1A�"O��ە*щm/���扂�tD�d"O����i�MA.Lc2˟% kJ ��"Oݫ!�4�(�q��D-JU^�j"Ox(z��F+OJ:����ѓv���Ya"OM�"Ì�Z�^7.��"�,�c�"O�ʷ�O�c�f)��M�r��"Ol0p�cXV�z1ce&K�8�X"Oh�c���qр(r#G�u10գ�"O,��_�)�8��хrzJ�9�"O�]�q�W�G8�mK���0o���"O�\q���Q�󢄮yX�<��"O���#獶��#"�)G��%"OE���3j� �f�0%<�4
u"O���𯎄/�J��l�/b94x�"O�9������N����?F��"O5���~�F�1�]���H�t"O�!��䘈M�j��`���v>���"O�`{	�>\���jɠu^f��"OJ,B�hġ#�t:��	%e"ī�"O,��m��O���p�Amf�]��"O�;��[�y��h�
P�bv�1!"O�I!�o�\�C��Z%|��6"O(��S�J�y�TacE�	PU���"O������w��%(�#_8X9j�"O�Mh�7,&�LSƢ݇V���"O������̥jS�2��	�%�yR͒���㫎��.@�`���y���WZ�<����9	ݢT*`�˪�y��Xa��!Qlӟ{,�1hwiL �y��؊4R"U��a��hˆg�yB�N)nUq�"2]�hM��F��y��/J�*�ٳ-IOl�x�@ؘ�y�#�?�iKK�2����Q��yb�#w
�� �F�?%#����K	�y�oӌM��� EM|��
G'��y�F�'�NE�qL�H�b�4&��y2���hxj�IY!pQ��""�ޑ�y���[��]��ɜ
n���(�o��y��^�/�lࡕ ]	b�Z�b���y`��m�B�yQ��VZ�ع��S��y�!p!E�pND�y���+RO���yb��(g�**�fH,\
Рk�,�y�O˵;���A��N~F��"�!�y�@�:o��1*$Z���hդ�y�A%W,<�B.�Nb(��+ހ�yB�A�Y�n`0�'�KY���hB��y�NF���8�.'MJ��E��y���?9yB & �7Ӗ��2!ڞ�y��,Ir��1p*��1�D*cE���yr�ӄiq4t0������\-�y�j�c�Z�2�H�c����э�y!��?��a2�(�1aY�����yr�܅��E#�
E�Z92]aSJ�y��=u
)�t��z�Ȑ8���y
� ��@d�!1h^���.-1U��7"O@�y�敪9��5�6-�+E8��"O�)3jN�\�@̖],B1i�"O�K���-&F`MM�V#��kS�'�����1!�k��1 ��\!v�q�:D���CI�#:���Y�*,,��m@8D�(���>Ð}i2k��e�z�A/*D����A1#֪��J��!F	H��$D�(���z�`��!-�Y�J'D�蘒 8z+�M�E+Pj9�\�&:D��SЬO?s��=8U�O�'����*9D�p	6k�A���Se��Ag&i9��6D�,E�2i�*���%�'�}&�5D���a�խ$h���aH|jM���'D���SH�-1��{B$ �D�2'� D�P:���0`y���6�4^�����<D�X�Jԝ,k����,��7�:D�P�v���6%8t�qG!Ob��{�5D��:s��q�а�5��2��P4D�`��չ`���*6Y�r��[E 1D��A	�:�I�ȗ4J�d���+D����k�lzCAA�9ܤZ�d(D��'fʑP����2b��G����w�2D�Tڔ�� Xz����?r܋"/D���f�Z�A����+3<�p���1D�p�C�xGn����83xXX��")D��b 	��� 9�A�9~%6��a�%D�����-7�`8'��o��E)$�"D��B��
�:�"O�?,�=�o"D�D���M&�U8��Mb�cH;D�8��d�XE�3�P�J|��!#$D���P�ר,v���f�x�0���#D��2��3*�]	Ц�9b�̸�"D�@���sh��@ܮm-���E�$D�\�#P(���hژ�F$D��)EN�+���	�ܞH�lC��"D���Q�~0��(�(Y�	ߖ4�w�>D�$"�.({s!{�ׁo����?D���WֈX��x,�DT,�0# D���Ǳ+β����.$qd	�3�<D�<����|	� *%y`��b��<D�Tjr�op
`�Qf�)4+rq�/D�L�D�3d��y�OӘj���8qf3D�p�Áм<C�`!��N���]�j0D� ��'e["��!@	�2��ఓ�,D�HR�r� ��O�H�Ȑ"�%5D���2�ܫt����
�Uh<��.D�$�#$��Nk����B�&f��p��+D�xڒ&��i�F� ��y�����)D�X��'Y�k�Aq�RS�(�F"D�X)��X�nY�m8��FN�N<D����F�$��m=o|���Q�$D�ؠ�HS�c�P��V�%fV�Y�K6D�0�a��Y���s���%*�>b�!��4RH��R�n[�V(^]�A^f�!����9�2g bqH"ֶE�!�DË��Ձ��,�}XG��!��!k���0�Y�^�P���	,4�!��Mp�1�OQ�X	`�E@�.~!�8tk��xU�_�j���� �!�dI �F�S�]>
�z����L?�!�dR�Z�	3�gD�(�)� ֧h�!�d�*]������9B�����XR!�0�|0!�Q�W�{�@H
!R!�� D���蒤vf@��c�4h����"O����!)&㺕P�l��-ޤ�*�"O*��㠙�@�L��۽++���"O��䍡tk�xji�
0 ��"O8�S��-,�H@HÛ �H�5"O>�BeB�'A�n	�$�C�M��d�R"O��ׅ&���b�Ʀf޲ip�"O~��ц�"@G�9�RAæ8��[�"O�Y��%E�tZTo^���y��"O2e#�r�0mӲ��"���g"OX���̴%l�K��B�t��O�O���Tj߱�M��O?�I<y�Xr&�H [@kN5��ś�-�=a�A&�$7��2��W�M���>�����"�L
i9� ���L7_>9мi�H��˒\�<! ��ħnH�#P�;��PnM��F�P�ЧL]�Iw`�Ӧ�A���OR�$�զ��{��M�o�J|��!T�Yz#�j?9���=�ߴC�@��#�֡#����V胊qLDy�oc�8�8�S��];C��%gt�s�mN�mBj���5��W�^�n�mCX�x#s�	3Ŝ\P���4�L�Y�d* yRHq���g��2��@G!�y+��3�D"<A�+�7� �g��L�ޔZf�-4�����H�}�w�I2Q��OH"<I��#~h��cG[^ �0��E�4L��>&H��~�d�(�������'wԥ���^!|{s҆�*���ēLHz���ۚ}��0	�eԧrR��tksӂqo�k�I�^*�I�<IӬ �&�hqfD!*�V���T/b�N��VJ���<��bڮ)�̚�D*��TL�6'ذ!"E78cj+�L�>�Z���=#?�e^8H�D��fR> ���2@�рc��<IR�?'��UJJA�9�ĩ�%�	Ft��n�(��� �3|b�c��''����M�����$�O��ʧ t,���b�"�����	4��ѦO��=���f�	<�.԰���7XH�����t?���i��\�p�L �M���ħP�n}�aϗk�݀�K��k��=���/��L�blȄ��@���Fi��\�k�fE�vC�?n�h��h @�~#=i�m@)M�nѣ7��{����N:x��	�o7R�Sm>A_��uT�������Oz��a�ߦ$ϱW��͊E�H�_����$�Ł�?I�ʟnc�8Kq-Z�21|�2膸a���h�.�Ox�oZ��MS�4V.:����xI�Kǌm�b�r@[�8���i7�dѰ%��t�勇D��!2�|�	{�/�h�xtp�l�6����*�q����wZ��o�'���(d�8E8۴{\<Q1�C[�-�ĭ��*�;>�x�F%1�����#�BŻ�!
M�L�BV-Ӧq{� �OF��ɦQ�IE��M�P	Z�@@�� ��2%�T�A�BS?�����>�C�R�c��๒�!s&z�G
O�'��6��Oj�?n��?�����G��0�Hbn4*�s(O����É����'D���N��sZ��%�ˀim��P�bT4���c^�mG�D�u@���
j<{��h'ˁU��i�����\��v��Dp�k� f���&�^���/�#| ��c,�3*RԨ$��Eܹ1��'�8���',7-�9��Y��Iz}�͟8S��1!��X�v�aB��p>	K<)�H�1��t�T?b!�]�t�6�Цa$�T�Oe�'��6�
� |  �   W   Ĵ���	��Z�JvI�*�� 3��H��R�
O�ظ2�>���& �ث�O�=�p@O�rh���EL�G��-`1��Ѧ��ߴ�?1��'\ʓ���iӞ�I�6��I���F�p��Ŏ�b��9��1���	:�ɺ1H�l[ǹi���نU��}���	\Q�(O�r3Jˌ_�&l0�\�l;Ю�;,�Y��¶>y%���S��p�J�:o B�2Qlɾۈ8�u��a���`�\�D"y!�xs�K�<!/K�ϲH%,�o��Sc�_��l���kuӴ�'S�$bW�1p���'I�Y��Ɋ+�Nq�;+ӄh�����;�|+���#���$��(w�=�'�Z|�A�K<{�8�
Q��>M�'��8Dx�l�h�'`��A�<�&9���T$F�/�{��"<�f��>��I�u��P�-[74�����\�$D6�O*�0�{R���fLC PD��g ��M�Ԍ?|�d"<Q�o��	�$�����l�Pyv':e&��>1�a1�D��n�,�g��K�N�BV��8p��'�.]Dx��Z�-X��eޯ7�D-:u�[�c�nY+�a:��#<A�B�O�%�L�@TA�F�i��i ��䒋�O6]�N<���Լ6�`1��)�l� 	�J?iC�,�Im��<1���L[����?vT���)R@��F}��?�	�`2`��1�p=z'h	P,�t��S4P(��)GX�@�L�p�O~4��Bٗgщ'��E�׋P�I�*Q���d� Y�OTL�O<����{��UcK>��,��=��O"J�K��A�8��PB-D����(   ���d�X�y"�
-�DC�B�j �u{dW�yi7)>� ��L�ge���S�0�y ɕ~�b�e^�\� ���y�(�<N�^HbE�E'Jv�}m��!�dP�!���V�w����@��
	�!��R����Q�Z�޸���
 �!�d��V A&o�!a�`ӆ��=a�~2ϘDH>�aU��p;��CW�K�F�l���[WL���S�? �U)��ATE�u�p��P�$Y���ɽ+�)��
�>j'?E���W+Ătb��_.�HѣJ"D� �d��3�T��F%�~���1f*�O�����lRL�ٷ��b� ��7,ǿP�nh
�	����́�Z��y"� ��ν+V�F�tJ�pcCʎ�cw0�gꜻcQd$d53��������K�	�9�,\�Ӂ� ���5F���1E�Z�EqO�L���Jcl^;DD�Ct��_v������_Âł�;A�2��5G�zX��(�zc�a��fЎZVZ�R�"?�fC�!����]k`�Z2��4Ь� È�.-)f��O	xġ���7��S�P��[	���c�`ǝH����Q�,T�>8��%O�|�~�*�j
�0`�"Ej�	P���Gl�/��"}Z�iW��[�`X$eV�b%�4!��È�D�?�H��G���OH���I��l$�$g�ŉ^�p�8���&bH u�L�ȱ��
���) �gH�M9BE�>V�Q��aB�.�p�d]!Sس�ڴJ�)�$>T*��E�!�DIt��Q�l��6c��N�6 �@}�8zE.V�>�Q	A�/)Jau,�Y�E��F�<�"ԐT������2Zf��I�)'Z!�lH�[�A+���ô�1uv|�Ȇb�(
r� �')r�B��>����� �L���ȅC\�4"as�ZX�~���L]Y4�}"��5�Y�5��|�O�x�o*=�6�Q`%N�hQ"�'+(���LCe�Qp�E��˝:*��T3�bVb��QĠV"s>�@�F�4A(R IU�ݟ@ vB'���kC��%�M5N���n�k`��R5D�[�(��$�՘\�u�v�+TB��'�IU�#�h���Aƥ��i�%^��Q�cԬQ`&��%��.Eµh>�O�c&�4�1�'ٜ7�⌈��'2lM1⬂vx��Y�n�	z��)K�C�%�>�!�'�4���'-��pcшT��r����Z?~d��	�]�x�5���/��t2O �E��C �8�͋�,�!�n�� ߦl0H���Y=��HE�45O4]Xf���Pk�X0'$�#�ʰy#�d_5gp@�0H �H����!�&�6�#���=T�5q$H	��A���<����e�D����7i�<����R!z�d��̍�Xe�u�f+�
X�"�O���|�0K��S�Ĕ���l�l�A�M�wQʈk��r���H�&�'����D݌u��Hp�HL>Z��dX�<�e%�@�ăe��#�Ý�v��\h6�h��xQ��iƕbs��뢤L̈͐r
��p>)J)Uz\�ɣol$��άv.\� ��
g�#on((�A�-	s$H�0���?E���J�Hhq�X<�l9��*�:wy��c��E"��Q�b�BJ�0:��t:�'���S��Rގ�	G��q�'��ܘ��!T�T8#s)� ��u���U��
����Ƹ6�q����(;�RY���:�ܛ�+�L���J*0I٦l4�P�\1gE:��)6<���ɞ�W�x) �(�%e�*C�I�!\��	�L�N?2����O%�"C�	*(`9B2	�^�$�!��^B�	�;P��ɸ����h���C�	�y9.\(�� B��K���&/���Ē @��CK<�Q���UDn���b�6T�t�aSB�]�<�F+̯�@�d�.	J�#��Y�MY�2��s�)��*v��DC�+1����H*��C�6`L�1�&|�d��%�_s�q�!�$}2E� ���}&�����]�\q|!�ũ��/��=�pC���'�&���D�N�^�q�ւ7�n�!j�]=a~���00y�AÉ�;+��J҄U��p<��%>�p�k)?���RmҐ��9u �ãk	T�<�!٣u����f�;>:nukƮi�č�tvl��vl �0|�/��P��r瀵5���0J�f�<�5c��C��ay����;�p��/�\4��*�[� ���_�Bvq��'`�pAE�#0]<�h5fĵQ(���'w���E?*�ib$�� .���45V�����'D ����%V��i�1Ȉ;s�2�S"M��x���! �V�a,
岁�v���G^%�x)PU��|�z��Eh2D�́�c����f

HZ�K�o-�L���7f^�=x�G�D�F�s̀�%���
H������y"�O�j�V����*��M�W/�,����������޽yb��?�'�-s�MZ!/�*�2eF��~��
�'SN�n�.}���I���y"2�N��촁�	���0>DA��	���+Pj����]���L���2Q,ƺ~vy�%3OB�@E&�-
�P��@$l����"O�,��O"�8"��p��$����^9u`��*�	����� �u戗;���:S�ˏ<֜�xF"O~c�"W�8I�� ��a�/13Af5b��>�H?�gyME�,�La+W��8�%�Q�ybB�^%ɶ�#1=����@U��Mc�@K"&ܾ�p�Y�tA��ڧJJ��:���v�$�Xj(xGP�TQ .�a��a��W<*C��[\!���0Y�0�ҵ�T"w���׉�K�!��B ����"c���b�EȞL�!�d�`���A��>c2����E�'�!� 	^���Sm�t���Û�t�!��F�PD��Q�ǒ'����DI�!��8 L�Pc�"|��a��N7�!��EqD��F�$~4rD�V�!�����YoI�>��r�+c�!�K�u��h�Ќ|�q���L}!���c�d[M��|S�)6!�^�u[�bT�+\�`�2"�j*!�d (Jz��ْ�T= `xM��L8x-!�Dʏe�.�)TFë6	,�s [0!�ĉ&XDf�{s!�'9�(<@)Y�L}!��K�y�d<�T�Q=|��ˣi�{!�D��	g&a�/��U����(Y[J!���$=m���7���j�a/o�!��K�lf���&� $�=x��_�Z�!��p˞ �$k�l���q��� �!�մ_�꼛㣍m�x��E�&�!��h ���F��x�x����V�>!�dN�C3>��É�h��dq�dw!�$	u!��q��z/�9��"�.�!���_q� A�'�D#Ea�FZ�R�!�D�70 ��h���?)6��[sD!�dX�$��A�Ɔ��s���+.2!���:v��%i͐�H��#<A=!�U���p7�_8G8	!d1M?!�M�	�f�9�l̈B����
��z�!��Z'8�!o�\�21r�H��T�!�B�`�\90�'K&��	��B�j�!�d����-��nʄ����Y &G!���<0�b�pa�9W� ���%^�h?!�d|��}`t�C�4�T5ɀ��A@!�d����PPT��)|&�z���h�!��I�w{����U�\l��\<�!�$J6��}H��UT�t�!�B۝E&!�$�$h|r��D0Fm��')]�!��/A���'�̎F/�P�Gʺf�!��@:�A�jػ@~�lp�R��!�d�/��z"�V N�<��1�֫F�!��-<Z��A�[�*��!�@��#b!�d\�)�ʘBB)F�f��P���P�:h!�D�ou���#�u����#_�yA!�$��P.���`���V����C��K�!򤓂9�.|�%�-N��ss(N�p�!�$�,_pZ	䉊�l�}��h��!�D�I���+ҢZ�j�.U׆�;t�!�ǅX�3�lȍ&����T�v!�J6=LaE� �&�4mp�o��D!�D�(yh�����<��=x�臭,!��\�����+	�w����F��+d�!򤎼:�A�PbZ=B�v�ZE�
0!�D�o��R�r��IFe?!�dП�| �OF�iunq�f��'m)!�G���@��H�,H�Y�bA'M!�	&V{L�9֏�:C:�����!�D�
@�ҎʈVG�6BW'F�!�� .M9p����޵hH¬-Ϡ�Д"O�m!Ň+LȐ��n3t��4	C"O
9 b�*v �#�+W�y*���"O,���&���`�9Z���"O����89��L�v)ǎ7�(��"O��t�L(��3%��RVKr"O&I;P��\���$��!��av"OL}xb�*A��s㘅tp|�"O�IR խw����5ቺs���0"O��3d��m��ѓ�� o��5"O�R��˭p4��#i˸s����"O��zG�άDϺ�r��J�e��T�"O��s�ϥ`�< f��UΤ��A"O���Tf����T�T�E�u�d��"O<$�Z;u��y���)�4���"Od}��M�^d��_�r`�@JD"O�a�g� p�Jܣ�,O*��z�"O�\2Bڞj��z��ܑ@�|k3"O~h
���U����<a�:�"O�����}���S5�P�^��B"OB4�M:}[>��L���l
R"O}���>�K!k6_�����"O��[2
.OÈ�����l��TK�"O�Q ��!�"����ʿZ'j��"OF-(QI�G�`5MH/#�5�"Oܨ�4F� )�=�1��C���#"O��j�9nD����.j��E�1"O�8��]52�z]�`��;�~�h"O��(�/h�=���N�:-y�"O���"Q�6����@�K�TES"O!�Ɖ�i�����jB�!r���"O2�3��W�9�삐�Ȇn��iZ�"O�y���N��$Ȃ�� �N��-j�"O\���&� J�Hi�᧞��iQ"O��7$
�.�N�($�!�pta�"O��0�O�w�(�D�ϣ	\rM��"O�5��	@P�tjٗC�:]�s"O��s�̭'���K�# G�E�E"Ot�+��p��A���?=32Y�C"O\M�%�w����lĊe5r`I�"Ojps������W,�.����"O��� �XM���KҰ�YV"O@�q��k@�h#@����C"O@̢cʀ�\k�t��J�&!�0�"O y�֣Y�P�t�[ �A8Rw��"Ov��@�(YQ�y�H�{j^%W"O�����p��q�F�CN��"OB���H/H�%£&E%z#¡�"O@���m�u�4����Q�B��2"O�˦'	R��Y1&���"Of�����%4�L�f��,\j��T"O�@3��˸r�������TJf��"O�)
���O��@TC2�=�"O:��q�,A�0��N	�!27"O�����S�8RU ��z�j-�5"O"���鍌bݴ�� %M���r"O�$h���+"�B�,x�C�"OpբbJ�?���㇩ʢo�x"OV���@5�T;ANZ�g�����"O��S��o�����'h���j�"OD�k�7Ll��T���[�X���"O.�+�k�&~E��9�B[e����"O���@�#G�a�'���Bv���"O�|�#�=Vx$��$OR�j�����"O� ��S��W?k`��v�4�����"O���0��%�����%_&Z��i�3"O�M�%M�u��d�ģ�=<}�Qy1�'UZă!�7��1B� �DD��/ly�ii�J�]<���Зa��CU��E�&��d*Fy�'v	�b,�0{�������N�+��,����n�th�d��y�Ə�I�]��f�.b	8�@�)�?��Q$j8��`ӊ6�fX��i�42:�11H�%g�d��P-�)}�"C䉈^!�ѩA�@��H�9�G�K
Μ�U"_ݦ(S��+1̀ȸ�I@X���d��?<�PG���}�BC $!���;�-�{J|b����O��9Ф�6,�hy�iS�m@���X��C$P�/�faرI3�O"�h�mz((A��J�(B��՘�T@��YPU�l�#
6NXy��D�ۢ����$a>����*_�<�xu*0�k�������i��P*��ζi�x8{0史$�bI*$�,܀d����2Y�+���J�!�b�7訟x0)��V�e�%K �׸pP� 2ړIH�A�u%Ex�b?�y�����Q�w#F���iU S�qg~���m�|?v|@@쌟S*�g�'G T�q�"E�$9kP��!%"Q�s$���2t�1L�S�!'(I����*�0"�Ԁc��	'ƕ"���	%�V%af-�O|LaWƍ��ݸ�*��
Kxyw9O�00���\h��$�������;5T��tAIo�t� �;���x����$aė���=�a�!Ar��H�58���K�$��|�!� Ѷy�*�O6@Q��N�`:�g��u�#�U ��`�A	I r�*�[��[p��}��X[fk�^	�b�2��0�����áv����Zޞ))[��'hhS��ԩdf]�G�����٨&�|��įIl�%�I�z��b�'��>�ɮ>��8 ��JXH��s!ɶ�"��c����"�0ɛ /��/��!3���+���S���)��i[3!x���)��,5�ĔA&�PCBO�c��{BB�4!�,h`6J�)��P��F#Oc.�Ă�:1���"O��c$GÝ��ѻ�n�>�>4�B��چ%S!G����H��0�d!�*4���B�,~��c2"O��� ϖZ��u���� L`��_��bՑuKg��-�g?�թ .yR���{{�2�_�<��@�Rv-��˺w�>\hbd��<!E'�\���s�i��bcl�*1]� ��)h�����I����R7Of���	�|�@a��I��U��q�"O��⤦E�
$�W�P>�Y"��y��
�g�:d��'�@4H1��m�-�y2+ʆ ��P��8��M��ȓ�Ny�._�L�$�yA���̘��r�f�`A�mZ��Q�ۂ0q���
lhc��M�ta!�@ɾFM���|�� �] i����(�>,��y��HI��ِ���uT�a Y�/D@��ȓ'�"��rlR��t)@Ƈi����ȓl����5�Ϟ8C��hBa��h8�牞9A��xR�x�+� #h�iR����ȃ��yr/�+~A Fl�$z�v���
�ēI�����K����S�z�J����g#�}�B��p؁�ȓʜ���1�T%�4��v�.\9��I�DP��A���L>�Uw��"��1]]Tu�_}(<���H�a&~1�0'��%�L�J1�$D��IƢ�w���ݯf���jE(�.���[1ܗ,s�x�ՠ	z�<��ED~�#��y��rPcP1���!���y�ե9>(*��І]���FT3��I!�$Z��L)dna�4NQ<d*H��K){�&�T��?�yb��%T�$���	�i����CV�@\HR�h�<q¯�_�>�O�D�geMC�����H�ABPz�
O&ტ��o�ȝ1񀐶Z�<�)�$�Arh���L��m��ɝn��ؐOӑm�$e	c�i���DþOA�}���L$}^�ɛ'x����)�1Ө`���ij�yH�'����w�^0B,��� V+j� 0�J<9��A-T��)06��;8�?!��_"���ht�v�I5,,D�hQ��@�FQ����({t|h���2u9T/�<���	�����	n�ٲ3�	!�i�B�NޘB�)� $�A@���*��c�57i�тvE0�	��S>�a|�CӂG�<�8��՜s.l��7i��p=ie	��e"T�k�|1 )��8Wt�K��Q�\)�Q;�(&D��A��8^謈&��!t{���D�+?�p`�S�#g�?���ÐX�p���ͻ��E�+<D��1t꜔�je��%\��H�bٚ@��QA��6}��s���d�f�D�R��z0�aY��Պu�!�d�RԢ��ň� =��A�d��V�Z2���'yޝZTj
�~�с�(����Zߓ8���8���>9_(&U�C�5@ oC%Lĝ��D�z=��lG��\A� �=�V�ȓ(��Bc�=qA�@��O�a�����:�ˉ>	�H��H�*q ���&�aT��y�*u��/�%@F�1��x��%q�OP�/�Y�� ��ȓTA���f)��
8�I�W��W�4���)q ���I�4�Μ��	ݭ)2�Ćȓ	pF��f��"Yf��{��M$"'���ȓX�~������8����Y�\,6$��MR��0"ȼA�����(NɄ�I��4{Bm�d�T�3��ՓO谄ȓv��\i"E�F�ԸK�G�kD���ȓ]q��S�障=��%�*EPf݄�o�8thoL�*`*iP�B��������À�YN�H��.�Q>�=��qǶ�ȓ��%�9�'EÕb1���Y@��eʫG���J��_ɨ݅�B����ʴft�qF��\9��P�޽�C(ZXzA�L �E]�8�ȓY�d��E�!�R���U/#,Y�ȓar\�1!�M �:3�ѷZ&���ob��Cɚ8p@��b	�BB���ȓN����]�8xC��֠2V8m�ȓ~�*9������kA�\�j��`���>�Z�-8v�
C �/�����4Y��N����T:�#N�����M���f�r��wx�Ņ�Hm�%�Hq���ZG�ϛ �DQ�ȓL6)J4� �uO���W�ܫ���ȓ\6�HXe���Xc%���"���ȓGĆ�;�kK�:��a�CǶ!���l ��
YT�P83��מ]h��ȓX�j�j&���Jv��7B�q{Z�ȓ-<�x�/��	zLu����o��a��T_��A`H�&.�7�_�#�f)��O�v����V��jb���I����ȓ_א�Ked�	V����	�(n��L��o��m�`�=$�*T�>a���ȓw����1�A*y��i�7�B��p��ȓ?�r�����os���-]W8��ȓy����Eܨ|"x9  �3Ip�Ȇȓ%�֨9�^'A�j���#_�c�dцȓ0�4)HAi�$tX�cQ�Pn����;&�� ��-$r�Q+�~��{�h���M�N]j��!��'��U�ȓl�Ȩ���ٓv�6�Ӗ�Q;G����Hy�[�J�qI�L3*��ȓQ<�Y��#z�P�Bt�E�ug(`�ȓ_�p -��	lH���c����g@,�b�����(�h��1�ji�ȓ\���
FN�W|�ũ�+�?3<ąȓZj@ah%n�*��M�Ub����ȓY��pa� 	f��pM׷6G��ȓu'��� ��vmx$���;�t���S�? tx[4)� B���!�=O���+"OP��)7Ha������d�be�R<O�L��F�+lt�3&ʗ�*�l�r�	p����5+��#�,1A�%)��B�I	��R3��@���Ưm0B��0NE]�4�ٮcm��F�D�&Y B䉷#��� tO����Yy�m���C䉆s��rR�S�Qn��r �� C�I)n��h��,�X%�$c��g��B�	i�h�`��lN4"��.tKdB��;!gHTy��GF�:�XA�Vw���	jx��?E�T�wJX��j6lk����*@V(8q���Hܓ��I#ʧ/f��5N�nޜy0�Y�y���r��^�	 y����ӂ� 5I��$�����TAI>y��G
�PI	ç]���"�J�+ P��@�Q���'%�H�bK� ���Ո��=91����[Cb¬w��T����r| �A;5%��7�0|ze�xf\="p��E?X�ƍ+wQt��w�c?����5o�����4��32"����	¹�NB3K2��6�  ��i�]��^>M#�i�t���[�Dn�\XƑ���I��^u�Ԅ�0��ަ�yçK�\�����
��q�����I:Ψ��ρۦ]�2�iza�4��<@*Wh��7'�]��`�9�~���#!�M{���>+>�1�O���J�F�(# m����z�����)�Mu$� � ��e"�a���z���b�P��U�Pl
��M[R�=5Y���J�;J�I���s�:��;"i���hT�ra:Ն�Ty�*�f_�x�4%HW�<I��Pm�J��	��5�3 ٚ�������"]� ��8�7��"4~tY��d>���.Bl�T���h�����fR�l�06��J����߷1��HF�,OHi��l�2���$F�i��P��i��i�B��"�ƌ�O?7I,
��͡$EޤC��rK��c!򤟋=�d��Go^0yȖ�$וUI!�D#`�L�5
�FP�<�Dc�0ld!�&[�(yX��[�GhTD9�#S�bc!�Y&�8���+�)ZX��p�^�Z^!��
���р�ѫe4x��䏭iY!�L9>���V�x`�)��i�!�D[�6^b4 �瓗YLX�`$� �!��Cǐ�#v,G`�:�]7g!�%�"�*ë�"��#�/͑�!�dE�zۖ�����b��$MpN!�$%L��Ѡ�Ŗf�I�Tnҁu]!��ű>Ң,!rd�!X}ꠊ�DJ!�տ1� �+�U�q�fI��hB!�$B�V���1���BЎ��­ǐ>-!�$I
Q���q�/�/��$��M#w�!��T��,ф*� ����-��u�!�&�ic��L�p�dC�{�!�d]1*�>M�ՍumFdɥ$ǻ�Py"cN��)8�eW�2'���j�y�@Q6P���,�z�P�gÅ�y⡒8��F0p���W��y��	�x|�"ٶ���
��yr$�-? 2� '��, ��B����yBAǫ�Rc
��t��Y������y�c��n�h�*��]�j^�Ɂ'�y�K�DR%DN��������>�y��1V1��i׈���@�Ѷ���y�BZ/1Y��A�Z�^�P�/P��y�䞫N@y�#�OS��q`u�
��y�\�r�ΔA�� ���gJ��yr�W�0rθ���зcC�]�&攢�yb�V�IX��۵%�[~	ӕ��y��^$@\ (����C�4�B�Ⱦ�y�_�8�isdPH�|��(��y�儀p�DA���38�`��1�(�y��4\<Q��̰)��s�⛠�y"	ݎ������0����p�F��y
� �LB�cŤbg~!rFSA
j�z�"ON����3!"�ř��nh�6"O8�P�Qf�b����0R�EKW"O�� +J�s\Lm`�-ȷZ@���"ORu�6M>O�a�+֯A?Ɛ[�"O�m�"/�?#v4��Q�M�M'n�C"ON��w@F�b�Reb��˷��hW"OD�� ���z�j��v�\Z���"O�����](i�* ���E\�)��"O8P�CJ�2�XdS���>��%s"O
�j@�A�X ��#�R>,�2	�G"Ou3�D_����ȍ8�2�x�"O�9�u�*LN�ي���42�(e��"O����<*ќ���ċ��V��"ORM����O(^���0�NI2�"O�[Q%�r����R���^�����"Op!x �qn���T�d��%�3"O
UK /J$V6b���	#�y�"O �b)F�0:
-*�Ú�F��� "O2�HQIG&?~q�2 �>�S�"O����+P�^�`������z �c"OJ`���#�"�n���0x�3�=D�c��U������z�P�'D����dT>G�q�P��)�0�G1D�Ly�(��dR��
�-=�=��E-D�L�C���H���bGY19r���j7D�$��.L�\	Ir�
��qW@yZv0D���� t�yP� [�,�q6@3D�8hC&��}��}�v�˽{����o/D��9E(F�cdF�j��
��`�&0D�L13Ϛ9Vp:X���C&U�j�b6�-D�`��N��k�T�e��oyp��(D��0%�R����6K �It��U	 D�i��I�(�
l!RÑ��3�0D�� s�s��ĩ�B_��9�/D�TJ�bͻ4��`�ebP�|�XaE*O��!@��5
�9�(�R��q!v"Oȁ�u���3
�@tFJ4�T�s2"OF�b�E)SnY;��ڂ;�R�A�"Oz �� �.Ql���n.S� xh�"O��bp,W�6�1Ѝ�:Wͮ5*�"OZ�(tȁ'N푆"�(�>�KW"OH��'@�5h���'�g`�{"On�i2Ă�7䙹�l�����@"O�l��,�K���c��ԋ:�a��"O< ��dֺ'�H�+S�҇��s�"O�R�IZ�t�z��ȣp<����"OR�z�)�۶�&��}8�� �"O��v�aC*�r!,��Z���"OH���c�|r�t���Z,B���"Of���]�}� ���iO�y�� ��"O�n��l��ĵA�(T��"O�}�6k �8�]�G�V
A��"O��Ӓj��[��xW�A�����"O������SԚ�i� ҔZK�!�"OPi��䄉<H���`́\Ԟm@�"O 0Ѕ�0*���6L�	z�-Ie"O�3V₀A�����M�D����"O�A�£�~պգ��A$@|5p0"Or�v�5h:�	У!�0Uj�]��"O<�`$���vzj��!�ʜ��QE"O<@��eD:%}��1QO������"O60rdHQ=2���0h�>$�f"OV�薇]2c��p����9��"O� ��%�����e)c+ԍv�$5�"Odr⡈8
g��1j��s�pi�"OẂ�xe���h�t��"O����@�$��K�R0���"O:���.�y��qq4DýV�9Q"O(\���%=�}y��Û	����"O��q��C�ɸo۞|���'�t)Db�i�Xq��(L7n
4a;�'Ӷ%�bE��W�q��(�lO╈�'�BXШ�2	�a�P�Y]=f0��'�)*ծG�G^�,5�K�[����'�d��ʜ�bpeЄQ�T@$�`�'9`+!ϑ�tEb��9T�r�c�'�� :b'W_����@�x��h�'����
&�����<0� ��'	r�3� ��#s��@F��:e��')�����
�eq�&ۥH�*qr�'](*���>	CMX��ݛ-B��
�'����&S�0�ct��-;I���
�'���¤H��T+l��S�:�x"�'���z�@8D�J��3���]��:�'�a��[?�fl@S&i�Pi[�';�J��5a�m8�)�,�Q��'���F�i%���3��+$�:�'�$ [�aG�W���Tb5*�Ƙr�'�Ni��+T#]�qATȐ�Y�lQ�'����n��C��0VmA�'Ǵ�˲��0aFp�Ue��)(�'b��놭$w�	��I/
^H@{�'�H�s�\�JvN���!A��I�'�8}���jMl}s4O<�ԍ��':}�C�����9c��
u��'*8�O�x�dpү�<3�����'�P�+2���f]AE���t����'���{��5	A��IՃD�dz\���'3�T�0�B
M���i��P�X�����'{��P��BN��]:sG�0�'�Lx�/�W� �HuE۳"w��@�'����R(�a��`B ��i:�'Z�8`A��$�.Y���,��'l��h\�V���Ӷ艠l�A��'*��
\�~��&�H�U��'\t �ɟ���(��F
��L�A�'ҤY�̄�:� C%Nӛ{�L
�'28���΀L�Xj�
�4z�"S�'�Мd�J"��!�ז��i��'!��u�ɫg�Ɓ���$��'ٖa�����B�|$���y�'n�`�녤#/�]0UL�76!��'d��T�^`k�&�}:%1�'�|���L�+��"sI�r=Fs�'C&���!�������E)_�i�'Xj��3Ñ�:	#q�S!J���'�r} ��I2���)�$E�;�*P��';>��p���ZL��(��4���	�''p��OV#Xq��j$&N
;;��#�'�t]�!��@���9�e؁72�'�x�B�D��HbPHč),�*�'9�j$GI	W�
��d�ݎ �d���'�ҁ�C�O�3(�D�T���6"5��'�	�W�"��VF�=�0l�׈"D��c�*��u��H�&?:т� D�t�dN��(����r�M�d�F"4D�����za)�d�v�F# ��y
� ���J�Q�vԻS�L�;fH�t"O��b���:rIJ�OA����"O� gցv�0���'O�(���`�"Otɳ�Θ`
'ԉ^�p�V"O�P���ՊeE�@��B�̸��"O��3�̄�q�x�,P$��A��"ORTpd�K*��ɳ�(^���"OP1�s�l��)�%�1_�:Y�"O��)!�W�!V��5
Qu� �y�"O�)��jB_#�)*�I_9ՂI�"OL ���-�:hs�R�o눸 "O,M���S@2D;R M=8y�˲"O���!aI�'ö,���s4�Y�"O ih���~r��#@�|zj�I"OV����$+�0x�LJ�.Aj��6"OXL+SJU�ʍ��kϽH7�a�a"OR���gWt�Z�W����R5"O�T�2h��iR]��H8ߊa��"OZ�H�'��]`R!PC���	vZd�A"O���GӃ^�|�FT�;�p�s"O�p ��d�.Q�v��Sc.�1"Oz)A��<p�B�X���A<|)+�"ON���-I��z��9tjTç"O�#ҡ�+�Ƞ��O�
���"O���'�R0�g��7�r$"O���+2@�"@���@O2!�A�!-�| �)��O�����M-.;!򤏁��M�q�Y7H~���Z��!��WCi�*��{k���4�;!�DAܴ�لF�Gcr���댝`�!�$����Ư W�]Ybi�7f!򄈈'� `  ��     P  �  �  j*  6  oA  �L  KX  �c  �n  iz  ��  0�  E�  ��  =�  D�  ��  ��  &�  k�  ��  ��  X�  ��  >�  ��  L�  � (
 � � % f# K* h1 �7 1@ OK �Q Z d �j �q �w +~ �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c"OV�Wc�6�:�3�	�C��:�"O�`y!�������3-�<�"O��!S��3C����ǇZ��\�C"O�V��vA����EE�@�J�yT"OtXa�Ǫ|�t�2&�ۥF<��BC"O�i�w��&dUj��+,1�4�"O���I�tͰ5���߷O�y9p"O��&�(w�̕Z���
P�C�"O1@ŏΞ
f�}KT��}�P�&��E����8�8��͜"U�^�p"�ߓS�!�d߅X����%.ͼ2�EO	n!�� D���f��Ik���!ڨ$I����
O�6�L)n4\Tb���>5����� M�!���r��� �� �6<r&��/C�ax�� ғV�1q-i����
"�F̅�xl�X`��+D�ez��%� ��\uj�0��R>ܲ%`��T�ȓ%z�d��� �l���;�.N:d�!��_}��i�铬�O$�����%�tm�P��3�<�9p�'$
��,������/"��( @_�EZ��p?y��g0�@җ�L�Xw2)��@�'P�}�uBC�ai}1.I^Ȓ���&�v�<لBޥ9�����d�U��0�cLLy"�)ʧD~R�W-M�|E���P�ÁST2؄�?�V-���d�����=f�05�ȓ`�ꕉa. N�И���,eL��Q��=(#�UX��|��.ýN�Q�ȓ1���vh�9��R7C�7���ȓ0��	�kS\58�qr��*����y�nU9��ٷ%@�g�j�� �ȓy0��&�C�cja*�ɜ-w�
���W}V��K�:�qi�X-+����ȓx6Н"tLt�r4� �_!S���%��!��	�_Pq�'���x⥇�z�`���F$m�,�:�!�(T�ȓ+d�a��ڀ�XQZ"L$$}�ȓ[�P�Q@�>�fM�h�c��h�������ɓjfD��3�??���b�L�e�
*��@���1&�Y�ȓu�\i��K�c,���ɏ>��̆ȓmv=Z�'��CWx�1�����5�ȓK'�� P�yN��WɉQmj݄ȓb�ƥ2ڟg�a񃊑+y����E��B�X�`��i��h]>�ԅȓm��́��:("ĉ�gvͅ�e2�q�
*Y�P+t�&�Nلȓ�F˖�]6AI�,[@� =o*Ȅ�b��|�1�р]���:CCS.TRT�ȓ�GϘ�1 ����l�(LjB��ȓ9�^��&"�$|.)��J�wN��:M��vHP&%z��b@%g���-z�!�7;L��7�����ȓ^��x��iI[�4	7o���x��i�!sA"� F^<�R$��	�q��0�yb� �Qi(P��	)j����jR� �uk�$�$�����j�p�ȓ=g�`7˛D�`��+ɨD*��ȓ�p�R�]�
>^������h�ȓ"�������\gـ�kQ�@T��De
��t�@$�� �,�e��=�r�3BΏ{ DIHF�ԌM�^ąȓg>x��e�hF<�m�`Mz�ȓkڸ�iӇN�R��@���yF5��"���ł!n&5�KՆ��ȓ�����G�1Y<�r4�Ŀ	'��������p/҄"� ��Z�< ��ȓ�Q�IWL���2чF8�Z��q���K�	J}�܋�ɓ	A����u����wP�|>h�#�G��x|�̄ȓL�̠�Ve�]��l��K&cD��ȓB�v��nӝd����ҡTh��ȓp"�Y3�Ϲ7�``���5����ȓH&�%H2�@�f�@ (Vc�:o���ȓYj��p�،=��-�%AƭJ�l��ȓNH0�
��"[~�x5*M4NB4��S�? ���09�45p!�Ђ�=��"OV͓&��!]>�j3��E���S"O�q� f�1&aL�Xb*͹	���H�"OH|P0ßb �9q�dhʤ�"O��S����@��B��:�f�'�b�'���'B�'���'XB�'�xH7H�3'HZ����N�0̺����'�R�'���'���'^��'�b�'������&@�1�aDA�V�#�'G��'}�'�"�'v�'���'IXݣ`�;48~�Hg�i�eq�'�R�'"�'���'.�'���'��	t��w�(��B�+b9�W�'HR�'���'���'~��'!��'F��Q�˥R�\��F�H����v�'�b�'���'P"�'�b�'���'�L:�#L����MB:p�0���'�r�'�R�'���'���'*��'`��r֥�Q�r��φc�d�t�'B�'z2�'�r�'�r�'�r�'�����uM���C&K�_�����'v�'�b�'�2�'�"�'�r�'x�<��B$1��Y���%a�|��!�'22�'���'���'b�'I��'�&8���<�.���eϫO*���s�'��'XB�'��'��'�r�'�<DR��9��h�� �����'�2�'�B�'��'��'���'�P�rr�;�MZBn^�y}Ju�4��O����O��O����Ol��	㦕�I˟hz�	̍Y�LP���l�h�W	��d�O4�S�g~Ҭz���!7�R�f f<Bl�/#4�a����BB�I��M���y��'= x�O^�M�����U<D���'�"�������'1r�D�~�%T�zP�!1u�h܎��b�\{��?�*O�}ڐ1�\$��LA*z�h�%U�,��6��Ę'�|mz��J.A^e�DC�"��p��ó���D�	�<�O1���ZT(Ӝ扆��JBH�M�F����ކ!�d�I�<�4�'K�iD{�O� É�JS�藲P3h51wHɌ�yr\��$�Z�4mOV��<���R�c�P�E���H2A��'c(��?���ybQ�$c)S�J�6=" �ҷ$P)hD�&?��A�\œШģA�^��'�?D�O�Z���ʁ$RFxsE%�
���<y�S��y򢗯Iu����a�E���3��۪�yb�sӘ�۰���ݴ����DNˑ<�1* a�F.�h���y��'R2�'�()�ѿi����|Z`�OF��Yd��9���B&M����1�ݟ�'W�i>}������	П@�		)���GIR/O�d�U�f&P��'s 6-�j�����O���矲�	�O���N1�DM�s>�|�D�߼VL��'
J7͗צ���)�H����1�S��a�6@�6L ��F���`Ա����eM͠	�Kr�I`y�L��U4ǎ�6���Aj�(>tu������	����i>��'��6���h��'�hA)��N< �`��#� ��85�'��6�<�	5����O�$�OBE�'��1N���je�+��[�(�,l46-$?��oբZ����K�������lף<e� ��"ΐ�6��`�p�8�IşH������D�b2EM�a���	�h�0�2dl �?����?�D�i�(	�O?r�s�$�OV���(�H�22��v�f��$%���Of�4�z
��c����h4� �����a�㭍�63D�Ivl����N�ICy��'<��'\�k�NX�<��7*����L!$���'X�I&�M+�AM'�?���?�.��-h��Zq��i�$ǱBq	�P��|ѫO�$�Ox�O��N:�h���H��bK�J�꤇N>x��o���4�����'��'��+�ᑠ5ά� s�ף*ؾ��'W��'HB���O�	,�M��GP8 �� OL��iQ�I;W�d�#���?���i��O*��'.7�	:<w&4�g3�]��ㄛ���oZ$�M�u���M��O*	X2D������<��.�9B>p(7k�4T�6&Q�<,O����O*�d�O\�D�O:�'K��d�0��Y�A�eO�)� t�v�i""�)s[�x�	e��<���w9��kG͔�{���q��i��1�KmӨ�nZ��Ş`�rݴ�yBhFv���2����P���_�y���s6��I/e�'2�	ٟp�I>��1Y���8�@H8!>lx�	՟,��՟��'J7팰G}����O��D<�X"�_E�D}HD�!7r�ګO�Qlڟ�M�x���Ff��T�:Q(�W�Y���$�st��xQ�3r�"����0��p�����Q?h�2I�^dPȂ&Z8j���d�O6���O��'�'�?7�����8�	�n�Ƀ� G�?	2�i�РP��'���vӒ��aQ��Sva�#���F,�.e4T͓oț��W؊7��Ch�7-*?�V,�!f&��
�E��!�V��O)�(��A��K�H�N>�/O����O����O����O�M�2�Ҫ90Dpiáh��f	�<��i��`V�`�II��,"G�n�JT���ԕ�܍xS"O����Z��]bشn���O��T���R�05��A��^� ��J�g(�C�W����,%RM�	ly�" �k���Y��X� 	�\
V.a8��'��'��O���M37İ�?y�#�>z�T̉�̑&U�Ȱ22i�+�?���i��O���'�7�@�9�ٴL���1JBF	���"6�rg$��M��O�����%�:F�9�	��� �=�4/؅	I<Y牬"�i�4:O����O��D�O��d�OJ�?��gJЙ:1��2)̊n���ܟ���럘�ڴ(� ��+O*�lZZ�ɞg��I˃)Lq����!��~���t~��'%��Owd��зi����g���8 �G��(���Ĝi��ܩ���b��b��Fy�O_��'7�B��K鲝�B� ����5�&bR�'l�I �M������?Q���?Q*�x	3S�سU*��t��k�L��!��x)�O̵n�M[��/���N�"��Ǌf�(A��M�LuAT,Y@U�b�����i>�t�' �'��X��ĭE0X �������*K�����ȟ����b>I�'vJ7Y�"Ξ4J�fã"�]Ivk� %\p1�<��io�O�]�'��6��
��1�5���8�yHf��!�ةl�;�Ms����M{�O�9z1jU&�bfĤ<Iw,�M�.I�����u� \p��K�<�,O��d�O��D�OB���O�˧R�`��7(pڝ�gF�>{�Hm;��i���C�'���'���yx��nݼ3^����(J�Sbn��������oZ�M���x�O����Oh�d趱i	�ĉ"CD���j͍,b�qz3
S�a���D�I��Ѐ�5���O���?��=�A���:=���SeU&a�X���?����?,O$Inڐa���'7B��.q �K��L�}�Ҥd��$(�O8)�'�7M�٦�BK<��f�5g��Xa4D�e�\���m~�h�`Z6�d/����OE4�����"L�	�b�����,j=JsLђ0���'z��'���S��婛�*w^�F�I�:���
�$�x�ش^D�4y,O�nu�Ӽ�Q�:��o�&B܀��B�+�yb�`Ӣo����H7O�Ǧ͓�?A�ƞ�R���z➹��P�rPБ�����bY��O>�)O�i�On��O.�D�O�9��/ʐB������5���btI�<�`�i��5���'���'Q��y�H^+Wt�bS�`S�m3G�Y����r^�6|�9'�b>�6m�#c32A�T鎱!at�����y��2f�vyBo�#�!����'&�	���D֝w�d����+]ˎ	�I�������i>�'I�6��v�\�$����=N",�LSM���'F�6M)�	�����	޴]��F�j���s��paj�=_vN�e�i���Hn|骵�O���'?����h�a�o�Z8���	����Ɵ���ԟ��Iǟ@��_�'_!t�JG��5(y�x�e�Ў2�t��-O��dަu �f'��i��'W���p�ߨ#ƹ��C��1E*���O�6=�*1�F�aӸ�)S.|���$FV�� ��6T����	W���
����4�����O���tx��� ̾y����Q���p���O��i���*J��y��'��Y>� ��t��!{d�_ Y��ċ4?�X�0��ӟ�'��~�V헱_ez���,�8J>�2A � h��D�ܴ��4����'8�'[�=���@
J��q�
�!������'���'�����O��I�M+tH�U[�Z2Cҥ{���h5�^�.8�'��7�5�������O�(����r[G�ģa�B��gG�O��d�,{�6-(?�%K4���>=h��2i��@�!�5,��8�)l� �'%b�'_��'x��'o��8FЫ���BR9C��Mwݪ�"�4.g|��,O(�$=���Of�oz�=��Θd�<a�]��(�$�ȣ�M��iںO1�fP�e�|��牎P_�Xa�g�/��,��K�5CX�F��8��'��y%�(�'_�'���c�y����"[k|�P��'r�'�R�H)ܴ� �y���?��}����F��fI���T�J�2(�>	��i�7m�R�Ɋ6wȘ9�)��b�6�g�� j���oŘl�DIT�������'@�V�$��?Q�/UV��;��V�wwUu�ʕ�?���?����?э���O���!e��@x�ħ%0j�(���O^1m�6��$��͟�ݴ���y7�T�D�l����ւD��A@�(Z9�yB�f�^�nZ.�M�MH�M�Oz9Æb�4�B��L�+�摢�Ύ�tv,���&Z }X�O&˓�?����?���?�q��t@�)ߟ#���j�! )8�-O��mZ�T	����IN�s���@dȞ�>}"���JYr� ���Ц��4jC���Ox9�NM�I�T�)�/�|J��Df�Ԡ�aX�8y@�G�tW�NGs�	Uy%	aVX�dቭKbV���Ԑl��'B��'-�OH�Ƀ�Mkf�6�?9�ϔ9$T�"bI�~<6��K�<q3�i��O�P�'�z6�����ߴ8����_+A5�H���C:3�¥��a$�M#�O�4ۓ��:���
9����r�� [��>�Iw��>1u"u�36O���O���O����O��?}х�KV ��`�laS֮Oן���ɟ(p�4z���*O�n�@�ɮO"uɶI��8�{����*&���L<�i��6���89@Fl�j������+�1��y��M�?=�������� s�'�t�&��'���'���'����vaۤ8��z��)~jιa��':�[��Hݴgu�p�)Ox��|���̉|C�q1!/�7W'<�a�J~ �>�u�i�z7��O��~J�""1afm\6��D�f@rj7���gMu~�O=h���8jm�'��)YF�P=���eo�2ATX;0�'�2�'�R���O��	/�M��G�(߀���!F�4U� `K�x�r��*Ol�n�D�N���͋P�of\�j���! ���c��<�M���+̪!�4��Ċ78�9�����3� ��g�};d��rL#�jt`�;O�ʓ�?Y��?����?����IK�8E�B�.��cJ&�F�UL0nڈ�������	T�s��[���k��Ք9i�Mp��Ju:���H�6	m��ġ<�|�DK0�M[�'�ڰ6NJ?9 �u��&Q6��'椬�s��֟ő|2P����@��ȟ��L���C @YHD��Lß��Iȟ4�	xygiӊ���!�O���O.̀�!�x���H�&Ìu��	���3�����$Ʀ�ٴ2�'p�(����n�`�ʢ%�(�V���'���,���ymEo8�	�?���'h���	�`3R}�,{T�k�mI����	۟����� ��t�O��EO��6"�Ԕ84؊`V��cӞ̀% �O��$Nߦ�?ͻ6(�LX@�$BJ�I*�˚�5vu͓EE�F`iӎ�nZ0�Pm�n~2,�35l��Ӟ	�\���&0W����Wol���|RR�D�I����Iڟl�I��dJ���(��%�2��P�v��C�jy�$cӎL)���OZ�$�O���$��(�\���b�\f���f�'5�6���]JK<�|�0K	�Z�s��82}<���/_���i�� E���Ͽ5P����Q��OV�a���U��&$Y8dǜ�;T�t[��?���?��|�/O�l��9��I���ԡV�ڳn�:B��:�ɔ�Mc����>	`�it�7��¦9��S&j�8���_�����[�N}�%�i����;CA���O~q��.��0����f�H���g�P�=��D�O����O2���O��$:�5�����1ڞ���!J�~�Y�I̟<����M� ��?��$٦�%����.6�R�c];�ޭ�ݿ�䓺?���|��Eٴ�M�O�	��:(�<0t��Zհ���ah����IG^�O���|2���?i�w@�J6kS5Im0��ۃB{:�	���?�-O��lZ�p|U�I�t�Ib����7ut@�J�,S�VΉ#� ��s�O�m���M���xʟ�qQ���^��i$G>�,y��@+,6a�[�L��i>ʠ�'���&�(H���d#��*r�1�FB^ş�������b>5�'HN7mOD3��*C���$��T�̔<&��&#�<���if�O<��'�z6mڡ
b�A N�/�x*�I8�nZ��Mӱ�)�M��ObxD����H?��RJ��܊�aP�)�T�@Ug�@�'8��'r�'���'哒/D��Ñ�4☳��D9(�N ��4,�<����?A���OϮ6=�q��IZ�FJ@9�¤�;BY;2������4Q���Or����iZ�dH9K�<�0��ԩ.C�|�eMV�T��DSWkz���Z���Op��?9��?ܜ!S� L�;�RD,�z����J��?q���?�����EЦ��� �ǟD�Iן��A��k��II��PD8r BY��@��� m����JY�����.C�.����L��by�'�J5b�+�1R�Ѻ��4J�ĺW�'>�@#��@gJ}ÃV1�@1'�'=��'R�'�>����Ezr�Q�{��r+ıe�}�	��M3���W~q���+�.�Z���k	����_�`V�ڟ��ҟ4rG&������?�c�??�>�S�:�0 ��3ɒT(&�`��S�IDy�O�'C�'�fP�mJ�g�X���8NR�I��MS�ς��?����?�����V����bmK�6byk�c~�`�Z�fv�x('�b>q`2LC�g��TkG���	v�ڝ@�My
]gy�&طkm��I)t��'i剜}�d��O
�U>i��˛�~f>��	����Iҟ��i>=�'�6�+����H�b�@�mt~UIRBI#�t��BȦ��?�aR�|��4���kr�l��-�,k��;���*~x��9n��E�t6�o� �	�=O�q���OӮ%�'��d�wI��8���1E�`!Jۜ(8�%k�'_b�'���'t��'x�9еM�X��pȓH��#<PTKu��O��d�O�qo����ڟ���4��]~��gK��Z&��QF��!�����x��fӄ�oz>}�$,Q���'���զ�H�ÕM��y�|bC��S�VI��9\��'��I䟔�	ϟ`�I�iTP�^4�20jM
wE��ԟ�'�6�	��d�O���|�#L(�)�m�N��z��O_~��>y��i6�6MSJ�)���/�>XB�[i�a"b�]^z��쑖D���,O�I�0�?��n�O���1k#o[�`�rP�#��DO�m	���?��?9�S��'\�	��M�F	z��Ņ�+(x�BS+�a|�`�������I��M�I>ͧXh�	�M����+�}���N�~��aa�эj���'��Az��i��Iv�<u��O��o�("���}ʗ��M�������O~���O����O����|D)��u츓�cE�
��{�J�`ڛVA��wb�'�����'�R7=��yu	�k�rlʶ�_���8b-	ߟ�lZ���?Y�S�?��dm�����b5���gN�&{���&���Γy�<hr7��O��hJ>A/O�i�O|�H��R�I��`�E�ݨV *Hb E�Ob��O��Ħ<���iL��*�'12�'f�̡q/�e��}��)�4�=C2��c}r�'FB�|�DŴؐA�Ǎ�<�D�0
�����y�L2�f}Ӟb>ݑ�O���J�h�����ej��q��)S.����O��$�O\�$.ڧ�?����?b@<@(s��d��3�IX��?!�ih恫�O��l�៤%��*i^�	� ˏ[� q��J�D�	��I��ȓ�/I��Γ�?��%Q�.���3� �@�����fD��� '
�{��dZ�k.�d�<ͧ�?y���?���?ٔ�S�Ht�uyF��i��趃֫��ڦ�JI ��8�I�8'?1��>qx8P��78�8ER4��!N�BE˩O��$�O
�O1�TTpr�WT>z��F�-m�
M�WN�+_��7�R]yBh®rl\������Ē�<��f*��c��L:6N(ro��d�O����O��4���;ݛ&	^-7���T J
q8�ASQ*~�P��<=��Fp�0�)�O����Or�D�H���Ⴌ5�l< d��y�y0f�a�r�7$f0f��?}%?]�];oP0�)ug�!5-��J⌃`;�I؟���0������	g��Z�b7ǌ=("Ԉ��v�`�s�'#��'�6��ޯ8��	
�ML>����59{� �၀�C�*����A�}��'�F�s�l�i�2;�6�y���I�_t�UQ&�ʟH^�=��O�G�CsF˓d%��q��RyR�'v��'�k9h�T	���Q�-�R*ŮX�r�'>�ɹ�M��Z��?���?-��=0���#Q��xĈ�A�,�`Й����O�lڣ�M���x�O��$(�Մ��T��97�(�oׇX��1�a��G�jt��W�H���*S�E�M�	�>���Y�8[�^D�&��b�<�	ҟ��I���)�wy"df��B*ƕ2���jEAЖC=�LÒ�I�l�h���OHqm�_�G[���(a��Zb�l�T�C�6���a
����ɩ䞜m�Y~򇖈?�$��'��D��.����˝�o�0�#��m��D�<����?���?���?�/� �Z�+�?$M�u�  D��(�ېI
���`�������	Ɵl$?�����M�;v�jM(���1��H�ԀM�6��a���?	K>ͧ�?���l��8ٴ�y
Qn*\�Q�Ѻ}���j���y�µs����䓸�D�O���ϨM�DI��N|�D�+��c����O��d�Ol˓��eG*|vB�'H����0~�� Kwv��3#��O2��'��'�'��@t��W�⼙&b�=E�P�a�O��y1Mǡ>��7�\z�SCy��O�X����/Yj�Ӟ�V����O0�D�OT��O��}B��l�Aw�DB�,�y���7E(`H9��P��F��1:��I��M��w���#��P�<�L�ڣb��XNaa�'�7��ɦ�Pڴ貄�ܴ��D�c����'~��者� gmN$3#f��7�`Ԫ�� ��<ͧ�?����?9���?�u�3W���[E�U�^H�N���$�Ǧ���g���蟴$?��]���afL	]��`��#�����-Or�Drӄ1$�����ۀO�2^���Hw�1��Q1V�5!�(C5��,�ci*|c�k_�kyb��U����*/Y �Rh�v,B�'�2�'��O�I�Ms��H�<��E۵gqZy��%U04�@��<ag�i��O���'��'�b�2-"�c'/�2s��b�j
�0�v�@�iE���O�M1��/��s�����]T�Z�	{< �&-Ay@��`�j��������러��ݟ����d)31K�-�X"(��L�<Y��?�Ƕi�v���OFxo�|�	f).���lD�*��g(L.@,%���	�@�� T: m�<i��!̞\Zwa׻/��-K B�$����;gz�	Z�	ry�O��'��a̘v%>Ȉ�jM� �rxi��׷e%��'��	��MKq��<���?A*��I;TO��+�ظ���K֜$Q��ĉ�O����O�O�S�IT��+�# 8j��l�S @�$c�n�Xhog~�Oh�q���*��\0F"�p���A��0WϨ�J��?���?�S�'��Ă��ձ�a�'Hn�M{�IM��A;�GU7R(�h�I����4��'�
�N����Չs~�����2����V`�+<~X7�O�#�F�����'x
9�S���?���T���w`߮ZR�RF�_�"%����di���'x��'�'�b�'���V��E���"z:t�%hV�qRdߴ8
\�p���?!����<���yw�����q��wU�U�#d�9��7���U�L<�|����M۞'D��0S�5g�	wR	��=0�'t0�Z����0���|�W����۟H��c�*������s�cJ�� �Iϟ���gy"�lӪ�H���O8�d�O\�Y������e �&8�11fM%�I��������شy�'H�%���x4ؠrHJ*z*���O`8PD�1ڼT"��B1�?����O�h�p*�'aP�*�&ԆI�dɛ �O��d�O��$�O*�}���j�ԓ䯚�'����g�(#�!���j����Q"�����A�?�;K�b���n،Sv&���@�)�VU��?9���?��/���M��O(�
�
N���ḋ(g��Ű"c�.�2�ZU`�!u��'��i>��Iߟ��ҟ��ɇ�<��j�%����hR)I+H�'

6�ȿE���O��D)�9O 8h�^?��1�qEK%P�r��"@EB}��'�"�|���n�c��l馡Ө�8��˜hM6�s@�it��.s���D�O6�O�ʓJ�Z�
V'�]��T�W5Ԭ<����?Q���?I��|J/O.�nZXS�I�:��AJ�*��o[2��Qe�	�Z��,�M���)�>��?���r`A�v��,!��Q�NQ& "���%"�M��O�X%�X�(���.l�xjC�A�ݲQySbY���Oj�D�O��D�Oz��"�Ӧ��191�L�.��1��C='��e�Iӟ��	�M+�f����֦$�,���>%��yF��$qT�V�Ƴ��㛖%z���B�Qr6�<?y�k�]�? Hh(��"C����d	�,� ���ǆ�?�	(�D�<�'�?����?A㇖3r8��9p�"��v�W�?�����R��ck���I��h�Om@��ڀ��{cG�l'�U��O���'G��'zɧ���'S$`򰇇�W=D���I"
qJÃ-�
l���:�����&�Y�O�P�ޔ{PFޱi�,h�jD��I������b>!�'�7�V�/��p��� z"�2�~�"��%?��iU�O=�'c�.��5ateΩ�@)�
�#�'��gFwG�V��Hc��9�q�����T�g
*���*K�R�*Q8OL��?��?���?����i	?I����H޾C���񃓶YX�n�#?�����0��Q�s������k�BW�	�	r'i�7o�NU�Fċ�&+�6�b����<�|�L�M;�'^f�Id��zL�ӧ/ V��A:�'3>8�ǆN��db�|�V��џ��$��2�R���n��LAjH�BӟL�I矸��iy	o�ZD�%��ON�$�Oָ
�H�\�F��-���|�2 ,�I��D�Ѧ��۴*2�'�*lA%F�^-��P�Ru`���''r&eP����V���d쟚d;��v^�E8	�$U/M���QJ@5��@��'���'��'�>��I�2�|���Y (..I�I��_��	�MqǏ%��d�ئu�?ͻ�f�c��%g��+��_�Q�|h�Vۛ��lӂ�lZ9���m�T~RDE�r�����)}��,���G��������o�~�Z��|�S�����	ޟx�I�4i��1u�"@bV�U!����m	Uy"MpӲ�BU��O��$�O,���$	�M�P�
D�R��I�PkЉ:ƌ�'c�i�L�O�O�T�aQ���l�E�vL�I#Șfq�轀�[��P�o?Z��}�	~y�b2b��fݹ:9<1�6�loR�'z��'9�OJ�	�M+�J6�?�3���>��E���� kA���<���i��O4��'��7�����شٔ%B��6]�x�� ��	��AQ�oZ��M��'LR�(/��S4l��I�?��?;�
IX1G���fX�`CKN���ğ,�	������,�IK��TP�
dRw]�D��"ś���Z-O��dB٦5��d6"��i�'�&�
E��%
�5���	`���Au)2�$ۦm�۴�zq���MK�'�i�P�((K�"]�~j�-bW��^> �)d�B���|rY���	����쟈�B��	",	��Y�-DB��I��,�'�6��r�����O^�d�H�I��`hB��-<���z#�W�D�O�ɖ'i2�i=�ʧk^d�jٗgv<�ygfڮG��慔�}�� �c�s~�O�V���'f��'���1�^!rx�݃ea �QR`p@�'A��'���O �ɭ�M�v�G*a�0�Ȇ,�/Y�)��5rz�.O$xmZN�Y�	��M�DDK��� �%<"�SC��/iF���'��	���iC�	��l���O�']BU��%���,9�ƀi(m�����OX�$�O��O��ħ|�2G#F5S6�ې17�ճ�@��楓(f���l��u��y�lX�?T�a�� 'e�&���G�<x��7��ꦁ��ny���#�4w��5O���ɑ�B1�'�X�*�T�I'<O�	���3�?ao5�D�<�'�?!��q�2ap˅�,"�����X��?A��?����D���Q(��şh��۟0���ٞ5e��iSa�&?�^,5�R��0��ɖ�MK�i��ON]0�Ǖ%k�R��vNRwbV�x���R��\�}�X{�,�{�S|��,��4"$a�*^ʘ�dN[�&�HK4C����	ʟ�	�`F���'����LػQ����f#�4_j�!�'�7�%��I��Ms��w�L:өHf�8���Vo$r�'=r�'B�Ħ��期D �������5f�b�E'!�>e��j��}3*�O2��|���?����?���: i#Ȓ��l8�*�fh+O�nZ�Z���؟���K�s�dKD�R1Pب��b��4���R֣�<��D�O���7����}��L�%�4X�0�cs�Z��fNd�v�@ �Cī��T$�8�'⅑p�ˑU�@�HO)k���g�'2�'�b����P���4m����F�P	N�K�lE8a��3�ZA̓4���dd}r�'���'����f�:��Z�h¤9zT�BAݠp��=O��dn�Kx|��y�O�7�,l&0�	�+�� ����/��yr�'�B�'��'w��I�h��ꂣM�6��l�/ ]p���O6��[¦qp��Ny�#qӲ�Ol� ��8xhL5��MxɴĈЃFp≖�M��ig��)ZʛF7O��D�0E�zPp�˟ �)�흮v���(ą�?)��8�d�<!��?��?���B�u��
_2���{�'
��?9���Y̦��U���\��Ο�O4\P v�֒x���	!8%�x��OH�'EB�'�ɧ��ޠMp؅�smH�y���a�fF�qG���G�f�\6�Ay�O*p$����<"~����&�dA�<o �5����?y���?��S�'��Dۦ�I��.|r�@��()�	�S���*i�	˟Zٴ��'�X꓃?�5����Y�B��txdxPRoT0�?9��'��8ܴ��Ā%"o����O�In�$�֊��E�ē�F²Z��Ky�'���'n��'��^>e"�A��H�fY�5'�xb��1��6�M�7̝��?���?�L~�m0��w���H��J�m���0��j�����'K��|���n�P��&=O� ��ŬS�+CC�4q�r�[V=OR�z3e��~�|W����۟`�F�N5��Y��Y�|;�E�5"�ȟ ��֟���Zy�Dz�ֵ�Ƭ�O����O�@㵍̷���iU���#�b��a,��&��������۴�'kȹ�W���
y�Ԍ
}��K�O��)N�pN�����?IF�Oְ��!��O�\|Y�I�5�ݱF�O ���O��$�O��}j���"�8RcX�J�4|�J��m4�5i�� {��%�o��ɂ�M+��w������ʬfr0��ʙ��d$��'��6M�Ʀ�z޴-�:�ߴ���3#���'9���+vL�D���p�%J�r�;!+�$�<�'�?Q���?���?�kB�c��P���/:�Պ�<����c�� ?q���Og�`2Ё�6Q�Z�{�[O���S�$�>I��?IM>�|b�,��\	���VL}��k�-O�X���4���Z��~yR�'��'�削������G�Kp4B��W�-�r�����h��䟈�i>�'��6MMw8^�^/ �$CB�&0}�L*PJզn)��d��9�?��X�������� �^��+[�:�T�d�M�;��sRZ���'T�|9b��w
M~�;)���哅@��N�d�̓�?	���?���?�����O!B���� 2j00j��|Pf̐C�'�b�'�7H1s���O�l�x�ɵj������I�O��z�tU'���ϟ��spm�I~b�Z�2����4�l@����e-���2Il?aN>�,O�t��D�Ob�$Vͦ<8En���Q��K�uQ\�d�O\�@`��!M?fv�	��O���厈H�D�"�3%��=z�ODD�'�R�'Rɧ�	�=\`M����1���3c\##F"���E��b�07�fy�O�6��������4%һ���A�`�Ö�?���?���?ͧ*��@����D���=�&�K?���ŏ��4�3�n�.������ �ٴ���|"�S���ڴ3za �iR3�h�P���#[Ფ�iKr�;��f��8�T��s����~�ǦY�0ZƁ{a�U�]�fvCn���D�Ob�D�O��$�O>�D�|�+�&`[�xoُB/��#J2Q�o�/b2�'t�^>��	���2���ǡCD�x�b�D�T���`Q� ��f}�@��<�|�2L���Mc�'�V��&�@�R���@
��q*6��'�
�!��QܟL��'��zy�O�¦���a�)�0v����m�-2R�D�OH��^$B� ��ei�(������5S�LqW�\$c*P�����k��x$���	���d����:޴�?�*O��kёF����n˶P64A@��(��ݭ߬�j�3�S%����؟p�4�Đ �J��%Z��R�g^�������IȟpG���'!@����;@��ek]�.Hh�'��7O<A�h˓��6�4�V�Y�A�gځK��9@8鱇8O�AmZ��MS�ta�Q��4���9K	|��'Y����G"Y<Zcҵ3�*��]�6�z�;��<�'�?���?��?�Wک��Hۆ��#�;U� ��$�ɦ]���|������L'?�I+q�;�h�3fr����ř��*�O����OؒO1���QL9��+b�('��e�V�ܑ,446�&?�WaF��IB��qy�Ҡb�ܘ�d) �Q�(�Q �N?
?��'���'�O��	3�M;q�ܱ�ɚGE$�R���R���^����ɫ�M��RH�>g�i�T6-M�I�����,�=�b("P��1�"�X�n�X~���+����Se��O��.�cn��� j�L4�֏�6�y��'�2�'���'~r���$4٘�%J�'��2�l\�T�
�$�O������q���ay��s� �O�qQPDS�:T��,2)ØE1�MXW�I2�Mc3���4Ś+"֛f���b��<6źy[��ݶ�>X��Nغ��k��'��i'�����D�'���'���bf��.%*(ȋ�NāmM��G�'DQ�<��4_�53��?	���i +8Nzicg�
+&2���I�������pݴ\ۉ��i�ny\Xb���b��eq�Ǵ8�N��'�?y� �����S3�R�t�ɀ}�����`�S���R	vd�����	�\�)�Sfy�v��yj�5T?<a3R�I5�F�JUC�#h�|���O�HoZi� ���ܟ�k�	�8XC �*�Id*���	��HlO~2$Ζ������Xp��p'h�_eX�+����(?��<i��?����?��?!*����1-^=sǦ�\v���S��ݦ#�fٟ�	�x'?��8�M�;Q4���&.F�@��b�IR�����?1I>�|�g���MS�'ǲ0xS�$ad\
�۸-�X]��'T�@&a�d?�L>�(O6�d�OʽQ�e J���'c\�_��5���O����O~��<��ip����'���'����!
QpDD:"��(�$�<�	���D�O��$��ߣD��s��ݝs4jsA"�:uX�ɻ;�h�#oM�ţM~JǾ���Iy�<�C��44z���;:�j��I��D�Iğ��	R��y��B*���i��ŉ.�:�JW�g�r�`�=�����ش���y���fZ�31O�)�fq�Sg���yb�'3��'�i����Y��Xфן|�(��,X�`8��@eY(��2�'�D�<�'�?!��?���?��e�-}��@�B ܋.\���c! ��D�Ҧ��a�e�P����@%?牓=��	�� 
�X(xZ��F+7ܐ�O����OL�O1�*��� �xs�N/�rQ�R@x'L����|���D,��%��'b.WhG�i_B�AV-�;��@�4�'���'�����T\�X;ڴy�`Γ���u�w����@LE�6bX�͓@����d�m}��'�b�'W�9�F�T;�ar�kT7-�D �_�Xכ����{ry�Q>U�]:.]E�5���V�<�B(�� ��	ğ$��՟��I���u�'�Hg�/ BH��D`i���?��K���K�����'uN6�3��ҙE�2��V"͌|. ����<!�.�O���O��FT�7�0?�tf�W�N�E 0�6�k�M��µh���$��'(��'��'9Zx��l��|���-�8mN����'�"R�0`ܴtA���?����i�.K�,�@eӬ:�jdr�m���I,����Op7MB�|�B�B(rT��/G*AV9˅a+TP�`3��#K�Z���G�ϟ� U�|���<\lHAMďr\^��U	��y��'�B�'����T����4Rb �� �&-�%;�gS�aKh��Wب��$�ߦ�?Y�W�p!�4DhL����8{����BL˂MD��B��i>�7-.��7M4?��l�8t����)�MN'Y,�#���SQ"���o�;�y�R�@�������Ο��Iџ@�O����̐@]n�Pt�P�#�ە�p� � ��O$���O����DFզ��<���{�),.�R�Ǒ�#�V�����MC��|J~چ`F��M�'� |b�4	$t��O��:A���'N`��`aB�����|Q�������W�\ό��b�n�4Zǆ�럤�����Idy��~���b5O ���O0<�B�)O�����B�4M:!E"�ɭ���O���#���s���Q�~$���' �}��	�8�HĐ�	I�9�|�0볟��ɏ �*٨F,�0�r�>C$�p��۟L����l��Y�O>�)�9*QrD�##�>z��
Bg��b�nӔ�QUo�<!�i�O�.N#Z�J8Q��
�)�F̰@�L!���O��$�OJe�q�"�3������?��R��\�lx`i�\h(P6	�\�	Vy2�' ��'|��'W�5��f�19]�x�$��F�Ɉ�M��ၨ�?���?)��d��1rAK��W�6\�!nY>I���"\�<�	՟@&�b>��A��c��<Cd�W5�]��E��� o�����J���\h�'��'N�`J��sg"Χ��)�j�F�������ßH�i>��'M�7�@��$����G�F\��r1*��V�,%�ls���D]}��'m��'"d�fh��5�����}�2p	$��:g����ʠ#P�Q>U�]�`�4d9�!�f
<��+����	֟x��ПL������IT��;�M�e�ԃ M�D�%J�.R�����?i���D�3w���M�O>�SN��d~̩� ��4�j"(P�>�'��7����XAnpnZf~ҧ�{��<R�.��1���A&h�T�,�ái��H3�|�Y���0���p�� 葯�zF=Rk����JyҌaӦ�8f��O^��O�']�݃�d��B4�����P(a�e�'�f�1��k��<%��6�Jui�I��6��XR" !D�\Hc/CE�$� w��O~�O��i�ɚ��'���p�*O	qh����2�`��W�'���'5b���Ow�I��M�F�����'��=_��yIt�ϳ!���(O0nb�Y��ɀ�M�`�Ɣ&��t�SKT:P�TYǘ�-t��D{ӐT3�w���&ڊusCK����O���)'��L�����Є$<lp�'�	Пx�	�l����h�	S��%�a
�ƃm1T��f�Na� 6�_9d���d�O��3�9O��mz���ER�ur&N%p�8���M�c�i��O1�*��q��	&"��1W��Ք���h֍6��s�H�y��'�f�$�����4�'^�葔i.'�XT�U�"L�.m��'�2�'�X� �޴
��b��?������S8I��xz��K�_�T�ۈR��>�1�i2�7m�W��*���b횇FzmZ#۵H������e��#���|:u��O�s��1-�����uv�mh ���*�!����?���?9��h����T�����3���dV$2��$U�!��A՟����M[��wL��b���Rin�YD�@6䀐�'�7-I�Y�ݴnc�H��4��DZ, �P�I�'~U.�*��۠
����a�Kj{�Y��+�d�<����?���?i��?!%`��FO��cԋ��/�ݱ�1�������ώ䟠�	��&?����C�<%G��R�8��P�ٛ|�60�O��n)�Mk��x���oRs�<�4������^)X�SC*����	k�z�x�'Ov�'�ܔ'��T(���7I�,܉s�ʄZ��]�A�'���'�B����^���(pvT�IqPD2Di��Ȳ��
=r�ɭ�M���ɰ>)��i��6�����dD�*�A{����|���	G�gT��lZK~�� s"�/B��Oh7O�-c\�pk�H� �F�PŭB �y��'�r�'��'���A�jT�óM�I�VD#&����?Q�i�X��ȟ�=oZZ��?A�ͣ��Jk�9B��� '��L<q��iP 6=���P1&sӤ�}�$���ŗIg0��←�W�|����P���/������O��$�O��d<[� =9�f#}�l�zu�ۤA�����O�ʓN�$R��?Q��?�.�L��
�)�6}��m.I��:�����(O~�D}ӤQ%��g�? � 3�H\>;󞈱cT ���B'2� �"H��9����|� ��O�|M>�w̏�,~҅��㕶r�����t<���i!�0Z���,�L�fD(��xy�*��I�M��rf�>���i㒹a��٫���`Eb2Tpq06y�~0oZ��p�nZs~��Y�����S2�I5,g�}�䢁 b5$)��%��D�8��vy��'�\��t�ЏcW��(#�P�\o���Al�.�y`l�O��D�O��?Y����ŢOè��5�
:l�0JP��.��!x�v�%�b>�獑禝�,��X@�2an�aK6]�m�5�6!�(��f�O�őL>�.O&˓nh��6#O$a�Qc�6\ą��I��M�T5��$�O�A�Qf�j>b ̘79j-B;�I+��dEݦE"�4b܉'@�8y�!]�#��q�@��|����OZ�3Pa�;� �A!�)��?�!�O�;r'��YY0f\Y�)��@�!��8�4��rFl	� hbfƄ/E����ߦ���ܟ���;�MÊ�wkļD�qV��B�Ɯp�d��<���i�6���S�������'���:o��?����@�z���+�|��Ē�c�'��X�'?�D$���Fi⇭�&��lI�O��o�~���'H�i=w�����/��1��:��,�'�6��7�OG�)��\%6�:�
_�n�����-D���:�Ϛ����'�MP�� �����|�[���SNC�`0��`��jj��tK���T�Iʟp�I۟��ay�oӺ�94��O�� �ĩ|��8����νR��Ol�n�a�����8�O(ml��M�W�i�\�F- 1HR(�aj��Aj�pbBߘdO������C�ɠ���F��ߍ��46��J�y�g/|�H������I���I�L��' �,~�����G+�.�	D&H��?����?�i��!�O�"Fo�(�OL��� »BH䰑�C��n�E3Ն�X≊�M�����G��F��� ���H�E��p�b!���3H�I���E�Jyb�'$"�'2�� ��}I�.&<~PA1���#(B�'��I�M��T
�?���?�+���
�b���hJ\.��Ib9O6��ZH}�loӰoZ&��S�4�R�CI���HĊB̢����CHG.9�j,D�`aX��S-l���Es�I#*(�1�ǃz�.�ȆA�d�BT��ܟ��˟��)�Oy�Lc��rE�%6�~Ҷ�\�l�$AA�!�V~��O��n�e��Ο�+�O���­ :���P�L�7�Iʔ�ޒ8����O��˅GnӠ�&��ԓC$�?��'��)��n1gl2�Rq��$`���'����`�	���	ޟ���F���-����@�"���K�%oM�7�/G����Ol�� ���OB�lz�)�DFA�	�xLi���8Vhx0e��?�ش(�ɧ�b�",	ܴ�y�81wuдOݏh��r����y2��!M�����-F�'���џ���2���k dׇkW��D�I{W�|�	��,�	�D�'��6m�!�*���O���N� ��0dBCF`�q�s���Ov���N}�'���|�i�-���D���ژ����?	4���"/j��]'?eѥ�O<�d�$��Y2��&9"\)	Z�^]���?A��?a���h��.׃:�j�J"���D(a�WȜ �j�d�������C�<��(�M�O>!�Ӽ���L������V�p�_�<����?I���ڴ���5+���O\v|���0F�&a3H�$|}:T�|2R�P�Iџ���Ο��Iß��f� 8�n�B"�*M�pa�q~yr�a����K�O����O����D]����	gO�!ݼ����@�y�'zd6̓ͦ��I<�|2�
�7ఱ���4��.=�P$h�YQ~�iZ�]f@��	�"��'d��;�<X�5�	Q
*���	O���Đ֦�s��Ɵ��(&�Y9j�940)�b�ΟZڴ��'����?Q��?᧥#�zz��
>��P�ҥ�#Ml�(�4���K�&��m	�O��O�g�֦0wt�z֙C�-Qu 
��yb�'/R�[�6��yZ�ϛ���ҥ�'�b�'� 7�L�h��,�M�M>q�Dl���x�� 4'�h�ğ.���?i��|"u�R��MK�O9�򣚈B<ܑ�d��S�O<���'y�'��	^��E��I�3b����#g�!4H�Fx��`�vŘ6	�O���O�ʧ���ZS.ױHk����]��'���m�ve�Ґ'��u��Ӎ�%;�nHA�ڥ8���kP'	k��u�IƮ��4�������@�O�w◆9.��M;?h�����O<��O���O1�Jʓ%���]9rDB��`gV<}��,�u�
^�t�*�'rb�m��⟰J�O��Dܗ'xZ���4{���{���*A����O�ܙ�k��v��aM�?��'�^��U�Ѱj� �b�
G1�9�'���\�	��@����0��E���*���Z�� �E�N��"#��¶6�K�p
����O|�1�9O0Xmz޹�Ӊ�*i�bl2KC�{�� �$J���MS3�i��O1��I	��l���2`[�T�F� 6�X��@�s��I_��xhS�'�'�t�����'�|X@�h�n5�pIшDfniXG�'q2�'��T��Hܴu��P����?A�5H�5�"���U���^v����b,�<���M㗐x
� �H���,�D�B�ۈc�Y
�����E�C/b!(��T�(�S�b)�����Mn\V͛#B@� E���֎*D�8Y��N�t�����ƃ�8�x��d�П`8�4�t|����?!òi�O��/��	�c
+hTД��'E2�D�Op�d�O�Ł�'k����%��ɱ?�xV��XX����
_ �t!S0�PY�IayB��0|�@�pc��9X z���TAj��R��F�6Sm�' "�i��E��!��^�r'Pi��	�;�5�'��7ͅզ5)L<�|�qMR�R�j��C^fu��A
S�Huz �����MTx�j��d,�Op�yO>\A����쭲� �n�����?!���?���|R,O"mڈz�\����6��<*�nݮY<��� ��z,: �	*�M�"��>I��i��7Mۦ�*�.1�Z)�#ɕ�2�m�v�U���mA~��W�L����V��O��K��"�*���-O�.�bE��y�'���'R�'�B��ܛ&X��W�#c������]'��d�O��¦���d>!�I��McN>Iইom�`�DO	(�6,�SIֈo�'�r���4��1���4pSO΅G����ٓk�ތ�@d�Y�h%�wmF0El�	�j�75�����s�Nt�@�Z����Nt��y��o�|�X�J%*GZ0�X_�"D�6H�]@�u*Q��<d�|ӤO_��zE�X�������,&a�$Q�M�Ih\x���
�J	��b��j���'��i�.��p蔰O+2(�F�ӭp�Ph16i��fY[t���y�V����}����E�^�;dD9eB�&8���"�b� ` o��I�������X}8u��@��d~tC���8^�~V
� �#D��>lvPpA�K�y�H���K٠zְ=j��	�+H$s�l2�����O���d���� �r�J$#C�o����/LC�i&�t�	��+����/v�c�������*�T�d����*ߠ<n�� �I!Y U�	��8���<�����i��b���oit�	��a-Rm�)o���O�X��J�r�1O���}3���8yz� /ŝq����F�iqg�'Ab�'���O��x��76*`���YF6�=��b:/�&6-M !Y�6���<�PE�jr�a6�F�n&j!����M����?q�'�4�,O��'�?1�'gpY�$�CVU�E�	&�:!��(�ɤEPz��O|*��?���k�I�RP�B+@(�G�>�*����iZ���e������O��Ok삝9�ܥCg��7|���
QiF�a@��*U
���Ihy2�'�B�'���>Q�j=!�	�wm��D!��)�)�֡��$�<Y����?Q��ty�<����0�T��ӡ��l���srH7���?���?+O��j���|�.�i[V-j䀒 ;�$�� F�є'|��'���;4��Ֆ6l��#��v�@�"�I���ҟ<�	ڟH�'�I�P �~��6�-c����t�Xk�l����YG�i���|��'�2��)d*qO @�h��w�� ɢNXe�IW�ip��'X�&������$�O��IO�vN�z f��q�0�C�E�Y"�$�d���x�� �I�����\�H��"p��F*�6ɘ�Mc+OԽsAI��m�	ڟ����?�ۮOklvvlV�z}�,��Le���ش�?����8���i��S8����PF�A�ƊC2Y��a����7M�O��d�O.���~}�]�X�a��1cw6���z80)�)�MK�GY��?�I>).�����3V�KnH&����҈�������M���?�\�0\X4]�Ȕ'9��Op!�!MI'a���u�܆3�I�0���!Z_(�O"�d�O^���42\�GK��^�k�(��v�:�n�˟H1���9���<�������Ěs��x�UA�I;xA�#�}��	�'R�'�[��B���Q�"Pyq�^�T�����I���O�˓�?yL>Q��?q���'qޙ�,�~��	!�Пe�0�H>����?�����$U<Q~F�ϧD8̙�e� 9d����H!=0|o�xy��'��'��'�����O����$��Et1�`JJZ��S�Z�(��џ4��ry2���F���9�VFD4 �>>֠�����IH�qy�O���~� EO8|�~�Bf�\��@�u�����ɟ��'l��"I<���OH���Dh@Ԡ> �"l�0�Ţ{k��j@�x�Q�8�	韬$?�i�-�Bͺh���`Ėh+P���B�f�D��i��맀?!�'��I�����Ѐ��f��ʘ%G"6͵<9���?Q��t���4a<| `U%H'mH���rA�!��4l--����ܴ�?���?��'������8I%D�W��Y&>h��N
��7��O��D�OޓO��<���;�\�Iժo���Z=��C�ia��'�b-T^��O���O4��,pl �F�NyhR�AQ���7-�OڒO^���y��'5��'-p; g 
D!��;���3\�4`���$�"Xf��&��S�'���%=_D8�D,U/r�+�-��L�,O��d�<����?������o�4��3�O�u�"m�A�,��XK^J�	�8�I|�IlyZw� ����u�t����9��T��4�?)*O��$�O����<qfߞ~�	X� ,`X��)wo
h����ȟ���l��Hy�O���b���Ι8���PG� \]���?)���?�*O�p�5CK�+b�J�{:pĊu�A"تz�08�ܴ�?YO>y.O�i�O�O(虚�.��p�\�r�ڀl�zH�ܴ�?�����0>���%>�	�?�8� ^��ƃ�Ha�C�"ҸXd�xRW� �	���&?�i�1��
��8�=!1������i�>���a=��H���?�-O&�	�<��Fh5��aV����/LaZ-l�ȟP���<R�r�3�)�ӷ��)���#I�Q�X��6M�7f2l���O����O���<�O��i�%ڤ$�,R&eZ�&�T!�e�j�đ�S�� :51O?���e�7h@(�!��	byv#����Ms���B$/��S��>�Ԯ@O�"��r��"gBDeЀ�$71ONLc@`[짌?��'��`��P�*Âa����f��5��4�?������
U��d�u�\i{��8�ٰ�g�,,����'����A"Y�Ø'��Q�����w�~p�e��x�ܠR�J
�|���Ggy��'/����O���W� td��N�4yĮ߹>�������p�����@���ܕ'uj� ��>��m8���0�y��s��>����?AL>�/O�yC ��O�m2��Y3�J3e��,Yn\`W��A}r�'}"�'�r=�,�I|���&{z��@V`�+RO��I4!�%4�f�'��'i�
f��!��h�	�6Ti���ԠVJ�:���E�+����'�RY�t��d��'�?������X�&rB�bF�»y��#LC}�'剷W�r��	C�X���"C�BcF�jp��ŠR@}��'�hL���'���'�Ol�iݡiu�A6.f���L�2�&����,���Ot�����Io1O���`y���r�8�J��R�s�)8`�i�>���Ev�H���O���f�&��s����n������S34º�Z�Ao�V�RQ��O��d�O2������g~�k�(o�H�:A�;,�c�C� ��6��O �$�O�<�DOX�i>y�I^?��o�)��=�ni������	Pye�+�`��<���?	��LX���� �<R�T@���T-�|s"�i�B��
P�ꓢ��O���?�1R`�IP�P��L=Kq����y�'B^|��'���'��'�"]�|��F�iW���@CV85���
�kU"�n���O���?�+O����O��dO.m����6C�.ܐ�v/��,F>O4�$�O��D�O��d�<	�O"vH�@9]x�ѡWɖ'*�0�"��:қ&[����Sy2�'�B�'�1{��5Ƈ�X��@�O>_P� �M��M���?����?*O��'Bo����5V�	TА#sb�U:���N��M3����$�Or���O`4��3ON�d����O�(	^
X��O���)�Ct�l���O�ʓ��\��Z?%�inZ�?�S�ò#QB� !lW�,X��v�	5����Op�$�O�t"'4Onʓ�?��OGȸ�sNG�.r���c�*[�*]�ܴ��D�9��n�埜�	՟��=����}�u�I�<Ud�/T����v�i���'�R-��'��'�q����r�:G��U�C�@y^��6�iR4�{ �h���$�O��D��T�'��ɘU&q���ҟ1��9�l�(8��hJ�4���ϓ�?	-O��?��I}�\ �'�2Z:�h�kզz?fLJݴ�?	��?YAO��5���ry��'x�D�8�5��)��Q�	�0�ȼm�ğ��	�� x��p��'�?����?ٰ�3\�Fȳ��@�O�i�Fj�fc���'F�-ap��>!.ON���<)����i|	���<pr��zF��n}�%���y��'oR�'2�'��	�%-����B�m6����&����BP�0�
�'v����X�'wb�'�r�Tb'.  ^�H��MS X�ı�	R�<�(O���O"�� �r����|���4�H�,�U"Ĺ�dP��'"P��I�d�I�7���0r��dM��$����<-O���On�$�O����<�1mЄ7��Sӟ�䮖�*F�@����;'�@2���M�����$�O��D�O6T{16O&�'��l��AH��I��,9~>�r�4�?y����$ָFYf��OR�'���L�2K�Ԁ�)@�/?@l�	F$^����?���?����<�,��d�?`D��*�( �u!��z����`ӊ�$HH�i��'���O�z�Ӻ�`�ـNk�L;�㏀K�����E�=��П��m~�����/�Ӻx��!Q�����`ԡH��6�]o��)nZ�����|�������<�A�׾��͋�d[�}C��zu��s��F�͵�y��'��	C�'�?1a� �$�6I��o�>Bx-ڑH�(F���'���'�藪�>�-O��D������=I��D�9"B1�f����<!4���<�OB�'���e�$(��h]!7��G��5n�R6��O�K�f}r_���	zyb��5f���f5����u4A!�Aú�M3�c�~}Γ��d�O����O��y��[t⎕b� ,`�O�#Ft�D�ձ9$�	yyb�'`�I�������9�&D)��X�%	M��:��$- �d�8�	şl��柨���T�'�hy By>��&薨
����oðrpl �v���?+O�d�O:���� �ѭ2�����Y�A����E�WI�ƕn������՟��xy�9G�r��?�1_v��soH�,�"������p�n��@�'���'���(�y"�'��ąG�~5CWF7)NH*bT�˛��'�2U�P0'悙��i�O����<!2��J�~b������X�P�Br}��'_r�'�@��'M�U�����6�զ��"�&�csL��9. 4m�Fy��cI�7�O$���O��)�u}Zwx�!�`F�-R<蓧��9���B�4�?��^�������O.`Ȋp���Rsp	S׀�'.j�yٴ]<��"b�i�r�'��O�J���DQD�? r��g� D�f��a�	�B�(�iwX%؛'<"P����hby`���; F�IѮR�=L`0��iP�'-� H��0OP�D�O^�	*s*�AЎ�2^� �CuNf6m%��ݏ+Þ�$>��I��,��6 |�x��޶)T���!K2�j�l��<3��
��ē�?q�����Cc�7Oښhg�#�ŀaA}R��y�\�T��ן��Iry�L��;�<pTB�7D>��7A���S1�,���O��D:���O��d
�;����N�!V�I��!��.������O���?����?�.O�}��j�|�D#N� �ذ"E�hR���� _}R�'HҞ|B�'I"������T ��ST�3� %�ŉ�#i���ݟ����L����٣��'Tle���S!J�h� H٧\�ܭ0�iRX�����@���}m<��o��� r|�RU�� l�@����H����'�T�0��@���'�?��'(r����m�?��D
E�*L�������?���1r�iϓ�䓽�$	�*�b�9Pŕl������8�M�/Ov�"V���}Ӭ���d��je�'���cתl�l8IE$]�D�HHܴ�?Q��,y"���䓧�i���Y��PfΑb�I%*PJ��n�j�������	ɟ �I�?9O<i�v��`S�·CU�@Ia�F\��a��i�
�;�'-�'m���N5 ���EK�2���Ʀ��ʥm�ҟl��ޟӐP���?!��~
(qXHp
�J:	�����' ӈyb�'V��'�0(Aum�9��P�F��iq"�'�Ӧ�d��^�0%$�X����$&���1Ndy�`dǆ"�*q�� �;���JS�N>A��?1������=jyv�#�ɂF�ҡ�6����2��a��ON�D:�d�OL��Bl�P�W� �԰;�
M�[�r���c�Op��?A���?�-O���.�|
����N0G��4o�1;�H~}"�'g��|2�'f�CX�Xh2��f1z<چ�ڴR҅Q\�[E��>���?Q�����Gt�'>���	�
u�pA���6L| ��ӊ�MS�����?Y�ĸ͓��ɍB�:�"��;@��ZP-քm�6��O����<��h!$��O���O�:���������F���a0��#F%��O"�d�]�`�D1�d�?��u��!C��dA�Za�dJSo`���=-��Rƶi�꧉?��'o��9)��!떬1a0E�b_<�>����O2��^��6+տoT �JgB�"oڥh7�i�*���jӄ���O����"Q%��S�Yb�7a�.����}�,�ѨOz��9�)�џ@��#C7%y��0�
<V��e��R��Ms��?���LD�f�x�O���&4�䦘>K��;ţ����LoH��ӉO�b�'"��)(�#W�J'ø�^�FȰ6M�O
���d�w�i>Gy£܋�ⱙ@�Ȅm�04�WM ���?�+O2�d�O��.Z0���T|*�(Q���_�X��� 3���QM<���hO�I�>�}�gF�'/ARC �[,=�6�O\ʓ�?Q�����O���7�?!��b�F�p�HSv��PEm�L���O��$ ���O��U�����[�V�I��@�Y,����&���O��D�O4�v*��Ē�T��9
��!��o�`�ȁӓ�6��OޓO8��:�C���G�g��a��:-ptm�џ��yҧ\�W������쟂Q�a!h�P��w[5SBًp$�^�I�����R��"<Q�Os.���]]����й$���:�4��DH6p�0(m����)�O��	\R~,U=LG~4��
+;D���f[��M���?���_i�'3q����V>@�R��'#���%�i7���Jc�*���Ob��쟲d�'N剁}Nr}8 �S�=W�
"���=��4q�~]��?�/O8�?��	�yv0�6�]t�	��)�`
�qڴ�?I���?!���FM�IHyR�'���Ý)H YJ�B ���2������'k"�'�������O����O� �&Eģ(]�5p҅0+�<t�fF榍��.�0�Odʓ�?�,Of���,�h�
A'Ɛ৥�;c�F��BZ��U�l��I՟��I՟p�	py��ïu8@�b�o�â4�d!�1�iSl�>9.O��d�<1���?��]�؊T*ŪC���*EC��v�@�<y,OT�d�Ob�ı<�țe}�I�#�:�k�f�n&t��NOb��T���	iy��'���'�Z�O� ��!�"JT'ͣD �a�i ��'���'��ɜ]�����n���*�X�/@r����0g	�[夤c�i*r_����؟����\�Im�ܴk���
J�: �5��H5KP�lZƟ��Iy"������'�?	���23�[�jS�\~Yb�fȿ:%��ҟ��I���j��d�����]�@&��G�,��$�t�Q����A�'�j�Z��j����O.����Qէu�t#H=�h6	�b`��̮�M���?Q1j_�<�M>َ���X~��1	f���z@Ƽa�F��M��{6�'d��'�� �>y+O����Շq"���GĆ�w�t�C��T����soa���	ny����O}p)$�T�4=6 9�dݦ��@y2n|-���i�O�ӥ_��(��?K��y��K'.	@��yr�[!������O���S�v��qz!�R,�v�0R��:n$F�mZ� ѣ�0���<)���$�Ok� &T������];R�ʒNގA�@T�؃z�d�'�"�'l�Y��q�٥d$L�A�]6x^�ـ�̊�+���Q�O�˓�?�+O����O|�d�<gO���ga�i�]c�A��q\IQT0OT���O��O��d�<	��U#Q�ɓ1=�i�3�ع\'
�[F�!N�&W�`�	Ny2�'}��'cl�p�'v��٢Α!Q|D��c�!���铯g�����O����O��&���qGQ?��I:Gn�QuH�/	��@P
�7�8�ٴ�?a-O����O���J<�O`���|��-�7��"��)�iPR�'��	�~|�k����$�Ox���3ú,ـi]�:�*u���J����'�B�'W�����y�^>�Ic��iݤ��Y�ǍO�)���Q��ަ��'u8}�o�p�D�O����P�էu'F�z���rK�IU�e �/��MK��?��k�<����?a���O�^(`�D��`xµh����q��ŋ۴A�I#�i "�'�2�O�����D�&uؙ�ڤ":��	$��\P�8��8;O��Oʓ��Ov��6u͜�\85*aB�u(�q�b |���d�ON��:H\���'��IƟ���&2��Ӷ%���8Tl�>:4LoƟt�'�M˘��)�Oh���?9B��&��qP���0Ӗ�C5Cwӈ�Iu��ʓ��S��(%� ���'���ۤ�Q:p2�9C�� ���U�'�2�'U�T���0G>Ԕ����'W����7'ƄZ*� �O<1���?�����'R��R�KҚ��К���S���Z�%���'���'���'+��O�%_�KR�g�Ҥ�e������ ��6��O����O"�O���<�O̦�锉E��8�^2N+����f�>y��?y������>��'>ib�d�T�r���{�F�I1���M3�����?9��~+΅�>qA ���`4M5&۴�L��a�IƟ��'\z�) �!�)�O��	��i��ha��2zX��jZ/TFʡ'�������c��6�����L�{�qk�+�]>j��eF��Mc.O�Ck�]�������6��'��)��Fٻ^��\PbJQ3ޙ@ܴ�?q�z#��ExB�)���I��h]�T34�IѪ�v���	�7��O���O>�I�b�Ο��k�>-���B�Y&�q���MSV��G��������s8N-���*�q0�nV-GP�l�������<A����M�$�'��d)R�ƅip���t	��M/>�lEx�,8���O���OJ���ǜ%1���	6��?�B�Sȑ����I�����O<ͧ�?1���In~��P�74�x��`-~�VqjQ�<���?���?a�j 2�Ƀ�@)�y�e�<xճ�l �?���?����?!K>���~r-L�z7�5�5��;�:��V(׀�M� �F~��'[��'��Ʌ2�p���O.���R��V(CCK������O��d�O��O��D�O�̃�Y�|C� �E�^��&�J�G&��B�>��?����ץ5��T%>5HTm�7������("�� p5C4�M�����?���|�$�>�3蕉V�*9��c�
DA�ٚ%NU٦��	����	��,�hP�P��ߟ���?�2�$�!6����ca/d��ًBH�6�ē�?�/O�L�S�i���抜� ^��*��.{�pa�bg�^�G��۱�iav�'�?��a8�I	*38�)
�V (���D�J�O��j�c3���?O��B��?Q-�B/ �$�}ɶ�ic�A�g�'	b�'���O��@�$�N�,K䀀���=� ��G(�m�>�{Fx����'_`��%�*%������5Oc��P�e�$�$�O��d��Z�$�8��Ɵ���:�����(/TD	R`IE�{K���>a�N�]��?���?V�@�
q��Y8�`�z�n��&9�6�'J�'N2�$�OV�D>��ư�a�BG�[�̥j�NӔD�RP�R\�PEg1�	��I�� �'�,!J��פ}{���'�-c�!zU��0t�zc��	|�؟��\� ��冘aCR�#�d�F�u�&��ԟ��	џ��'k,Yu(t>�c��W���uK&�Eo�*$YƋ3�d�OȓO��D�O�]��X����'
s����e�e�T��a�>���?������Ѷ�`A$>鉢	�)���3�IH�	)� ��M������?���� �>�����g��ˀ�T<>�w�_��a��Ƛ�'Ɗ�J`&+���O��ɓ�*r<HD��{�hH2P�
)G�>&���	՟�@��,����e� W\����Tt��t�w	���M,O�@Q��L��Qy��b�$�>��'�6a#�
%(��wEHP<�cڴ�?����4�Ex����=Q�t� �ڹC�L����>�M�1LC�6���'���' �T	#�I�=� J�L�)�����BC>�M��ɜh�'����$[c�}�DM�^5l4J�FK�=8�m�|�I�<A��fy�]>���b?a�B�K�BU���ٛ �>;v, �I����J|���?y��EK�(�7��	@j���c��J��]Z�i��b W]t�Q����	e�[5L��y���81����%/E�'}�'���',�'_���.��5��@�e��G��DIbp�'�r�'��'��'��O��XN��$���+�:��P"�i4>��N��5%�X���
�Z�@cb��4� �gm*����@#ˮ�b�L�y
� �-ᤤ[p�be��Ót&��1��M:�z�(�lH% ֊���+Y���-T�<Ү�CԀ ��q�R�#���AK/*l](A��kep��(� �Fٚ,HT����]�7[Hi+�L5u��i����zɐT��<f }yB�1$��p)�G)r�`#ʚ�+�l��q��<��]�7��	��Q��B�e�d)��ԍk^ <�����B�'��au�O�MA�|XS+�e��d�sYVr)�����CE����]	>QPkő>9ӈ�!%��(�(A�zq��T9,�p%*��~������T�W�:�J���B�D��XR��'��>}���	?�|��\4% �K�E�3��C�	�5�.�h�NT9SА�%h�����d�'�$���W�j�)�D.XiK�>!���?Y�QA�����?I���?ͻ �����G
$���b�B����{cH"��SxJ �'	@�g��)"���է�$�hl���m��!�# �!h�ɀ��4��|�-�B?��	#h����V�Ґ��S1�O�)'�@w*b�N�K�=�b��=9�U�ȓx�#g$�4PGnU(�0��'�"=�OI割dp�:��N�)�Т��k1�@)�%�>�4�����	П:]wr�'P󩎍F� ��/� /Eh̀T$,"������ ���� �ʗ|+|���E1M���,B�I�+ք6T�@�Q9�Mb��oެ��d�9�Z��~��ȹ@��A� q��'h��Ic�Lܸ��.,Th1�m�- ��ȓ��	1��߇ #N(��!S�?]PT�<yA^���'�xа�l�����O�1dƏ_;�c��[1Nq@���OF��/����O,�hW��$7��Tosd����	�yΒm����	�x�
��,���*��}��)��ց+�2e��$YuT���+��=k����	^;uOz�Ey�$�?)L>��b�-h�6�YEA�!qq��AD)�Z�<%_�����G�]�7�Z��I�z<��i�� ��I�-'�T�"�=hM�Qىy�+�6FI�6-�O��d�|j�d��?&.R3K0�ԃ���m��Ȕ"�?1��Iz�����蘧򙟜�f��MLPT��-�6���u�0}B�V1�O��(
U���<���C��&ԥBV�>Iqc�����<�@h�:]���C�ςq�(<��h�i�<���c��:���/?�=�P�Ld����$
�t�ɢ�K3@H$!�����)瘟nZ̟ ���<i�	S<T����I՟���ן��!����ف{N|lcd�@ =Ҹ�<Y�'MHx���Ы�/p�����g�9�n�B/�I�p[J��$^���S*S�8vz-ʴ�Kw�c�0괅�Oq��'���toʉ%�n$ ŝ/_�q�	�'�4	�Q啃.jU��m)	>�y�O*�Ez��)&#�*`/�tm�"�H%U}`�aU-y�P���Op��Oլ��?����T�Bش=p�BPv� ��7/�dl��	�M_�pZ�}�R0P����O
d�e���\��!`��
I�}��	{�Ļ�	��!+��d(�.u�����?�!��e�r}�O݄�f�R��CF�<�󅋭7�����F,d�t²��C̓S��O��b�ƦM��ٟ8��ɐ\�\�2��]0tNhЪ�E�̟X�	%,�)���Lͧ�����r�ɬ��Y�7wלu[�i��R����;v0�Oba�u�^�)�����É[8$٪A�'�2�����r�&����	0��D��'�1_��ȓ?<�� ��#Y����u��,E�P��@Û�h�}�tQ���P�,��po԰Ԙ'r�UO�>����)��0�ğu�l�F�*f�*TOZ)i�����O��E˳u�x������T>M�O%^-�6\��j3��<l�
J�� �A˂N�ڑ9ŀH0����p ����m���ؔƋ����6�>��)Mޟ��	R�O|ҧ	/c��}��O��H���'D�@B�ɹ݈��⮋�@3VL[R�"����[i�'�B���A=b��)��C �Yd�����OB�Žk�(� �E�O[nן��i�E�T��ND�jR����2�c��d�&����ɼN�R1�G�9$`$@y �F�qz� 锥?<OD��s$	@�Jh�մOE`��)5�	�ME���|R&�2Hs��ڑj�
3�1i�&��yR"�=0�F)�N�`�B숥Eט���CC���ر���@�R�,,"���?���p�&2vSD����OF��O�D ������?�O��86��yt�ӤO�6@B���xBg��ڼ��E�D�R͋�G��q
�'�Ҽ����ش���CZ,�ȡdGD�?i	�S�? Z�0�A��@ѴT1t�wl
��f"O,��s�K?�,�VBݻ]zJ�)q�D�f�A��i��'"t�&/�r4�(�PꝒKN�Y��'��
�2�'?�I\�H �q���3�dɇv?���s�[�nڀPɂSt�x2X�^�` �x��V�b�H�I�MŹ(4����+���p<�&�៴�	iy�� -J*1!��o�ZY��I��y��'���ᓿ[����P�/�>�0������C�I �M#p�π+��Er�*�_T�9R�S�<1+O"��d�=��ӟH�Og*�i��'��چf�*08qx�N_f�h ��'bۜ�r�T>�vg�S�W6�p�2
*��9�O^��Q�)�J'�1��)�Rgx�u���N�'���0��˘��O�^�I�j��-[.�S��G1�8j�'..u��c� u�AJ1H�)#Ó[�ĳ@�J��Rýe�l�˖N5D��iqLM�N1�Y��vf���(D�!5<)VP8p%A�iUyZň%D�����o&�q���C�5]R|��'D��J��_+^����ÿ7s6ȸBB%D��	#HĦ}F���wA������ D��6��f�\!ЃN��8
8-1�=D�ī�=�@8�.F�F>��7D���C/%�rd8$'�-H�i��0D���զƤ�fM��j�!{bD����"D�pYH<����ơ(�"�;�D5D�А3k�z����,H0[��	`�=D��� �Z�!�rUy��K�![����-D����k�!0�й�򋋘�� �-D�
3�XnbiN*(||�f8D�J�)�ZGbtK3b�<`�X����7D�,J�m��'�p���5| :ѩ6D��FiQ�	N�Z7Ȇ�����2D�p��.�UZM9c�y4��+q�1D�� �#�袱��ݾo�5��n1D��JG��+;��9[����B�OlF�B�*���k��4X��S#M�B�I'u�̓S�
�f�&iK�>L C�	�h��];�ɃQߎe�Zp�p�&-D�<��fJ/j9\8dX�#� �$,D�l��3����E[�W%�<yW�7D�T��
	�=�q���C|���5D���VKM�#@@���2#h@�5D�!7�{o��H�Dҽ
���@s`-D�,�u��q���ӇI�.\�z�3 �,D�<;C��0TQ��	Ho���ܳ7�� P���Ot�V	װ<B��B��$u`<�A"O\HHd�R%��%YE(^���O:� �.�(�0>	�iǌ]�e���741 ��}8������W��d��hD��p����׀д<�!�䍄}� <��M��/�ɉd�ǘQ���`ጆ����=�eGś.?����U�}U�$a�"Opa!��.XTS��R
����V&蜭��y����c�X�@E�7c�r��
�4D��8W�Z�i� ��P	�|	;���O��ن�f�|Ҁ����E*���F��p�t ����=)�O���"ƜeJ�"\�C�T*�U�!��p�ȓ<���{��Q�A�0X��bߦ
z��?�4@@�Pq�qG���y��ɹ7�K�l��QK�.��y��\�����W:��q�cCX7P �U��{��h���X�A�H�h�Ǎ�<?ڈxp��!��q���%F��"��p.юR�	\jh��:��hт�z9���M��(㤑��51޲���'����d�		1�ׂhF�!#�' H�Qǅ�,r�"��uE�J6<1Fy��!w(X�~�cmS&7$����1�X�$�c�<� j��کd�p8��5~͈b��<(��
�}���'�&��g��I����(g�@	�'mXyp�-H=�[r�I*3�����'I:ȡ�g<�Ov��b�l�.���DZ���T#��'���Ɔx�020��0fcd���(�Qg�"<O��#��h�NA�$���F�NRܹ��<�>B䉞4�}i���$\b)PTO�0(�x�Or	�O�2����O*�-ɱi=V��do�9��0)
�'8�m[��R�.���H���2�b��<R����Ol���ʄTTZ�	P
�	H�M��OJ�9 �� �RP)��4T��1C/]�G	"XJ��+��
�A,mz4J�E&�옇�	�25
�N<IqaG%E�<"� Z�
��EQ���y�<yg�_*=� ���*E�E���@#d�m�<ɦjBBh��@2ዽQ������A~�<�u'ݞR�X�Q`�Z�֎4�um�p�<��E�s&Q��A@4x�'E�<iV�L I�,�!`,<Dxd��eGD�<�B�$?;�q �&��q����`�3CP��>�萛w��y����L9�5��e	{����cZ��$,���z��R	I��I��D�=�!�6`�A5*<b�L�K���=��O`�g�I�O�D�;EZo�4���C4Ee�|�
�'�J�p'��PՠU;!�\,>d%�ѯ�
#y�Oz�}�JHI9�O�X<�hX Mۢ�^	��_�������'Y�(3ng
m�f��0�O���h�m�S�i��(��E�X"W��8�
�r�!���| q���ܛ.��xADB�6ܞ1*@1�	u��~Ba��.��͂��&��9Ra�=�y���ǒ�rdI�@H闂�?��,.C��}��P�R,��kq�ʖD�JX�B���=	T��7% �	�u����uJ6E��x��
����B�I�b?���
=?!�[T�]�h"<I O>�2kF#��0� ��G
j<(c�#D�D@�bJ�qۈՠ��ާ8G��b!D��s��.4i���X �sEn2D��Q��Y����`�+K�X:m�g%<D� ���zV~�!"��"q�� >D�ܩ���Z�uRҎ0%�Z�g)D�D�#��"�X�Ǻ8�+� )D�(�Pe�D�xkbeK���щDC%D���d&َ8�VQC��G(hޖ� AC$D�  '5���ae��T`��5D�`�w�_ u*RKC7a>��	 D�h� :T@�h�#`|
l��H1D�����09R� �p�P5��u2�-3D�L��S�h�洺�,���A ��,D�<��*�8��\���ݒg�BaDA*D�Ac�D�N�����⚾Q�$���F)D��b���aТ��UA�,5�성�(=D��
���2y>�D���	�&���`��9D���t�&l��Łc挵C�,L�'�9D��7�O�Qi>\�h ��,B$B6D�� �Η��|8GeÎ��( !D�,��/\�6�6���M� ��I�=4��3V�?{��e���JU[�Ə1gmч���]�ć&q������-+�����$u���<�g�����:��H;6����B$Po�<�f�!",����5tBx0��m�7pJh�?�}z��DZP�Ö.T�r���#�@f�<9�%K�t���ڇ!O���e�th�J��h�	Ó5N�Q�o^�puzL	`�S�4�Ɠ=���)�D�bHxbd�31ߪ�q�:�xb	D�?9r���JI*,���y
� 2�a![�as�Ż�g��Ӥ"Ot��A!�@h��)T��e�i�e"O�qj��4�i�0!<v��A�����L��	2���a�B�2H�Ѓb��$�"���2#D�>���hV��'���5I��ژ(�wn�55;H��ϓ҈��n�7���/>i��c��G\�8�O�D�1O\�:�G�����O^���	�?Qj�i�㟪`6 M2K>)A㞨d>mrçizP3U��:`�R��s��צٙ�7�ɣ+S�#|�'zp�E�Q��T*�!�bfX d����fvx`��ܴ]�8��!F�Q��ڕ�L�;�ܩ0VK��$T��O�I�5��8/�9k�H
# z��x#H�e�te�t���B�yrʋ�B�@�ϙ�w$�rFFtb��R=R^P�h#C� ���ax�p�6h!G� �'.��H1J50�"T��ae�@Л'#�AS�_U	R�$y���
��iہ,�r$�䎐1�!sQ�+m�=�2+�<�D�*��E�T6O���C6 *�Hf�^�{Yʵ� 9,EA&�Q�$��D�/��K�3�ŀ�y��m�DP��oݹU�
����c��ِϓ
��T��9����U<������	�l �7 �0>�^t�g!�s�'�������|�I2�l�K��3`�|]�4��-4�#>�EΈ�3I�bD��k�����|�T�/H���i��f��4�Lwܓo��,Z��ڦ~�h#~
���#"V&Z��҈���"A��?!fm�,,�
�H��5I��a̧D#�;T���a��] '��,ȳaq]�-%�N"�%�O����
[?�C�ùc�$m:W��;�Ձ�o�x�*�:rAä3�\�WJ=X~6��ãҋ�Fx��[-}����!̊�>t	�ϓ<ެ��W�ѽҌ��O�X�!�ƃ;�8�[�CΧn��x��?O�qZ+��*L���ҩ�q1��0�FL��k�Q���Ǝӫ�Qq@6O��?+Z�#�Ą�?��̘U���<���b�L鸕@׾=��\c�ɿ �v����m>�0��#o hxRD�.D�Щ�,�	 z��C�F݂=�?E��?��r�  �H�vhP��\�A_�A�&��yrn�Q�LeYvɥ~B[�3���0�2�0�p��,;�b��W6u�@tB# ���x��?ҧ��s��Ђn|5��$��/®��ť2L����N�o��]�$�*�M���e��it1�Ӫ[�P	D��%��G)��1���8F�!�� ��I�p�ѐ}� -��TY�U���?h��22��b
%[�/(X��D.2���P	[��������I��I�*���aܗe�IY��%m�u��B+je[qi 22ȝ�Y�f�0T��1����Q��Z�<1v��	(��9	�) �h�tЖ�������F��P� 9�P5	���&>o�F�4�*�:OM8U��6b��m�p,�9��)`Q�'�
-�v��h�P�*B�߁/Ff�:�ԝVì}��B4|�flV�S����% �">����X�,C��*H���:�l�u�'��x[� �Kj��)��ؓ-V"-;E �Z_�+�	�(/����/��!�$�m+��+�K
 �b���f��I�T���CS�C3X����e�2EQ>yX�_�6�V�9Ш�Q@���4D����.U�c����R��0�^��g� ,KlR�:Ҁ��?	��E����>�O�*�&��CA�'	��
�,��!��,ke�����@	o���7+��!�d�%��ȓ�
�l�*Qc��-�!�ĉ�MW�QYD�D)n�y��bՆ*�!�$GH�6|iP�ë�(����J-g!�ˍԌ}S��)o�d��뇡Va!��@f6в0'ڱf�J�7+$D!�D^!�ܐ�B�138U3SjR@!�ȧ)V�L��Z����r�У%S!���9�	��:hrz�h�옃e�!�W��3��הS( J�iۈj�!�C�_�<��TaH@�Ԫ�;'�!�
y�!;u��f02E�@N$y�!�d3p
s�9&PB�ڤm�!��L�pG��q�ņ���9�ʖ�!��ӕd�0�XAG�B�)�԰;�!��
i�	�%��U�6c	e!�Ą<�m��C�/$�@y��g/!�(��c�.9�=F�	gy!�$ҏI>K6iA3��ck�Ar!��N ;��xgn�;|�В�J\?@T!�$Ǔ�ZDc����<�&�!*�D�!�؝ �����J�E�}s�&z�!�� 6�J��C2~�&�j"F0B�D#�"O����D�\�vA�#e�(O�f@��"O���Ѯ�'*%���D
��f}ɗ"O��c�#�:m�t��$�9�(�"O|Q:@�D� _��jUcI�n���+�"O����È�.Y�J@S�9*�:W"O����	�<����e	�bҔ�r "O���&Q�HW0�3&�J4V�����"O:��˒k��m����p��8"O�L����-���a���,9"O�t�\�g�he(�������"OF�8�f_�~����0�ĕ��"O �y�N%v��3�,S@�HL�0"OhڇC,��$Kǈi3���E"O�iq�H]���J���	o$lB"O�x���]!�<�sW��CB(�F"Oj4�G��9F8�A+Öv;r�("O�A1'��~o0;��3%�ū""Oq ��l�q"C��(�"O�ИLD�]����q�Gp���x�"O�fLK��8�6��F��8�G"OHqbt��>rqL�RF�?*f��I�"Of��`O,A�U�Vbԥ$n�x�"O6����ܒ`�R]�^�%I�"OȬ����/g�=1�FQ��0"O��wS)^崤�f�%��q�f"Ol)���F��䫃�}�N�Q�"OD��hC�
�ڤb4�Hlj\{"O\\�GOؠ-5>Q�B4e.M��"O��s̐,Gt����R5-��V"Oz� U�D(v��mX#�_�1r�"O�MH托Z����̡O��$"O�E�A��wv�i�E�A�M�µ�D"O�}�'�iRNp�SH?H����"O�����;D��Ԁ�I�z�T���"OZ�J�E�w���HM2M�x���"O�|b��i<��i�<�3f"O|٨�/dS��d�4\�Ih�"O�Ah��z�ڑ1��>jhv]�D"Ot�Q+�,��4s��W�
�
&"Of 0���<��,[�%	<)�����'À��4'�S��jbJ��X�P�	�'n����/�(v�0|I"e�,O�RR�'����piD!9�0qrT��{����'*���4�V	1߾�:�H�@��'�8�'��jF�T�@��N�4B�'1꽁�J�*�(�#��A�ii�'s���bI�u�ѪWBW5�fQ��'�H�Btj��h �9�!�&4	+
�'ڞD�M%k�F���R�;8�!�'CV5��V$��a
�@>r��i�'�.�xь�7X��|!kJ�s�F!��'�܀R.�K|�A�Ō���H}��'���Ej="�* 5��
����'��X��=4�q�R9-)@��	�'�MYTf�.*�tI���=<�6�#�'̠����L�[6BI�Ul��J���8�'7�I�ć�$&�� թC�BI�'�<( �_�lBL�g ��9r��s�'�4�Q��#|�mkw�4�b��'OTLA`)�q`x���!B$-��)��'Q����Nݡ0\��ID�0�@Ѳ�'z�ғꊩ=�`0�yby�	�'Q���#�ԙl��J g��oǬ$s	��� �,[�"�*pQ�-Q�!m����'�'����'�D9	�D �t�$����7i/2�(�'&�=h��*��a
��֚0�T5��[<&(#za`Ф��,X��V�Q�(�7'J~�<)�\l|�'�ò6`j�h��"�b�ȋ���O@��� ٩`�H��@+=0���"O�T# .ڣG�����J�& F"O�m��Q�<`��
�@�?v��Yf"O�I G��:@ʄ���Q���S"O�M���G��� ���I#o�|��"O��c#��&
���ऀ1?T09��"O���2"B�P{a![�g�0���"O�|���.�
X�e�-��J3"O|`�bNިJ�m��-ۈ[�؅!���6�S��OE���R=�i��+Qk�!�$.6��$��*�bU��R�A��!�J�2e���݄DO2		w
Q�b�!��A�FɚM�$)(G<�R�� !�䘿.����H�H.T�� ��v_!��"9M&-Qör$�\@/"!�ȹeը�Б��7*
 ��$&�/5�!��čoL�[���$3���G�!���1E�J�I�鄱V�rQ˔ �!��e���+`m�RP��膊�)T!�d��YA풍+7����D�UQ!�$�=;.fy!�eM9q(*F�dH!�d�1~�T)2oE��j��P�@�!�$�$��"AY]��13w`D>�!�$	�F�b�A�VoYҝ+!�"V�!�$�'u�(��3	@*�=3��/�!��I���i�	�&&v��w ��6!�D/��8��C\�C�U�樌#=!򤇬S�"H�"@�&\t��?�!�G�{#@��@I�=B<A���5u!�D^!~s q
��΀qk���Ɲ�g!�P�l"�Yf&��A.\C�%��n�!��fyر�FKV�4(W��b�!�D��;]�� d���s��$�rcQ�!���c��jǊ�:+���D�E�b}!��!6%���w-�+n��t	�LQd!��ۓp��Z���a�v���(R�!��6r��������	ǘ=�!��\JX�t��8��=&8!�5�Z9��� L�P�M !򤙁_�i�.O�X���:$�ޭ0G!��O���зcʦy#��ˆ&�-I*!���o�N�d�Y�%7`}s�	�g�!�$G>��@�s�[�o����C���!�dA�mo���FX�z��z'B[� r!�#9$<�����+g��y�@ ��!�D�=|��E1W�SA��3�!�x�+$,J<ar��PX��	]�O�8�1�� -1��W�.�j�':���	�5*Բ7k�B���i�' �Ԩ���.-RV���)͒
J���'9b�� G�6;��SB�.� \a�'�Z�+�H�L\�m
�ϟ�"��D�
�'w�e����f�v5K�fH�e6����'C�,c�+bc`�W%_aq��I�'�r��d�E�}�1���҅Y��+�'ib�Q4#����kߒdMظ�
�'�jT��B�:_3��i�e�5c��D[
�'g��b/϶MH����䛃[<���'� q�!iD*H��B�c�N����� ��j��ڮ�0�Kv@�*�(��"O.�P,��%�S�NW�\�eYb"O���E[i�@��QM�<��"O���%CaR �+VSv���"Od�hd�X!���b� Ui� �r"O�<�E��=2����j�TL��%"O��`N�t2-(��ئ'�Ô"Ox�#��әA�(���;V��x��"O��d'K2������p�&q�"OA�SF�>3�D���N���h�*g"O�!i�C){ǈ���Vl���A"O��*�F�P#��.��8F*:�!򤎏*�T%�u�Տ�B��Ei�E�!�d b¸��3��"M���fF!�B
I��yQS�Y$0�0h��NȻG9!��>��� �藱h�<�I�-��D!��ŏ.Em��M�"��,I@g_,!�ĕ(�N=��ԾTè4��e\�!��:���D�7��bd�!W!�d�K���rf�r�6���LW�K!�dR�A�4�ط��j��hе�g=!�$Y�H |�,H K���*��#(!�;m96U�V��#Cr%�R־e�!�E�t�t��6�˹J�2�q���!���M� ��bw��
��!�dB1zpP���)
q�T &�-�!�d���Z�f�R4�`�[�?���ȓ0P&Rס�<�<�[tkĘSZH��W\"Th���-LX����"��'���PZ�!x��U�A�U=,c������q�wDƍW��ېߺS��C�r�^�Z��7��Ja&�!R:D���N%a�.U���kH�%��N9��L���11J-U.~1��K��Ry�Ms&a1D����o��!�x��o�Q��J1D���Td *3챐���,���f(=D��2�?1T�}�� *vِr:D�� u�Lp��Ӥ"�
�dI�K8D�� �@_'TT���^������2D�����Y�hѐ�![ ��m��J2D��`K4�|��s��/v2����.D���'�[d��m����� >����� D��3ܷ"��`"eG�v5�u">D�x{�-�Һ��U�.Q`^��>D�����%�D@C�	$p�<�	QJ6D�����ͬ�����N�4�0��1D�4;�
�{d(�h���"����j.D��)0�;&�0�y��:Z��VE:D���梜�)T�P�Q�V�"��rK6D���!��Nh0s*ă �
Fm9D�|�0�ـ)��)) 0�]��!;D��J`H�9�L�z�ݭY���VO7D�Drvf����(6����2�� �4D���tn�U��84��"(�5H.D�����:O��(�Mϱ,�:u�V@+D�X�&ʀ�V��Q fJ�x�H�g�,D��0���B?��B��A�H��!i6D�(rgk+8a�3,΃T�� 0�i/D�<�'��NY��� )�`�g�'D��aJ<y իf�J({��y�#D�lӒ��	�p�;�j�� Ġ-�d?D��
щ�,�dL��瓣�:�	��1D�<�"+)K�0+Ta:$�(m�b	:D�L�CFf]PѮa����#c6D�� ���B��6���3E^%9��df"O.�ʃ��`{� `
�$�""Obd�p� i*�jFB� �60h5"O(�AA�Q�7��X��A�;��|�"O��(W�@,�B ��$`#�%=�Py���E*�8�FΊIւ��F��\�<�fK�&&���M�;����p.�t�<�Rl��n�\�� �Y�9�OOK�<�#ĩ�Ԙ�h/�
yՍ�D�<���
6:�܃�حT���ơG�<���]�u��lhw��)������B�<��;̤l��*�I�a�[G�<i��>>%���U�ڈcP1%l�C�<dƍt�n��w�T!�ҭ#Nf�<�d�B$+��E�"W�$
�<�+�[�<�%�@��)��j�Z��ƉY�<��T	�yZ��΄^�`�0�	K�<q��)q�B2bF�l������J�<����%i���k�Ȕ4ٚ����C�<�@ͤ@}Z|�ï�'�jU�Q��G�<I�͝5�:T0����(�i��GL�<�FеJ_�hC���vW2�Bo�N�<a���FF�a���H1o(:�i�K�<�f�Db�����Z�!_�\��iB�<it醧N*\��eZ#�>��FPv�<�Cg~����Y�:�,�!�p�<�AI	�
��ĩ�9���`A�o�<�7�čh98p!� @�~�B��C�<cF��喙*#��w��=��o�@�<9%`@�|�"`�V��:@t��NJ�<Q��QR�Ţg.��O`��PuMQz�<9��ʎ��	R	ւn,Nu�z�<.�0g��Ɔ6vh��K��^�<ytϟBƂ!� 0ZEpţ�O�<��cW�M��h#�2%�ʈ�1�M�<��Y�?��j�W�+.�{R.b�<�bkԀ��,xW��	�N=A�_�<A .�U�nhz�ސ.4��b`h[�<�a������kQ2��I��U�<�(����Y	��Y-I�z�1���M�<�f�\��$�ņ.E��J�@�<i/ʍd�L1I�h�-T
Q@'ÈR�<Ѣ�����kH)�}@���K�<Q�B�	7�Y�'�"<K�ab�n�<1���$�6����LE��]��lk�<!1eM#<�V���D@+g�Q� l�<1jC�-��� ���H�&��R̈~�<�q� �X0L�Ign������@���<I��Q�5�X,�r���E�XAa��{�<�.u��̨���:Y�`�֍�w�<)�-[� ,�u�E�š	�U3«k�<ybǔ���Dj� �2j'�s���h�<Y�(�"��XH,�%���ら[�<YVM��l�4T+�@�;s��`x�X�<�歜�x'����iB7�N��#MWk�<q�,:u���ۑCǅ.Ў}CV��j�<qA	Ps�:���?(���E��~�<9�N�**���Є;~��,)!a�P�<��A��^kb��&U�&�$�&��A�<	բN
X�)�OV2=e��x�l�B�<��l����LQ�"�Z=pu+��_@�<��M*!>�j1˚�Lm��3�&�{�<`�:7�pwAT @ 	�_�<�gm��A�1�0k��v��d;g�^�<� �T�jR'�ֈ:�kO�\��� "O0�ن�B*,2�tcԋ
>� XY'"O�9�vd�gk`|;�dMZ�P�!�"OFt*�e[�L���F��p ޑ�"O)*�_�~���'&5n�S�"Oj�{A�*|��sG�hk��3"O�]#3ᙉCFȉ�)�>|>�E��"O�h���!>�jQi�hɀI�D��G"O���%�E�4
��1�Z�G��Y�"O�pH�ɚ#|W�٪�̟��(� "OV%bìŜD��zc���u��	"�"O@�RQ�A�w>�J�I��9��"O���@�oW���ݶ^��|K2"Oh%��=-���GN��}K&��b"O��{���8%)�c��E�g;4��"Od�b�Qy(X���` 0dQg"O�E���Z( Zp��s-QtLq"O� �oZ+
վ8
��S�q{����"O���#	�K�]�r!�gB\�"O��s�M� �(9���G#�ѣ�"OB�`���*0�\QrE��ui��C�"O($�ѫ��]���,߄Wr�R"O���!`ُ�b� �O�lh("O �	�d�2ː�h��t,H�<-L����o۬� at(�I�x���F����8��X���ny�ȓ?,�:����o�Z���L��L�N���5F�0 5*]P���{Z�y�I�ȓq(��0��A�*���I���(E�t���r�RqQ".S&{I�A@��~�0�ȓRVu�q͇)J��3U��?R֐�ȓY���	�2/l�+a��_ސ�ȓF�ؘ{�GE"{������7c�x��O�5�5b��r���c�䑺dUh�ȓG) ,���4EZB�K㢓�;� ܆�s���穋$����hT&2܆�n6���F\�D�qdP3L ��J� � ����Gf���2J�6��}���AԁL�^Ej��DF
�1�ȓI���� J�p���K���fxb<�ȓ!
@u�.��P�u�'��>�RI�ȓ��'�W�XDY��F�,� �ȓgI�$�b!�\�Z�0f+�&k����ȓc�����	�=���S�B��ȓTŘ���F�/m̽c�K>Fΰل�!����ծXF���`�S
U�u��z�����*�%;�y���ȓʀSaD։�P(�d���BD��LS�Ъ��U�F=Li���[3Z:p��x"� ��Cw܌1P�'Kj��ȓ�^,��@�7a(�]��$�u�ȓH�H��c闚m;��f��3��H��0dr�#C���X#Q#�?LdI�ȓU��aB�D�!D�i3�
$it��i�h�Ԏ� |���cb�q ��',\�[1fƢeM��;��TM�.܆�s����焩��-�sBL�U�ȓ:��	���-.�� �@�uEb�ȓtO4@��d��W�����H��
܆�Zʑj���`̒����@�Z��ȓK��x���P���n��R�\���N1{5����LY���8���ȓs�.yk@�3)�i��)�[�
t�ȓm��RFc��,�a!�m3M @݆�S�? ��U�طI���ě��.�[G"O~��T�� )��BC߁Ē���"O��KgF�݂9Ģ��O��x�"O0����Sbˀ��a�6���F"O 8��Û7z���)e�I ���I�"O��	�� >�}�mT�(��R"O.d��bV�w��@��+=J �"O��j�eI�0$.�V��_
f�C`"O 8�!Bh�.�` J��K��K�"O0�yaH�l�P�( @���R"O^Y{��Fb��u��M�9ڍBe"Or\��ő�+���
�'X�AߦHS"O,��Sw�^��$e�;p�n]h�"OQ��<+|����?J����w"O�2�� F�b��I6Pp|Z�"ON�аCK�GY�\3���g�9��"O�j��ʰQ&���#%�2&W
x�"O�p���M�����%\�*��W"O�m����nL��z��Srz�
"O�!�%�1
�@�2�̌S�	:�"Ot|����G,��%鄝,xb�z��	ҟ���F�'aŀ��܀Lb2��A�~fJ��ȓJ0���˸�Z�A%�;����_6ؤ9���#�	"eD޲\K­�ȓi����@�h���Y3��.*�6�F{��'!��Hn��Lb�B�m�$Tn��	�'6r"GM���1�`�>nH�	�'~L�SEe)8$e�D&��9�\,�ߓ��'��}Y�:K��IST�ǉ?����'s��ّ.�X�4�QGj�b���'F�}끧�sH�a����YkJ�"�'��ty��u�� !��� F�x8�'�\���W��ء�HQ� �4H�'�\U���u��}�A	�B�>qb�')b�AIAo0��`َ3�� S��D�O��$.��]�R�� M�&oa
4�F�X�WS<B�	�S�X�x�%W����n���C�I�Do��ڦ�B�d�,�PE���C�	�OَL��4{�U1���qp2C�ɹj� Ī���N�Qj�o^,L��C�	4Jx���hN$wڄ��b��C�I�3$tP��bt����0/��B�	>`���L�}�MC��	j��B�I23(�ɚc�W��M�Ҭ��#���=�
ç:0RůRu?�F�+ 숼�ȓlJ�����,}�\0��M�=��d$�`��I�(��]�+ܔ�iGu!B�I(��Usuk�b��9��|�PB��lr��Q2�ٻɎ\H4����C��B�@�[D?pX��.^.�B�	9K/H�0%�ކdl��M��|��B�	�M��l�V�S#=��p*��MEnB䉭Ui�P�w�ЛzJ,���-y�0��?�\��M�@�U�A8ȸ���q����ȓ��)�,c�dtҕ(�M��ȓQ���A���qTq ��D�"]��V�^m�AG�8>*����OR��H�ȓgTy���� h0<��F�nD�ȓ(���"@�	'�Xa�����h,L����<I���� N�$H���a�d�Q�'�T�<��R�a�2�!Ҫ� r���oZO�<��E�3���!J8���H �f�<"��~���D<JX(�@���b�<�D�)S��!�`�8j�$�� '�\�<� ~�0槃�q�xq�&H3%Aۡ"O��bgε&�D��w��?
<X�O�()�"��v�h�#��0CYB�#�(D��8U���n¨� Ԡ �l���u�'D��*4#Ӊ[�(ѫBʵ���B`$D�pА �]����1J�#Q?��+G�!D�<�`K4f��KE9sC2���;D��	w��C����O��L���:ړ�0|"e��;+�vX�Mɖ*l�qiV}�<I.A�T��x�KS7>{��ㆧQv�<�bn�����E���;w�\pQ+�J�<	�'�)\�a90�Q�\�6=(� H�<���!R�����I4'+p�&�C�<y�$��N��EX��T�6�����I?D�`���ܒ]����I�7x��݁AN;D�`����"C&jeQ�Ӱ,�}�a�<����(�����N�	J��˵=H�EZT"O�Q#!�ʨz�8�E�h9���"O���1e��%��9� ��j0bp�f"O���i�i��O1Y'N�cG"OF�p���=�蕛CF�`�hk�"O|1[Ĭ��e�Z���e�0��AbO��E	[U���ǬϜl��  �K'�&�S�'c��Y�'C��6K0�i1N�sH<�ȓY�&��u��u(��6�H<q���ȓo��Zf� R�8�d̆�g�F�ȓ��]q�jвn��,�vH�7HZ���
i�oU=EFq�7E�Q�ȓ�vx�c*�v��e�9L���ȓQ�>���,��@A���<5N��ȓ-�n��R@�&OS(RSeS�9<|��0�͉����dņ�!2
�$$�Z8��m�<�ز,+B������!E�� �ȓ~0D�P�)R{>ܰvGR<#2-��	a~�D�lN6�6��Fxn ���ς��'�ў�M�LqC��K%ĜQ���1t�`�;�'������Ǿ�@�r[�~HK`l�Rh<!�C��z�t�r�`_�ddѐ�����yBB[�v���S\\;�F��y��78�B!��k��D"����� �y�d��.Ar��F+�:�а*���yb��1[#��a�O)�q�0�!�y��R[��- �� �Z K�0�y"��&5�8�Bo��;����V��y��G:�Y�� �!4�P\"��yҍE�1�JɒĒ�6 �]J�>�yn�3��ە쓾��]Y%�F5�y�ڍ_<@�p$x x���i̩�y��K]xi)���dg�hqP�5�hO���� <����
H���
�`�)r!�@ A���D����!�µBf!�O�c�zI�a��iP�xL�@H!�d܏=�>uاe��(ՋѢN�B/!�D�,R���NS*\b@ G����!�䌌]��Hh�bS
;֐�3�|!�d0mde�U�ˑJ�`��f]�Jw!�G�-���a0O�!+޲�R$ƗDs!������Į�i5�`;r@�J��yb�ɥm�rѢ��ӑ 8H�#���9M#$B䉥-w�H1�H>��\Z�cB�I���řG�S��x����.P�C�I $&��R	_�T����y�C䉱(�|�b$�2%F��6�,�C�Iq��<� i��ݲ���?F}�C�)� 1
c$F(w�H�bMU*{Teaq�'*ў"~2�Ŕ0-q����-e�-�6����'OazI���8d�@*(�8�S&ҳ�y�&G�>A���-	��q!�J��yR*�6���Z�M�1�����E��y"�C�BC�%3���y�D�{�� �yb�I�O�����j��U� f�?q����'��=��J��vv���3׃YZ��G{��I�<qt�P�8���k� �O���kf��Z�<��!��I�e���
1�L�"��HS!�
�W4�����K!���.�=D!�D�R4���V��#h� �F/�!��L]����n�D-
�,Φ]�!�M�1A�%�=J�����B,+���)�'F�
�k�%R:G2�t0�A�.Y�*����hO?��F��.JP�Y#��
-#���G��e�<�'�� w���5�v�~u��_�<1Vg=��9-@�H� ��B�`�<��ɵ�(h���>$�ʄ����^�<9��\.���k���6"̀�[� �Zx� Gx��~R(��2��|��������y�O@�K�� :�N)u� I�j!J>����)&
����0���UKO�9�!�$�7G�b`H�Q�hP)Jտn!���*�N����9F@���(�@b!�,G�5��1V���gĻ-V!����9ۢ��� ���!�LFFџ0F���I�`�f`c5�ԇ-��������y"�$A�%	��P8+��� ���?�S�O���6�R�p���-�]�
�J�'2�5r�f�
Ci�<BR��W����'D+$�Z�Veb���њK�����'���@ש|��9�mL�Q���B�'l$��O��5��u�;YdH��'��Ӈ�Y5su��ҕᅩe����'���jH�@5AĂM�Z�DI����hO��̓x��� �T&�>�!s�.J��5�ȓx�F̐0�H�?Vy��Y�3<H�ȓD��`.�D�p�ȖD�"���ȓ+�,��_
i��9�/̟�(����<�cɖ�#2΁�! �)v���o�N�'�?E��ɞId��J���7��S�l*D�x�/�$4(��[�(h��P�G�'4�(�A��g��Q�.tgrQqD��J�<�b���0Lr�)�jm
q SD�<2i��]O,�SŞ�t�Ĥ��,E�<)d��]�ŠC�:Lzp���C�<iV�òER�����*��lz�Їȓ@�8��EO�W�z��0g���^)�ȓF�n�*��Z ���W$�YM�D���}Y����7.�7f�.L�6B�ɧ#7�-2֮ڽ$��ԙ�DF/fB��<G�ֈ"��K�-�0	��aZB�	1w�����L�i��:ƍ��|@B�ɓ�8=ȗ�θWitB���Y
�=��'6>�qP`8'D����A��5��1˂��-�C��� 4k(/!N���^�t�Ռ͸[Ͱ4ʆM�:Z��؅�]ސ)�b	�A.Q���<2��ȓ_�xE�V6�;��ڸge&؄ȓ[m�՚��\@�x�W�Q8�U�ȓd����1IZ$f�&��'ֿ<��ć�:�꜁&���'�FU9g�I�u� ���؍�S��q�$�өU�m�tA��S�?  �zB�4jX������t	6�q"O��k�kC�`,�	Hp�X�$�Ne8�"Oh���OX;Uj�Q��o�F�N�Qb"O\q	bjπ d�c��ڂgd
T�B"O P�2�֖s�!�f�x��"O���g�ٻv��cc@80zBE��"O�ȓ!�Q+��j��Pbxj��a�	L>��L՘=��	�u�t� �bh7D����Fֵx�Fy�!��X�4!���6D����+�@��@�P,|v�lR��2D�`�!�ח"�Z`I�
�'o0�p:��/D����!G&�@��,ũ2�H�۔�8D�t�#�	yK@|��E�n@hȠ�(,�$(�S�'�����`׌bMb���P�RuEB�%|�LC#�5�� �cℎ:�fB�	�6�<sA�D�n���c3���C䉤{��i�TH]5F�m�.#]� B�	";�:}Ӓ͋�0ѺpI �ҊR���=YL>����b��gw�� ,�5"{r���i�y��k���5!�5L�����yb�;x�`� �釔�Hbeh��y�f�@Z��ǁ'kf4��Uᙘ�yr�-)�i0eh��q�e�C��?
�'�#���4����%V�:I�	�'۰���l�>@[jL��P=nf�ۉ�$)�n�W)�d���*5�J<2C���e�'��П���Oj�ɪC?$���d��E�b7N_#snC��0p!�Ihb��e@Y[��� N˓�0?Q%��*Md�ػ�IR={IP�R�Th�<!u��6�`�rS۴�2Oe�<�A�6~L���DF�D��4��j�<5N��iB4 J0�?ɖ%��g�<ٕ�!�R�)C���X���J�`y�'��|��������+�;!��aKF+A��B��>d��A�v��P�X�*����O����D�=�8 ��;��D�&�٠R0�)�c�ܥ���C+��C&��$�f��'����WgVl�P����_�����'�T(��ƃ�r�d`���\@���'�A{1A �Q0�ͲfiA�X���+�'?�=�5�>Yi5A�"ӆRU���
�'���'#]�&�<DrV`ٗ~����	�'��IS��Q����	�"+'�Z���'��� ���(���!?�Ҥ L!�Č�D����1ӚMX����1!�Dٳj����h�z��}
pK�
/!��^���r����NT�״d���'�(�@�Y�6Q0t��'+��}��'���T �ˈ�CZA�!9���C�'�a�ԡ]�(���-�&3�%HA:��>����?ّa�2C��C���h��g����y�f@!} FM��σ� �݀�Fˤ�yrٰ[BH�J���T��ȶ�2�y2b(o4LʧS�@r1CJ��y�BD/vW�5����69� �Ѵ�ٟ�yB�^�\/�y	��ԯG*�e�g�F����?I���� 
xN��3A$�8�0r�`�1�?��'y2l3�^�iw.�2C���/�?i
�'�����4r��y�c
P��Ih	�'^��x�K�m=���B��HR������hO?=�b�F�F��yU~`ޡ9�F�<�%h�!P�,�!��2�����S@�<�Q!L�;6č2coӉP���s_t�<!�ɔ�$F����ވ	�´��K՟H��S�? ����ےR�]+"�%Jmpѫd"O4��2�K�e�&��G���>�����"Oࢆ̵�2�	�φ���=�1�'�������
�&�h+�1��<��q�œ�m������!��\(��ȓ�<]�Њ�����5 8�>]�ȓg�0\ؕ���9Kf���
j���L<�Ā:D���$L�$Av=!s�F�<��'O�`@�AK�Μz���^K�<irF57������-"Ԝl�d̚I����<2l^�:�hB�A�$;I�`�p�G�Il��$�Uݬ� 玬o.Pt���!D���b�Ȇ6<b�!'& �x����I;�OZ�o�*R���;%��C%A�'9X���ȓ#�`e*U�Ymb�0v��� Y�ȓL}��X��X:+�r	Q.o��ȓ@t���uMɿb�HUP���Ow���(d<��HzH9U�X*�����'�����ך]jDI�����h?PA��'?ı��J_!5�0���e��= �'Z�,¤!��Z&�T�b�L�V�ΤK�'�"YR%�$�hb�,�b ^a��'�>X����T��)c�!�	��d�	�'�5�/
�"���ܲ����hO?y���7S#���6�*YRL�� x�<����==*����2iZ��{�@�}�<��j��/j��t���~�.MѲ/y�<��l׿}3Аy�c
|�� Ф��s���0=��M�/E�0p�&�
`�p� � r�<YC�$��<�f�;V.i��H�<�# E8�*�Ab�H>{<�a&Hy"�)�'l~p��� ��KG��0D̰�ȓ.�<�䄁::��k�-�%����n���E&Tvo�[F�ޢ.p2}�����'�fx���l�6�,A�p�����'��>��$@�Ļ�dJ�O) =H1��� �I�ȓ]^�P 5�;E-�P�r��6��4�ȓ�^�q�'��+8�8��c�F@������R��#g���1N��P���U0�� �o�8u�Q�0*�ұ�ȓ�\9�Ft�,�뇨�<��q��=��K��=f���D�R�c܆,��i��	@KZ����ӄH=H�pІȓri��-c�	:�aI,Wَ�Õ"ON�Za��L T�t��Q�����IG�Op~]cg��-Nj� @��X�4y�
�' ���C�5~X�w��P�j;	�'����%R�B�^S"C�G�`���'�f,�p�&yg���g[�>� ��'!�Œ�d �E{-*ᄙ�9����'U���`��i�X�r �G��j���'&L`�I?�!�4�^MY�q�'���ӕ�س%���H�m�t.�K�'˼����!]TdӠ_�q�� �'���	P�ʇ*��)RU��j��1����?qpφL[��ӎ��J�����y"#_�T[�g��Q��]���y2c�]�r��bK�H^��O^��yB��!
9��e�E;9��������yB�ɭ'����ČfﶝH2��6�ybC��S�	��nBV�Ġ�Ѩٞ�y�&Â(=j��snԮO��)ԉ���x��y�L�Oǳ?���5Օ��Op��2&M�pZ=�e�ٶ*_��"O� ����"�@p�RG�ޭ^�#�"Oh5���D�uH҅��`@�_h�i �"OJ��@H�;�t5�A/K�neZ�"s"O����KmH$(3u�ބL��a"O���n������D ѿ':���S"O�q�6ş�=?`%3c	�<4f�p'�|��)n��1 �,I�w�yeŇ,�C䉹<�����8[�0"2�XC�ɊM��i@���9�� X�J�n��B䉋K��d�ԺJ���C��~��B��x��ʃ�&7�F�a�]�h,C䉫P�>�:Q 6�$+�㐉#.(C䉒'�
�@7��4,P���C�\�R��?A��OI1O��	�� 	<�a+%`ȇx�=��"O��`"��t�XU�¬ưn�Qڠ"O�0��1N3 �x� ��2w�xhp"O��� NFR�f�#g"�>uk��k�"O~ݩ4c��;u�l!ōvV�0$"O�yYqK�K�>��/P*EP�U�"O.�1c%�t����-ɃOG���'z!�Ĉ��C�B<%�TQ�ABQ����!�'�A��LP�j���l"b ��'~ҭ��.��X��|�(�Q��)��$4��dF��/ojYD$A�"�i2"O��!��E ?\�吃�S�'����W"O�8�S-1�=:e��T#B	�"Oʽ�3�=4T� �T5dn�m�E"OB�� �1Z��Ĳ�&!iv�R"O�݊�[�Kv������VZj}z"O(���C#c8#�U2=XN�q�|��)�B.qD@�=p=�b�Ų"b�C䉍La.HBd��*"�������4p��B�	�
�<J�ycŏ��n�xC�	�u�F��Ħ��B0ΔaU�W�/�FC�	z:Jl�S`�NN�d�R䖁�>C�Iy��٩�@��p\$ u��	iC�
����3�Nvw���K,Y`�B�I5���ʕ��)��7�ɸ_h�B�	�wiY�	0p���8�'�2*=�B䉳Ob�M����x|�D���X��B�I�d�*Ѹ1c@�&s� ��:6ٖB��b��)��NW�5V�b����6�C�I�%�������7%>�9�d�o���Ɩ7h�0�')ɶ#�LuH�l݀d�!�d'��tr�A
L���`�3`yў�����R��Q�܌[�*�y��U�!��B�/BIJ��KS�����ZF�B�T�&���&��l�ܠ1�Y:>[�C�	#`Vi!֥ 3'�
�|��C��
u�$�O�'��ҧb�I1�C�	%�Ơ��ʓ6��A��">�(C��Kz��R�٬Y��͹!N9'�=i�'p8X��U�Hzzcw��	Lp�ȓ3���.<}F��
u���oq�Ʌ�)���*bӟac 5�7㍸&r�Ņȓ4,�����1\+��Ġ�2k�|�ȓ$���0OÀq����L�FL��ȓ}?R��%Ċc^1��.q-�ȓI���5Ν���k(I.L*�D{��O�r=�I�HQ��[����^Ƙ��'�,q1+E��5�a/MA�p��'g�a��m�|V�A��%�C+ �S�'|X��u☛W@z%�0��0J�)�'������.p��=J�f�-#_I�
��� z�J&k�:"����F����� "O�"�ݐ����d�P{�|���	]>I��������dHe�� 9��<D�@��(��N���bӌ�M�� Q,9D��r0F3"�Pq��
)#Fq!G�9D�Q�)@�\��Sq��Cp}i�#,D�0{�(��"��	�r�z�w,D���B��	ᐱ���Ԑq�LQ	%�.�O����@_����	wH(�{��W`"�=y�'gf^��0��y���f�\�M��C�~�c���8�2pа��!n���WR�\i�F*Hj4��m4'�i�ȓ q���V;��L� jZ2 �d���[7�T"�@Q�y����1�Q�ȓ�Ĥ���Z��j�cd*}�X��I�<�r�L�Fj�H�����̑ђ%RV�<�/� g0���@��橕y�<���#+v��D\��>r��~�<b� F�6Y��ɐ�Q�8�	C��@�<�������d��j���i���z�<��dίU��) �b��(Nh�0j�z�<�fτED�]9jћ2��� "��w�<qT@�5~T�Y�3�]f�0�Eb_L�<!QKp�8@���E��x��'N�<����I��30)�o����gH�F�<��K}����!ڬO0hU��[�<)QG�)K�5pg�=8'��ba�_�<!Q���)��i
�ϋ��8PA��C�<����Moͳ�ꎚp��p���Cx��Ex�n��h�E�^1��۵Đ��y���o�����O3Y��5����y���yZ@�3���:�5�tF�yb��2't��"�܄��}�$���yR�W�5�0H��n�����ʣ�E�y�L[�qCjp��B��,��� �ybEA;��NX�
|}��']����hOq�����n�*H�m��W.(�T��"Od���/�;@���9a�x�9���'�!��
����E�}��L�aoߴ-b!�$E�X�z��ChӺZ���c�,DH!��0$lq����^����]/@!���&]��p�Lͪ9��|(���U-!�#UI\�x�HD(;��I�B^.K�'4ў�>-�Q��X�L�A↔�Z��h;P�+�����B���c<!��jB��\�<9�Ϥ]�dp����+W$��a��b�<�Dٳ�\��ĎN��ܡ{1�N]�<���Es  ����8`?N���+V\�<a��Hyj�Qb˶`~�d@& �T�< 	��D��cG=�x�F��xy2�)ʧ�.9Ç��4Ndy�$����<��t�,�Bw�S7"W5#0g�6�a��/\�t��N�(y"\B/�"9���r$�`���60N$m��?u� ���
���G�Ki�E7���*@��ȓ?�D���N,,���i��2By���JA�B�&h_�=�`�	1*ƾ,E{��Ou����ޚM@>�"ǜ�kP r�b�'Q�>��f}��w�Mx�X:4)�:Y�",��]�h�p//)��Ղ0+ҵBUh0��xI�1(`��2s]�<Z���af0�ȓ"���w)X6�v����ƭo���:��q�"��OX�ٖaM}=���X���h�C]蕰��'�����b���	0�)� �䈖�_�Uo6ћ�@ЌM�~I30���O�=1�'��|�7/M)*�	��&ùE�H���'W��59}�v1t�T��
�'�Ti�`H�.on�œ��_h�B�I�P`�P���"����qMݯ>�B�	�(��p��pO8��S��6|�.C��(9�P�X�㍳f,AᝇS"C�I:;F*�[a��<|ʴ�PKN��>���<I/7�D�@�C\;$xDCCJ#�y��F
 H��j��͆ߪ���y�"K�E�.���
	x��)�1�y�DD!]�m� ի8� ��G��yr��uDd�` 2:K�\��Q��yr�GR �I�6��!�q��@_��y2%�k�@�K��2%
���?a�H|P�SU��j/�zU@�;3��z�'��Mp�D�&�ru�d�Z_|��'�^��a�U�<�VmۤHѵ��4 ���<�̈�	>=G�T���LP �"Ov�� �D�"{��d��V�J�*!"O0�(�Y*�]s�A�%Q\Q+!"O"�P҄VOg���v)���!�"O�@�l�62&
c�����ɨ��|�'�azb/�|6n̊�"�=�"AB��-�y2��9^��7-W�.}.�kf�O��yb��*f�}q�*])�څ0���y2�R(p�)�v,O���Η�yB�B���Bs/B���i�R �y2-XT�hh�0v������yK�7y����H[� ���MK���'�azR��b���ш�}h����
��y�F�zc�SU�خ"�B�&���?��������FM�03�2�JFN�.��@��I~�<��&H�p_V�1�ރUd��C)\v�<��M�3pv�(ہ�RX����4Br�<I�Q�54q ��?��1����c�<�P��+BҌ�VT�4���j�mZe���0=iA#W�YDh<H�J͍ \Z,
�k�<y�nO�}ѲmPt/�f�b}!��h�<Y�o��$0�0J��@"`�$�b�<��'Қi���d��D��! �[�<��+�p�~�dd�e�,"�J�C�<��)I���u�M��T�<�u�T=^x�0��,,�K֋N�IF�@��Ǆ-@ٵ��6X(��Y��&D����l����a���ޒ,V��{u$D�4�3�_�_b�*���~�T�� �?D�4Z�dR��[�ےx� ,�'�=D���vB
3\N��r m�;fN�{&�:D��
��L.c% �Q�@��V�>�`7D��Zuf�$��ĊU�A��X���5D�hN̓pd6	�a
�U�4��a7D�4�#̷+�F�(��&z�Q�
4D����@%�~Y��H1��	�2D���Af��v7�����-���p�!$D�ȱ��7r��q� d@&d��УB�-D� ��A��%��<)I<>�V��D-��W���ӊ,�X;�ØR����6㗥HB䉞I��X+t��M_�]C�'$~�B�	)�Zh"�G�X���W�BR�B䉍Ta��{�� �{����B�I*`���->	�(5�a.��B�I�s�( PbI)oQ:���N��B�I�8���9��x�@9��&�e�f�O��G�� �
�H�+|�4y�g]�"��y5"O��{�MC#���(!l^��ax "O(�
�ꑶT�|q��Ӯ?{��q�"O��PSd��Y��%qpiգ=c���"OV���b�u�Z��0�N!I���0"O^�d����1��&c84��"OL�:�f�1j�x����
(ݐ�"O �������Nr��v"O¸  ÁK��� td2���"Oް� �W,@��G@b-\D�Q"OB�k� (Jo���ce;u���"O2�����6/�>YC���6V�`��"O����,O5"�pu���w�����"O �x�)�*
+4d�P��c��q��"Ol�SU$#y��2"_u��%��V�d��	�>���mN  8����v�B�IFAz�iR�ÿ]�@$㒠�0�,B�I�4>Hԛt��mE�C�6O@B�I�0m�ps�T�C�^ J`��/;jB�	4��IS��aJH* ����C䉧	���u��:Aj&h��g��,C�ɣo�ƈ����'��*�*`oZB�I$ ߂�a�5��1�bt�.B�	����홸~w���W(��B�.UDl3ԡ�n~�YP$�$�B������ODr����JU8B�ɭs��)#-�& ����p"�i��B�6�`UH���G�\)�H�]ȊB�	�gT2�¤J�z|��\�@LB�	�a��A�AA�,\&� ���>��B�I�+}LؕG� ?�Z��6�B���j]0����1°�V>?�B䉱b��%���CV>j=�rg��=D�@�g��z�lɩ���E�Ja!.D�x гh�Ƭ�7K�)�p��SM+D����ǁq�D¹�yt�:��B�I�!r��b��?m�0I��N}�xB�I�O�0$J�J�4�4D�f�U�"B�IeL��WH�!(��1�c��C�	6Ȥ��s���OX!6E��|�B�I�y�d���D�X��Ő��^�*C�I�Z`�4AS9�z�ȃ(Y��C�	�JdF<H�(ю ��az��R n<�B�I�5��ᖦ*r����p��C�I�2ƀlyh�HfrD��ꚙ7�HB�I/3��KI	]r2�X�5��B�ɩKET���1���`�|B�I���`�! ���"�Z!Y
�B�I�l��9)�FM7�8@�L�b�B�%fn��B�.�u�D��
DC�ɞ(�xQ��]�b�t�s7�ZL]<C�	U|&\I�ㄺF39ҦMԏ`�0C䉲: Ѡ��ԙ<�����'# �C�I9z4yAB�B�]+�hҺ]�C�	7\�֐��EJ?IY��VD��>�tB�I(Y*�e�Q���6�V\%���D�B䉘)� T��b�*&��dl��[�C�ɤ�b5�Е�F�b��ww�C䉅��mP5�D2e10jVd�	 �C��&aG��@��^/������ l�C�ɶ$s�!��$&(r��Ў,UHC�	�|w������=�ĺ�P�2~B��e?,]ѧ��B��H �W��B�I+�pʒ��Q��qb��( ApB�)� L`����5^(�� �J�QS
@"O�����M�v���B�����b"O���� ��S�2�@�䔱Rq"Oh�q�@�&B��"QE��Z�n�Z�"O�X�F`���6���C�x�]Ц"O�E���]`+��!"u�1�c"OF�gJ�i>�H1�ǅ�m扲p"O�eR6���F{<a���e��e �"O  �� J?;�vl;ԯ=?�����"O�q���=@�5�g���T�q"O��h�턍� ����7x1� �E"O�)`�=���ԥ2:Α�B"O�DG�g�D���K��`,� "O6|�⏝T@�S��`�R��"Oi��䔸#��E�0�Q�<�NU�"OTma�kO.f�p�s�ʄQ���X'"OB͛w!_7"1��[���"O�P��f$(҈�F�G;J(.ű�"O�A `*�.9��k �C/&�|�p�"O���QE�@�$u�s,� kC��"O|�;�a^3����O�:S���T"O~,Xtf�/ JJuYc���]5��1�"O���C�R�L�\��&�@�3zia�"O�}�� � X��K�aUl�"O"!��̫�b0˓#"�"O��ˆ�1dz�X�+r% �"O��8 �`�rL�D�c}M���S�<��J��>��<�cT [�Y�L�<	����(�����!>)yHp�E�c�<��	�2��|b�ܱh�>��ե�a�<1�X�[6>�B)J�v�ҤQ#D \�<9C%����jp��&���A���Q�<�ÀN� !���_�q9hYqc#SO�<qg��,|�Lp�V��=�}�u,KV�<Q1 �!�v��q`��<��P��N�<�`GȖ#_�8 ���
8�L��k�U�<I6��Z���w�}�����gU�<��N\�R�Aψ'��A�I
y�<�q��8~�TE1�m�5�@����x�<���R��J	@w�T�B��E��F�t�<�V�S� �e؅-� v�l�s��[�<��>Wvz�I�E��p^^Qq)JY�<���1dLlM�t޻r��6E�R�<�'�J��j#���=5��x�<��Q�d���GFWҨ���t�<��	E@� ��hƖ �L�CQ%�r�<�0	C�M�(�"���<YY����h�g�<�e��4d�,�ZdF�&���\k�<aa�1Yp �fC�%���V�SQ�<I�G˪��T�E��y�P&Dt�<��A7'����U�M�����3�!�$�	Oo��ɤ���UU�y����4�!�D�1в�`��� 9�u�Pl
:�!��W�Q�L ǚ�2�\(�ʼ".!���uc�p7��$0�����E!��&(6�C �'����g
�.Z!�$Ǣ��K�;pn�I ��B!�DW7`�s�( Q0z�e� 8!�DH=-y��`�U1������]�!��noR�	�<�&����ׄ0�!��V�v���c�b`J�!`���Q�!�# U����uXt5��mZ�x�!�U8���� �_C�и�L\�Z�!�$-�٣�B$vZ�P�
��3!�� L$RUC�6V�(�*g&Щ~\1Jf"O���ұq�0����ksHѠU"OL5J��];�d�c_=rࠐ�"O%qvL y���aײn@�ըd"OT���b%[���:�V�8n���"O�e�p��ba� ��NƎt��,K�"O���χJ��qz ��Y���Ib"OBQ�0��Sf��eA9?�$�Q"Ol���I�.I�i[��\I��ӳ"O�:�-�e�ĸ�c>|�"O��id�ȸN����Ϙ�YS�ЋT"OF��׮�~�4��h��FS8D"Od=!��\�qq��E)�LJ�x�S"O0�t�ur$Yc6�]� �$�"O�1v�˝>�ZXe*���x�U"OX�k%��J�k��j	#���?�y�茵*��T!ˆ�Vb��°����y2��@A�H§��U�<�����y�L��h�J�z��I�I�"�Щ�y�`K26�<�DH-CO.��b�چ�y2m�9�������@Lj 	R�$�yrFM�\�D����͎��{anދ�y�� H6+�VPh8�U,�yR�N+\� HW� �I6�0�a�'�y�,HS�D�� �Ev�@�'^��y�Ė%M�M�s	˞|���Sv���y⦈:�h@�QI�$;©���խ�y��~H!ȵ'S�d����쀀�y�.^�V�"=d
��}J��;�y2E\��\RF��46�@I���̪�yҡ�d���7A�a��#&C�	�y���457�xZ��^��pYd���y⨔� ��xv��y����L�:�y�i ���gA�Bю���/«�yRD͈\{8 �d��&&��Q�ݒ�y��Ѷ@Hd���ݭ醔1�Df�y��2>��]ɴ�	��&ᘷ�yB�<
K\ڰ$ƫ@je8���;�y�
��tĀJ��^�&�"b晌�y�'�xJju�c��jp���"�M��y��� v�svJ\9a"��	�풗�ybW*�-��@_-p�B�zTH��y��*3jUc5j�;bK6i�SeǗ�y�# �YO�iQʋ T��M����y��Rvx�i�'K4�j�־�y��LN�yb�E18�yy�h���yg��8�*��+�-� 	��y��6�&��c�1y0��c�yO������2z� �A`O�0���ȓ�e@�(��)H�`	0��1W\�4��Q���ƮS[X�ct���Mָ��q�=a��-G����b�*X��h�ȓ}Tn�i��D�Fp`�b[$,ez��/d� 
��
=[d��f��%�Jp��5�Lj��)VQb��ٺ��ȓ|=@�S�4TBhcU���C��X��6XD��ˡ*��z�dۓZ��8��i��K��#�f�:@&D�>(5�ȓ�8���A�,I���2`]�t@\��ʓ?K����F"�
Q{�KJ�}�C�	����ۈy��8��	�T��C��$\@ApSj���81��MjG�C��g���Q�_�e���fL�G�tC�I�2��9� �[4t0B���2�ZC�)� ��3B��9t�H#�M:=f Q�"O�(�C$C7wRE�F��Vl�Љ�"On�j�hT6���0�� ^�eC�"Oj�p��qoRa��0��S��'�ў"~�&��*]�K�D};6�9PRL��Ua%�7�_Y��lCUj�:{T|�ȓx8��	��ɻ|x�!�m6Ȇ�I��DO?GƤڷ'[�na9��#�!�A�,�n5B6j˂i�Й!�!�!�Dŵo�fe!gB\�Lެ	  �U�ўl��ɥ����4�T�z���H-��|>��:�S�O��zǄ$N8�
��.�"OBy��
�H2w�K�Y����"O��u�H+8��;��ڴ�d��Q�MCH<�2@էB����٘t�y@�O}�<A���-�����)p3����d�<�F��8��܉s�ߪ�����J�<ɧIY'"�� �c�&��C�j\k}�)ҧb2P9�k؂��IZ��I6'k���'��~��:L�H���dW�F�$J��6��:�O4k����KR��H��$�4 ��"O�\A�F�_f`lcC%Y�]l�Y��'D�'uհ�-M��ha{�aJ�W�.���'i�d�_�z��d���� H�h-)��
6�S�T��K��x�窑6ċ�G�!�y"�g�\đ5����������y"��J�l-�E�D'Č�Ғ����=�y�cp
���h�,C���I [pzC�I� d>|���5��x%��h����ĝR���u��3dƅ��N���Մ�[*�qDO�#�84�S ���zT��~����S�ORn�"�A��hPqC��--" ��'�D3`Ō�(4��^r7��N���'Y����	T����m3.ʨ��G�KS�C�Tk��H�@�H����ب!J�C�	�;	����[�m;��0A�Ҵm	JB䉘��ӱjB�/�� �p Ҕ�6�?)����!���1��"l���q�]�!��:8��1zV�z㊽BM/May2�
X�\h�#��	ĮY*6� B�I�~(X	�	�� ʾ�¡�/�:���'�O?��W�D����<�c�^� �!�U�Dl����+]�ȕjJQ8/��'�ў�=��	C���u��hzj� $�`��'��`���"r,��/C'J�N���!-D�$9�%ǆ�z�H��Z	x�6�5����	������2�M�1��hzB�	�{dBAX�N�;�t���m�
6�h�=�~�N|��O�$R^{��D���"�<Q��ʛ[���A3��}JƼ�ծz��e��=�'e�H�)�%^��:�'�"�za�'$~!�=9]�\�� ��WjE�W�= �
Q�#�x9O�}��W�:<k�Cj��E�է��jJ������YB�X���`��I�����	"�a�Ƅ�q3�r,*}����Ă�7��O�23艓F�z���h�<a�\ ���I�P8����L��tZPq)c$=��"��$�ƨ�vl���z@|����A!^&��D"O��Г�˚p��P�W�=M���<Ov�'��z�Y�h�� ��^�jw��FE���O>i����?����u�1(���5�1��B�	\�ƹ�F�]�Q`l�s F7 �ꓔM���ᓟq�*�J���I`���f{�F|!
���'�4���\d|QK䢓���+ٴ�hO�,�S�? X)�a^�hF̋�B��1�P|�p"O*��`�3��UbsB�|�j	��"OX}:��KD?{��˾"���0�D8�S��vlV3U�¬Tv(M#��T�L��a�����x��+�?#���b�1��9��	h8�<hreH/����PJ�.A�&ZWX�x�'꾙�u�ҼYԠP&�2:S��'�ax��d/>�hHY��-�0D`��V� Tў���~��ɟ[��0�"�XXt�� �DD�O�=%>�t��d����O�'\��1VM(�	a��ħ��y��WG�C��7u8d�=��'H�x�JCqp)�mC�e	ܨ��	�OZk+OR�<�$�3zԒ���_6ܝq���_���=����A���Y�@�4*j��C�¦�������X��Ӛ}�!��Xo���3Q�"�,@#~j�Γ	Z�r<:'GJ-<
��h`�v̓�?���|"�B��6ݳ�Ѿ_nxlq�ؔ�y��2j�@-J��������'#-e���^ �`�B֤��(N�X�Ŏ�2+�!�D Z$B��t���U�
Q�1
Ҹ1����P��s�E��sJ �C��	���'���D��,�C��8a����j��YZ!f���yRF��L_�Ȣ��6\[�UI�GΚ���hOD㞨&F�z�4��ǣU�
L�� �9D��3��ѨG_�q��ϒ#pP�����8����0=q&Z�j������	T�L��3#�py��|�?�JC��;��}���T(*��5D�,i�W�d���-7,J�����K$��d=CL���U�O�~�HlB"k��H�a|ғ|2׍5�pl)����u���Y2�y��'@NQ�bGI��sE��F�0��I<	������Oh�䙱�L"�>�;�g$��!	�'�}!6�c����D��
�N�3���i�"~� �&��wlBc=����^�A̲,�ȓ@���p�;N`Y$-J��P���s� �Ń� &�L��㜺
����#��0|z�͎�P�"�Y���m�B�K�<aK>A�4�O�S
RŌ��J��:�B�S�MW"�T�X��)�e�	�,��I�P�U\��{�MʔB����:�S�OÆ�Xq�/{*b$څ��	|AHbr"OĽj4c������M.^��A�<)Ó?�D�'�=�T���mV�e�B� :���	�'��ph��B����sj�-/d쳋}��Od����",.�������i��Y�'��?��ׅ��v�Y�����ԁy�j��W�)��<�CT5!�L4Rb�"� T�^��G{���iQ��A� ͱ`n�p��*Bb@�ܴ�~��'��y��"ĵ� 4crNT��T��OV��$^*F�Lg�?:�ԩF#N �!��=��Q#�KO3U4�ȗ$���!�$�%BR�� ��2Hj���:�Q�,F{*�4�&�̠\'��BA�22�h3"Ofp��*�Y`\��U��a�(OL�D��ORE�r�.�ʖʏ�*�Ѱ�"O�ɻvd�Ą�X0�B�]�&�"O��9�	�}*8��%a�?�v 1&�Iw�O>���BO�� �H@���7[S>e:
�'�U"���z˞���[W���ə'qў"~�MX�*��ͣq̑i��rug�F8���~��*edzH����5y��9�T�1�y��	���%�ٸvO.�p����HO|7m&�R� �'��"9S��z�6��������ቯ]%�i#�)ݾ^�标��4"##	W)�E+�h
�7�f���S�? �,@�E�}"<`��M�Q�����"O�\B��@�Z�ҹ4��*� X��"O~�p�Y��zq0�'�Z�ȩ�"O^H��S>����N'KV5�"O�r�nēC�`��.Y<cb$�w"O��
q��an�S�+V(	J�0"OrMkf�k�yb笏(9�-��"O����L�Q`�������W"O���̍cX���P��W���G"O�$�'�
f� X�D B� �Aa"Ob���*ԑ$�<H�4m]�E�z�;�"O�x��c��Bfn<��V�B�U�"Oj�b�(2#��̹�d�B� ��"O�	�'����е ���"O�D׭
a�d,	bk��t;�"O���p��7�X���ٽt�9�"O6��f��?;�0	w��}�&�p�"Op�9U(c"����29��	8V"O��j��M�,�	#`D��|[�"O���q�i3
8�b��;jH�Z"O>����_�Q{w�L� bL�"O��ɷᝄK�[3s H +R��A"O�q��\z�(��H�;@f�:"O�ɛD�@?[*�)9��
�W#N�a0"OvP�H�=G�l�� �i��MJ$"O�l�MR\. RQ� �H��"O�8��f)p4�3��-�"u��"O�S�cĔVf��Xg��G��u��"O�B�,9��[����U"O:1�Tf݃#
1� F׷$-z$"O�)A`ԽN/ y%C�3���y6*OV�Y3�+g�8ly�+�=r��
�'!��ئ��/^l܉�F�?Si蜺	�'b4irbP&K��U
Da�R�[	�'f����
#qQ��ό�;�`a��'�F��D&����z��w�����h�<���I��T-* )�:_��YJpPc�<)�NE/#Y���&�ڰạ���^�<	!�B|z�o�a%�<CፓO�<�t�מ6Qb=�Pj�)H�AQ �Q�<�c3���Ú|�1I��K�<�A�:�V��#'��8�Z���f���� �D�:}L���M�M���;qM��4� �b��wj�ԛE�&D�8��.[?	b<��Ӭ$��<�a'D��0����-���p��E��V�"�E%D�l[�+�5	�l��Z�a��/D��+�FS�F��I��v�,D�$�*D�� P�m.�r��S�N�FԁF#(D�$r���S��!b�G�q��D f)D�<���u%��{����dAA&D���d38b�ѾR���i�)D���5��@Q�5xUF@�Y�p�c1D��!���"x����)I���I;D����"��hR��A͎8�6M��"8D�`1T遂|+4�!}�
�ۆ 8D���7�_,!SX�+H'V�6D�PJ�<��(��ǩ7븐�n D�T`�,͎@F�,aG+ŘB�����%D�x��	�)2	�)2�B�LpZ��B D�l8�U�C�@|��a�:%-L��G�2D��00�H�@��#����M�T�Ī2D�L����$G݊@rD b��]��N"D�|��A5�� ��~���:�K!D�L#G3Wt�hɰ�	8���H�M:D�� 
�f��4/���(�ܔBr��u"Oh!լD�d� ��EW"O��s�"O��󢎑P�
ĺ��͏BH(�2w9O����,�p>���0
�j|ӳ�?r�ƨ�5�]���3���XW���.�h��4Dq�2�2U�V�/ؘh�ȓJ�d�i�m� m�L*�K��B&��>�FJh$!��-ڧ1d���' �xlj�.hn�A�ȓ��=ql�c����3\�h��|i�\b�j�(N��ي�Y���"�C#r�����!d��4��.)D�D�צY]�ҸCݴwx���T�{�� S+^q".���/PNlB���i~ �c�5蘇�u+��9��ǜq\���,��L��m��b�@����y��B)s��Չ���3P
��!ᭈ��'rBd{�G�)��aF�T�ۗr|]��iȇ�������y#��AUF�R�KF�n� V .7��H�e�+w��?X�>�p��� �8��+`��S�ظ�ȓ?~�w��;,^<��R][���o #��H��uY�{"Q/;�֙Z��/w���IƯF6��=y��f�bl�'�f�P�cJ2���b��J"Z�'}lՠ�G��ڬ0�e*۰L8V� ��$G
��Т��I� @��G��W4R�0i��{�!�DL�(���G(��.!lQS�����!���RwPy�5T�V�0����/{!��"����ʵ ��A�wkB�M}!��ԮM1���d
��"$�[�WR!�DS�	�mx2"]�K㈄aԉK�|L���Z+����w�Ͼu� ���%��y�.tZU"���E��E��+K��y�c�%%g`� �����ӑ�Ɔ�y'\6�X�{Vhq \��F��y�ƚ7xh(�
��~D(
6���y��I�z���BiI�h�ҹ�����yb!==������D-c�Zh��:�yR�ƯlV��3��͊ieJ���y�D�!�b�q�>lz�,���y�+N��)5Z�XE��"%K_�y�NQ�D4��A�I�:\�\d�C���yR뎩&a������Bk��3F�Q;!�D�_��/{��M�dk��=�!�DJ,6��g�V}��ivK/D��AY|L��
�������'$'����1Lx~��I����್Xf~
�U���RcNL .���QM�~�<1'g�,}*����ڠr�✳P`Q�s� �>rs�?y����Hex!�VA] ��=�u�=D�`ZE�A�raֱ����	����Vˈ�P�48O�l1�S�g��ȺR�u�)��s�p�!6}
��J�RW��`0 >3JNe�d+@-P��aեO 	��#����?3HJm�L<i1�R�6��� ��o �	�g��@x��(a�)h��GZ���	��-WMQ W,=�$�'<�$��$]p�iBo6��iM�X�c#mٔ*��y����;��'��e�&e�8���&?}�ƥK;��)�>^k�0;g^����DG���ϟ/��I�M1|����|����L9��Y"2���&� $^ ����C?}B�P N�d�	'񉚡�l)��㓫z�.YP���v���'�GZ��w�Ӓq�����c5��
c.�*Q����&Xf�'V�d#�'L��  l��\d�����5&��h�'[@1hA��65z4] �e�:v.�ӓ=�&��b�;��$U$�X�R��Q2y��Y��-��
,PM�p/U*w���'}�~����>��ҵI��� Aџ8��qW:?�6�G�������a䈅r*O�e��N�*��S�
�V2 �xrB�"hY2=b%��Д���g��& B�'0�5C1��JJ�D|�I͑xex��BL��b�|��[���c�\S`�ڿ"��4���ƙ*��8N?�r�԰�8ِ��ʃ=B��Tl[Z%���K�a~�"Ҁ^+q���C�D��'�*&':%�u�%
3"t0���>~G���O�<Y���Bc����'9�=��t�LU9�˕r/�h+
�':x�{T-�+K;�[؝c�m�!r�+���(N1 �Y#o�;cӊR�x�ޫuì��O�5��m̈3Q�41�( �v����'S�(a���+%�x���_��� �q�I �v���&�)b��D+c#�5��'��L;Cc_X�'cJ����F.,
��Y�#9*��I>�!Y�&3>��a��-z�r@bP ��O��@��pǒ�����%�Y�	�'��|�D$K��`pI�q�0(L�J�j�a�����e�1���O=�ɵ3������Va��'샋m+rC�	�&s�-��¤p���'^106�yr���"�,H��/hz�s�'�2雃"_Z\x��W(�oݎ�ד������O�	ۄ/N�K�t�!	�	`�ؕ��D,�l��'�vܡe�\, �,(�h^�c��:��Ď-A�h�E� �ӫ:��9`�!Y�S%&X�wDٞf��C�I��TmG	"���Js(�"B���ɧk>F�E��BX�S�O�J4C*5�=��"�|D��'�4H��sM���%�"j'9�M�lC�KE-@�^ R��'��:�ʑ.X������ۈcl�	+
��zǄ<`j�;?*�ڑ	�/���@�*2t�˓�2�D�i�W���Q����rvႧf$��1�/X�fJ�c>́"�W�}/�`d�ߞu�<�ku�%D��qg�O�NWĤJ�o�
=���s7��|�RfT�x�B��ԗ>E�䣊<M���P�şh(D,�sM�9�yRh�5r\H��^(o,R(�Ӯ����	�R�H� ��q�ax�C9�D�3���owl���Ν�p?�S��~�j����	6�D({�e3���b���;[bC�I']�4����V�B����A�y�|�M>�����{�֝!Lg�}���BB�i��W�?�����! �{�G$��J�)��|8a�2!0=����OX���N͆�n(s1BS3ɸ�(����G$;Bj�ӣ��n� Xi5�I�]�Q������O]��c�Fؐ	hX�e��9՚#�'�t�+Ʈ	}�\�!Jk+O�IC��6y><mPp�-����L�Tf����ˈ��g"O|�V/^'|���`�'"� (����.c��� ���b`�|�3�I�h=,�:�~�8׋��X�A�����p`
�!ưl�6-�#	L5�q쉓w��$B��'�O@4����Ś<���� ���_��$����	Z���=��KA,�ά�4GXT�����o��kHt��e�ϳJC��*)u����x"�*VV�$z#�	���TS�0R�w�n���,�P��ӥ�DX��2O1+^��� �E	;W~��A/���(ȥŞ�aQZua&�)CҰ�Y��@�|����%Ud���
-�>q����/��<e��iرO@ݡ���{Ȑ�����9!��0hT��J�0܀��I�xZ��;��E�DՉ��y̘���I8"��(X�'��)��
L�c���fm��0�[�F��H�4a�:5/�b�D��NL	>��� �C�nk��|��aq�^�%���שb�:u�Wi��VR�sR�^����1}��O�*+��a���=�D��O���P�HU4M޽����Ce̒Oک�0C�Ei�t�	��PM��]��ħ�a�oV1 �D ��"p����qa	�d�dD�)��J'-ϭ�u��O#�Y�VƑ9oup��-��A*��,f>y�eI�S�X�bq��&+�˓$ @���ܴP�F�*�͜7RU� �88��y���?4�Q1�U$�����*ѝ%�|����?Bu�@��y�Q�
�! ��i
�țb/hH��N���� Ͻ��	 >��c-��~[�]����hT���  �%�2�+G��+G�=��� 
8lҺt�B��"�>�I�n� �W ̈́�������7�5�I� ��0�r�x!��jSLѦ
i�P�+���؇"�.4�U&�6�|���L%���J"]<���-�q%���R��.�m!�B�O���7�Zz�EX�I�2{{
��!/��}u�5�G���D���g'�;����O�Up�I�0~p���w�`�K��N�#o���$�/g��5p���96���O��K�����[���N��*��F��� �ݨ64x��E���X�-��	�̑�`��R���j���'����Тk�V5ѥ�B5Ul�q�
�0n�%�vM5��4c�j9�m)!��q�&j�,=kV]+�m�2/��4��J0���x�,I#fY��WȜn�b���S�.���:%n�(����$�Ă�����bG�UBt��b�(�8/z�h�!���#ˆj��ф'Й؋A h~��ȓW4H�� G=L�2�;�͈����"�Uu����ӻuچ�@,U6�S&f�Ѕ��t�n��WO �bj�$�թ�A�T��$܎+	L�:� ��DptQx%�F���P		����Bķ�N��"�?o�0HBƼq����	�$���s`�^��pvoQ���$�@]J�y����>�:0�a^#�?���X�-Y*=Z��? �l8C�O$g�`��R%Ӡ3F��;!�'�tP�aW/n��9��A�*��G�wx��6��"�aY��Ρr�rX�!W.m��Q B�B��w��P�d��&^*�{��F2m	����'5p���
I�xqK!o���6×��ލ�t�V5#Jq��AJ�n7r�갌�Ȧٺ6����0Ty��ƛ��W+lU��6 8΀I�fC��=�v`�5��@�e�]�8-<�ZBX�)@��hSoԗEZ�zӵi�LCseH�lb�H*Zj�l���q��� �!r1eQ��,�K�> 0���s�d�5�찻v�D/B��$C-c���#۟��JC��O��=�#�!2�tp;�۩5vȵ�d�?�O�)�ǩ߷J���e,�4:��( Se�{��Q�4�PX�@��L2Q�>���'��)��:)^V�� ��.gfM;	�'��9�#��tD�M����) �љR<��yஇ�rݛ�!ѷ������ C
��g�
&a2�3�c�U
a|���8�v�B�'��3�bϓN�\:#���U|� 
�'������M��,q��˦&�& ��'�~���ɂyk8�,�����'���zf��m'�l!M��l��'7܌���>G7c4G^� e���'ޮ|{���?<�1@c�	�|���'O�(�#�C$$d>]j3�ҹw�,�A�'ǌ!�t�J&
�T��Ӫ�/Q����'0d�a욘W�A#��DB�
�'��1@hw��E�V��̴�
�'�z�R��"�4��kK��l
�'����c"�O��8[fG�(¡��'�� �&�)q�^4%=�4��'��� ��kMl��l�& ,��
�'Κ����ʑ,c��D�:|��$�	�'`�-+�e]�h��HC&�Y�T 	�'G&�1��?sw�����E�U�<�	�'��ũM+n�>�"!D����'���v��Ö�ҐA� -h���'�ވȄ�	�d���GkB�K)0�@�'[f�b�ö3�d(�w�œC�����'ӺP�ө�!�ȳ�#B>,�@�'L� �#c+Ь�bvO��<���
�'"�z����=E�D�&��DS�i	�'0h��.�J�r�:ņ�#Kk�s	�'���KA �%dk���W-M��Q��';��H���r�.͓�@րM!na[�'\��[��92P�zgeW�v&���'���iv�qj�QswIٞ&��P�
�'(d ��[��+��P�aO�yr��zE�䋂�	LPa!�?�y`N�ʹ�Гx#�0��yb�	?^�u ���hv�a�"���y2!H�~�1H$ː��J�	A��ybɂ�{��%��挵 ��\Cნ��y�AW?�и�%�֭t��س�%�y��X�J�h11�&N1`s��c�8�y���<l%" 5G�dn�d�b��yb`B�	�0E�Sf�4)���'�H��y��	-��(�c�=K���6����y�=u�Y�㔡I��0�0 Ə�y2�P5=��#�C�q�Fy  *Q��y���VM����턬j�L�W-̹�y2�<Ubx��I:]�20C�j�=�y��A*�s0��WϢ%F���y�GK���SS�W/bX�eI��yb�-Hz)p�.�D�ɘdn_��yR� @s�]�$��)�9"wE��yB�I�H���5���,�]u�=�y��'�M�r���T(V�D
�yr,ĵ,�X8*��d�*L�T+���y�JK�t��@m�e�NAJ�&�&�yb�-uN,u��	�K�RXQ����y"%�/�M	2/�Lc�oI?�y���8O�pT�WN��(:�9�Q��4�yB��g��SŅ�tz�`-O	�yr�#7�`���O�l���!��y2j�*Jڐ<�
�u�^!�����y
� ҜZ�H�<Y�I�
/MP8�w"O���FW�2���ꎉ l�R"O��G�e���3I�1I
��"O�I �ζOn*�@���,V
&Ia�"O�H9C��+Y/V�k"�V�@x
�"Ob�� E/GR��2ȅ4"��@��"O���A�sʆ�k�C+=�� �0O�(�,?�p>A�����pYA 	J���C&ǂ���(�l�fv(�ϓ{�M�j��+��T8��
�\T��DxT����
 he�CL�9&օ�>3�v&�yU�*ڧ �UXR� u:�3���h/6��-���q�1$��AD7���,"�d	#I�����Y�jP�M#fl)�� ǁu����� D��3pcS�7 ���@��q
��I��m�jxRP����<���jl�A��L�y�M�K�>9��<5h��.@�aZ��'��V�^�Q� +§r�@	�'T��+v�ܒP.`Qu.�$Q�L�Y�}�8V{�a�wXE�O�yp@՟�`�[eDW�^�Xբ
�'���h��Ѵq:�<˓,�U�a��
�3PU;��>a��>)���;"G�d��G�_�\]� *�N�<��(^�>�C�aK ]��!Y��;& �u�<x��'�r�@�c�70T0�B1;��<�ߓ3�( ��HM��yR֓l��UB�)U�2>"�
�lߝ�y�Nӷ ����̆Z�����A��O�(, �a��I��Mlz����1D\D��eńi`!�db�vEy��4?1�X����T!�$_5��۵압	6�E��YY!򤐩J�=��)��/q�)����x�!�r�(l��0on�|���T�%�!�Ч��}A	Lu�(;���8�!�ϩ�yP5&E�#�dŪ�.�*M�!��Z���Ώnܨ���#J�!�T�1ܐP�ek�"�$J0�O�r�!�d� e��g@�x)��q��H�8p!�ħI�
x	B��S%n���E!���-�,�Ӈ%=b.Eٶ�<@!���I�:6�Ҥ?�h�rЉÙH(!���Lh��s������c��!�D8l�� 1���C�P�����q�!��"�,�A|���[ы�?F�!�dPsW��6K	��a��A7��d��L�d��eQ@��4G�	�yR-�Y �Ⱥ�@�v\��S��
�y��;}-��� �����K�,�!H<����
��0?qQ��b����6�^�D�<�Q��b��|��X�ؔ'��a��
b�E�c�0p(�=��'�X��eG�?F�ai3.�5{�,��L>a�
�x�"��$�%�'�Y��3-D���E��N����ȓrhi�c�O�Ɗ��䄻SE�q{��'?��v���G�L�kB�J�z7�m
3��+g�pY{�;4�PIs�W:�u��)J�M� �Qd�66`�(e�Xi��d6NS�dzM<���2�BXP$
f5��qx�PxTJ�j))�U��b�S������GBz�bAD(���*��(���Pq��($)�,&X��� V)�'$R���S.�$?��'�`��2���Z���Ev��eT�0!��d��0ȢYV�"�3���#�ub�C�'p �D�E1(xIyr��g��L�`N��2dPb��(���eȡ	5he�7qd�q(g��KF�E��cЃR`y���lt�8��!ޑT@���]4U��X�O�����O�ա�-N�p4�+�"�l���O����MȈIW�M!��ұq�'�"��V��^�剕}��& Ʋ'���Jg�ֲ`��]ɷ��k
t;�JX)pLx#��>}RU�W��z6��?"$Ω^	8� BXA0H�%�=�I�! ��^� 0 ,���P���C��݉4F�/{2��c��?*�\�҈��Naz�OP|�b%Y������.'�h&@�=/�A*X	M��'�YC�j�H�TP�"��c����~Ҁ%D\J	!V(ҹ���F��O��a�a�&��� 
��&U<+z��3 ��C�Z(�)�+mJ��҇X:N���	�G��	�?��(/M!���V?6��X!�]�KR��A��G2==����%��"�^5�4y��M3x� D��!�!}!樺Ń�c���I 񤇑#��9v/�����béj�P�����ND�@d�!<OT�۷��HN�\:A�8 .d����Rn\�0��7��0�VhI�)8�O�8�v(���O&��/R�0D��%ثrQ�d(f�|"�X�v[�Lh��2�[A�,R1��)k!�I-k^�ҷ��q�v�*�"Oh|c�@Ɲc�|� �U�w�hh�k6E`�)� 	6�Vjg����N�?u�0� ��e_J-�*@L��ȓ(�*���!� lmt���aX b5��B)�<: ��f�)|�vc,O:uӠ)�7=��I�JX�d.� ���'��6c�˟���&T� I��'!�mRՆ� �~�QO�I�bђ2��H)&�T1�d��	������
qܧt�n���Q<@,�=� �Q�����ȓ��B�D�J�)���_�P%��'x"M�E���2d�ҧh�z�Ν$pE��zE�4=~H�"O6�!aC\5;8|*C)�9C�>��8FC�J(O���''?�")�3h�f.<��W�'��I�7���<�VLZ�IZ$��l��1�d�AoCA<�%vw���5j[�B8j�HS MX�'S(\0�'8\��m�|���U,�%:,hw)�V�<is�ڍ'T����L���)�I?i�F%h�P�-0}���݂w�h�+'���|wVx1�Ψ!�d��*��n�~~FX�%D� ��K��RLJ�kE���$ͤS`8����ʰvy2���d��=��~r%ϻ7�@���.*k<e����H���@��N<y�F����FƢ��L3�p���{uFtzt�|�	zwB|�;(v��)����Ӻ"I<�$�F䈾-���k)�k<�S���(�F-E�nD�GlD�b�t21��h�P�qQ��4{�qOQ>=�nv��z����=i�9��-�EVB�ْًY����ϟ�,�F@X8�옲�KT��8�"O�pb�����2#O^
�s�T�$8V�K�9(Qi�N�R>� W!
�Y܁iB�U�J�BB$#D�$ ��l�d�����$gŀsD\��H8 �����g�2	�Hɖ��1�,�����>x����ɀ0�x�ר5I|�3���%�^�;qn}�Ta�aW|�'�$�Kr�U��T�	(�I����"B)��J�?����x�@@CL�Di@��h��$��
XT��l 6)���K��`rJߝ+~b�p2�
.t��&@3�'b/�eI��<HS�)��l3�r 	��L��T%i���y�.�S�Og��h�'��Y�1k�C[��H�5?�!h^$���(�U��a���M�g~"�%��D,L�<��up�ֺ~B��p�� K����3�in��W��&�ўHK#�� -"�D`�T���"A�6�%����&�D�}��.U�.�k�$o��X��H��g�� ;D��_.H3��z�~�R���0ÈO�� a�o*D�S&OP��趁��
��L�An�J��H@�/�$��I��x �m�x��lL���L|JD��,<�L,��`�r�Y�Ɉ.��PٲњB��i1����0DI��
�5������0��!M�]剌'\���O85�So$?m��K5J�
>D �`R�=�>hʃ��>�q�H������S�*�b&��^z���8O_)�)�.`�9���'|O6U �m]�hȬP(gA�hq(L�"NC���F,�w.8�>��!]����AG��y�d�>"F&���NJ�y(��D�=��<����;z <̒P_�=I"�w��%"�c�z�x�kJ���p�@���:-'yr��	R�~�T)P'H�c�H����Z=A_�'�L���$Z?DU4�ۗ	5�'5m"�1�h��I�l
ÅI4κ1y���a�4�'i�eK���!�GN�}�F! ��Ey�pL]}�(�'-TB?�S�Xaﱟ�'�\� �d C�`����H�=��%c�1LR T-6|Ok�L��YI$�X�Z����0\.|�A�XG�J%��%�O��!K�6 ��0 B�V^er��'�L��*BJai�齟���� �\���F?<�����#D�d{��.���ge��4�(�2�>}�o
de�a��l<nm�?mc���*��q�a��7+[0��ש?D�� W�Y�Yqt����H#�X1�F�t/�a�-O0�[e������|��X�W9a��Q��"mi���?Q��͙98�(��ᓟ%4xQ�� ɓG~~�B��A�yB��&�)�G�NX�P�u�Z{�٣v�ʩL����ʴYPD�ŧ�<���T����?o����t�ϫ��� j�J�H��Q�����qZ0��"O�=�r�ÄT�<,�BVg�Y��iW@P�0�T`�N̊���Xʤs.O��Q�.�^?Y8�cA�2>�0@Ç��,0ea{�gфo��<���ͼ�MSf��u���F_��I9 i�g��XO���2�������Ia���BA��/J2E�Wa����>�UB�F42�9���E�O��U���"˜m��#��<KXL�5�J�0��'�ȭR�ŒV	�S������(@�J�1%1?���>����B�V9�ď�r�&�"/}�<�$ϡtC�,��ƚ^Q�%��E���bGd�[j�M��w<�C�ׁ)��Aa�OZ�_�����~֌�5}�RU�Z�B������w��E�F-:D��7��<%��=B���[1N-)uN5D�@�$C!�}����I����?D�tPW�#90��ۤcגŁ�(=D� )�N˳â��n�<*D�ũ9D�0�`\4e��% ̭rg�ڣK8D��bR��+v���0u(��aH�d 2D��跮4K��q{�˳$��,2h=D���sh� �Q�gӶd�2M���,D���t�	�@�$uٷ���"�x�IRM$D��)��ѕ6LP�{rbY�8�HU��g$D�dSQ�Z'O�t�pu��	� AI6�%D����(�qׂ	�_���c$D���F�]O2i�1(�+��,hwM6D����U
^���TMԡ�Bd���5D�L"�]:p����6J���?D�xK�b��}��qwoB�XHl[�;D��9�T8P�Z�t��*��4vB�	H�u3�I=W�%xq��:~�4B䉗H�ֽrpm	3+fi+g�ԜG6RC�	�.��@m�,}Z��v�ӂk�
C�ɣn���K�-��]�:X�-���B䉷�8ŰG��~��CE��j�B�;U�p��v	!�ՁT�T�`B��%�p$)Ӣ��.{ڀ�$� *Q�C�I�ZU�<(��b���Ӱ�̙w��C䉢O��YH#��c�)xt�K��C�	�{�F]���Q�#N��[c�[u�rC�Ii|u���2L��8�$L:dn>B�I�A��h�	�9)��c�,Px��C���n�	p� 3�X�2�3|��C�	 �\mP���|J\h��˒�7�B��_�`q���:m��}�3�E�-��B�IM�\��#��V2�M	�oC�r6NB�	����[�.��"㬽v	.C����,6����q+V5'e-&G��$"OB�S` ��4ގ ie� L�	 5"O�lx�I�!l�Z���:;�ձG"O&��]$#�R]���Q$���ӕ"OԼie����҉�U�ʭ� �Q9���AY�(�V� ��'��!B���,l\���[�d�6Ł
�'�xU�0,�0eR����Q��	�'H8%���9,�p��#ڊ:��,��'0��q�G�{֕XSOM�.q�Y��'^:�`��8n��ū����'����3��0�BjF)���z�'sޔ���T�;t)k�81�,�r�'HXġ�A
�B���cI  &E�Ի�'��ճ�Ќf�0 �X�r���Y�'a2�J � �]%���Ͽ`_�Y�'���J�OɊ�.�XV�ёU�4�h�'ʜ<KRNT�T��� ��q��
�'�����ߟD�,2����,Y��'i��1$A�<c2L�
���
���
��� =[F��(b!�p���ڎv.F���"OBtҡ�ްg5�8���E���q�'��	sF�>9���M3�ӎM�l����5B3ּ��B�z��iS_<��'�����O*(MIW�T�Z<T�z���=k�(Ტ2}�{�"<Yҕ?�X�����o�kv'��N�����~(,��v`8fv ���ʔ�]OB��S
j�W��b��U���� 8��H���n�V�(�pT�F�a~����0|2b�_�mzٓ+S�7� e
p�@�#W�1�'n&E�����On�OO�I8�D���`�9S�N?c^�:H�Ġc�Vĸ�e�O,�P�7�D~�jר	�*`�4��O
$�3`;FLQ%� Fx�/@ЂB԰W0^a3ÃK��y�Ɛ9�:9R�::b�`��y"�4���	��"-	N9{����y��=������%��DX��V��yB��8���S�ȍ"�:Y���_��y҉^}�,�ě�FCS��y҈)�⍻������W�y�N��+MӃZ�����Ɉ�y"��@���b?H�rTzp��y"�#K�������8��`�t�֨�y��� ��,qd.�")28���ĸ�y�=:�$]����4�{�뎌�y�S�Ɛ�e>��=Q���y҈��/X����Y��,�Hm��y(�8//J�Ѧ� �@t�#�yB��Pe�p1�[�s3������y2"��p`���
K�A��)i��݅�y%O�ZK�tl�#lDcc���yR���	�R�Kp�T(�fX�yrJ�2Uީ��EE�ZMD�yB$<W����W�QLx�C�ء�yr�Uu*��FH8�XS���y¯��H֬�SOH+=��$8�O^��y�`����GN�9O~����Q��yb!^8��@˃�3/|�eR�M)�y�D��ѶN�(��dQX=�yb�?d���ŵf(@PeQ��y�h�p����P������y"-��p������7G@�՚����y�]�=���s��(CkT{��X��y2�7dj�i�,ǚ	��Z�j�4�y�ŗl�5i��ƕO{��귈���y��9��3���}���2h��ybnľR늴�&Q8?� qQC)�y��X�|��]��m	�0w d��S��yB�ʱp�em�X� �*�&�yR BU����wBM���w���yr��r��h�q�3}u(d�QK�4�yr�Ĳ� hD/��	��� �c��y.��eR��˝��ɹ�IZ��y�I��[HbL��
�*���q�ݫ�y�� ���"(�,���)'`ƴ�y�� iP�!��B�&�̬����+�y��B3Bs����FL!l����)�y���6�`�U��-���a*Ϋ�y��ɧiV将;*�>a� �E<�y�M�?�AX�̚�
�<9�-��y�����f芻M����Eԏ�y"m��?:�M*4*�F�`�7M9�y�ɓ��z$���H�>����W)V��y�n��llHQ��H�7�H�`���y(�,M�`§df	
���6�y��H-u�}U�ϳj�pk��B��y�'W.~����N�h��p�T�+�y���*\д�"�Wp"���;�y
� ʸa.ճ��Y�)ܫ#����"O�H�ĸ`E�`&��(*q8%�"O�\r��� �b���V�"O�3Gg�?p[ �pth�A'�e[�"O�t�P�	`un�zHȊ �Q�t"O��" {���2���~�V��"O@�6�\�FɒQ��GW8q�M�c"O�1D�W�-4z�j�K�B�ٲQ�!�Ę71wd\�3��F��#���{�!�"f:�P�ߩ�X�!�V�b�!�D@!116�a⑘(�\�VbP�o�!�dT>-�Ե�d�](b&�Q�#՛m�!�䟣2%u��-ِ=��k�@��T]!��l�,A�kӖe�1�Y�V!�D��K�J�`��� A�^Z�-��X#!����x���Z��\ȡM�!�Dߍ"V��0O�a��г����Y�!���2��h�2��O�x��Y�x�!�ČvX���0f�PR��H_!�D��!xr�sū1���Nʍ[A!�dߢm�D$��AH�m�t�`���:!�/'�4�΢ZzQ� "�<!�$��T��(�Z��81�6"^�^ !�G=T0(ѮS.h��)�G!X8N!�D�-;:Q�H�u���	��!�Dʐv4j9Ӓb�8|d�6�8 !� 3k6m�c/�H�1!�^�dN!��$a�bE�	�]���J�gN;.M!�d]�u��E�%U�j	�A۟rZ!��>iP�
�@ث8�abGG!���Np��f�ƹ� 
�wW!�D,7�&e�m�?/y�u�tE��!�d��H���;t�N�(N�䂦D��,�!򤊴��H��ץB���(!D��/!��Q'mJ���J��8��}��җp-!�K0bb�s@�z�VI�+K|!�䂢'����Dvݖ�#��W$
a!�d̿K��ɀ�%�/*��0؀e�4 !�d�6*��a{���8�r<I��̫<�!��f<�+�{�vCtiK�4�!�d�=%��;a�D�zMx�����!�DU�;½���(�J��î@�z�!�̃6�$���B�	�Ų�E��!��#PN�Ԁ��Tk΁S��Hu!��#X�J��ĕg^�V<x�!�ф5�Q��]A%�h��i°^!!�G�@/��뒁�6p2�)�1��R
!�ڭL��t�"��<G��s%C�L*!���TX���`�$2^��(/#!�;B��P��L"t��6���Q!�Ć:N
J1,�cd�,!3�$(�!�?�
p��^xTH���!��Y3*̔��j�@?�{���T�!� -�I�4�%<2���މ:�!��9>ѐKe)@�d�VA*���o!�D�X�|H�pA�?k�b���.�
!��]h�)�A�o������5!�B8i���1�ʝ'"[�ŉ�i�%!�$�Qz$�b�
��E���8"!�d~���0�%U>������D\��'!��JR��{�l͠V�X�:���r�'2���Z��t#6LϷ6A�Ș�'"��ځc�=���o�"����'\�}�����x>�c?�֘H	��� �H�kڀH���S��.5L\��"O�i �L+}���	�i�g���b"O
d���Q%t���qH����I�$"O
]S�-C)Q^�ِ�Pl2�y�"Or�lވ(z��ּs:��� "O�)7F�1(�p��C�RO�2s"O�I���	�F=�8r�K�$`�y� "O�E�2�׆�+�j�7}#��z�"O2����6{��:c�	
�� �"O����X�./�qq�Ƌ6�t�b�"O�0��V:?�&�Y�*.(����"OJ�A n^=Ic��l��}��"O�8�3f"Sr��x��$:�켱�"O�0�D������FR����ge/D����O�d�Hnت>0�q/D��E�����*V�T�{�H�$�.D��a�CO�3�̭�t����eB�+D����k�D�H��kQ2J�a �(D���1+����rf���X�AI!�'D�4����_Az��!Z�ԙ��+!D�<�$`�)t�\-`B熇Ϛ�9�#D��ÀA@�;�5�_�un!�q�5D����@�-yh�*4�ɥ:�09k�N0D��z@��\�va�a��7i��
@0D�l�0��+2}N}��D@4U*>�ȵ�#D�<pqC3u����_j�RyPC%D��*�ꏐU�Rew.�^ak�o5D�p���[�${l�;�&A�]�(��� D��(�I��J@V�)��ԄJ�D$3!A>D�(I�"չ}�~}���ϔR�@ i�<D��YwA�9b��u�RɊ��~��-:D�Pc!�ؓl�=�kP^���7D�H�0M�/I:����ܻut<�#�7D�H���Ϗ0�|:Q+��%��\��e4D���2�Q�kحHab�r���"3�3D�T��/S�����&12d�94�#D���v*̑�`��5�� %�Eh�&D� "é�; |�Mk�C%?N}[ņ0D�������c@UZ��m��̭��y��,\F	��_�GO�����^��yB�]�[�Va ENU�v����B��%�y�+*�<�cЉe��� "��yz7�l���-_@K!��3�<C�	W�H0�BZ���o�R?C��-Lo|����@��)��N��C䉔]9��"C��v���0xέ�"O�؃R��1x�P���c�$�`)�"O,��R�Ȑ)�X�Ã��:�2h�"O�qCg\�.��x�[�\ϐ%hF"OT�Ä_�Z�����n;�L��"O���@��:3�:�Éײ8����3"Oh]�	E!|t�Rp�&�֨{6"O�����q@�PR��O�1��ea�"O�Z����u#�P�G+*m<<9��"OjXғ@�_zj�J�(�7'��b�"O�Qq�ٜ-u@iQS���W��x�"O&�&�G�Qߌ�e�E'S�l=r�"O>����>b!Z�j��D,�8h�""O
�� ��<]A6H�����"O��!r��G�r)��&f�$��"O$���I��GV�r3(�$4je"O�[�閆z����d&O�3�4P�V"O�b�*�}@���R����"O���7+˃{��8���=]��4�1"O� ܀9��H�B����;Q��C"Of4�7	R�q,!�ʛA5���"Oz�*6�˿��̢�\LRhq�G"O�l����g���8d�H�z�(H��"O�)��!��j�}��CLkf�"O�!�C���:�v�Cq�&$WBa3"O�j"A�g�}�GQ��^��d"O$4:��������7��}4"Oةi�.��>�`���I���"O�;0��	�Q�I��y�c"O���p#C�p�~��HE�mP�1�"O�t!x���F�'=6�]*"O^�	"f�-"ek�T҄� "O�z$oݰ4.�#Љ�b��(�"O��g�*9>�]� ���C<h��"O*�8�   ��     r  �  �  )*  j5  �@  SL  �U  '^  �g  �o  7v  �|  ł  �  J�  ʕ  +�  ��  ٨  2�  ~�  ��  ��  B�  ��  ��  ��  *�  m�  Q�  ��  5�  9 n ] � �" �(  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��l���_�a�)�Y�!��-�	W<)���&M���#� Z�kY��3���p�<ɒ�`H���p�ݎNLJ��m�l�<)C+��5���k��n�d<V�o�<�Aa]�K|-���J�ș:C�t�<��E<�	��I�����n�<��K�
Z6ͣR��3�&�Y��T�<	�F��l<�p뒔g�zhz��˓Pn!��AbM�#& W"C&)ӧ�ܡn�!��;
L���WQ%�=k*�,�!�DǨ0�4���jR�[ �&�Wa{2�dF)�bUY�C�,_+�	i�E�xH!�$,&Ttx"���C��yuk�'[�Ȣ=E��'����BAA�9��m�F��o�@��'ζ��1Ǘ����E��^��N����2 UkW�^	&J��*pjѳw@��=����y�ÆF`R�ʵ��%Pq@DJͷ���0�Oh8�ugL	Vm�E@�M*Kx�[�'#��P����'?����*m@�X`!�;D�$�j�Sľ��"�R47�����8}�[��'��?�+W^^-V�уI��zG*2"1D�� �`�ckۧ%�>����B��$�R��iQ�'��)��|"�	(KHA�gMկ��R�\��Px��iDH�ş�`����#��Db�'.�QS�$+4D��I�<;���D�h�`�n�;�����`��U�!�֛�J]��eE7E�l���	)4�!�d�v�Z蹠k�Ck�)�����O!�䈫T0��c�j�? E�4��	^�c�!�$*n��\����5�uQBbJ03!��P┨��$vd� ��o�!���d $���A��IpoC�y!�DD+���A���3"� u�3l�".�!�DO�*��؀B�:�|�q!V"l�!��,<xСY����oI4�!��F'��!��F�f��#�n95�!��ztX)���>7v��`K�U!��w�N!�b(U3/����Ȕ�[�!��*Gb��Uo]�L"&��L��!�D�7+�2<�6*_N���I�!�6�(9���Q�lL�3goݥ?�!��N�dx��XU0�y��9Q�!�� ��8�O�7\�xM[�b!��<�"�)�XF�C�!�D��/�z��	Y6=���P�F01�!�dI�U�}�C>Y�(gۚ0�!�$ťH~�%T�qZ҅G��!�D(=Ŗ��̏Wg|I���Ǒ?
!�DǏq�Z\q��&nH��K�.�!!�DR,Z~���4g�R�XSn!��;%��0&���@��8�4�'4!�d����I�jE:�\�f�D�T!�;`����s�W=EF8�!��`j!��#���U�M-�T��a�@�!���nJ��`u|�BN�"�!�Ĉ�^�
u�E҆9b�-�b!���D�x�T�N��e�D��/=p!���g�]Ʉo
4_�Α#���G�!�d��Q7 �����)L9Q�!��,
�,T�����mڔ*%��3�!�K9
�X�V�e�T��,�	�!�$�\���S�/Q���Y{!�d(��a#�]K2���K�<�!�d�6]��z��8���s�]<�!�D�[Mj�ifFR9l�<���@�Wu!�$�/$�p��v��=nT���b�M� E��^��H���8e��2S	
4+�n�3U�$�O&�'�`��T���y?�3���e^Tb�'C���6�ďy����6��?bȦ@p�'Ҥ\+�cZ6���� B�6X^`��'#>��0��H�`���~�TR�'NB �� �-������v��i�'Z�Y��C:e�sQKª����'vL�b�MňE
���H�������IR��EJT�V� d���.H��B�	#"��+�`սt�^�"7�У=y�'$�P�ՠT?9�P��@�Zd�N���O&������H�^���J�>���ȓv�lt�s�J37�.`� �Յ~ �EyB�|�d�?� �v��<nF�(6��b}B�'����j��9y�	��߲|�'�<H��g%Qx�dڂJX�]�x�'�bQ�l�� d���ۆ����D(��Y�ӎ��E�Bi��!4Ph h�"O�#�-[�h��U���C��Q�"O� n�0 ��c�6 9�n���T���"O�"�&�!bB�%
Z?��*��Gy}�'I^hP��V)
+�Dc$�Z$0�~|3	��hOf|��.Z#_Dv$!w�δ#�����"O`�q��!�(Պ��U�n���O��D�@�Y:�L�G@©�F���|!�$��#򬺀jHf&ν E���!�ҠY���K\�-�a���r���"O��ٖ��cVf@S������"OvA�&!_ ������"�b��Iz���I�#y����	;f����'W&�!��K�l(S�M�=��"�$%�0�Fy2���0��(�p�w�Μ�$=$�\#�#5 yY���!��1V���j١�ҡrP���7O*
�y��>�Q��'y<=�|��c�=� �J� �$�z��Z�<�2DM)q(l�����TUx 1�c�U�<�W�FfTY���%��$�rDS�<��M״Q�&8  )�91��Ny2�'��R�K�_���b��IG�`	�'#ك�+1EJ=a�(,����'�쉫3iy&����-�����'L-�W'�&��$�ێ�l���'o|�1t/C3Y������C+{�58
�'
�8u�$Q�l��R��n���x�'r�$�Dl��a��8@3M�+l�b�a�'�p�ì��.: r��c ��r�'���$��>�Ωp�EH�ո�'Qvj�e�5iz��;�U �:`�'�b���d۠)�9�CLƔ�����'�Bሰ�W4[����E2s,�Q�'ɂQ����==�0KC�q����'~ ���K>\@�5C��:��-��'d��Á<����v��.6�r���'�h���e��?���V�ֹ^�>�	�'Ѽd9��
9�d1FA܇ I�\S�'�y���(PY��;�(ղe'J���'D�R�Y�y��i�PY�88P�'v:�HFD��bJ%�B��4Nm�d	�'�܈Q�"{�y���z�& ��'*��{�d��J�YCT=jr,��'�Ze8��B&/=����c)�LZ�'±3E�0*���C�[�`-�y�'ِlx��N�<|�tJ4.^��@�'���1�!i{j��<A�H��y∟�DUy��L�3���9��0�y�\#G�eр���I�Aq"�I��yr�D>�:�HV�ن>%h�Ӕ+,�y"玪7M��u�L>&6�P�"�2�y����o_�mP��Ņ,�.�b��ǎ�yR�<�6*T�Uy�%K/�y����
����6Lt� W'݈�y�M@�[�<9�Fn�( �*6/$�y����y�r��0j���H��\<�yBʋn�	�g�5>P�iU�I'�y2j�J��ѣh֔+Wd�2r ��y�lǨXc�4s���	��Y�fb��y���2.<94 ��b��%�1���y��Z�t?�C�@�.?�|���y2�C�4 �&D��aE��K��P��y� B�:(j&ř$�ܵ�Шׁ�y�HT�i8>�	!�)� Ԉ���y�)W��� ���ݢ6������y�YB�X��]�;P���I��y
� ����b�z��`��M7���!"O�)��B4$wP,�E
g4��C�"O�H؄��#@���P�\~(�ȣV"O��0��M�2�˱MQ�Dh��d"Ot�ѐK�(#5�d ���/3��Ȱ�'���'���'�b�' ��'X��'�^H�nrR��Cb0I�\i��'�r�'m��'��'D�'��'�n�	d�V�,�� #��V�ڢ�U�'T��'���'�r�'���'���''x}��+̑B����B��&*�B�cf�'���'�2�'�B�'���'�R�'�DeB��_)Y�e�F^�7�.%[��'�2�'���'���'r�'���'����T/ÍZ��,�X�PA�w�'���'���'���'���'��'�R�릯�7WH��2D�V� E��'�2�'��'72�'(��'���'�Ʃq �H�N�*�S���BĔ����'"�'#�'L��'���'��'�*���2TZ�a��ÖR%�康�'gr�'��'|"�'���'/�'i~Es��20��Xqg�@�W!8+S�'��'�B�'b��'��'+��'q��5,�	�}(&�� �y�'���'�R�'g��'�B�'
��'� 8`�ZU�v$8q*�F�R����')��'���'��'��'�2�''"�Ң[�$%hRo �}�ZS�'�R�'���'���'v�D`Ӽ�$�O��R(R O�N�S��%d�F̲�DNy"�'��)�3?��i�N�j���.5w�d)4$̫Z�����4��d�ܦm�?��<���C1Ҩ1V�Y�j9��Q�ś�;���?�a���M��O����N?ٹqE�9ZT�I{���(yT|���%��x�'��>�x�M�0cWص2�h�ܒ�o��M�d�F{̓��O/�7=��թM ��^����Գ2f���k�O��Dw�4ק�O!4XzӲi�B�T�t���L%��"��C�R���f��Y��2K8�=�'�?�6b���!)J5f�U����<�)O��O�nZ�(۪c�t���K�e�٠d�4���3.G�{i�I۟���<Y�OF-�d�*k
|1�'	� �����$���Y~y�5o.�*Y"o��H�"jK?a���;E�$dt�)��TyR_���)��<�R
�0M��!�6� @m����f��<��i�&%�O��nw��|�1m˂ho�|H��D1���#T�<����?���↩��4��do>� �'-H�©E�:\)	E	�)C�4�d�<�'�?���?����?��	�0~8~T`'��<�,�σ���DޟPp�D�O���Oܓ��QB02qRL�� 4�P!�$6�(��'���'�ɧ�O�}��;C��!���X(|>X8EM>h�+�Ox�� J@��?qW�1��<yՍ���Vu� 	 3+&M��	�$�?y��?Y��?ͧ��AĦA`�A럸ZGcI��u���1(&��6��H�ٴ��'
^��?����?)D��C،����E�%ϹM2؅�/V�M�'�6q`��LI�O�G%$I�R9�2KY,Vty3��V��y�'���'���'�����'!b,B�#�>\�tD ������'���'p6m��WV���'2�ɜ㖤1�
2x�(q`F�� �>b��������&x�r�o��<��9-�-���	�v�a���:R&��$gу)���D������O����O��	�Xbj��T�ǡ[���`o��3T|���OHʓf<�fJ��1"�'�bX>�X%�E:c�����ܜu�m��#?i�R����՟�'��Qd��*!H
�T>�)1���:� �	E©� �Y�_:��4�`�:�{��Op q%��i�&P�M]S��[B��O����O����O�)�OʭS��<�#�i>�=$옂HZ�ͫc]�4�0�s���"A��ɽ�M�O>�����Ο�P�LP�\�����]���0�- ٟ��ɴT��mZ�<��43P@}sa#��?	�'V��Y`���.�Z�`��O-*�H���<�*O:���O"���O��$�O6�'`3��
ϐ!V�fp�c� �6��3��iq�:�Z���	s��V%��w����r#Ϫg�H`y�I��xQ\Pv�'��|��ԣ
Ow��6O�9�v듦 mD�Cwf��l�hL��0O:i���F��?���/�Ħ<���?Y��@F�ѻ��T�C%@5;����?����?����$���u�c���t�I���`�JTx�J��Ҩ#ŬD%�J��$�������ON�O�E��C^<�D�A,�0��"��4B7�ƨX�@��%>�-X�b%��I���jL\����
0�`�Ο��	ԟ�������r���?�dÛE�Y�&蟅5m�ɢ�,�,�?I�iJ:���'��f�O,�4��T��k�0d��-r?�C�:O��$�O�8W�6m~���ɉ[�~ ���O9��I��>��ͬ���§��oF&�$���'#�'���''��'�b�sUܒ5�m�F鑙j�̩�[����4�lPS���?������<�5�ϹB����n��o
Xt���	����	a�)�Sp����_�3����ꖸHL��J�N[�y5��p�8����O~xaM>�-O1&離1@0	4*˺*2��#L�O����O����O��<�i�U��'��Svj�PJ@�
w !��'4P7M*�	���$�O����O��8`NRA���kQß�5�0����$ ɔ7m'?����g8�|"�{�?  �P�悟
�nY�,�x���t8O,���OZ�$�O���OV�?���W 	!�"]$,��Xy��^yB�'��6��[�	�O �n�u�I4C��iI@��>N�5�#��.�,d'�4�����S#F�UlP~�P"}��0��*@�<$�� .�P�y��ҟ���|�[��ß4����X1A%	�v��Y��ߒ!�����ٟ4��]yb�p��0���O����O��'b�\��g�J��,j��A ��q�'��?!���S�4"S-|�bw+����t��f"2�3��ճl��ƈ�<�'$����� �'48P[0���a!�@@��+��'Vr�'�R���O���MK��W:"T`9vHӠ6�R1p�Y�0?��;*O��o�A�3��I��8���v�ֵ3�R�*�̑�0��@���,�oZQ~���u�NM�}�������xAO�%�K�� �<	)O�D�O��D�Od�$�O(�'w����0���
�M
x#Qi���M��e���?Q��?yO~�f>��w#��b%I��~�~t8T'�B�z�b6�'2Ҝ|���Y�L���6O���N-vl���

�b�8�;O��A�"�6�?�
&���<�'�?�" 6uȔ19�;4��J��,�?���?�����$���)�u�]֟��I矠@` ��l�p��
@���(�ccTK�in�������h��-a��҆c��=����-��Z���~{��
��q����O~����O����g�H�c�h�
��e#�KŬmҦM��?���?���h����	���M���f�J�KKl֎�DU�I؆,Y�`�	��MC��w`��#E��h0ɐ��1K�t1��'�P� Ib�Ʀm�'>ų�
W�?���Э)qzIq�}�h� �.�qF�'���џ$��ܟ���������b�L5��M���!��ΉL���'!<6��LwD�D�O��-�i�O��Y����w��-���̫[d��2�]}��''��|�����93)����I�U'�`��E�&��L���i�L˓(r4i梟�'�0�'u��"dP6z����dԠ#i��B��'Jr�'������W���ܴXo�%���jZ�����k��X"f�ˊ=��̓;���~}B�'�'�����ǅ}'R�Y4�:^Ɛ�Sk��J"����pCKίm�������]S3�`p�,b��V�[��d��4O*���OH�$�O����O��?Qrd'�F�́b�Y ������ߟx@�4hG�e�,O�nE�I�s���T�á3�x��&�T�*��]&�,�I��S�h&h�n�g~Zw����C�X�z���Ks�C)���i<SR�o��Ky��'I2�'2�ŊS��u�����;���#�A��'��	%�Mc!녩�?����?�.��+w�
�(�h�;���:mo^Ñ����O^��0�)�h ����A�U;	"p����
�jp	ԯ�1DT9�*O��?�?y�d"����<�;��)?�	�I�>�
�$�O����O���i�<Ľi��iQ`�3�D�0���M6��2�M�� �'W�7�'��3����O�`���H:݄ UVp�,Y�pA�O����/4
7m%?)�NO7+	J��wy�F� XS@H�1�� db�]�$��y"U����ٟ��	ߟ��IӟH�OW�t��)WlZ�ˏ5&x�ȢAi�\|#���O~���O�����ܦ�ݷ]=��Ph�.D��Q!FCƷYj����ҟ�&�b>qʅ L���͓}�"MA�
FN�`[��R"Z���U���I���O>�(J>A,O�I�O�`�oä�4���V)Y*�O��d�O���<a��i{��x6�'���'����F���H��,y�ڐ�e�$�_}��'���|��ң	��3ǫ! }��r'������Wj@����H/1�����~��	��QQ��e:D�`'DO��d�O���O��$.�'�?I��(NW
)��D��=���?�ֶi����@P�D��4���y���_�dzF#׉{n��#̝�y��'T��'d(��p�i�I��|� #�Ox|R�eS��=���Ȓgt᪁a��Sy�O���'qR�'��dM�d�n4@eL̾�Rl3�D|x�	 �Mc%�ȡ�?���?a��Ԉ߂;��T��B��#��#ckK$C�듵?���S�';��}X�+�%2`�B�#��6X�P�%�>��'l���kD�� ��'���ny�h�J�S��dj1���E�<���'�"�'�O��	��M�v*��?iB�j@����'��L�ҙ0�i�<2�i��O��'�b�'E�L���)#LB>@�,5!��[�'�P�҂�i���n5�
��O�q��nY*x��px1 �5��Z�ሱ6�D,�O&����VX	i��H��<!��@&�v���)Ŧ&��P�m�{�HUd'�_��;P�O�����i>����ۦ)�uw��r��b�8g#x�6�Y�n�^�2pf����s��|"V���?�G��)r���1/+0�S��R�'2^6-X�tF�ʓ�?�+��]#6&F>V��lZ�G�����[���C�O�D�Of�O�S^�P��Ǌ<_ږ=H�E�2�UV$��Qy�O$P��64�'C��s�P�A���s�
	��z��'B�'I����Oh�I�M�p��b�"���!Pz���	x$:.O��oZZ�|���ܟ��G`�%}g֑#�A[�Yi�س���H�I�O��lj~Iߍu��x��X�� D���N�T,�2��@�>�X�I�1O�ʓ�?Q���?����?1����̬#�b@ �&�'m%R�8Q��33@$nZ�@���	˟8�	X�S˟t�����-�::� 3�W:R�ZY�d"���?����Sܧw�2�nZ�<!$n�H~u��+�#����`��<�$R�/���IF�Vyʟ�b�@�@}�V�R Tq8|�p�'v�7��w�&��?-8����`�Hْ�j��~��4�R�>���?yJ>��aR�<z��I򌈢%V� ���Z~��E��-2ÉUd7�O��1��d~�Ȏj�zhi�==���C�Z���'D�'���쟸�5Ꮥox�tqSN��+���3M���L(ߴJ���?1�;���4�V#��Ͳ���TFL1�e<O��$�OZ�Đ&x�7�2?aU@��T�r�i[�4�(S�Ӧ_>��QT@Ԉ{p qBK>Y,O��OH���O����O��ȧ��6��90hIH#�� �i�<�D�i�� A�'��'���yrG̃�ъ���<;����pO�L����?�����S�'[����L��B�'l[w�X�cG	�[��]�'���@��ӟȻd�|RV���AP<#�&	ps%N�0�YҁĈџ��П������py�e�>t�pd�O���1���b�7��E&�@[6O`m�l��MK�	����	��.׹BK&���J'L{N<��dJ����nl~�ȗ�)�B��SP�'Կ[F/Q�9�np�C+*uz5��O�<���?���?Q��?���$Dǿ?��]9�mX��T�h���*@B�'���O��"T���4��s�f, C_:�AZV���U@D<�d�O:�4��l�p`m�f�r��,Hp̍ U@!��P!m�D�p�N�%���D��䓎�4�����OR�$�ei��iv���l\7}.���H�O����<)2�iF 9C��'���'�ӛX�����
�j�فJ2/����	ʟ<�?�O�����N�vR�Q�F��5���X-F�`)�"]?��i>))��'T��'��ABA�n����+z*���n]՟p��㟤��şb>i�'%�7�`�R5��A+w�b�C� p�:9$��O��T����?�_�t�ɠ��uH�L�F�"%�����C�X��ǟp�`Ӧ�'0RE�t�,O�(y�L��JXd�*���*d�:5��1O�˓�?A���?���?����U91���/�>h�v���	�h�}o�1d�m���P��j�s� ����cq��L� qެ&
�U�9�?���Ş:Q�ěߴ�yR��>rK�/WZ�c5��4�yb�C!�����9V��'��i>��	e�Ty�сY52KB v@�T1DI��۟�	͟��'(6톾'�`��O���=*��9zP.�c|��zf(�!� ⟄��O��$!�	�j�p�hÌU���ق�Q7������Q`"
 M$
�!L~*@��O �i�w�x4Kp�hGDC�w��!���?����?���h�>�D��=��Px�i����+S�Ǵ94~��˦�y��������M[��w�Y�EL�r�8�Z�=i`�Q�'��'I�N%n��F���ݏ=}d���[�V	A�I�"�t=:U�#;�r�0ӛ|Q���I����ɟ���⟬Z�'W�
:�LI�,�$:)��G`yRab�����O�$�O����d�+J��"O�U"x8��A��\�'8��' ɧ�Oh�����6\���rm��΁[A��Yyx�q�O2������?��+�d�<I��܄O����I������hٳ�?����?!���?�'��D�঍���YßDAE�Ӡ^kvS^�j�+�K՟I���Ă�)�?q�[����ڟH�ɋ7�Z4ⱭE�L���pAa�r�2A3�#��9�'=��ʴ�M�?Ekњ���w�$�F�F�E�H	#���G�4=�'5��';��'��'���mR,��#F���LR�M,P��s*�O���O�]o�g6L�S՟�Y�4��h)�5��/[:{���*r�EHR ��N>)��?ͧY ���4��$Z
HM�5I�ř)O@~ب��� �Q�o��~b�|b^���	ПD�����	��4R<x;d��2� �(Qԟ���{y�h�
]�PB�O����O��'k���Җbҽd���D����� 0?��Z�4��՟`'��'d(��oz�=�O�+�� ��%�8���;��4����B�ƓO�YR�m^<jI$\�pK�s����T��O���O~�d�O1�T˓M��fN�9�����˥
Q�4
�b֖	JP^�p��4��'��?y�Үu����#U�h�$2Sh���?��Z˞m��4��D\��b�P����x��	�h�0, �"����yRY��������韈��ǟĖO�HP	���.���0 �԰#!.��`�cӚ���a�O�D�OJ��
�$��睽*���� E�H(7�����Im�ŞT�@ʦ�Γv4%𵤟�2���C	^���ϓ_K��c�h�O2��O>y+O����O@2��'1Ĭ�G��gv k1��OT���Ov�d�<ac�iY����'.��'� iP�H�mx<r7��/:�d)W�D�V}�'��OR�Ҁ��,��� V�P89�҅A���!�����e*L;i��O����	:i�BH�:��� e�h־<Cue�����'t��'q�������@��J�|�r�����
�؟(zݴ_�n�����?�G�i��O�N��O"Ĩ��W'�Lm*�-�"��$�O����Oʁ�Ja�J�R�Jm��?� |�@,F$Ӱ��T'2�YT�.�d�<����?Y���?���?1��L"�0�-��O((���.E,��P���!�����I�4'?��	�
��x����N:6O��Y(�0ҩO�d�O̒O1�f�#ծ�
DfL�jgӯFu܀ʇ
N�] جT����U����i��_y�ň+8�B�Q�@�8��&�vn2�'2��'Y�O�割�MˣOE��?1d �*�akuׁ:	
�����?	F�i��O���'5��'�fD�6r@�Q��T����ݎ{���:�i)��2w{��ڟ쓟����59��;�BX~����Í�1��O����O���O���=���- POU�8��9�.�e�t����I��M�6f@��c�v�OzT��J�7k���7ķh6p��'�d�O��4�꽐S�u� �Uf�#V��<E�CF��H�����iT�	m�	tyR�'���'�r�ϰbk��C�ץR�v��g�D�uQb�'|�	(�M��1�?���?9/�Dq�!�2Z�<	��^�Tߎ��g��T�O��D$�)���3,�~Y	���By�[�5~-�1�3�˅]j�j.O�	O��?���0�$=Q넨�!hJ�U�N��C w�p��O����Ot��<y�i�,l9� �Yy��AA8h��v��1#
�	��M���>9�/�Fku�]�:=�)��
V�����?�6�Ɨ�MS�OH�˖O���M?���g
�%2�l�eL�)}�rx��nt���'��'���'���'�S�9ټ�%���رxT�Ėd�Hڴ5�D�R��?������<���y�!�q����E�pv��@�ԪD�2�'Zɧ�O�	��i*�dM ���)���lע�E���$��D��
ZR�]8���B�G?s�ܫA�a3j��A��&�P���e�6?�0p�b� =����s����N��Q�,zLYK�,���y�R�M���O,-/wP�%���B�G���� B���$�
��{�k�
8Km*��R�� ��Ҿy�� �%ԭt5F�ѥ+;u�0����'4NK J�S����k�\"�@�dK�:܌y�&-%I���ie��\��
�L��
M�S��v`fΌ� ���+��1�Rq0Q�JV�,�������� �Z,mhL���M��?Um�	ClXH�[刌�dϐ*>�&�'h�'U2�'j�l(T����l����J��'��ѱ�l�!#���'��T��"�C���I�On�d���I�TƱ;%RT8��B�Fޙ1�U\�Iş����+>6��?i�Om<�#4��m�ܝAI�$�x�ߴ���ۺ[cn-m˟��I�\�����Ƥe�WLY�W؍�e�St��R�i���'���p��7��~�4܊��O��C�/��7�E�H��mZ��@�������0����<!��/FT��
e�Ȉb� �$���I囆c�F��O�?���,*er��`��!d��Ճ��\ۆ i�4�?���?���D��Iwy2�'���Ƽ{���i�J��m��Z��O�=[��6��Oj���O�E��.�ff���/6a"����A��.-��1�O���?yO>��e��kӊ�C�$�� � ̤}�'+��Jw�|��'�'剴HIԥa�.T68^>�`-F>VΊ���f]����<y����?q�y\�U˅a��%��i���(���#���?���?(O9��|�螮�R��W`�B����� զɗ'�b�|��'�B�Im��C-Mx4�e��%d�¤��P
4H�����	՟��'3��b�~j��-Mp��̝	<���h�Q�t{,��i~��|B�'�ʃ��'�x!��\~At��!��m�Njڴ�?�����u	l�O2�'7�䇐|�^٠F`)��C%I�e}0OP�d�O~�%��On�O����g>��!�!DDK��Y�/R"6�<AL�2͛f�';�'���ʹ>��ּ�Z�׿R��aV�I�.~J(l�����	p_� �?Y��D�0��QZ���U��M;6@��(�v�'���'��4n�>1.O��Q�@�2�D���ƚ5Q������y���i����O����9�� ���<9K�ݪ�EË�7-�O�D�O��I�bJb}�X�H�	\?2�[!Ҹ�g�L_���C��E� u�}�I>����?9�sp�i��P
Je�7�)>jv(a"�i���:L�O��O>ʓ�?�%��'����Ϫ{��1t$6A��'��Z�8��ޟ���jyr��JF��""]24�e�E-�FoI�D4���O\���OF��?y�O�R��5&��OG�YY�hH>#4\#�4�?i,O��da��'W�������N_5&��)ޜo�<j�.��y�F�'�����O>�n��o�B,�W�Dfp�<�Pe&!r�OP�$�<���b|(4�+����
-�]J3�I��p��mXؾ6M9�I��,�'sT�BK<qg윔R��hd�P�zڹ2S�NҦ��	Yy��'�&�:f^>y�I����s���GDg�0��g�25oA�NC�'|�U��6(&�Ӻ�s�Ҹp#ҹ���Ө[�dAʴ͗O}��'>�;v�'���'���O��i��V��I>C�D�<>��SVmg�H��<�
GM��ħQ%�)��2< ݂妉�6��ulZ'��	�\�	����hyʟ�)�q���VЕѤ�ȧ[8�1�E�E}rAS��O1���$ʻ[<���$�/jl�����DD��1lɟ��I�0za,����|j��?)�� !2�%�
F�HS��[�aI<I���'�Y��r���˧�?�燎 �� A�K+y�
�sd·(	�|pb�i7"��t��	��i*�I	"3�@C�*a~\IH�D��1|)O<igVW̓�?9-O����>�,�i����C�~E{�M��h��"�<)���?ى��':��צ\PU���5�-�@lF�]��fn����O����O<ʓx����28�µ2A&�2C�ޑۧO]+T���Q�������}yB�'����4 K4�V̸Q���r������?�����D[�=tt�'>M�]�'ez���c&[����Y��MC��?�,Op�$�|�����B8�k��Zp�l��)ޗ8��6��OB��<	��]!hf���l�I�?�(��E�"f�i�Ś[5`��S^�����O��d�O���4OԒO��ӳ �I �gכ$"��ˍ��7-�<aȞ3m���')��'{��ɭ>�;rz�pn
ml�1 @j͘Jc4%oϟ(�I�<���If�~�')Ŧ1��*��ے��r��n��C#�@;ܴ�?���?Q�'��	Vy���
o$ � =R��=C�˃�*�7-6C�d�Ov���O�2E p.)�J�Aו@�dqd�o�����O ��Q�i����'�����4��)��A)��!��J&����>�mZUy�'�,5������O �d�O��qQFi���0fy\i��E��M��Q����OJ��?+OH�������˘p<X{v�,d&LJ]���{�Ԕ'���'�BS���q�ؿ���c�&�4"Α�b� �O ˓�?�(O"�D�O|���Q� ��]�b��(܈sG� ���<����?������J�=^̧?�B�Ԧ�-YE&i�`���\nZjy"�'��	�P�����x# v��:���;gHH���z�������Ms��?I��?i+OD����G�d��5V��:.Qb�r���0�������M[���$�O$�D�O2�0�=Oj�'�i d�*k:���2���F��u�ڴ�?����÷IDZ9�O�2�'D�T�����
Q �R��$"�DΩjp���?9���?).��<H>��O���kg�_, xQ�@��(n�ɐ�4���K�LӨHm�ٟ��	����������G� ~��)�*Z�;<♁�i���'��yb�'��a�'Y�~�y��K�Ii`Aj��� ۰n��r�۴�?����?1��<a��]yr�-$��ӗcQ�d�����o�6-�, ���O���ON�?Y�I)q�#���#4�|j3mZ� ��Hݴ�?���?��V�o��	Ty��'����l��Q#A�Y!sN�q!�L
-����'&剧H��)����?a�O���剙]�B�..рl8�LN����1��^y��'P��ޟ֘k��,Q�T�`~4Sd�D�&�p�Jq���?����?i��?,O��a�S%-J��P�
\k�)X2�P)Vg�X�'����Е'�2�'��E�+����A<��h�
@<S�R�(�'���'��'��X�HZD�������6�>q�B`ܴM��
�̓�M3-Od�D�<9���?��TE���Or���۵.=�j�-Şq�N���4�?���?a����U9;���'>�'+�#5(��QbKo��lG�L�Ms���D�O����O��F��O��'c4yz��M�@��W�ڙyVu��4�?���;��0%>��	�?9z�MH��"l�<��a����ē�?��Gh� ��䓟�mU,*��1���K��Yq����M�-OƸ@�Hʦ�*����d��'(ڔ���김�i�17R|�۴�?���`͓�䓗�O����iۿb�T����(>���۴��ika�i�"�'9R�OՊOx��L	�%J3�х~ƞ�	�eZ�C{fl�@H`�	r��v�'�?a�HX*L�3wY��\8a�����F�'�"�'T��z�>�I͟���>��U+�/(��X3Ș� ���=�$�k�������Od�]��������i�ɂ�(_
T,Ho���[�� ���'��|Zc��|�4��:J���$�,Un��O�ks��Of��?y��?�-O΀`� �3:���0�E�;u��̠�Ь3P5�>	�����?��	��,�ɗl^|q�U�s2�Ӗ ��?�.O��d�O��Ļ<��9
�)\4��]�aE�V�z�#$ǅ�t���Ο4�Ie�Ο0��0���ɛg��		���y[�Y����	^�.5��O��D�O����<1rK6?��OF�թ4뉾A�Z��2%�z���s��rӤ��9���O����=hO�$3}��׺0��))d�&�(��d�ˁ�M����?�*Ob��k�X�Sٟ��Ӿ0���8p�ƈS^��ʁ'-Eq֙�L<9���?風�F�'��Ɋ\c|�R��d͞��'F3 ���[��Cd
���MC�X?9���?y�O@�iC��=�4���Sbvȳ�il��'�R���'z�'q�Taf%Un���㳇�1HT(�b�i�& #r'p�p�$�O��D��	&�4��2+Ya��$��,��0�S��x�ڴ��d������O�b��'4��%ϝ�&�҄h G>7M�O��D�O�8���g�����{?����S�h���/����AÏ��%�re�x��'�?���?��W-IT�$��� 65��i�+q��6�'��H�o"�	���'���| ��)Ti�;kJ!�O��_ˈ�A�����O����O��T^�|s��+{i�h`�7Js����7k�'���'��'���'o����V������P�Ĕ�yrY���	��x��ey��V�%�F�3� ��"�!1ͨ\cS���cbZ�B�W���IK�',����@DC2�FГ�'�Y�!�T���$�O6���O��>n� �V�����@s>�g�;8+NaUe^2.7M&ړ��$�O��'-�$1�ńM���d�pmn�I�Í����<����O��&�ҕ$��H��M$�3�"O�y��
��!��(N�1㥘&cv�� ��T�.�j@�9J�Ҧ�ٍ
�"A)�jǡ\5L�pb��,w^i�p�SS#HTH��I�s�N\Z����2s����K�n=tZTjɠ����^gK�4��B�_���P♁&[&Ɋ�5i\ zbk��X6�1����@�:u'���`�$QF���a�O���O2�����wd>#�9�䠛�V1R��<K!� � d�i����I�jHˏ�t�(}���:`܌�H�(ۈmz(����H��,C��p�|�x5aա�65���D,�A�r��Y���i�f1���l��y�g��O����E�i>�E{Zȉ*Fe��R}<%��C_�P2�'h���*A�5Z�0K�E���*� �OJ�Fzʟ.�??mɰ��( 8��%gFz<8,G�],����?9���?����p�d�ON�ӵn[J,f��)(�J�2�
�H]XD�ʯq�p@��	�E�NP�'�F�l!���Z��	2��%9<��	�%9��2e��r���k��Le���f/�O����O��D�<i���'ۀT�0G��R��X�F'�b�Vb�'�(u���J�$��Ma�ͩYu()�y�o�>�+OL%"���D}b�'qČ�TA̎^�Z=�0E�"Z` <� �'2�ϭB�'@�I�d�"d���٪|ܸ�Pm8��ԯ_:��X� Å�i[h��I+Ia:d�`���dը�'�z�Xu� `�� 7eF�H浑Ǔu�]�I؟Ĕ'jP ���R��� �m].,��y��'F\EH�j�y�y��M�6jƊD��'��6͙u$��R!b�$'�d�*UN��E��Ĭ<A���!l����'g�Z>IK���x��aW�"o�Y��\�v5�]��b��D�I�8)*��N�	U�dU��+�� ��]a�䕦x̮���5}�0z�R��u�׷A�*ᆓ%�Ll�k��k�Ũ%hB 	wn� ���X�'�����?�c�i5��I�1~������0`�@B-��Gr�D�<�����d(�L�]�v�҄&T�U��/����ۦ�Jش�?!��i�r�O�Dc�)�c�$�ҵłX�6�O����O����'O?S�����O��$�O��n�R����7� `i	��;CZX*��҄�����*Q�i#�|�蕖'�8ݙ7+�}�$���LR�7���O�E}R�U��<�}&�<2��-L������/UH�t�Cb�,QH��)�3�Ɵ`jX�se ;�V�8 C�O
!���r5�t�-;���6���;��ɼ�HO>�A�&ˑOr=As��*f:���цhUP��PH�ӟ��I��,���uW�'��9�,� �#�g�.%���!�X��7J�I]!��Q�`�K#��+�j�+��x�X���xrk_R�H,�V䐦?���%�ĳ"J�T ���?9ʵl�py���:<B����G�<A�o��2y��p���#�Lx�HZC�sܱO� Ǝ\����ϟxT�	`榝c��[ `]Dm��Rџ���16��)�I���̧C�~�b#�S}����OfԨ���+s�؅�bcMl�
�ʁ�'�C��#�#������c:��ц�Y��9O����'�'������Kb�mqMK��$ �'�(� �b7�6�AB�|�p1�'.�6M9^r�a"�ȣ=����n�6L1O��N�˦��Iߟp�O+\mb�'wH�!�+�:6'�0��H��fK� J��'�r�¸}���T>����&�;D�I����JI�Y�Ot�w�)���Il��u�/3-�C��9\F�'aR8�������Ovh�Ie�S�.�rSG�88~�H�'�J4b�CƧGo2=Ks��?��HYÓ`͑���7�a������I�`��Cwh_(�M���?Y��D{CǏZ��?����?��Ӽ�A��F�%�ceޏ(M���"J[���'hQQq�'���4&(`%���D,�).h,=ʌ{���ay�~�Pi�EҴ?��qd��=���'Y��G���,O����
S�Dj7ßfx��k�V�Y��C�ɂ��	�$8ҪA
�&U�n��7����O��#nV���Ƙqg.HPc�QY�B�	�x	��`oXy$��F\I��B�	�h?X����1,�����VV�B�I�\c�(d��>Rv�ґ�Q�#��B�8lk��#�ېh5��8�D";�B�)� �๓j�b%ʈ�`�>8P��"O<����*�B��Wdh �"OH�Ä����QQ"�'|�!�"Ovy����b!�ܻU�_^h剕"Oj	ӥځ�h���m@1ZNn	�!"Oll�����3�~i�`�ذ&���"Of���
G	C'V�qD, 5���:�"O�p��D�P�JŃ�dN&�SG"O���НG��ص"F�c�-��"Oz%u-)c؈��S��M��q"Oz�`�V��Dd[Ǯ�F�&���"Or�B�;�pC�����q"O�H{猓'��-�l?���b"O`P��
<L˦-c�Č�B�ظ��"O�9��eҖ4�Ζ:���d#��y�J�'�r-Z�*]�^�y�ǚ2�yR�D1.�: �aƑ��dt���y2�ƂN|MUL��;"�@�N��yI*f�P�J&p�QbSEQ�y�W �n��ī�>4C�Ԅ�y�
�;<_���j�@:9k���'�yd
}w�	ʤ��KJ&�rªI,�yr��e%�Ł�@eH�aEՖ�yb�	S��aAsσ3�]�
��y�IC,Q<!I��Ϋ��y a����ybF�#~Z0횰�Q	EbΨ��դ�y� ��bx����?�x陑Cȍ�y"�^<{���d�K:U�� ϱ�y�d�5��P#7
�c �ز�y��Ԣ�Ωa�^%"ЃR#���y¤�j \��P�I�uQ��y2IU'Q��p��D֮v����iM1�yb�0$�HM�V��;j�0��%��yBkCO���0�]�|���G��y"*�8$���#�"TF�A ���y���;�dڷ��6 �� P͎��y���4g�^]Ckx<�pS�B'�?qB��$0�d5� uЖ���`X�]qE��.Hy�.��L��9�f�c ױY��xJCJV��H�7a�.�M;2#G0�H�H�h
	��d'�$⮰���XF���j��#��]��I�9(�Y8v��%db�����5=�5RkX'��h�"lH�[��@R��Me0�t@�iY�l��a�2�Li�������>���SB��d���q�X�0�)�Wy��BO�!�#M�A0�pW,��%A�\���.���m�b㰘ۂ��/���"��	^��+2��m�L��N<%>q�3�Hp�7E<Z���������"O.���D>pg�X�Ξ�]��-z��|�Ǝ���,x�ᒟ=�@�sN����'N&9z�kT�D�,�����S���ϓt,�����6%���l��Wrn�3�D�<
�q�&�&z\ɲ'�Cϴ�q��	�:�Ri��I�$��1f�O� ���G�A��O ���O�c�UHv�M�&�!#�;*��YVG�:���c�x�E{҆K-g���Q "��t0$�,,�;�b��G���bUHX'Қ��޴!�Z�'��OJԹ�w'Ψ
f*̥Y+bP; �Hȵ���d��|�5"�w��������h�%群��o�|o��2�c�8��ɲcx���a��̺k0㐲3���ۋ{Zuk*{�퀮>�~I���<�&ʓ�ꈻ�!��r�qO��ДIT<�
LBFf]�=^��u�=P���@mΙH�P9����p�a�Y�HT�#>y��(��3
y��$�!Q��� �ǜ/T� b���ό+ ��]"Z���f�<��]mҤ����:Lݸu����F�4#>�0�L�p�y�I��q��Ѳ����FP�0�ݜ���K�`�y�dIC�̗��O���݆ng�9�˲�j�R˖�#�C�	'G�M�.�+t9�7k�\�qp(OT����όY�2q�[w;L�&�~��c������4�z4��+�"_�4\��I�f�xZ�Î�kGTsQ�7�pơB�d��-Z&l�$�p���!�*�J��'��h�TkR���l���Y�\Y�r�}+G6#\��aB�	��`�I�6���O\� )���-aź-q!j_T��|���� 8U�E��;�pU�P���P��C����i� �{5"Uy���+t����k�p��Hc�]4a��\P)4D�P&��4I�Ս�5��A�� ���IW`��W����)'tb�@@�g�]��sG��SEvػ�"�O�\����j��Ii�!�\�$�8�T�b&��\`�T��r���r���x�B���<�`0���|џ��w��+}�� ���N��,B���v�Fq�dW�0�������V����65�\P��s�x!�D�( �)�<!�T�h��(bW+�%�Т|�s��� �w`P�"�X��Ee�i�<yU��^���j󁜍��TE���*��q�
�v���I�j�4#|�'�4Qy�B�3T��0:��֪|�����'��tA"��7"\xh�-{�b��[7dr�Ir'ʕ�v_�@��	
HZ����_�v]5���U=����V�n	�{�^AP�B�B�\
��9��Al���!��H�!�dB�o$0�T
�&\|�X�F�� �1O|�Z�N��@&��B*��(�YA���P��P �m�,]F��"O��p���EF���DU��rQm/3���S`,L��~B.�����I'~v̭aP͜�M�J�+�0F�bB�	,�|�c6M�m,��끏�o�B����"[D��ª��^x�zB`�3-C�
�ʷx�����^-�0=q�K8k�(�b�Bc�hadJ�=P�r�[�	�7{f�0 �g�<A�L�<�x��I[�$��.�`̓	ۮ�g&�$n�yɰ�#ʧHH���G�h�E��<c�$��ȓK~��"u�	�`�BU�%�;m
H�`�����	�&��hQtH+�g~�/L��*A��wl�|�gGE7�y��>nMT�I$�%,� XQVß!vH����Lż�,Q�6�u����#��x�vM���9�|! �#7LO�L��<:>�ٕ�X鸅"��vޒ�c�N�J�b�s�"O��k&��#Q�5�0�"B�j�����h�Y�&��8���M�&�L���És0����o�~�!��X2��}Ip�˦\)l�yq�T0q��$�U�ε@��m��'&���O���pU>�\6�Y�����9 �
��0l��	�P�F�'}HH4
�|jzp�	9���[׏�4��<�zr�ʞi���x�P00���,�=c �\X3a;�	�O�M���@?��$�#��]Z7i���u7χ���D 0MN�ـ�Ȧ�Py���VZ������U�1�"g׻hP (�i����$���e���i�ۼsugI'�0P'։0�I�0��|�<	�)W�$kb�C����2F�)&�߁ ��0"�PK
�(-O�.O�@��<��#Z�'*�i�ύ)%9��y��z؞�2�(��\/8}B��'�|@@��ԅD��	��� ����'�L\J@E�@8��2��R;�`ؘAn�t���
�$:�I~�$����*��	�4���ܟ�%8�HM��D� M>L4�� �"O8�$���C�g+�Q��!�j�������<�E�R/N�8�?U�wFv�zR�@p���ШP�^�J�[
�'���Sn�98n
wē�Uچ�xv%�*�6����iݩ�Ub�q�'~d@�p��D��;�C����
�����G��=|�D �(�v-��Ň� i$ܛ��Y�X�dǒ(�|y�P�&�%D�>�4�����UV�g�`��I�ek��!Ɣaq���/eӦ6mъK+��ݘ4 Z�7��y��9���#3��B�	D��}� L��Lt��ߤ]	�yB��߮S7�3�M���B��!����$!��ʧ�
x��{^�p���/f`u��c�8y�@Q��'�|� /�sy�˽3o�����C �x�	WA��y�"���<0d�W�0uz�۝s�R�FyB�%�M���:��͂�-yy�>�OKL����ѫ�V����,�����c.�S:D\����RM�t,<}f�2	��u�g�~��� a��9��ە�J7���1�n�'���i[hy�7�>�*���}pl͛��Q�7"����"O�A�O�3C�lMї/�b!F,�^py2MO�8누�'}�91@æ|��[�C�G\�^��e����)�x�#!��G<a{i/8� ��'-���"A���2I�0�����Z��
V̵	j���SDM��Dg!ʓ{ߪ̘3F	���"ұs	��>�p�L"���?�ɗj�>�� A$�����
6K@�%lm�(�V��	d4$|��$E��Չ��6Z[�ACBK҇|�HP� I�x�.`��}R_�ͻ/�P\�� +@߮�b��R�M�I�ȓ��HC����$�� w�ʤ$�T�5��D�(xEJ*0W�MHvB���&� r���.<�HAA��Y�oq8��W�'(�<i�%�{|��20�	�\��B�ϐn��L����Vn��ú��7-B.GlZ�C�U W*��Ey�ȝ<�rl������:=�S��7��'��*�7rȵE�#?�~	�H<�[^`�0���m��,�$���j�����.�.�q�N���E�����E~��&�=Gm��� N$iY�=�{?Y�8��E�ac\;�� D'���H�e"O@�cb/� �<��eCQ��0��Q�X�L�_w��$�ȇ�Z<l)(њ>ID�8$!�S���n� Q�S/A؞p��E J���"���X"&�&�)�T(9�%]F� 3'jR B��0�C��s��$c�C0,O왱�Q# [D��9	���u�D^"b�~\�c�V��m���`��h����oQ�?lDQ��������'6���`�pF	�u��}A�`�ri�)K�vPci� 8��9}J~=���KA�gz�K�jF�_ۀ���"O4�b#͹N&�0�'��N�h���NSQ�D�;D�Ђ��m�A���LS���=�!�#:~��WK��HĹx��`���+�L���^ �%㙳i����Bܴ ��Ũ�#Ә�rgۑz��L	f�@�J��G8���`B朽'��S�3��< g��0����Ō�;�*E)��<��ߊKf��W�>��l��B
�yBG��v�X ����~t�Љ�w�MiӁ",���C�}�S�@tn�.�%��7옽w�nzCYI�!�Ĕ��|(Ռ�4O�q���A�dB�&�p���Q�Q�B��U�ڧMhM�c!�Ƀ��xB�F�{�|�K�>k���򄆭w���� J<V�y4���I �eƦ�	 :I��C�1�r؛ �K!�J�r���]�a{R��{D���%0 ip̊�#���� ����W }m�|f��px��?�ҵE ��a��,\!md@qTF;D�TY�@P�řAb��im�xU|T]�@R�չ���ke	�8�|c?O,)��-z��l���H1\�Oʴ�aO�L�(UY�`C�cV4\J&��XvD����B��6�8bM�E��H�r�a�-z� (�<{��+<O�,x�1h+=y���hW�}k��E�DY��݆ `���� +D���AE������� �XQ2l'D���׃�Mk�d�ӧ�
OEQB*O�e��j�͑!w���X�"O4�Y�L��
d���چ� ��w"O�@�ҭ�=�{�KC�G��,h�"O���L�4��V ��y"O �+��^�y�
H�R��6���#4"O,�1Ѵ�.0�DS-�m�ܐA"O�(� �0���q`޵�ƅ�g"O�Q{�kր'����d�θ%��!�"O�ɪ#زP$­�c��
���R�"O���L%�F���˄�2�l4�"O�p�0�З����k��� �*�"O�Ha7��t��2�
J���3"O��"�͔C<\���_ c�|�ز"Ob\x�. �_�`����1�h��"O�hcѮ^L��G��*-�����"O�̀��ɨ Kr4R�ɉ�^����"O��g�0��}��I8`���"O8qRsg�-n�5A`��F�2d0�"O M!r'�\Ɛ9����0t�UZ"O�)�Pc�	dQɧ��oqRE)P"Ojp8e�S��ęP3-z�Jq�$D�`9�i�<=��	QAS�7 ���e�?D� �5�F:nOV������!%��>D�0;�Kĺ ��,3&BL6dμ:1�<D�`3���x��]t�0�4�=D���Otnr�a%��l��bK/D���j1���5h˰~_0IS+#D��1�TV����A����釉 D�XC"J��!�r(�Fo� 	������?D�$�%���?z�3�n�9I����7D��iD!�,�����:}cz)�A)8D��Ԏ�2��+��i	P��4a9D�� �h&���_\�* ���a��R"O�XR�%k���b�e�2X�v"O���v�)��� �ɐr���%"O��
�+�#~�xq!.VvX��Q"O�`�c)l�n�[�̖�FZF|�"O��$��(^'Y�6���B;�m�"O�Pʴ*��x�����6=��"OT ��jп]�����!�S��g�<饪����!��F�	�f�R�]d�<1�/�� [�Y�g�@�5�p�Rs�X�<�3��M� yHD>�Z�r��S�<	�a$�	@)�9]�HQDS�<	Х�9V*j��2� �B648�dPu�<A�)u��"B�и��*v��n�<��.�,���x$$�26�H$����j�<�P�R�,X�@�I�|GHx6o�g�<)�K�__���,j:�ų�aa�<�f��P�I¦	B��y�0� h�<ACA�oوm9���Y�L�� hc�<AG��$B�h��S�0JJE;��D�<Y@�B!C5�z�'�
�����)Ik�<��+��2��. �z�$��! A�<9���Uz��b��A�a���"���z�<yt�_���*w��ev ���� D�VA�aO��#�� X/f�A$����y�nuU�)� ��7W6����	I
B�	4�q� J
�(�R�8�G���C�	\Hघ',H�A���	"�K�C�ɰlT�#d�G(Y���p�ϦX��C�I�g�F�H�N�u΀Zm��;  C�ɩk�X���^ ]$�[`�:��B�QVj�b�ڬ4���3n���C�I#�ԕ@�͕�E�=&
 )��C�I�Ih��C��-q!,,`#.޻z�C䉭,v�m�s��-\�\*!��C�IG�l9;�)�~#HY`�[8ck�C�	�|Ғ��oμeۄ�(�G�2!!�$� `cL�[3jc�aV3v�!��3I��@6���17�1G�\G�!��ح^N0s�W�wE(���W(w!�]-�¹�qNF<}+0�����Ad!�D�n����q���>�n�C�ŨmK!�d��}��L��߭�ƽQI�rF��!�O��(=KU@i��LH�~2�Q�"O6�t͓�|i\�hA+~u���"O~��f�Ol-���8̸Q0"Ov���sQ��b�N�GN9jq"O��p&�Γ<�z�LP/cd���"O�8�� Cb5�4^'���p"O��QoR�aG�x��é8�	�4"OD� Q*��YA�H�XW��pp"O��`�(�FĀ43CHV� 黣"O��`Q��2���{0�������"Ov��#.��c�ZD���&gE���"Otx�I.Ƽ!��9[#>X0�"O̩�,:,~�s��c����6O��=%>��OX|Ag��A>�r'eX�j�܄97"O")P+O�I�R �hMyg"O���!m�$5���P���'"O�͊c!>2)5�УRZx��t�'�'%��"e��0�+۔�:���B�	����w��(�d/	�0�7"O"�
��@.�.DӀ�#v[��s&"O� �P�F�@�A�6^&�Y���
}����
� 0A�v��%pR��/ۤ?����"Ob�9*[#z��҇싮�`��C"O�Ka�
t�!�+Τ����"O���FE�c1�d߳Q�RYy�"O�����X�{e��<J����b"O��,mk^���k ��"O4M��P�-�$daG!�Z�p���"O���#�����/1OF)�� ]��y�&�q���z���w������yb-�E2d*AUtr�ё#���y"'E�<��p��.l���Ɂ ���yRa�U�4�۪Qp� ����y���:c����'ΣQ���r���y� �?3��As�D* �\�8sO�5�y��2
ƈ"t���r��щ�/�y"J	9Xg p�����\򁐑&B3�y"	K=�J���ˉ�R`���L��y-��x�h8�F�VX֨�ɢg *�yB���D�1q���]Q�ȒBT��y$�pH�d�^�W��%2뇄�y��,��Kh�2\�(�0f���yB�G�RL.0F�<
`V�C�m�9���F���O��QY�h�-N`J)p*K�H5�Y)�'������?�B���YC�-��'aN��w�/P��ˁ<>f]�	�'��Tॅ	��l���,ݲ���'ᔰK%�*n�\�����)EDZ�'�ƌ3��Z�@ ����Gւ(8t�'O��U�z��HY���%
׈�!�'��`��e�P1>��Ӫ&����'^�I����;Dc�-�F�@�}�0U �'�2��0B
&X$%�va��If&�+	�'r��b�C��S��}?<����\�<#�[�����G�~VE*��Z�<A�C���@FN�"� �ۧ%�T�<i筇0#�0�Qu���{&
���M�<90�@-�X)�aˢ-	L��c�YO�<��c�!�0�W�%5�����I�<Q �8o^m�vADD����B�<�G��9�q&F�4����ti}�<Q�iR�KZ��'j��K��RPoy�<i�/�=�v`�gEen�U��.Eq�<q�[�L�� ���-:���d�Un�<9����v$�	i������Ypb�t�<�aU-@R�@k@�ڰtD8��kEp�<�e� ������o~���/	e�<�v��o�E��.Ł7˪��@]�<�u�Wz�NP�D��XV<d���t�<�o�&]p�	�`J�*"b�x�!�o�<�� �2aqnX9��էB�j�JnDT��hO1�H��W��iv�eZȈAy8}��"O�}"���4Dm��'�
#/�J-h�"O8Y�3f�(%����s�!����"O��q	̳N"���gɆVV>�p"Od��F$M�/��+��jO�KB"OU�q#W�u�r��Ӈ�{Cx`�v"O)Z ���E�V0��J|1���q"O�p���ƞ��E���s\ ��"O���"9�L�1�/|\�ica"O1�Dh�*h�`aƥYW�1�"Or��&�4�!�#��lx�"O�١�l͢Mg�tH0�Rz�^pq4"O�����0]�D�zF'*�[�"Op)1��:S^�}S���9�r�i�"O� �� �^;t�������c'.� "O�1�G�˔v��뎱h�R�"O��IA��:���d���P���"ONaB-O�&�A��P�F��(�p"O�y$��:M'���ugz��mb�"ON�*S.ϛY�>���
�$�5"O���t.�	P �D�4)���B���"O�+gJ��_�����"�����"O��34M^�:s� '�ħ�5Ҥ"O��X��bLiEF�JM���5"O�����q#]�R�A�{�)�G"O����/J���t&�&�=�7"O�xb��1t�P]��D,F`d@�"Ov�Q#GLq֩PqX��E�"O41k��Z�IG��(�	�~�l�"Oư�`'	(hx):a �W���&"O���͖8|'�Sq��<R�"O�����T905��f	q�S�x����T�U��y���{�h�'_z!��0J�֬���]++���"�˂�!���<	_�����!1��� $�!�d3qZ��c�m/!��`K.
P{!����N���g��v����l2[�!�D@�%wF��A@�A�\���8�!򤃃>��\����'l��顫W�!�dNk���Aq+MF�@=)T����!�䅐p�Q�#�GlֺH	�آ*}!�$=)��!"H�?B�|0��I-j!�$Z�E�x}z@JO�c����E���"E!���xR�e{diE�Pj�A��'�!�dl���h�>C&�s�P*2!�U�-��pwG�
��)�ï:�!� !>�p�՘@�2dB���2�!�ֻ�RL���6~.���@<"!�S�X�����b|z�|����d!�ӑxٔ�D�dm(̋�&Y�jS!���]�>�+&-�)Q����� 5!�D��h"t蒅^����!(E�2�!��<n�����N7b�J�r ǋ�j�!�$2)#~��Pc�A�Zh�E��&�!�;$�xhE��0��C�'��`2!����*u5�B�P.ZV�|?��ȓU��0���ťU�@��e�S,���ȓ=�"q��:M4a@�h��O�L�ȓy��𠊸v��X��^����W��ò(�����FF�.fRɇ�9�N@@v[�-�h�W G-6�
��LrQ�w��]}N%:d��0,�b�ȓ���k�- z��	�e�4=�ȓFd�1m։ƙ��"تڰ�ȓ��h�s�A�P��S�,=����ex ���T.5�A��d�8z���LXpX8Q �b��*��b�-�Q�<�K�j�5�p ,)3��I�gKN�<q�eF~=��K2�E'y�EQ��J�<����dْ�#7.O$z���p}�<	g�ʀnm�[S��I��Br�<y�o^����1gH��
+��� �y���!~��2��W"U�tY!R͎��y�$ND<��[��Ғ@��>��e�&�c��"s��1+���2#�漆ȓ-���t�̤W�z]Y�M%w�R������Ckԓ(;"���T�.j85��x�n�QF�(�� ���6'�6p��S�? D񵎈8D��s�n}���"O@qH��L�^�X�q��_�>D��"OĘ���E���q���  �D�	G"O�����4YU*,	��{�����"O,�
c2�2�F��<M$�f"Oa{Ճʶ>�-���9��=Y&"O�@e�+"\ q���&���"OxM�DI�"�rx( �-h���"OZH%��OYx��	#j�H�"O~Q���͢�J��ǰ4Wz@x�"O��(b�I�<��Ԑ$�C�Z"O�x
��ƍ'�,يRÙ(E;�\I�"O 0���ŭl�Zd��Z5"21Q�"O$-zd��B�����&�J5"O��r���T��u�C��$bZ��H�"Oj�����(`B��osR�I�"O��u���H�1u"؟F���K�"O4,A%1�j��w��N��}iE"O$:2�\����&	jh&|�7"Oֹ(�"ݩNd`��� �,�C"O���#�f3()3%�/-h� �"O
-�#�X�p����"�p:9�"O~9���L�CV���1���K�8��"Oδ:rfѽs���/��D-FM�"OxXs3��?-����T�85qA"O*i�� 1j���hB�zt��"Ov%�'�b�ԭ���ԟ�֤K�"Oء��],bh (��?��]A�"O����*C1a���;��Z(c�h��"Or\�Q�?m�4ъ��;��\��"O4�Z'��7x���)�ԥ�D"O��;�-	?Ђ��t��wP(�S"O�X��
;-4��b�g?�V�{�<�҇�	j����K@��8�q�w�<�v��{	��ҫ�lNZ* \�<���C={W�����X�z#�=�d�[Y�<��]+yƨX�nUb���1��[�<�$KZ?R������j��I���o�<)��FV-��I�C�!̬��@��o�<	��^�9G��h# ��D�Y	&w�<9"�}����O�"I0��#P�n�<)��ߨ]R4���	dRn`����P�<���ԡ@:��˂ m����&PL�<a��:x�<��튞 p:BŗG�<�P�v��&�]E��qq��A�<���̰[��A�&��w$�]{�Rf�<ᑋ��G�(!�@BH�$�KT�Vd�<�Չ��2w���s��(�V]����_�<���3}n8zW�C;,X��3��g�<)�cV �t�`�2-BiQ�/�{�<Q�L�oZt<!�-	c��$t�<iF���ё��r<�@1�ȓ#"z�Sĩ��N�lX�cfQ�|N܆�@Sl�H�G\ \2�m2T-G*Ȃ���paP10�c�B��*�NM�pr:���~࢘+����l
���,M1dU�ȓ7DJ؀��΢����C�/դ	��=�ͩ��û%.�1`!F�	"�4��b�|��Ӈ�����U�E��ȓ\mZ]Xe���<�~X*�B�T��E�ȓ5�D��əu��
V�R=}����4��Є4P�����e9'��͆ȓ%~uSf`�'VQ*�	 �/Z܄�z8�Q��J�i�B�9���&�<p��S�? 4YJ��
���йS��@sN @�"OX	�׏S/j��a9�}S�4��"OJ��'
�%����*�QPفv"O�@�$LD�~}���e`�;|2"O���%\�H�	d�ɣ���Pq"O�E����@�o Y_����"O��!�"�{p��@�af,A"O.�s'��X�h��5.p��C"O�5���DS�!�F4<&�7"ON\��1|����P�B����"O�`�`� x0����@;[q\P"O"}�e`W�q���Z�e�_t ���"Oj�RC� !!�"�"4i.%��"O �2�l��_�$���N����rc"O���P$k(�D�D�#�l��"O<�R�Æ'�%��CßH��dr"O��ІJ_�-���A@|$�*�"O0 ����:��T)U���;R@I R"O�}�!l#��F/����ru"O��!A�ܷ�Pqtnˌ}~��S�"O�Y	w��
D�x|����!yL�ّ"OV��#�+�J b�$q�<��"O�4��h����W��'j$%"O֨���0B)��`��M|\䑫�"O�س�U�,��8��@\1n\ `��"O���KΖ;�F@Oԋ{;����"OZebd�m�a�&G�
L�"O���P��B��xK���6�Z0�	�'$��Z��W�]�����d�@z�]��'����_I8��%��9V2@Y�'?\��w�e2┐@e;�
q��'�4��^�5�&E�BC_)+�2���'��p���ZuL<����:ZTr�'8Fi�A��98Ԩ�$��_Ҍ��'�"w��[�N����0
(����'t�iC�kݡDp��  W%����'����C�m} �0��d2�'�lB�!>jt���
�%�@H�'C.���C�/n������C /:}��'�>��!E�8��ZPaU���,��'�!`�'�72��-8R��lMĄ��Z�$��H�)�ƕ��?)����VpK��w���"W�� F&��R�`x
�,�*J|��@!�@.$U�ȓi�hc@U�|9�mXJn��ȓ&f�8u�:�m(�$��b�I�ȓ,�+풶|��)���_Yc "O���a���fD�IB�=jx	��"O�:6BNO�aY���:\I[C"O���AՔm�=����3�U�"O.d�1�N<�|4�0�%
�(`P"O�E��&7$p!j��ܠ�@Y�	�'{��[� /�v�S�'td��;�'p,�kv�\�w�z�!O�lg�$�'O�� �c֦� \�<[k����'3<��'!u
9�`�$XWBy��'�<����7Us|�!A��O�����'���&�A�4LD��l#pJ~(��'��܊��z�! f�+:���8�'�`@3��K�(�����9���ߓԘ'u��&�U�G��IS��B����'M�,c�-�)j{��q������	�'��8�T�Y<y�H�پbˤ�	�'�
4xFh��>>�)Q]BP A7�VH�<� �����N�����b 6t�"O*�ipꟀ{�ʀ� S��0"O�뒦[iz��gcz�v����'Fў"~J�n���f�c�	��;�~`Q�f��y�&� "񇇙,=�5S��ً�hO�����&r��CLք=,�hʓ�!!�$W�_�p�3
�r9L��h�;;!�N-}�p81ɇ5#vd��! �4�!�$E�:&z�F�=R+�@xy!�D�,0�x��kB�Up hML�X���b��(�����<o�P�o�8�J�"O,�`Ώ�q&Q��� ô�h�"OD8�0'�n���%D�o�����"OF���T�	!�D#F�P�i���B"O��X��+X����Xqz"��"O�e�T���\x\��tʗ2Uo ��"O�`g��$i�����.в��'�ў"~2f�\�[�N�١���XTΰ u�7�ybK�`k��Z��HF���MO�y�J �E6���8r��4�Ulޖ�y�g���*�i�?^�e���  �y���Iɒ�U�7T�Ը��J|�<I�#L�_R���d��Y�X��SE�<�p���{�9j0C9)Yܕ�d�M[�<)���Fu@��/||(YkǢK]�<��D�����Iu�+E�c��hO�Te��z�DW Q�M�Psr��'Wa~� G��|��O�&K�f�k�I ��8�O��vCǖlp�����͙c����"O>�Ě I��_.\oz���"O@�H�+l"��F�9je�q�"O��WoΌOl�q�N�(Xr"O�N��D��m3�ꞏo�\t���'�!�dRs� �C��9.���p䊞�!�Ώ��.1�x�1��_��@�'3��a�˜�4����p�ʱ6�z��	�'`<��Fw�&��6g�_P�!�'ߎQIU,���x��UǄ�Q�8�(�'
]"$��%�(�bƥؗM�h,Ɏ��6�d"X���G�1��x�+��9�������	ؽKF�-��j�0g7긗'�ў�|��5R��i��e�.�����y�<���ڀ���ތw-�/Lo�<1���4;Rm��
�Rdj�X���i�<a�g{5pmz�
ɊBDZl�ӧg�<���=��y�Ί�)1�T���j�<1��O<.�H�QI?RZ�:W�Qh�<I0+�|X[��F�<��J��m�<���(k�n�H�7�h�[���b�<�pED�sk��pʐ>{V�ؚ�c�b�<	7`l����da�%1��`U`�<����+&��.���Q�!g�q�<1 ⛴�"��d#H7}m�:���ly�|b�O�hb"@�;e~�%�1�]06�x;
�':���WF9&\ވ�a�QQ���
�'.>�r�;,�}!  �A��1�J>ɉ��	�"*~B�	%�J���\h�GY�X!!�)�y!�$7R�Qd�!��$@� �q�V�H�xz��Ęt��yR�Ih6����TiĖы��'����2扔Wc2�0�.� l��`�D�SF~�=����hO2<��.�Ḏ�ޚ4�\�PeA$D��P0���x��X�pW�O�R�x��%D�0Kf��$�B�:'��t���� D�� �xy5��Ovxu� ���`+�<:�"O�m0�/U	SG�1
�G� �p`�O�8��ؿ�,�hl�"8��m�'�;�O����E�J��uؠ��iф�W��B��Q��EB5YH2�@�� lړO��=�}:S)K�O|��O�!�X5��H�x�<A�CT�J!��TEL?6д0�k�s�<)�bE,kR=��^�L�"j�!�D�<1bK	;L�I9"��->�@&�{�<���Ѡ#���Q�(ۀW�>T���Fm�<�rC�K�T�sv.��/��)e�T�I}�x�a!@�6��|�G�]�o�I0%D�`��n��;2�[�W���
�!D�TBciH �:��殘,K�{7�<D�<��,�>"�^q��
 �n�[�j/D�h�$� |�V�أZ�4��N(<O�"<���� ��P�tX�oR���vD�A�<!uB�$b��H��WM���5��|���0=)Q�;�����w����̝M�<��j �>Lj&�FI ,1��@n�<!5�%v3P��w��]de��-�g�<�ы�`W(A �	X�F���I�<�qo�(+��01KX�wî\�p�B]�<�Ɋ;q�>i�c�	�M�B���&�V�<a�,Y���D��-[�a"�SQ�<�Ɓ�%�8 ���0n4nұe�L�<�8S��,�C)ɓ���I�gG�<��Iՙh"tu[�lr���!�Ey�<�ҥŰT�\q�H�<$kT��i�<�C�I%.��%��F��,����Pf�<1���M�AZb��"B�Z�RS$�^�<yӇ��@N�a�{/,D�g�P�<%c�6<d� u��//���P�M�O�<��,��p�N�Jp�!���`�N�<����g�2l�Fk�@Ȣ`r��H�<171�de��XVHђuLHj�<Q��_�@����LEq+�³�g�<��]�0�Kʖ�$�5JGf�<a�k�8Ea�%ܒ_t�5���Re�<�`A��J8�	s	�$H"�zAF�<�q嗉N禍�4���PWڙz�I�g�<���4�4�u�ׅ?��]�$�d�<q��R!m0̩��(�"$@�Ƀ�[�<��-J
+�x�cP�zƽ�d�GV�<�G�SR�ޔ�* 
 ��`1eeCR�<e͗�R�0�*�#�	s�Hq` �֟�F{��I��pP�e�bdڢ�%%׌#=����"OrP��� ~$��&���)Q)�yb�A	hr��ҧ��*����E͗�yBL�
�4��N�N���r(T��y��ڭ+�^T%	
��VA�w���yrnH�Y{�6�Cmz�!"
-D��c���
QזiI@!��\�`6L�<����S�I��D�W��Z�hXh��E�pC�	r���+�.�Xx�r��;�>C�		�R����Ţ�H\�`GE�F��C�I�u���D�(>��@�B�7��C��&�r	���I6n�q��T��C�Ɏ-F�e�4���L�I#��Ɇ��C䉢n�&��'�0FN�$Pt�2�(�=I�Z4�xJ��M�>yHT���kP�̆�`[�1�	V��
�����6 ��9��:�4ړ�BZl�� ��m�<��ȓO��\���� ��y��D8q����S�? �&�F:'�BhJd�ǨiԼ�1B"OʨhǩɺV�����0A�$A�V"Oby���"�	�z�c�"O�U#�/��H���&>��r�"O��Z0h�H��T�F�L�)�p	��"O��[�@�W��P��hM��Iq�"O^1 �fӾ_��i�X31�d(�"O���N##��%�a��?��1;�"O��d����ӖԊ�j�)�"O6�+��'4o�����Q�t�:��	z>��@X4E�����?��C�1rc�Q�6�;0���*�C\�e��C�?m�踠�����:׈[�Jf�C�	w��%#�e��bb�����&C�	<L��t�D��Gn�R&*lC�Ɂb��RFՓ�x����,����4	��r ���]:�U)3J@�\=�O�=��´8 ��]��%���%	���q�"O������n�*����C����V"O��r�L����Ep��4"O��Θ�tٴt��F�7�5['"O��gGJ�J����+�1O�Fp��"O��RagI� ��q�k;9��z�"O^Mq�+pG�4a���82����d/���d[�m�vi .]kn���!�dG�X�`q��? >��� �o�!�d_+c^"d�f!K$�y�#��!w2!�֪,v^H���
e�t��(ѻy!�$��8Q!�gB gx
�[s��+m!�d�6m_�d���O��5��T+_^!��pМ�n["F����j�4�'�a|rf�>m�tus���,�jİ��ɢ�yR�G�jC��ӆ�"]���
3�H��y�U�R�RU��#�DF�;��P	�y�iZ�:�b�k�Nˊ;��8k&��&�yRM�)[� ��2EׂHMrò�ӟ�yb��d^d�s�K�2�4Q��y�M��D�ܓ��Ы9=�0�%���y�-�l���E�d(�p1�j���yR#]�|޸���X�.���]0�y���8.d����� 1����ߛ�y"(
0R�`=H����`ʐZՏO�y�`�K��q��
1e���T�5�y�茍1�āY`��tADis�n�5�y2�w@���i���������hOq�b��v���?I�)6�*0�(+�"O��� 7t�+�J�T�D�ӵ"O>��k)(�jԪ�)�:q�pq��"O�,����;� q��cN !�L���*O��{���	fq�A��DrO��j�'z�L�7j��5����E�Z.y�'��0&��e��|9p�H�l�x3�'��xPD�*TJd�xw,O:R�����'~��F�)Z���F@�T�j;�'�(�`A��k�f���a�?�{�'���o]�H-:�q��
+Daj�'��U�
N�qq��`aj
��Tr
�'���ش.̺��$�p	ˢH�,@
�'s A�2J߸$'�l3!�O�*�e�'��y0���b��,����y��L0�6��Wi�V�� s� M(�yb��2\��3,ɊV}1���y�[����C2��7V���0����yR�%#�}�&#�K�x�(r�5�y
� �H��H^��!�3�!\��(�"O��Y��A>�0řv�c%���"O�s���y<�]�uϨ<0�t"O2�����"���r�B�w�!Ca"O�pv���p#��
���T"OV��5��4y9��:�2C�شa�"Ol����_�\ӂF�{�p�3�"O5 ��#� �֣�6"���#"O	�m�7���@BȷP���C�Iu������h�"�0�-�x�|�g�
�}�!��D-G-�D���@��)h�� �Q�!�_#G�LD[Ef�3b�"�P�o�"jc!��L�����U�g�m2DOͨ?P!�ތ<��3��ԑh�b��&�!��'OV��E�(Z�z�R�I�8H�!�]�ņQdmCX��u��+�6�!�D����ôD9[���Q*�a�!�d�=�ځ�R�-1"��BJ¹�!��I��̤˔)	$<m� h�/A�!�Ě�0Oz�A�M'&缨�B>N!�$�2�>k4*_�E��o�)p!��
��`-��x����+Y����%"Oz�$�;Uwࠒ1-�P�f��>ړ����*�ڙ���Q����kU�݉,�!����sDh�&z�|�j�U�d�!�r+gD�ї)\�x�9����!򤐙,�� �"zP ��Aw!�Z8]�|z���tiހ�a�'<�!�D��m���@�Ij�]b!�YG�!��aS�\j�G�;!�n����Gl�U��(�e�a���;+H�@��M!t}����"O�Lk����cI$tj�h�"OZɀ@S�7��LRvG
�Go�E{�"O��:��,(�.��g��NY4P��"O�ҁ�ݼ~��:���yR&���"OQ1 e�.�41��UQ0D�3"O���3kr�<�*2 x�X"O֨��f  Xn�"`�yp"O2Qh�'C\(��Cl&MT�U"O(9�a(�9;�8���Ou�]�"O
́ Kˀ^z�q�
v�Ĵ� "O�#�1 x�׌]���"Ojqi�D�TZ��X!�ݪ���"O��1�^5=���	B*V$i|6т�"O�5�1�؉���`S(��@UB�"O��zo��A�6Y���k���V"O�9���ڱC�q���L�gir��g"O^�h���	�fD��b��D"O�I2�BQ�b�@��фΎ T�}
"Oʄ�q� ��<\�u�"%@�Z�"O��^�	q&���S'Vx�G�'���7_-h�y3� �8>4T� ��Y�!�d������
�:Q������G�!�!Q���P ʩ\�Q�EFK��!��ף]��B�6e�z�C(ֲQ�!�DN j�ЍAE,]
�l���i�!�XᎸ��R�1k�y!�Y-t\ ���&?:dxZd��> !��U� �Vq�+ߌ未r爌p�!�d�#)�� � ��:�2%�����9/!��,/��Y��K�a��]	D�2H!���Es��V�c�����E*C�!��zqXMô�B�{�X��Ӥ��T!�$@?��v�O�[M����.��$R�}��� �:g�7Ŵ5�� P�Hiʐ�'ў"~�qJL4;�J�J��ӻm��X����y�Ћu�2q ��b���)@�U�y�N��lQH���%P�|��Oƴ�y��
\�؃F�=Qبػ��
�y"�ȣ1Y(�Æ$��H	�@ ��y���N8�T)-_D��$
/�y�l_�WL�=ѥ��ZXb0�e��	�y�`��{�:�)U�ӂCΩ�T�ĥ��7�O����`�&���B'S6e�HZ�"O�I+��H�T�MK���]H�e)&"O2`s��Ɂ-NE�����i��qAP"O�@� ��+3��H�� �n��ps"O �ZŁ׻g�����ݿ`�z�� "Oh◦	�C���4D�;Ix�Y�"O\�34&�:.~$�J��Rd�Bpɥ"O,yChI�:�RM9��Qr��4hW"O�@�䟐��hs وK���hT"O��R;~d�c�IÌ<^X@�p"O=x�(K�X$���ӯX'\�@{�"O�$�*�0j1�@�E ޽i���"Ol"�!�A���R���9�f�z��|��'�x�����,�p���!dZ8��'�����~�F�v��F��	@�'�xQ��oH�����](8�N���'>�����"�z���o͚/"���'� c�+�t���s�&O�c�De��'����En��\���W`��_-��'�ڝ҃�O�"���$����P+O���	���YU�EL>������>�!�R��j���	�`9�����D�!�D�g]؝�s�ˋK)�1K%�B�!���[��(�C�^2���ʲv�!�Ad=�	��e]#:��
��f�!��o��K�A¶-yT j%��;v�!�[���@��V�A��hZ���na�O�=��Z)��'�� wt��n�r�!;0"O~�''�-~��$�\�5Z
JG"O(,9��:=Vj "�@�9V,��"O��1�?A�D@"��8T���"O����IR��1*��ܶg�2գ"O��x���=>z!�d�т5x�3W"OFuBl׽?h��2�2i�(v"O89��B�B��̓+m���"O��
M�N�
U�u��{l�q�G"O�*$�GK���g�B
w`&Dص"Op`��^�+�4�)��-fB��3"O#n	0y6��F�A�2�	�"O����B�b_R��`�����a�'��I�4i~�QnD�+�l��t���7|XB�	���\�lO�.2I��+�( *B�	�L�p*��L� y� �L��C䉀b���Em݂5T$-���rB䉏E��h��Ƀ/��;�+����C�AH��[�	V��cFG�	�C�I e͌�����yA���$"�#aC�k��H�Ȓ=�t2�.��FC�ɊY<.$c4��R��52CgL�u^B�I${YT�yh%S�IrB�+c��[-�.u2��2��T��C�I���ϒ*^���ई�6C�Iw�:0#Pa�N�J!9��"^C䉺v�l�BV��IE��76��B�	�]�ܴIs�.|ۤ�*��'l�B�)� ~�p(ޥU���qR�D)b�ek�"O \[�፨�5�T+	��>Y�0"OyB���b4J�����B��K3"Ot�f(V,<���(��
�����P"O����C�Z�;��ہs%F�xr"O�$ѤʕB�8u�N+i�"O���mI�q��p�'f[�.)F`�@"O�E�S��;Kۖ0Y��+R/�8��"OL�{�Gǡ,=N��������r�"OB����Z�8��/�,����"Op�0&�
�y�j}�/���"O|XEI�C	���`�� �"Oju�3�I"�npi%�
�@�8Du�'�1O֌B'o�K;�=�n�7b�:��B�|r�)`J�i񦅙��R�;cw�C��:�~pR��1G�Š�JЪ+~�C�I�7����E$m��k0�"��C�	YZ�8xb�@�*�Y�h�"�dB��4:�Z �԰Jt{b�P�5+�B�	�C����k�&�8̐��P�~B䉪 mH���B[����eǌ�n)XB�	�Zp�J��o��P�&����VB�I�4�RJ'x��K�+�55�C�	�v\qHS?Q�̋��י2�$C�	�::�r�1������e�C�I!F�sU�/yEn�ɷ�� 9�C��?g��Rd��p�<�SuN���$C�I�\hT��Ũ�`��/A ;��B�I�7��`�#B4��SFd�j�zB�	.,�e����<:¸���.#u3bB�ɯt��ܫt��1m*��z�����"B�ɹ4��%"S�ưl3�艅[-L&,C��#��I�@����C��.b�B�	�*�����M9�ƜB`�Y�O�B䉅5[Nx�u�N�U�<�'��W\�B�	9"�����t[�����@�cI�B�	�0A�%RZ�&"i�RE_	G��B�	�K�&!(�.�c"�D˕��a��C�I�'���14�A�(�����e\���C�I�6� ��]49��}!R%�4aB�I�%98p�B�����@Qf{�C�I�CM�mY����6����Q�c:�C�	�~��$��#E�pu��f��C�ɭ/�@�Ŏ0��c���%��C��46��+��O�Kp���	WJB�	2j���SH�+ ��#��	'B�ɽ5���g�P4 p�0��J�.B�I�#�P50��/�0Dh�DP4#�B�&$rb�s�_�l�R�$��0r� B�1 tr���wE[�-ͬ �$B�ɥ"U�5���	?��Y�#L�L��C�ɇSBV��礕�Ks�$�r�/�C�It�B����	]��z��/;i�C䉿A������T(��dU5f�&B�	7J���1��&;|<�
�g��Yi�C��J�qc�W-m���F��lh4B� [�8������}j���e-Y'u$B�$�ѱ�A�=X�Ț��cddB�	p��0���s��c�
Wb��B�ɜ1 $d�GL�4,�u[r%� QHB䉫d�ɰ,��1�)kWK���$� �[Έ'�Mhg腍i!�ۿf�6X� ��c������>$!����q�=e��)V!3G!�� ���uF�+O�9����e�*���"O��B._	8�%�@��{�ґ9"O乡c�-��۰#R�j���"O�	��ՙd`Δ�$�Q�hu�PC"O���Ӎo� gaV a.�02F*V�y�O�z����fcAX�fH��Q�y���(\`ZI�dH�;�a�I��y��՜;����Wǘ5)8s��9�yBhٻ2�LE$L5/�\�@h���y�Ɓ�*9�@ł(J���^�y�g�E�v�q��\'|�h�&@�yB��h��@��g� 7X}���9�y��3q9�i�qG�% |(��M��y�F�c�6@�AX�ҽI�T��y�Y�,�A�k�u����3�Q(�y�;�Dcԁ�;b�섚��J�y���D&��YeZ�m��a�.ս�y��Q"3h� 䇕n����G���y�O�]��pү�:czl`�'�R��y�b��&�D= �ŗa���Q'�ܻ�y-^Wg�j�'�^���1eٗ�y�ì#wa�4'�U�p��nY��y��9*�V�ئn�Ku�sd�W�y�͚������l��$�H���y��_�da��v�Y;3��#u$C�	 1/�r�]���$"Se�C�I`ծ�yDJ�u�Ʊ�� �KՔC�	�k�\��S��V��%��n�B�C�	.}���J��P�ZR�K7~��B�,N<������]Y֮��z�B�	�.l����S
E��m8N;�B�	�)�܍3͔9P�$4!����B�ɺ���K	������ !#�B䉙,�I�K��H�'ZC��B�-9�b�ZH��ゃ�lC�yQ�b)D����]Kʴ���p!�A��K:D��Qa!Z�h�B��#�ؠ
����9D��R$�3冬�Q��6��a"6D��X�&8F���p� ����)�� D�$��!��M���|��e��� D�0��$�!_�h��-б"\��CA�=D�X;uF��Y��*���[��e
#H=D�l�VŞ�R�2�ǯ%$��i�+!D���R�WQ:��ɔ�I�|�Qa+D�Dw�\=]��a�ȈM�5b��6D���sc�5�3��0K|1с�6D����AN�4Ҽ�  ��h\u���5D�����
�Xز0A�nđ�L4D�����,+Q��w�dc�&�l�!�DţkHv�
ႎ9���o�23�!�Y��ʡ{@��7��(���,]!��2H�n��E��x��8qH��dI!��2}�i�$�9�hT�Y�'D�8��NCq�#�/v�J��7�0D���$N�9@^� �I�V�>�[�./D�DH��
vܤ��Q'TY"y(e-D�Ԃ��^�':�"q���L���?D�`���)����#��(!F�>D���'�Y>Z�q�3���|�n��4#'D�t��P%-��x����`(B*1D��xa)_�Y<��KQ��)f�12��9D�,��!ڋ<�`�� ����K9D�# �/l�H!pъ�0i����Tg1D��#�f��@Ej� ��/(�щ�0D�� &�a�&�3׊�X��8k�L�3"O���gd�OU<	��g@���D"O��P��J�T�b �	i�@� �"O��AQ�U�jnP�q&��5�4]9�"O� [BGC�]��8P�ޤyI��3"O�t���Y� If��
Nd\�c�"O�:t��	&AN�0���CL�y��"O�@��f	�VM­!�L�~� $"O�Rd45BD9��ŤHz���"O�$Ct�$d��ءÇ�A>�Y�"O*pH�eлb䂉{��!�@90#"O���%O��e86�Q�,{��@"Ol�W	&f<t�Q� S$gn�Ӏ"Od��%*�(v�FoE%[�y�"O64��gC#k1ȉ()_����"O{�BS~���H�f$Z�"O:�X4E�m���U%�dN�lA"O<�0�C�35C"D�u�X�AM��Qe"O 8���RV%�Fmi�	���yr$G���0��w���ؒ		��y҆�,�`1c�j�.�т�E��y�ȇ&V\�ފ`�x@BoW:�y���Co`�*�Ɯ�Y�&����Û�yb�˒w��0IĄ�8c�28X�"�y����ȝ��@R�rR�Ywh�2�y��)���c��f���)����y��V1x�n�ӔL�2Y�6i��
�y�"�2,#����׀Xq*�23�y�Ë�!����ȭIl�Lꂫ:�y­U�Z1��qF
�I&�I�k��y2�V�V�<���9��I�0����yҭ̫=p���Ah'~��FS�<���įt��u�,c�2��cSd�<���(Wd�S�d �FLh`K�x�<)��F���e��\�d�p`�|�<���ι�uͲg�5zuN_t�<�wa�;&� �rɑ�Y[v<�'�o�<�G˔�4�UQ4E�����*h�<�n��b¨m�&'�+Gv�[�Go�<!1,ۢqyu�a!���Ne���n�<A��;w�����kܰ`�j��¦�O�<QE��\,���Z�g�e�AL�M�<���έR$�9�d��#���D�S�<�����b�� �le숻�de�<ٵ�UӶm`���c�� �!�Pc�<i�.͡.��
 � n��䊑k�c�<���S�P��\"ٞ�a'��: n'T��`'"O#c��Z4K�`�pK-D�p׬ɛjI���&	�)$��h_�y"$�� ��h��q�Z�3�	��y2 F*q��H�ނ�m�(l���F�yRm";�0�IA�D�N}Hi�a��+�y"�X�u�h��6;A�R�i!hC��y�'�f�@ u����ua���!�y"F��xzy��óUV�����J"�yr�W�c�#��:��<�����y��ؚ��XG	�f��0 ��<�yB�K�7cj����T#�T;�@V��y�-y*T�$Nѝ�JM�5�#�yr t@`P0�%�<}�dH�)�y�-�RB�\I�-MS:�Z���5�y�Y97y�L�� $8& �B����yR*�a���" �3/��U{
M��yz���i�<�n1!B��
_�9��S�? X��֕3=H����M�5�@Ag"Ov-KG�(3���WKW�r��"OJ�&F�p�e�0�^�]���Q�"O���s�e*`����<�(s�'�1O����K���zDK�0�Πh"OFdi#�\t�I@��䆜c�"O�aӥ��KvP��(�ݶQ8"O��0S*.��T�"��{2��`"O��96'Z2�(��a�B�̬<��"O���ʠ.c���@/ɑI�4"O,��iȰPl��R `�%��Y
�"O��'��h?��㡩�3���"O����=A��r%	��l�|��"O�Y�Ģ*S����Az�d|��"O��B����c�<]Õ���E꒥��"O��R�Ұ(O�j���7��!�"ORԲ&F_qd� �#	�$�"O��3���!.�00oÐ
oI�T"O~�{���,:�u�f́k���f"O<���dݛ,r�T0��4iRHa��"O�!�v 
�[����al<��f"O���0
O�@% 8X���}WPU`�"O�\q�Å�R����Itf��"O�l85�
�0e=�φ!U4J�"OD���F�*4쁹���&@ص�"Op��oA�M�1 ��ަB>���g"ON�yq*ׇv�PK!MN A�y"O��P�i�_�j,�1!,4�N�*�"O I��H�=�BH�c�`��%�!"O^}��g�@-B��4�ٶI�=:�"O�mF���f<�DO��xs"O�8YpK�34P���a.�� ØU{�"O��3iB?T��@JAn��1�� �3"O�� C��2\�m�3�Ҍ-zTh�"O=c�T�Rdxi�&�9�p�`�"O8���%"J�`����"OҠ"Q��<�H���g�/7��p�"O��+PS�2�Y�iUl�A�R"Oj�±���n+pXB7�Ç �~�"O ��([y�҅hö^Ţ��"O�h`@��i�hd��2��(a"O�jF�G���1�f��b�N�2�"O���R�B�H�K�3^�t=b�"O��3�(� ZW����5!�BxR�"Oڍ!Ó�tX��ǘ4"O@@�cZ}*%q摉O�$	1�"OTDI0��IW�]���n��l(g"O��� �~A�d���f��X1�"O,�8WHU$H�(9�/=�Ru f"O�<���Y�{.$0G�ͺ��u"O������b%R�[ ��		B"O^���Ԭ|��F#%� �w"On����\�.���Iae_�݌d��"O�I{@�Y�h���Ú�AԖT��"O�1��;]�.�b���5T�pɀ�"O��s�C�m�إ)��g�h� "O؅Y#�F3:D2�Ǧk���"O@i�ߢyo�T��E�C�쨳�"O��8!���0��J'@z���"O
, `���p�P�D\1A#D��v"ORQ�BI &i� �dcJ8i:�M(�"O�
$2D�=�L\�3II�Nb!��)/z1�N6<q��I0�K=uG!�d�9�4C�լSR�YS�E�m>!�� �Z���5�a�sM��NN򴚓"O��2���-F���UY�)�\�"O:�2$�LL� Y�(�8cpV�@�"Opu2�@W7���ڡ�O'r�,�"O�.}�.E�.A=;��h�$ݜ�y�M��+�Dاm�7E&E�Ć��yb�ގ,,A¡�˚B5�aN��y���<~�\�$����s�ƅ�yr	ȫt%�"��MZ�p�j����y�P�!dȰ �κU� �q���yBL=v��U��U)���.���y��]�@�b�K�`�k�c5�yB ˂t�P���y�U�o3�y���E�8���ːz���`����y��7Z�jU8�\n|�P� 1�y�I��m�V�b�lG<e�a놀	�y�9��ܺR��Y�����H��yN�0�P��̈z5�T)!��>�y�*ĊhJH1G�;'�@�e�I;�y���(e{P�)'S�/j�"�Mʰ�y"&��ߠ �u�L"���;�m^��y⏙�t��a'n�%��o���y&�����Q:	F�):b����y�*Ӯ=�\H�lؓ{� ۢ%[�y��7
g�� "ɂ-\�%�	�'���[C��C	�-b��")3\�i�'9�M3
��s��8��� ��S�'�5�o��E5�ܫud�	�le�	�'��
PN׎�$y�!� Y�v���'�l�ϛ{a
����+V2 �'+f̐E&��=��iY��ӘSԤ�q
�'~$�)&�"^�;T�I�6���'�8|j%
T��Dg�9�����'s��R��п@\��he@�+��+
�'"u8uDƽ��1��N�ӆMX	�'�8�3T.�$S��1V����'B�I��ƛV)C�턉,�N		�'Lԕ��	�V����R�ޮm48,�'�ȩ�sd\�H��2b�k�z�Z�'i9���D���rN_78#�%B�'_͊ׄ�y �Q��U�0E�!;�'H����M�H���2���/���'���s�ف_�N1*gC&�� �
�'��\�էQ/4:4pX$$��"9�R
�'���7�$.34�H��e�h�X	�'#|Hhu@ƠR�@+�1*��m��'�&q��0E�BأF��qnT �'$`Y��)�x�YF��)�
�'��欂0#򱘶��3x���'��@��31�a�%L��Z�
�'2��5��[�j�8���;�h�p
�'�N��fM,Ӻ��fl�y��'H�"@�IW|  �ݒ(���'y�i�vfC��+��Y(X��:D����  _��J#Ώ�o�r��8D�pp��"Iq��R�c�6��x�`,D�l�"kܩc�R�ؠ���zWv9s7i*D�T�
K�5�f�X�� ���'D��K�"���\�!h�*
��1�-#D���AG�w���h�v�R�Z�"D�ȀW�A:|��a!w&!x��s��-D��H'	4Q*����
$OX��x��*D�ܐ�L���<I����U���3D�4s)L�nx� �@Ɓ-G@Mڷ(3D�� P ��d�~�Y��*4���cU"Od���U?BuP4`�@�/t����6"O�|␮X�U�l�1���$�*�"O�%"�+ɉ���iCK�+K�ZѐE"O�a���")f<8��*������"O2\!���b�j���ճB�"�0�"O(T��MQ3ԥ�d�V�vz!jc"O�Q;���Yo���#"3�01�R"O���(�d����E���3�ސ �"O���G4#�\��CN?5�r���"O�X"�'�$��	��B$B�
�R!"O�t��ϐS�%�����#BHB�"O��㛨���u�	��)��"O�|�C)K$:����&M?Q��Q�"OJ\b gϸ8�X\��N��X,�y�B1��,�F�F�p^�X�!&��y��]*Rz�9����<E ��p ���y*l7��� �/>굨����y�K!S�`����,/�u"R��y� Q����6�@���e'�yB�[�(�+�W��=�1��y��F�=c^��`��	��A�����y�O��n��	9��l�N<�@��$�yd�	bb轋��c�ir *�yr#�8�.y*޸R21yc/͉	!�D-%w��ENڡ�j��(*!�Ĉ�tx�%��"^�\	-��!�D3$+�e����2�����}�!�Ď 4t��*7�N�^=���ug!�DK�A� �9�h�ٔ� F�U)P!��<	����QbF%a�G�k!�Ý5dRr�$`f�*��UX`!�$ʞj悥�V@��}9���6K�8Q!򤏚�|���-ŐYq�$V$9!򤛽9���05�	5-�<��&�A10!��2%(�2���UG(�K��� !�$��t���Q�5	'He��%�q!�<��(� ��b
��P3EI�*!�$�����_xM0Ĉ�F�!�ա/�p,	6�:yV�� "G�!��XBFI`T�	%��B�@�7�!��o��5B� ��fۤ��6�!��˛T���0`˦7�T��FA�8�!��f�j�1���	���"o�e�!�d �>��91�^(6�޼���^�!�䍒a�<��'\�):|�����(%!�DF�&��|���@=5 �e�t/��0!���9:4��{e��'s*`3ɫ.��_��(�ʔ�D�[<+��9�'�>~S���q"O�Ca���y���d��0<�|@"OP#o�5,��zZȕbJ30k!򄗣6�ԓf��C]�s� ��@Y��~�����Æ&
�>%�	��B1d�� �r"Or��@��#֊𥢃P@`�PR"O���g�S@D4���<���"O$�0�J
�0= N�:;#ԠBu"O@���-O�u0&�
�I��ѫ&�II�O����$�:*Hɸ�Ᏹt� XB�'f4�!�����Ȁ&��=F}��Ob�=E�DO��0y�(��KŢ}8N�*DM��0<1���M�#�>�2�A%zH>5V���=(�e~"�i�ў��Ϊ�r2��V�%���щ;�(��hO�~~� �5zr�c�� h�mChC��?	�A'�S�O��q��"�%�$@Y��Y�j��"O� �1yk��>V���CO��ќ>aÓ��ɇEmd�`�RZ��1�.���J���ɱ"}�?��#O5G���U��D��r�"��hO��W�И�f��Cv � �`
���ay�Z��?c��@�/��m��ZE��s�&ђ�`84�<��Q��N,rӄ�82Jx�c@�0��$�S�O����V*$���P`��nrlp�7��OLdJ�����YK�/�J{��	��'��ĈФ�{Q��=L�0�e��=,�!���"s�����N�2�嚛'!���*Y̚"O��Cv�X�	!򤔑7Qx��Ó5� T�!�R -!��J��� ��f�2��֕1�!�d�x*P�b,
wBlQ�c��6��';ў�>y�3���"����#�F���N6D��'.�>�<(�H�j$(P�`j�>A����dT��Q���!�"�!��2v#<�z``5D�X�s��`�*,����Y�I��/�%�S��v��Օx\
��q͋�|)vu�ȓ�ZEҖ����b��J�Y�.��ȓ�8����V��cĞ�MK��ȓ"@Z]qV�N ���H���8��Ot���͔k��m`��֦.�cS�Њ@!��+��,�P="�@yt�!B�!�D��	�\�+F�Q�T ��,�X�!�M�Z�:i�5�ҍ8�Ly����
"�!�̐v]�0B�(w}�`B�
�a!�X�bl�xc��]�>o�cjEW!�$��G��Y�abJ8 u 9�(	�vT�d"�O��סB�^vP�R��C�����'��'�p�cB�\wWQ�cE1��Ex�'����#�/Y�v(r��={�� ��'D0}y���{�ʜ`D ��)���
�'L �S#��YU|m���[u�AY��������d؍.���A�V�;�6=Z"�CFQ!��(�^���!57帬�mB.3�!�L�-7,9���,�<t�l��an!���O�i�g�"������	f�x�7"O,��%���G:��0�	�lG��"OL�bĔwt ���[�v<���'8�'�F͉����C{�q�SA�b�ء��'
:P����K�@��:����y��)�5C��\б�7>�ukt��c~�C�I�`�ɻw�/G
�(��Q�gP�"<�ϓ7������s$>�Y. �=��������"�K�a�\�@�X�	[�HE~b��8R����Ms��(饊O(?1t�� ���'ْh"�q�4�-��$����hO�>�*!�;O�L�x睐'6�DX��=D��.�3�V� ��'6�PS@):D��a�M���FЀ�! n��Q@�O��d5�)§�y�.��i�>ȉf��d&�0n��xB�'T^ �	?\�UA�fZ89�ı�4���>���T?��J�sӾ@b�T8wd�*ab"D�HY�@Ӵ8ݾD�����	(��StM~��=E��4+�T���)i�N0��:8���ȓN�={rT�6���I7�S���0�ȓp(���V�:1c���Y���l�Z���O���& u� {&�6�^��U!O,�B�+ߖ�*1m^<V$�A,T�k��B�ɵ`�@%�2T���{ �ռ}U�B䉠{�鰠e��*pm���?pB�	Z�B�@)�$�f o�PB�IB�������'A2��FџwE
B�)� ��"��$&ݠ��s�ݝ,]�Đ "O,8���t�d��$f^�CU ¶"Oي�c̗|���`Ǐ�0Q��ؓ"Od�2,����U1�ޖT� �1"O�E�͈#��A�S��\M��%"O4��&����b��4�F�+��@'"O��� ��v��t��Beιy�"O0�$��ic�%��kX(n]�X�"O���c�w
R�	!�>2��2�"OĬ �&��P��yP
�,8�i�C�'�ў"~r�%Ҷ$B�zs7N���kסO>�y2�'+f���DI&*ұ�G�/�?���M��A��d	O����س@I|i�ȓE��EIdG�n]D$3� �/���ȓR(��K�k�"U�$ "�ԅ�� 9��&ֳ"��	cs�
e�4e�ȓ{�8�"׎U<Gr���c�cG���ȓE��H��V(�V�p� �E�ꈅ�����O�B�Hs*��1"ȼ#��Z�J!�d�)�5B�"H�:�@�c!�ҿ
]!��]��PiQ"�fr�`cD�ʚ�!�ĎL�e���=0�` cX��ay�I7c�:�"GO=/�����Ů'��B�I�`
�ɻ�pX��x��31uz�h��(�S�ӑc̄H��^�`F��B?juPC�I�4̆,��ĠH���#H��|�C��4�p��L�p��\+7왥O=8����<�$I�Q9�'Jh�ْ�L�<����>N�>��U�Ԍ .��ׁ�m�<�@ܝG�Ȥ��jG�&��A��Z�<!�@*o�(����w2~���w�<)ѭ�/��L{�(�GCj�8ԩ�G�<y�N��2�:�Sa�\��h�3I�Z�<I��i��,�Bkΐ��`��kA}�<��F����#AM�[���'�^�<)��!�)���=��ً��NW�<��H�<Ad�S��K�{��mS�+
z�<�f=6���j�cB�/��h�$��w~R�'�F��Ù))F�r�b�)T��9����ɝy]$�B�֥6'I���O�#��B�#�U ���s�Dk#�?75x���U0GE�?��5������=x�0T�2D��yo��"��1��18~,d�`��M��)�S�O�$��ǿ#��h�
�Hr$"O�Q��1F��	j���9��Q�"O��1C�"%7��� h	5Ԑh1"O� �n�2!&ݫ���j�h"ODEs�
�������%0�Z�x%"Ob��GF٭X�lDY6'BM�Pd��"One�D�A�@:��'�	���I�"O<�"ĪOU$u��(Ό	���T"O�c4�C�00�b��$L"�c�"O� s�IH(HH �HL�hn��U"Oi����<W/�H��gD�i��§"O� ���!8DLhp�[;3a�x�"O*i�b 	��,!$+��}��"Ov=�C��D��Q(aё7G��i"O��r��D>;/�%�Tͅ$b>��x�"O
}��Ж9����tkH�n&��PB"O��P*�0X�Fi�p������^�!�DØ���$�
�_��e��+J��!�$�؍s��N�s�R!�Jٳ:!���[�.��Q����-��C
!�$��cBh�r���a�[+_!�� �L����w�h��#,�����"On��ȼ��l
��7PcP��"O�(A7
	���IO*4���"Obq1PbҪ?9<�@�S;ND�a�"O����
Z�½V$L�ҡ���yi�"m�\I��"Q�f,�af ��y�+�w7�h�GD L��8f�_��ybGQxG �����4CH�ݸ�l��y�Ǔ�D���RH	)sV�����T	�y�a�FGf�"4""��ɰ���y�	\,]�]�0>@���y��.7��ԋs��lj�G��y��/Рej -S	K�p�6�yrjU<w�|"�f�:*�5� DN1�y�gC&}K���k�})���5�y")I&u�(āǱ_#��a X��y��J�2�9� �֮ uV���%J��y���4? 8k�#/7Pp�V%�y���tܘ�`�	��P�FL[��y�-A�>1:�X�J�0��d�v��y�#G�+GZ�"�0 �,�F.Q��yB���=�HL!��\75�!{e�L��yR��%@��Kf��|!�q+�>�yb/�7m�tU"◇t�@�T��9�y�ťe���u�@�u�Z]"u�U �y��҃Jj��� �a��2���yR��sg*`�Qdx�]��ʃ�y2g	��	�'al���[��yr�Q�G�$��c̆[z�pPC���y��\�C��-yb`U^;�zo�m��')�)�vL�� @��!U*���'�D $�*z� �[����pA��'��k M����8B$�G4�p�'��b��M#�H@����M�yC	�'M�1��厩�N�s(Q%G�z5y�'tܰ��nu�� e�2r`aB
�'�ص�ƒ-�P�P�$��-�����'B��s���E$�8#b⛙!^���'.yڡ���oY������s	����'�9�FaY�:{�)!to��tl��Q�'��t	�hE*I��4�9c�P�'G�!�7$H�4hD-�K��P���
�'�t)�v"�6	��q���ŨT�����'G�Uq�P�%H�r��Ұ 4�
	�'�����D��}�Τ�TA�Y6�pH�'���jSA�8a�R%����$`u�U��'*\�V�S!e��Ę�+7jŸ�(�'jA2UV�`
Z!+��]�;����'�D��k�}0	��l�" `��	�'����1fN?r<�� £*	�'�r-Hac�	J|b!���:N:u��'�n����?$L�P��3�v���'�<��EI�B�`�[�z�`���'�^Tc�i·N{ར�k�M��d��'��ZE엒Z�4Z3��+'R�R�'�H��`b�7�y���I���(	�'�VEp���=z�aaӇ۳a\ri	�'�9I��X4r`�����d��x �'٠9h��Q	+�֨Jr��$gu���
�'U�dg��O�
��A-TX�@a�	�'��1�Q��=�
�q��%Wd.e��'�m�"M�2zgj�sT̍�M	B���'�J��!X�?��� '�'i�$���'������Z��*�dH$p�b1���� �-����$U��M05�ޚ8��r"O<�da�m�nኲ���D۞�H�"OVX�`��z@�I"ċ���F��B"O�l�kW�9ֽ��J��j���{�"O�=��� (��d�$H���D{�"OV-K!AW�]�(��GH�)V��7"Od�BG(�-W�%� ��-+���"OTc�+Қ/��訧&I3F,4-X!"OP�z5���i�UA/��E��"g"Oȁ��̠*N���ư$$�W���y�����I�E'�W���j����y2
��(MI�X�Q���3ʚ �yb�M%o{d�"a�8p�`&;�yb�U!u��|�2�C�a��a2�[6�y��X�lP�y ��	A������yď"y����`IJZhx�#K��yb�@1H�h(�`��V9 ��B,�0�yb��<6���'e�,�<ģ�枤�y&ۉ}LM��ǈ�	��
@��;�y�iF-=Θ�
6�SY���Gχ�y�M�5G�i����L�Z岧-\��y�,TP�0�1����XI'�@2�ybD�6UA�a��R�t(�l�!I5�yR�F�flI��uy��Y�a���y�J
�7	��GF��xs�(�<�y�M��|�:Up�����,��"��y�DSTڼ�"���C���h�	��y�f\�tJ���NU�O�������yG�#<�\u8��?��T���8��'@��r�9�\�O#
��C	I�&���qC$R�^9
	 �'��ᚗ��RF�V�(U<\�egL�{��Br��Qyb�������$s$�0�%ַD(J�၁,�B�ɤdD^�@k��K+����M8,	^�Y$��7�ze�Ģܾ[sڀ�鉠t��y*Cf��Xf���%�	���$��[n�W��oFH�w�],w�Tc7��� �as�"�5��)#bO�,L$<�V$����+ue0T@�@�B3kDB�W[�1ń�A�.(�d�]�kp���3�T�_��p�U�T�R�鉯ft2т��y���2D�"�9ʐ}����S8�	��E�+fi��L�'dP��L� ��"�.n���#�̾�v�zc�5�$L>�x�B �����fA�7��
���%)��r]f�Y�gS})���m��Z��Hw�ƚ԰<�pG_!u����d@S�d�ha*%}�rי>��T ��	]' �������U�$e�O�|�t��Qh��Zpl�Ӳl*P������}�pX3�]<���$�ڎ>�V�q��޴2�����ᎨK����#�E�D��QG����T�(��2n��T�`B
��0<�W` gc�A;��ÄP�ɭ]Q$����@,]�5��D��t��U��:��*PeY��M�֯��?Mp'��X�3?q�HL�&��hf́ �䍁U/�fy���2 `���W�	��(�O`��-�Y�6lΧ.fVi�sC+*�^D�J�}>�$�r&�<5���"(������'	�3w��9LE���TZ��V�4 A?pC��I'X�D�@Wjߣ�3��O8ŲbG�Q�18�ܻc�Θs�X*&��3rg��U%����u��aa/޼����.�mn2a*�����ˑ�j���֡���/�=�蹖.:�D�>z���c��a�t�%�0Dn~P����!���p�ֵ<����yO�0�@��?��p(7jJ�HmT��� �q8���p�����K���3dH(���#�삾v��m�'�n���Ͱ�н2��O�e#<zl�}�WN�8/��"����t(�馁��
.�y2f����H+ĵj;���!ŁgR�Ԧ��b
��+C� �N��ڏC.6X����(�Dk�'H2(��[�A�PX�'��<�4+\�%hr���+w��P��B?3
�1b&�:��jU;ci�pXAh���4i�K�~BK>�D
�(��$��$� ��2OP<����^���=C�4�w-�S�V��A�	�Ny:��Đ}�0h��D�.���'���<�7��;O��25�X2b!�b,�@�DL�e�F  �O�0��+Ԛf�`��I�i��v�:=��fN�E���#�/U��C��4p4|`��J��
�C�����8	"��F0_&���·�/e�Q����KCg�H`၉,�e�Ê��yBG�>&v�P��E�h�Ĝ���Y	?x��g��{Z�)̨[������|
� By��.� mI���I6��:�O@u0���[jV�����!������Ӟj[а��	 �Rߨ|�>���$J�v���$4.��a��<^ax�C�'��Q��mJBr��ɲ��%m,�qs�D�3$qS�ړ?3!	�O�Q���ޛ`�Μs�gK9uo:��ѐ>)�@��q��P�U�@=��[#,>�'Z<��Ɣ8J�4�ѵ��ijA�<�si,)�p]���4&�h�6=����2ɗ�)Y��A� ��4�||�}&�L9��ۊP�pAO�X�� c;$���f��HԨxx�,O�<Śy��҆fRT��$mJ$�� �̉Q��Ģ���}`j"�S� �NzӢ;,O����&
D� �F��[�v�KgⅠA=҈���#?�<c�mXl�<�T�ӡ���Y#�4�0A@-�h�I�4�6M`V�)M_*5z ��^�O�����/0N��KU�8x�Nr�'�>�@p	�!x�������v�~����Î��)��
ɮ�~�\~����3vb�w*ȝ>��Q��"
!��T��d��̛9�Ҙ1�P����&Zɨ�+pnL�Q�azBOW0�"d�@a�q:�8�����p>q�`�)Yw���EG̲V��R���}+1��%c�'9�M�W`Z<i�F�yT��+�������81�e�נ�k�B��}b�,�G�p����t�� u�^�<�2ϟ�qgZ� 1�ŕhÜ�U�
.��=(F�T@�f��P?E��"F�2;,i"���R��0�ȓ*�%(�&�i�8��U�5$zj��'XX��i�w����'O�;�M'T�F�rH�i.�����'/�����ݳ5�J$���LE24�[���:3赚dᅃ�!�d@�HI�A�D�Q���];���Q�,���L��C���I���']����`��#�!�p<�xQ��ͅS��$��	����3��e�!hAA�O�>�b¢YBݒ,B�}o2�2e(D� Z�i�C���aZ.�ҥc�*"}�C�X6����D�,�bR9|���p��7�y��K$�Ox�:�@�	J!���$:��My�*ˉG|V�y2�ğC!���#[�(�1m�a*�	��zG���Ȓ�	4r$�m�}�cC�3��Tp��ԟ��Q���Y�<�ÄF%ѦA��Cܙ ���iJZymNpe��=E��n��}-��F�C��M�c�.�y���{�X��	Q�sm�p+3'�y�mq*�q�'��B�������yr�F1c'�E
rHY6���d�y��ׅYF�8��r�HM	g�݀�y�����y��hM�s�r�C���?�ycM�R�P`�-Ȋu� ����yr���\�h��@��lG$d��.�y�e�$Sfҙ3��Y&0�Ѫ�y��!��c�6T�<��i��y��>9��@k֭eP�T
�)��y�lS�q��TrG �DŸ�M��y���%=�"@����z�pؑ��yR��c@H؃HM.o��l��㘧�yB���t�	����Z��)�3���yB��N�9�1ɓ�,H��q����y�;�IA���]Ya��y"* ����)�"�$��}��lV��yB���	L�2���?F]0s���y�M@* \N,��J�vX��2�Χ�y�A��`�Z�-vzAx����y����h� H��^}X*�x�g�'�y��K�<�|A�S)��Y�}"@�Z��ybJ[5@����\
m�:ĩ֎�y�
0u������?�4)@gFT+�y2bMM�p �b���<@�<�6L���yB�5��Y�nO2��t�fӡ�y�)�WE�Cs�G�6�*%a1��y2���B��򮕁)|�� �_�y
� ���6�ٝs�
�C���
a����"O�yщ�%Eo�)�q�
�T�$ٲ�"O�Um�O7���g��6�`t"Ofl��eٰ@{*E�P�d��В�"O(� � E��ҡ�D��]`�"Od8x�n��"F0�@V�H�`�I�"O@��T�˱x�.��kD��>q�T"O(Uc��0�V3G�X�z�Ū "O�L�����3�\ �/�-?��i�""OPl�"U�z���)PiB�[�"OB=�ʃ,���i�FBE�ܚ2"OHL�BY�4(�!҅`8mHY�"O�����O�Mj��9�o��J�[C"OBT�ªg"n�A�u�q�"O��"��M�:����U��0P�І"Op�ʕL ���u�3�S�a�d��"OJ��5������(�MM���s"O0��)��fh"�R�����P	�"O�y�g	T8fW�0�V�2)��T��"O�����7����X�*Q�"OHљ��7*X���)@* i��;�"OFT0Ce���(7�? X��#"O�P �'
6�Đg��#At��d"O��#��'hJv�� �2<֙��"O�l�qC10�|��F�D-�9��"O�u��jQ�1���b��Cׂ6D���$I�2���9��[<Ĥ��a0D�8SM�/L)qGo�%pa�`�Cn D�ؐ���.�@X��%�3B��s%� D��Z cÓEH�e�`B�$ZBw�?D���n\�y�d�Y�&�;�|�vF/D���'�U�@t�+�K^�o78T3t'.D����fO�����u�^#}�����N+D��Zq��1���D�Q���	Ad$D�������Y��9� �#��Z��'D���GED�(i�q#Vm��0� D��(r��l�R9��Z�
9�1�>D�L�"_�t��	{��C� � \��:D�`b �	�w5�<����#j���9D���/X��xgdI�k��-J�O#D��A�GɃB5fY����,t
b%D����ڨ.g��3T
��B��-@>D��9%M������g�$_���*D�d6��ZO�q(�̇�<��!q��&D��� �J����=+3����'D��sD�� �>I��2	���S��%D��to�!d�)�#IѧyEΩ��'D���f掣f�Ё��mE�/y���%8D����&�#C\�
�,�
>��5C�( D�|�ԿrϤ���G�r���% D�@��E��n��Y[�#�1G˲����$D�\����d܎@ '��㐼pWM?D���#	 >�&9pDl	�$V����?D���I@m;�5p��� � c5�?D��H��Υ��m a��7�$�@�<D��B�֒]��hi�䔒q�4T��6D���B�$F����ӟ_Z:��@$&D���Ṕ	B|�A�ʹ`��=���'D��j�ώ�KP"��a��鲡�Ʃ7D��J���/v��&`ϵq؞��'o?D��R ��e���@�fM�5HY��?D�l�V�Ȟ���2Z1%�%�T�Կ�y��ס�xh24�F�rj��ƒ�y���Q��ɺ�A.�Qh�a�%�y
� ����$4�(�2�H	�|�&"OrL��c��J�\p�wA��	��hau"O���G�eg�PF@S������"O,����%7�����ǳ[p5*�"O$T��g��gvh\�1恦a�5CQ"O�P�a�<���	4o�4Ie�\2V"O��s��n�`�؆H|�q�"O�}�p��.�-;qLW+b����"O�]�� +Ai��`D+�b��"O1wAؓK,D��`�=5VЙʅ"O�}��i�$MF�X�BQ�6$S"O�հ$Ȅ Y��q��׵%^��Q7"O�m�����Vp���0[�t�"O4}+ǒv�ڰ��Ȧ	|H�A�"O�Dn8$!�L-3�`��Q"O�"d�:9��"J��L����V"O ��Q/_Ib� ���QdZѕ"O��ӷJ̧30ї"߀9881{�"O��t!��Zi�4`I�S%�DK�"O5+��sYb���M[!H+�9Y�"O���_�61�tL->���"O��¬�)| �upw�W�T��ʦ"O�����,G�)�c�B&"��
�"O���pX�j����K �1�"O��I�@Ǎ �=C�L�%�+�"O�h[���	*ʂq*����f�a�"OJ��7KA%C_��C ϋx�Q�"O��p��.m��(g� �GB��Z�"O�A�lFy�&���W(=4"��Q"O"��g.~�F�!�� j��"O�Y�g�%%*�qr��0V�as"O�����X����6
0 X�Pu"O�=�c��}(�8�@	�1}�������xrB�c��A�����`K'�E�P^�ҡ��$�<�"c"O����,�l��|27N^t�����ڈI�����Ϩ<Y�n�v����I��H�x1�O6
�>��*��:š�DN`$l�7�ҳnR�*���"R`:��d�~$!�F�#^���O|��� U��08����B�_�yr1<���Y[ ���7��<�А�@ Q
J{�����O�xC�I&Do5��`
��T�I�dJԦгK��D)JO8���O@�Bg!������O�4H��J�4��
ㄒ�2착�M@�Y�ҙ��DFR�t��I�V��"��D�zDA����� �f���(7e�y�g��I�A'��R�B�oH�(����')��'I�<��"&*��D�T�	]&e���K('=�C�䄾%�r��E�S�"��;QMD���	�&b��f��}	���@�;�BY:����+t &��O��M�"$"p#%NA�S���I�̝%H�����jҫ��)m��Q��'�(I�v�S�Y��Y�Ƣ�>)ɘr��k`(�u._�h.�E�âQ*0�Ղ��)�w�&\1�δ��/,M	��'*�0�چPK`�(0)�>��B��_#� Y�Z:7k-(���K(���U��:��NMڦ�Y�)0�g~�H&~C*�b�/S�t�ҝ�4J����>�僚�v�^y����Q�O��L� `��l�4,&� �|�����*L R�ۦ�C#b���׊+,O6P�/�l�X�-]�6ݤ �r-�1�����o���E���g?ɂ�
6O���u�W7����$��BȒ��.۰?�5P�4"�	$��O|�10�P�CR� �ScG0���7���bE8�{��z|�I���t��1Hum_GV2�E2�M�[s��+����c�'TP�$�
G� �!�%CO,����p��p��`YfQ���ǭz�L��'9�yɅ-!���#��O��-�t���j����F�y�6 ��'�|�bCC5<C�a����~�0��b�7}���$I����{"��%I�h���J>X@9�C��?dL�Jw伛FO�ςJ�=!L�g�Kipꤳfo1�O��U��+~����w� .�@�c��'�X�S�l���'@pMi!"¤r3�AQ� 1�l1��'��p�cP-q
Vղ��,/���)N���E��8X_qO�� ��2�9�}!v��+Z$ ��"O�)�f��(PO����Y�l�"Њ�"O�dC���.(CO�n��P��"O�{��Y1:=��
��Z"R�ta�"O ���P���2E���h��"O��Q�B�I&H}G��`��m�w�<��:����@��5(
QC�J��<9�����s�)��Q��Z1@�A�<y�k��Kl���Y?0@Ấ��E�<ydβ�x ���M a�0U*$��h�<'��{	���U&ߜDl�������ڹ[dqO?8��\Qw(L��i`�@�q��{�<�FȒh����r&T
�D3�C�u}�L�1��@��'�T���/��UB�S5��|A�M��R�	G��',1`�J16�B-�*&/�l��6D������W�|��`�JYjlC@1�e�.Z֠�R���!Y3��)D�.�f��d�
4��B��c�T�	���h	~�A�D�� 4!V�řF���Ơ'}���'�J�y�UJ�d2�x�B�r�'"�
���w���SM�%t�(\{�'��eΞmE$���IKeRȠ�B��D���*�pjL��T+WؙQ5'�)��s�m@R���q�z��Y ��?$���6/�Z�t s�B	�!c�隠1ʓ��ۖo�Y�~0c��	B������$X��S��!�$ӭ*�@�C��)D�IB��%=`2ٺb��=��j0��%����O �����#�J�4�Ë[�tQA"O��ô�<0�
ٸw.��d2TU���h��p���3擠�0<�2-���xB�	4(Gf@�GE�yx�D�g�8-�:�!�jNO�M�����l����3G�쬅��`.��WA�,O�9�c�ӇP���F}¢�xJ����Çi|xR2��18�ha4b�=;�4%��G*H��7O�?Oޠ��E�u8>E��xGJ�2��?*ҧh��l��U%K<t䂡#C"y�@��"O��$��@Y�"�B�9"���F�>a��vNdc�,O�	i�CV�,�px�GĸO���Pu�'9PI�VDY�"ᢆ4_8&Y���6?=���n�P<!�%+u��U)�F���1�Im�'�L�C�կK q�����g�����o��Pҗ"O@ĻРK�^">�+t��)���Z����P�wqOQ>i
�!�$��$�A��k�T�؄�3D�Ě"�,M��d�kİi>X+.D�l�B�	�;�x�H$�-`�:D�肶��d��=�'%�0�ujf�-D���C�Uo�S�e�<]hF�Bg�-D��D�O0:�i'D���rK)D�����8hWpxه�M6�����)%D���0-�R���5*��9!�i�r�?D��r�B��lE��Q�';�Q!�n'D�phv��R��e�e�=3tIh�M%D����ŬQ� ��$�["IV]Hw.D�����Y���X��-�JZtp��
-D���$.��(T�K�iv6�; )D����]RlV��
�1�蝈t�%D��8���E0́�FoIf��}�� D��9��Q�yk�d�e�H2l�y���;D��"ƃT�)�0|A`�8[��C��6D��`�FL�1���XAg�8X���"�7D��ZE �S�~�.$�)P�!g�B��ib��rÚ��$�XP*�-LC�I��dC�&Y��A+v�˱Y�$C�ɡ\��	򊉦k����t�ڳl��C�I�Xed`˧/�.	�ܘ���/�B�	_�F��5X���e$��sNC�I��r�Sq�4]��XAlN	L�C�)� �����'Ƚ�!�ը���"OŒW�ӭ7F���A�aB�($"O$�����	��<r�̆'k���f"O�<� ��
b�d$��#Ź@��@�"O愫E�ݤ!oq��!F��"O��R��
<.DA��U*q� 	�"O� �@��T8e$�F=4�$�C"O�mك�\�D���`�T�D�jq"On��D�p2<m:C'ßv�6�("O��	�K�F��(������@�"O LH�Ѱ|�[��P�I~�a�"ODŇ�����K�)`���"O�@����+��	�Æ�no��F"OX!W�Ɲe��ED$l��+"O���� �%s�D٣��J�l`�"O0(²I�o¨�r��ͱ)0�|�U"OށQ�GE���$�	̜f5l�q�"OR� E�O�~��(����3I$<9� "O@01v�æjF*,D�[K㖠�"O���VL���@�"��#�D��"O�l,IFR|܋���x|"���"O����Ίb� ����A% x	"O���MR��B���.�"��d"O��X6�T�.Xpxӭ�i����D"O �����r�B�V��n��eq�"O0l(��*^,
�	��b���`�"OkEIʩq�z�H����p'"O����㐚?����M�,���R"O`E��-�i�vpXק��Q���r"Ox�ӱ���*Bt���\eF�: "O�`�[A��)ã�`n��8�"Ola
��Bj�ȥC"�ųr��Y9"O����H�+Tx�"������'>Q���H��|����V
��`qg:n�F�0�Wk�v�O-��ӯCm��u��5�*���يO���2��
�YF��L�]�Txz�\>�E�'�1`G@��n[36�@Yzâ��q���)�1k�+�%7-��ç5\��C#o�`�׋��\����y�
 ��M8^��
T� ��A��X�|i9�O��
hR��[�J��Y���s����q�O��.�'a����cD(�HhydkA�P�����>�B�!���<5jA_>��P��$1�j�J1*��XY�\رĚdLӏ6?��C�u>��ՏŗAP���c.E8QV����Y�Z�O���"4�����ǋ&H�y0� @�>���hV�|�  >���`F�OeN������"Z�eI�`��vҸ��-O�l��A�ؓOQ>��T�*"nR�{v� 5F�ő#)�Oj�*�U<g
�IQ>ͭ��h��e�O�F�䒿JŎ`+�f]'\G�p��IT]?!f$�4�8���^�V �c�ٹF��M�r/޷$�8�'���&�jӼ!y�'pwn!J�/��*����-B�Z�h���.��?`��A�FK�<%?7�F��MKT���2Z�1R��E�Q�4��Gp�����-��b��覵��iGa�dA�rv~�R�IK�\��D�"�vu wǇ��M�Kp�8��%���S �VT�6#M�_	P݁���J'L�	�Le�d�A�A*;��<JA��I>}s�P�Qt���w�S�-��a)~�� ��3^��u"��#.���S�&����(�6w
6e�փi�qcb��j��m{�@��Mk� Mt>�z�iV}����-��_^ :�F[/W�d����|Ӵ�Z��D��l�� h�� �0�dջ��AG슽	P�vӆ�A�,z6T= �q>�$�wlչPKB�Ef�thdx���M#:hM�I�"ʕa�	O�x��V�^)s~<03�Z/\T��$�G���>!�N-0JFHό�1���
m�<I�C�Kut��Ec�)q~]3CnD�<�"I�:T�����j��ఎ&T���I]�Eb�e�2l��
vC�*z!򄜇}��0@��	�A���c�4c~!��՞tV��@E��\�'-��>m!�$^?p�U�0,K�f=�#l�h!��}�<�2C�G�f�����k��
�!�� ��eH�X-p��E�3 ���h�"OZ��r��!]�i���}t�(2"O�]�vDˤ
�@�`�IIt�<�#"O4�ۣ$�BN��G�2vl��ɵ"O:�" ��w�u��ǚ%XW\���"OX�r֨�Wo.$����+E(�
p"O
���*аߚ���	H<@^~	��"O^@���;�i� ���t"O8(rd�)�&�Q�,m8����"OP��!�T��Aә!x|�"O���CL�(��-SfN��(�E"O�${�B�'t��h���!-����7"O��QS)�J�T�G,�:$�W"O2����M�"/B��%��"�ĩ�'"O��+Ubbx20�ש w��@�"Ob�a��>x���{A�:my���"OX�u��>%�XP&�!el$�2"O�Ph'�1�p4C2���Y��CV"O�-��E�F��j�Μ �Q�G"O�,p0�D�2@pբ�+��B"O��t�NGF^�v��r�����"O6��e#ع
�<J��_�x�<U�"O2Z@iI5tF�H����Mʶ풕"O޵�i�!k��d�$a�i��y�_�<ON�JQ)6M��\�� �>�y��˼D߄�)��C4@���a���yrh	�~��)�C��-B1!��yBHܶXƜ !� �9R���Q�y��<9"`���Ɓ\�0����y��3� b �
.M�	��J�y"�X�i�ƽ�5�^%>'ĩR��-�y����-#�Pp�M�^�n��!B	��y2�J�X"�M��T�L�Ґr��+�y`Y�y�=SA��H�N1(�ʎ6�y���,�r}���.�lR��y�h�
�t�rch֩��	$�y�aݽjjj`cl�+���a�넸�y�È)+��X��\l0懭�y��\(A�rh2��+M%xIb �L��ya�d>q�#�8[#�(�LU��yrOHg��wᗝX5��vD�%�y�M�3&%L���H�&�2IJ��yrA�v��]s���V���H�h��y�O��q����{����镧�y��D"l�j�E�ɣr.&<!��[��yb	wJ����^9mж�@�`D	�y"�ȥHߪ	�w�g��0�ѷ�y� \$��HP' ��	��نc���y�W&z�����E1`,�Rq��y"{�|l��G��.�@��E���G�!�$�%^��	�/	��A�� �!�$�,)>Dҧd÷5�}سƁ=u�!�Z&*��@1��/���$&@�\�!�d��0J>t�5f
�z��	9u�o�!�$ +�vxK�-�t@�O�D\!򤓴i��pC�C^ܘc5NMnJ!�$^�c]α�3@]y��-w�!�D�.s����
� ��Sl�P�!�d�,s�`�t��4	l��z�-Y{�!򤒔fz�ɪ��E�t_puy�!c�!�b,(K$oM=�L䫒�@�)o!��P�)1���'܍s�����*a!�7<tD�A�D�7r���B�0�!�Če�zabt#0��4)�ܧ
	!�� z��tF[>l������"���� "O:��0C�n�re1@��)eI�؁`"O��Ɓ�?)��P���4��"Ox���T
@��88���GT]y�"O�@j4��%l�4���C-=�<�#"O����ŶZ
���q�����	4"O�j�g�]r�dK��ׯlX�x"O�HS��2+>X��b�̩{<j�K�"OB��L��J�9%��+pYh�"O�	��P]�i��݃I��a�"ORy�[�"\L�e��EBc7"O$@6�J-'�Tɗ�K�8T�"O�E�3 IR@.�B�n�.J�T�d"O��A���#yc�0CoI�I�y�v"O^��Z�T઱����$"O 9X���7k�9C�P�P�F"O�Yр�JN���C�� ��"O�\���i_(if��E���:S"O�DS3!S"+)&D�aMX�Z�Dňs"O�0Q��/^���a�lI%"O���R!A-iP��%V�&�H\�"O6���f�IuY�����U�*a�v"O��r��d��i�7n��p�
�8"O^$��D��#�X��L֬��"O$�`�V�pJPp��1����"OF��NN=�&haf���>��"OΙ�QHJ;�6}:��d2lT�"O��*V������7B3�"O1%��:��� S܂E��9w"O�yB���yj%y�oF��@��"OD�I`ܒM���fa\;X)�|x�"O�b �����N�S���#�"O���3̙�M���j#��3�B"O����'Z�[��7��!�`Z%"OZ �,�1,���U��\�21	�"OH�â�TT̍���ʤu�`���"O���ㅞ8F!�1ȤE�^>��0""O��D�H.�Q�
�-A����"O���7LOm�4�V�U0@�Y�"O��4!�;ԶjC�Ax��Qr"O�ta@ �R�ti"�J��u�"O��A(�
_�n��	�{�:��E"O^�"c�<;�{3S��UIu"O�հ"K�tn�`c�ذ{���8�"O����\�*�&G�T�.8\"P"O�%��H�"5 ��DKř�ĉ�@"O
1����t\H�**rF��SR"O���Ё��A�h����6Tr��3"O�p�B��uQ����`ȃ[μ�b"O�xS��@3�f���%�f� }h�"Oj�b$/�!���DT�l�"O�J醃w�(���D<��80�"O|�bRf�{b���3�E ��8""O�00��6=�Ĺ��*�r�
�"O��S�k]�&<���͐K�R �"O���LD�WY�� d�ey~���"O� A��Q�{ �\�2�T�[y��{u"O`���U)"/|��0M�&FN�HH�"O����')�]@�	Լd����"OJ��)O���=�!�4�F���"O$�3�,ۘ&dڜ�֫[���Ļ�"O ��Y�N��� S� +���"O�	�j��a���`��S�C�2�y3"O��Jb� &S����'�<��p��"O� T\pBf	�bN��x�ȭM����"O�}Ҥ瑜�RH��+@I�ru��"OLE��hW+�����S���"O��#l��IB�T↢z�0��"O�i��#˜@��c��K
Vr�|J"OJ�a�e��*]�8P)�:Wd�X��"O��A4ď�I^@���~A�`2�"O�	
E�\Vv�$�V���f.B@C�"O,m��B.S?6{ㅓ%"�\s�"O�p��ʏ�k�q[�B�dH d��"O0���9Z9&��wCJ:=RvM""O$�A�>jr��bu,�y[�"OR���
u��8�J�)��*g"O����z[JI �!X�B���r"Op
�fT�j���� 3o\N�Jt"O���0''8�<��&�+kU�0[7"O���to�J����&�HRx "O(�S��8^TjҥB��`+R"O�,���8z�ވ�QE͏Px>�rB"O�t��NaVt��MWϖ@�"Oȸ	��1:�0@s&����d�"O��* ��S�P%Jx$Iz"O�� �z�J��	�Tw8p+�"O0����M%��k��ͨ?X"��"O�ģ��Ք/g0�� @�M_��[r"O�$��'fb��nF�O$�%X�"O���p�ZP Ss��P��#R"O�����a��pᄬѣ#�ؠq"OĜp��Ih�"eK��=�BL�g"O��D	��=��Iz�e��"O���F �z`����Z#_l\�V"O����w����_2�n4Z2"O�Ȋrݠ)(�������1��a0"Ob0�K8JA��ƪ�p� "OV)�3��*̡֨#�5�@P"O6Q�c�ݨE�P˳�Ѕ,��0"OnXX��ǉF5v<맍Q"<��tys"O�qIBC������r�гjJ�9��"O�9� *��%,W�2He�a"OH!	�� �D�P��:���"Of ۴
@�H;����i�?@�T��"O�B�K�"�R��Q 9$���"Oܡ�"T&f�,X�dn�q��d��"O����o�`�K��c��!C�"O��F%"y�1�5i�c�64��"O
�A��`�>�!r�JKv�df"O8�W�A��H岳�1.]v�	s"O�Y�m�?@��%�].6��H�"O�D���Ƹ)�V���&�}�"O����_�"��X6�?QbQ��"O,HH�����i;�Y=(�:�c"Ob�� ]);�8H#4� �RQ��
0"O��RQ@���͈���'?.mH�"O�Y�cF�>�>|*�j�
G̮Tp"O�a�.? ̎��'_�]�"�@#"O������lhPeg�_��۷"O<�;�ΰ;���"��"��@"O6L�B��a����ǩgǈ��"O���n�� Q�	
(��b""O��D�ګ�v�x��R�n�fA�`"O$X�   ��   �  8  �  �  �)  5  �@  
L  �W  �_  g  "q  ew  �}  ��  >�  ��  і  3�  ��  �  Y�  ��  ��  O�  ��  ��  �  ��  ]�  ��  ��  ��  �  h 2 � @ �# �) $-  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(�"Ov�M�{�Ҵ�U���F�T��"O� ��M�g��l�a��8{�Y*7"O�Z��іh��8`�tm�`�"O&ESS��M�,ɠ��b��b$"O,y0GD�!�<�Y#dYF��c0O��=E��Xj�z9��&�
W��b����yR��tR�D��A�(�,5�4�1�yR+��9�s�B��LsӬ���yb�Q�j���s6$���w��y"��#}�i�hK*?2�X����y��
�+U�y�VI�����y�kS}�Mh��+F<�M��F���$9�S�O>(nR�xЄ)0�"ǈ^f^���'�$+uP�+���Ũ�\k:��'M� �7���.�di��. W�0���'!|�QB�9K�Tj�F".�0��� ~}��.ު��S,	�Q >A���'ў ��̗+Y�*�yf���c5D��ˡ�ΩI/�Iy�e�b{����=?���)�'6P���B"e�rE�g��3"��Ɠ��a�U�^�[��%F��2oy�Tc�'�d���ᅝ#�fЈA�?��a����	}�-+IҰ���؉$NVA�� B�[�B䉉~]2(��^�"s��LL�"<q���?Ms�@,X��#p#A p�4Tx�(9�OZL+۴S��p����n	p�b�` 8���)��<i⦓c����	�9Q�:l�i8�4hg�	�i��C%���e8���@ɆZ�"C��x���I���=Y�$�[��'�ў�?i2(�hd� ��k�6"�H�(�H)D���c%�)�0�;��¦Q�P���f'��y���p��F??!��B�J��$%��+� �E�O��0�b^=.���d�(�(O?Ab��+><󳢝� ��j�t�<�7!2���X�	'WEx��S#�o�D=�O� (�Έ�b ���N'G��j%�IA��	�oQ�$r��X�R���"1D���:}��	r�U3�>� 
.D�8:ƫOO�)X5c�;v*�*�c,D��0!�V
A���j�Qz�&D���i����]�U�A�K��T��%2D���q�ϷHjx�UD��}��E0D��g�G�x�pD�R�PL��za+D��c�\����4���1y���3�4D��u)SB��	J� �n����3D�����y$Ԡ;�]�e�2D�(I�%.E�H�
�ȐYXz%��<D��@7��mA�aS4 ��U{�6D���6MJ�I� 9�C��(+��R��!D�2����dic+I"�vtKԆ D��㑼q���dG�	=P4a D��(�ɑ2ZE0��FPf�0��!D�ZS�8�
���S�T`^E�խ!D���C�X8�y�rGR=^�:1�C"D�lB�ǘ��Ba��d�E��Db?D�8�#&�'iT&;#$	@]��ؓ�>D��j�W�9����K0�c��<D�$z��N�<�D�R+�� ��W�;D�0��������"��1�K��%D�8����I���DJ�{Ƞ�.D����ę}� �;�L[�-q�h�0�+D���$`
�j���*SNK�
�p:�#(D�P���^��h�Q��[�����!2D�{b�]�0�<�j3���.�(�B�2D�@Juj�dk0l�$ӱ{a�t��;D��1��Kk����Zx|3@�9D�@�E��/�(���Ϡ3������#D�<� ��4�t0 aNQ
RX���$D����ܯS΀�1.ћMҌ%��#D���&�x� ʅ��3#phu�C"D�$"70'0B�{2�N��Z��P(!D��Sf��jXZ����k��H��?D��!�X f�U�c��(ٜ ��2D��(4�A�-�R�c��HCQp���/,D�4����V�L4�$"�m*�'D���0�\g-�D�nɂp@��31F(D�4�6	L�a�R�&D�W���VB�I�4�D=z��B�w%��h�:�DB�I�U�(m�`�ǃk� �� ,+B�IC�:Qr`)�;{�����]C�C�)� �Q��tY��3����x����v"OP �� 3GTdIX���7L�(y��"O�X*0��K|((і�P0C�0u�6"O���GĺCN<���a�`0�"O�b���;\�h[A56{ڙ��'���'d��'��'R��'q"�'���m�r�P"nR�RucP�'���'��'�2�'�B�'"��'��a���ü4Q��#M�g����v�'�b�'��'@2�'=��'���'���a!J����]2���_ˌ���'���'ar�'f��'���'��'�	c �;Hآ�J7�ŤmK���t�'��'�R�'h2�'���'Z��'�)r&	_�B��P�c�C$%& x
��'���'�2�'���'���'R�'�<�3���0\6��I�)����'���'���'��'R��'"�'��q�c�B������M�0�N��?����?����?��?���?����?�&��kuʁ�&��Ja�DJ�.N��?A���?q��?!���?q���?���?1��;�x�Ȃ1W�R��У�?A��?����?����?i��?���?1��(-��1���I#�{2AH2�?y���?A��?���?���?)��?	#��U|�Ѱm�!ZP�"�I-�?����?����?)���?a��?q��?�Մҥ7,)��*�Тg
ɝf.�l�	ğ��ğ��	ǟT�	П\�ش�?��i���I��ԫGG��aVa^'�9�E[��	Ey���OMoZ�[����s`U!J$�yr���F�*�I??��ie�O�9O��D��$���{㬖�\��t��쀤~�����OzC&km�X�������ONp�bH�Y!p��c�\NEb�y��'��a�O�6��*��w��$�N`���hu��� �7�S�M�;-dؒ��;1���ŧa�������?��'��)���@]o�<��gQ9W d�a��@�ЖB��<�'����@��hO���O8�+�/4
�)��߲:T8x�6O�˓��v��VE��'t(�#���ް�����l^�C�d�d}�'��6O"��r�b�/K��y���,4���'<2��h}��y��4�R���yb�'���gE +|�����0dQ����^���'P��9O
a�i��p�����"���*2<OimV�v�Pț&�4���Ȇ��n�Q��F!|���� ;OJ���OB�$�~ˈ7�7?i�O�>�	6~{t Z�����0���.�p��O>)-O�i�OB���O����O 0�-3):�[Cg %��(�ͣ<a�i#�8��U����F���ܵ�2h�%��$#%�N�ҀZ���	��%�b>��% Ҏ310mX�C� q�|��"	(��l�~��ˀh&���䓍��>�2��M�C@����KG8}DR��O����O$�4���֛殃�"�r�k���Q��4@�a�@i�yBCiӄ�DЪO&���O��ğ���ı/Q#:�PT`�M>BJ	���k�.�6��7&�'����.R~\��A({���!e[�<)��?i��?����?ɏ���_V�!jdW�N�2������_���'J�(eӄ���;���d�&���rmH5G�ZH���e��d��	n��۟d�i>�H��٦M�'��\��S ,y�HS	*��J`�2M�X`�����$�O����O���ːsm`���"0A�L��b�12����O �Y��@06��Iҟ$�O����%��JK��0t��_���`�O���'W�'Zɧ�� s_�|��I�2��9�d��F������	��(C�M�<�'sy*�D����#����#Po��!sN��6rȠ���?Q��?�S�'��Ď��a�Ckܣa���{�!ȫIA`�#M&c��-����ܴ��'�&��?�R�R�l�vMP��II�f0� 䗄�?��}v�Iܴ�����M�m�r0�*O��{���aP|b���R�>H�Q=O&ʓ�?��?a��?������0Wo]YR�
5�B���(�	�l�o&K>h��	�T��a�s��#���{���/@���ب_k���	б�?!����S�'P�����4�yb���lN�a��1P�.X1��2�y�$`���������Ol��T-o�.Q:q�ʑD�`��f� ���O���O��{���OW#A�b�'�B�l̨������5�����X;�OJ��'���'��'�Pq0rEDJ&h�GH�:dDm��ON�@�o�-u{�6�'�S[����O��z'��IE�|yl�$h8Ij0��O����O$�$�O��}*��t�1�4�w��$���x�Dq ��Qӛ��D�"�'��7�4�i�Y���[��n����*640��V@g����ٟ��	&	� on~Zwn0��&�O&��3Q@�4r6-��@J �&ݢ��m��ayr�'���'�"�'��,ި~�~8�5D�$�@Ǔ�0�� �MS��N��?���?�M~���I؂\ز��ozI�H��u�Ι��\���Iʟ�'�b>A����*}.$P[��ɭ� �w�-Q���nZ��$мK�J�g?�N>-OT�J� /=x��ՁD�h�8d�'�n6�T!P7�D�Oը���/&���S�)&��Tɦ�?	TS�t��ןD�	�-ܤ�`�.�8�DD �>&�*h#P�צY�'�����"��?��������� ����l&����\'C�^�KB6O�����'��
pE�[�P=@' ׋Av@���OH�D�Ϧ�yg�.jпi��'�����"K�`���)p�@i�|��'��O� D�i��	+}���T�Q�&( x��oPY6��qB��	@���"��<����?!���?�q��9W{�@*�����%���?����$��5#�����	ɟЖO���)WfH L��\j�IF.T2�I��O���'���'aɧ��V[c^��b�X�b�1%j�>J�l07F�2T������ӔP`�L�	q��d��N���a �jiDy�	��������)�kyR@z��9����\	���,֮U����w��2@��$�O2�nZv�^��IϟAR��
�F@6S�~��%	�;,��$�O|���s���Ӻ�¶��%	�<��BS��$��AE*<"�L��<�(O�D�O����O���O��'+F����eة���!S#�8c�i�~`2��'9��'^�O;2hf���^�JH*a	1�Qq+��`�J'=�l���O
�O1����en�^��%v�|H3B�"NI~Ak"��V�P片4����'(�<$����t�'\�Ñ�%(ᘴH2��0a��x1�'�'2T����4h-� A��?��y `s@F	N�@DHRa��X<b��B��>q��?	J>��ؖL�JY1r���zN�<v�	]~r���r��O��	�	TҬߤ��%�T�}	*Ar&L�y2���!���w-��!dF�1�c
S�r!mӎ�$�Ox�ĜŦA�?�;<�|�p��?$�\�P��B-����?A��y2J �M[�O�I'���~R����O�!(DT KG�?PUʅ�M>a/Oh���O����On���O<���CR�R@�|rA��a�N}�g�<��is`�;7�'��'b�O	�B�dT]:��I!E켱���
]	d꓌?a���S�'��Ѓ�3�8d �6{>lpRK+>��Mp)O��`�iǌ�?7�,�ħ<�T��z��A7�ÉN����k���?1���?����?�'������l��ti�
�y�n��U�H�k��P;f�ן��4��'_���?���?�4/Ǹ7��A�#�xh�Yi3k�=I�����4���ͬd����'9a ��"���^��$����<���7d��~2�'L��'���'����j3�a�G�G4T�@�Q,��d�Of�D����s�A{>%�I��M�L>9�E��"@�ьi��Dc�h�n̓�?a,O�� }Ө�C[�!���~��!��		w�JP�J,����������O@�D�O��$��i�aWAR�=,X<BF+�(4���Ol�4[��4AR�' �U>}P����:�0�C�ƒ��@g)?3P����ןh$��'}mڷ/�
up~����5�~�7A�&FcP}޴�i>q��O��O���5	�,�DߵE���;��O���O0���O1�X�nC��啳o�y:"]�R�)�7��8�-��'"�Gxӎ�d��O0���9Nl��FL[�t�J�q�N�09��Xq, s�4��^�wĠ}b��u�d�p��)�
�'Zۦ(�����JJ����O��d�O`���O�Ļ|�ď��d��E�����^@2��Ư���<H��Iß`���y�B>|�����@J@Y*��O7Y,��'ɧ�O/v(g�i��dVU`ęs�L%o��`e����$F�.��P��''�'k�i>�	�{�Z�� c��F��A�ަ$��I̟��ǟ��' @6M�kd6���O�睅}�|Ǭ[&Ws�q�dY�Z��⟸k�O����O��O�\���YY�6u�%Apd�����d�dH8d�~t����D�S<e�"�֟��n�.� ��-ʦ�J�CaX��|�I͟��	㟜G�d�'��<Qပ���{�BY':j�}ye�'(n6�G�b.X�d�O\�mZH�Ӽ�@�?g��k`F��=������<q���?��q�\��ڴ����K� ����c��%~���!7��n3$���Ư�����Ov�d�O<���OF��I�R�<Ȃ!-��d��A�()R��`R��IًF�"�'ҟ��'��%�➞
��(�UA�M�*��j�>����?�L>�|� i�2<UZ��F"z5�er���d2��R�9��	4*��E���V䢒O�˓#��m1Fm΃u3>��	Q
��L���?1��?���|�,Ov�nZB9��	.">�(��4;�$��d��o�l��ɂ�M��⢨>Y���?��B�P ��[�Yd!`���x��b�B�M3�O>|`�������w-F��cB!^>L���8J��''��'�"�'6"�'E��"ga	�I���to�*H�P�%�O��$�OVln�@���ӟd��4��z�x��3RT�j@a�v��ճO>i��?ͧH����ٴ����F��u�rj@�	0����d�<kP�d� �����O����O�̅m�FXB*��|�ڝ����Ӝ�$�O&ʓ���G�7J�R�'��S>5P�/�!o�:���K=^"����6?Q@Z���I�8&��gs�@g��=
L��->�Qr6gL .�℩�4��4�����'��'|&	�SAP�4��닱��Ux��'E��'�����O��I��M3#˜5����(ߵt�(EA,s�z�H���?�i��O���'f�S;�p��!%
gz*�� �F�|���'��؈��iq�	+[jt��O&�g�? �iP�i�l(!E-k���P>Oʓ�?����?I���?I���_�P�w�
�+����eO�)ɚ�l*#��E�I����}�S�|���{!;94�t	2��;Ab2�&ͧ�?�����Ş��d@�4�yM�t'�!A�k'��ۇ�ӧ�yb�4���������O
�d
�&�jA�7� yFX)���_9����OL�$�O�˓h`��c��#���'mЁ#8ҵE�$�B �f�:k��Of��'���'��'-X! �b��U	'Hq��4��O8+�4�
m9P�S�?iP��O�4 �LS'wc�=[XA|%�)G��'�B�'k��ߟ��&��5m�V�b�)�.WR	��MCܟ�S�4��i���?���i��O�nR�3�2�3�ON; ZV�n��M�$�Od���O����tӜ�����3��ڤJqH_4�qےl� �4Ja��%����4����O��D�O��ʈl:�P�C2N%�W�>�~�kV����4������?���䧱?��ǖn��u�@�Z�(D:sIW�;o���D��[�)�ӆQ�8 ��&�G��\��	
��|Ci�ݦ��'&(T�S-�d?yK>�.O��Ĺ�P��T:;�X!�G
X� ���O�D�O��4�:˓f�,ݥ]��lJ�Y��u�P��Bt���],�rӠ㟈C�Oh�$�O�Η0F��ۖ!�Idd�('��fia�#w���9���R�矢e�I~���t��'*6u ��h��˒g�^�Γ�?y���?Q���?����O2Z���GX�f/�V̬,ڶ�҆�Ly2�'��6mQ2b���OLm�`�-b(M�a�?@ 8)$�I%<�*�&�8�I՟�S�m�Y~B�XJ��)�!� J��֢Ǌ'N�R%������|Y��Sܟ@�I�p��T�	�а�B���Ys�Y�EJ������wyr"p�-�B��O����O8ʧ��@�|����O�Ո�(<?�0[�T�Iҟ�%��{���N��6�RGEΖ=D�� E
l�R�
ٴ��4��UR�'��'�b�eD;Hĸ�5gK�'�Ԋ��'s�'"�O%�	��M�@�U+3w�!T��uQx@��L�1uV��"���?�i��O�E�'�� B�TP���Ra�YH���Yn��'TB�zղi�I>�h����O�'�6lq���
�J��ϔUmNe���-|O�cG$�-<��p�뀨&�h�1������ �ԟ����<�r���y7# � -��LSp���w�\S"�'�ɧ�O�l�1�iE�2*d`ؚSc<�x�C#��.�$��5��c�'��'��	埔��0;N8���=�2�2@oN4#�����������'�d7m�O��˓�?)��D1`�)�膤G��@���'� ��?)����3U���a�ܩ�r��F�ݜz�-�'�5"���#�0�c��d��⟠ca�'�V�H��M�OM6��e���~�`���'��'{��'��>Q��$G��I�Ĥ�7'Kx1�4��"_�"|�i56����$�Olyn�X�Ӽ���P���$kD�rf)`�ˈ�<	��?i���v� ܴ����Y
F���k�t��T`R�%�f��j_=v�Y�o'��<ͧ�?���?Q����oT�E�$�d�,I����F� ��$�ߦ)�������	���'?��	��H؊@���m�&���lK�p�ۨOT�$4�)�Ӟ��@��B�*���cw��<`�<h�ԛ8(��'�-�0៴(ט|]��	�/YpPis���
��ES���џ��I��L�����SVy"�d�|\�f��O�sW K5Je航qHB�b�z|� �O�o_��)������I������_�8���Y mS���Fُ.m�~~�"Pe-,�E�D�w���WL\'���K��%a�0� �'�2�'�b�'�b�'���x�%略%0x3`k 1&�^%Q� �OT���Op�o�D��'-�7M&�DT�+W�k�K�	���0I R�@�O��D�O�	�8@�F6M3?���|�ѡY�l�s��!A\.9�@I���'�L�'�R�'���'���!6^\Q捛�֜��G�蟰�IRy�ab�<�h4�O����O@ʧUƔZEAQM=� ��L�8i���'�Z��?Y����S���_�b��G@I/S��b�
��3O�+�	�cF��
�\��"{�+�a�G�")C�� @\���׈a�T,�	����	����)��pyr�w�@������[,�|2�HP4>��GD�W�d�OVoy�G��	�$�k�QJ ���:0I�lV��I�a�T}l�~�C�@*8p��E�I 'ˮ�Y#N��m�����üaR�<����?���?���?�*�<��+�#7%H)H��ˋ�M+�,��?����?�H~Γ9��wc2]�%˜=��C�O�0\2�-[7�'���|��4�[ wv��8O�)Bn[�
=�����~��!�F=O�u��#���~"�|rW��Sџ���[}���@.Ӗ��A�ʖ��X�IԟP�IXyrFy��d��)�O����O��Q'-4 �����H�o�֩Y�(=��3��$�OD�-��
/�5 ū�4�-��D�9�	�i��5�&�����H~�tͤ�X��7I��1ˢ=Ƭ="r/�4
s���	��4���P��U�Ot�猐tm�L�hĊ.�L�˳lV�#w��l�҅���O����ݦq�?�;2n�DI�"�gB�*gϜU��E͓�?q���?!&��M��O���1��1��� ԭ��]��ZY���ƃqh���c4���<���?����?I��?��ށ��.C&Z� �$e����ѐ��䟤�����&?�� Z6�Q���G�)�T(`��?�"�O��D�O�O1����ʙ�������E����-�"�9�����C��Z8���r�Ipy�@�!fp����ѐ��L��N�;Z;��'2�'��OA剨�M�Y��?q��9�x�R��V�-��Y����?1Ѹii�Ot�'���'O��/���*�I�L�����1�����i��?��hjt�O�ʘ'?)��� 5h@��7)Q�JX�f������D�I���������IN�'�.%�����٘��Òx�fis���?���#�,�����C�%��'�R�~�b�#��:nm\d
�(=��ڟd�'۪P�i�	�p4*��V�H�D����K�6$ �̚j��H�j�\y��'���'!�+�?*�,�hШ�9"��H�ǀ�7f��'��I�M�wEW��?Y��?A(�<��U�肬�p��-<��%j���٩OF��<�)bg��>�Z%�1����RI2Ä�vv��1�j�4=�R�+O�	�*�?aQH'�DX�]��Ū4Q,L,͂֨�(r[2�d�O����'N���\�̫�4)�j�J��9f.$�c.�eO ��N��?��)�����y}b�'|���� ġ;���$?R�H�[�$x�\����'Bĺsn��?�c�Q�Q��-��5kAG�#��!H�ov�ؕ'	��'br�'���'(�1�p�Ӈ(�0 ��L���"T�ܓش'�����?9����'�?qC��yGfՍO�LU�c���\ �@Bg�%G��'�ɧ�OeD�P��i��D��r��h���Hj0sm�;El���~Vݪ�6�D�O^��|��Q��K`h�$*a���C�����?y���?i+O6�n�$�U��ڟ����2pt�\���K
Z	�e�)�	"���O��|$�U�Smy*��[,lo�8�0:?�T��!)���ܭ��'+��d�-�?	6㟿4�p�z���6�깃��&�?���?����?���I�OM�CN�C�$�:�n�/pqI�O��n��=����I���ش���y�<i,.��ELߑ#�p�����y��'DR�'K��rT�i��	5\�i��ҟ�,c��A�2�Ȕq[h�"W�>�'Z�	ğ8����l�	��D���%���М6�%�"�_�5�h�'B.6-XW����O��.���O�8�v����L2a�×
�x(c�W}b�'~B�|��hZ��Ji����>LTs��I#�։�!���A�6F"�;��O(˓Y����Շ��N�HX�ɁNKp�8���?)��?!��|,Oνn�}�F���;+l��ђŉ >�
��cb�@�.����M[��G�>Q��?ͻ"�.]��
ͭSEv�� ч�\���K���M��Ov��g*�?�s�=�	��:���DD^��L�kŏ!�L�R7OF��DJqm���W�V��Q�K*fk����O�����5˰N-�C�i��' �TӣF��o� aĂ˼V�z��!�|��'K�O��)Ƿi��i�=��-�3	����CmǓ1�L8
��F!���;��'��	矬��ǟH�I;\�\��M=9���RF�VM�H�Iߟ4�'V87M�/��d�OJ�$�|�B-G<�|�����!"r��Tc�@~�i�>����?�I>�O�\qEjV�KTnÕ�Y6�6d��h�Wɖ�3d�Ʋ��4��)���`�p�Ofܣ�*ss�x�&A[(Z/�QW�������0�	�b>U�'�7mL�dqu
�r��(��Gغ+`>��D�O�����!�?��\���� tm6�`��ؾ�a�Ͻ(�����Ο(�	��m�uw�
��ď�oy�iL)N� *�m�o���S�ژ�y^���	��x�I�d����L�O
��)�kD9e��H:C׿D[��:��xӐ�H�l�O����O�?������F 
��@!iZ�S�J]Ql��?����S�'p}X�ݴ�yb�J�~Ԩdh���
�n�����yb�J�V����	�q[�'��i>��	6"^� C�i��?,Lъ�G�"��	�T�	�� �'�07��������O��$�(Fsh����h�ySc�T�4���O����Ol�O�l03�Γi�=z�g�c20zG�� zTOO(Bj0aTnZI�-C�n۟�k6)֑B����͎�B��2��\�Iퟬ�I���F���'�"��� C>m���:s���'8���';R6W�ef����Ohn�O�Ӽˆ�U;H����S
_z�3�e�<���?���1֚�y�4��ߗv�q���RU p��o�Z����#B��0莚Q�0�(����N�@P�ͷ�������t�v�)���)��K�ꉔM�x��\�+w�XA����7�}�T��PN�0��
f`���'�F��N�Gb��;��V�^ ]��*��?��-�4G�8$�@E
���b�zx��ٙUG�Y�3�S�J<p�Aw)��#�.d����C~�K%D�"AiQhM9w�0Xwf��^V|���@��������oS��
�F �68L��kJ7k�;c��)^ ��+&ߪ�| �wfЦ�p��F����4�?����?��'^���ZB�
҈�5��㆘�o����4�?���WEp)���iX%x��5#�?pG��ʂ,+t���2k`6��O����O��i�L}�U�[���=؈}�#mQ,#f�HqE���M{W�(�?)O>�����'3�T��FTD�9�g�<��䪱�a�F���O��Ė�O4F0�'���͟ ����-����e_��u��1�H-�>	�S����?����?ٷ� 9@qŒ�����є%�0�i)@O=A}R���$�O��Ok,T7A��)�� T�}Z5�qa(;���6��'���	Ο�	Oy��ԥV�T���l�����K�-h��b�#�>�,O��#���O
��\�_|����-� ��ģ����u y���)���O4���O0˓fIz�A�=������}�{'.��\���is�۟�$����۟1�N?Q��B����G�4~m�����TE}��'uB�'��Ife�����D���1�Jt�aܩ��-���g��l�'��I�d��sܓSzx�P%$$Ĳ��J�B˄4m�ş8��Dy��E 	պ맋?�����͈b°5Pl�+hK:�Q��Q�L�'���'P�1��ġ?�b#!��eW����4Ezl)$�z�&�$�����i�r�'V�O1z���cG�6֤�"���1���Hg��m����  5��ޟt'�|�}
ѧN�LN�Q1v�;ia�%�Ea��53�뉙�MK���?����rEU�8�'D�Q�'��%��s!eY����tӠ�[�#$�IX���?�BgC���{P�#2��`������&�'R�'$��:γ>q(OJ�D��0٦cL�^м��3�Q�3�`�2Dp�v�O���" (�D�O��$�OkLZ�2�`qB N�/��@D כF�'����Ҏ%�4� ��=������4i�. �.-kƢw'T8�x�'��I埼�I���'L��c�"1+X$��]��:,��(�/� O����O��O��Ӻc�c!����ʍ3f���#�ꦵ��uyR�'r�'��ɗ$G�K�O+��Cac��:� �#�!O���O*���O��O(��|
�g(Fax$�P1?,슦�#��AW�x��'��<�vFt�$�'�$�cq#�A� �QEeR��[i���D��]y����ē}L�I�e�*��@*`F��d4o�ğ̗'���ǥ&]�؟����?ט#b�|�X���"DR�!��AϜB�O����<��m��uwfD�_eD@��e
& XS /	���$z��S`�O�d�O�����Ӻ��ֺ/��H����"bľ�CѦ��	[y��O�Oh:��Ј��i)�F�tt�����`by��ğ���˟���GyʟvͰ6I^�^R0$jZ/3y�@[S�_r}b�_��O1���DV�f��5[Ď lfX�Z�iE�Bh>�n柴��˟�c�+ͽ���|���?�Ԭ��/�X����D'I����\��F�'��S�Pڬ�<˧�?��'6�E�'b��@R2OñQv�9��4�?q1�
��]����?t"�������ZC�"B9�L%�HB�9?q���?�������-O����P�aO�7���i�f^2N��'����쟜�I@y"�'����	8�(u�����$��҅ߒ~���'�՟��Ih�'��SR�`>e`��
�r����S*
���6b�>����?�N>�-O���O�T�S̛�
�#���d��q��s}��'\��'��I3+&F����l�$�,L��qc�	\�����:�Qm�џ��'�"�'F�I��y�Y>7�\��:v��mh��p��3WS���'��]�|��\���I�O�������V-_F�Y��T).h��S}r�'�R�'����'p�s����A�@��]�޴�Dɓ���l�CyR���z�6��O���Oj�)�S}Zw���2�`fl��Q/����4�?���F,�LΓ��̸OW$�Ç�_8�x�SdF�z�N�k�4.	��c4�i���'���Ot����>I5VQ�o�9C�����f_t�z�lZ�F5��	ܟ�'���$�kLPS�OW�3��#��B<Al�˟������!Ad����D�<q���~2(ʻk�A�l Jv��4�-�Mc����DA�qi�?���֟P���RT�r���~��$��.T�9�j���4�?!M�x���myR�'����X7Y����M(Y�*=DΗ�Y�l�_X"��<a��?�����")�Z �T�{J�1��T�5G�i���a}�W���IKy��'�"�'���P��٥HZ��f
=J�P�ą��y��'n2�'u��'� /y��j�O�dКSH
2X�hI`!D��1����4��d�O:ʓ�?I���n�	��扯9>���/�4�� �'��XV��4�?Q��?1���&x����O�Zc*�Q��ϝ�7f�\Xp�� N6�k޴�?)-O�d�O��$]�?m��|n�$����b͛x��=9qn��b�h7��O.�d�<Q��3���柘���?y��'�3q��r ��l��]H������d�O����O�\��'��s���'>�.1v(E/�2�����/T�l�Ey��#/��6M�O<��O���\}ZwC�D�ubZ�O_�%& 94�1�4�?��<�(�����OR�����=@�J��ՐU����4F�TԻ1�i���'�B�O� 듡򤈰R���{��/��
�D#O�mv	f"<1����'n�=�7�V8����I�:v^���nlӬ���O4�����*��'��I���1K6X�1,W>K3 PQ�H�!��	mZƟ��'�����	�O���O4X�"��%?@�a¢��[��X8���Φ��	Z6x��O
ʓ�?i.O���X�����0)c�K�d���H�~}b��yb�'{��'R�'��I�fK�#��%*���0J�2�����!����$�<������O��O�]����
sv8�5��4x�huarO�JT�D�O��d�Ot�D�Of�q2���=�� Vh tG��`�R`���z�͂�i���ڟ��'���'j+��y���:d�ݹ�E$�V���ڨ?Ē��?���?).O��)��j���'��[��K�nb�(Jw� !$:���%x�\�$�<����?y��'���Γ��i�T����&<h��c��ڨ��c�����O�˓U0���Y?��I���)N�:h1tH¯Jǎx!׆�2��4�O|���O��D�J*�D7�ĩ?� �ôR�L;�B\'D�sG�~�ʓl�h<I�iR��'��OQD�Ӻ{&�ܫ?-�Řd��5{�N�3j�����	��Dzc�u��&�|�}�`.\	Mf�C"h��{� q�alI�-w����M3���?Q����_�@�'�"����J�9�D�Z���8T�i'x�fE#�6O����<����'����q�<�(�0?p��)��tӬ���O���6��'��I�����	P��"��@��"�K1Ϝ��>�!�f��?I��?I%+x�Nȉ��װ-5�d�U��?-��'���6ʦ>�*O���<���a 
���Z���2p�k�~}b�����O����O6�$�<��W�a��`��C�48�wG��7���Y�x�'�R�|�	��<�	>;�4<�gDގ,���QbaV4]�@ZP/n����ޟ��I�����Oy���/x擟Tn\yR@M�/5�ucF�,V6ͬ<������O ���O�`I�6Ok���h����Vf(ѳJÝq�<��۴�?A���?����$[�2D��O����9��p�qf��_�.�"6H�6��O���?I��?��Ǒ�<9/���!Ȯt0j�2���}b4 UK��M���?)O�`� d�z���'b�O��m�� x�-!@
�<�ܑ��'�>����?���|��)���9O���;1g�Ź���B6��!�؁k�6ͬ<9/V�Ǜ��'n��'o�t��>�;�<1���:S�|�9%��0O��9m����	�Y�	>����Oz�>�j M=2��U��m0C=lZ'Kd�FxU���1�I͟����?�j�Oz�u��\�7QL��yU ���iH,�'�RR� �:�7٬pslܘ}�MW�. P�0)��iQ��'�����&�0O��$�OX�If
8YuD�3��qآ*�HE6m!���9��?=���4���{�p�Sʆ�	�*�s�,�}ش�?����Of�$ ��Ʋф��#C�&6�Ͼa0z�H�>��%�<�(O>���O��D�<VE�7s��=��B"`�PY�`�2��y����O�O���O,=�b�,C�\���^�0T����G�%e�D�<y���?����D��]{�y�'2����U!e>����&'���'���'��'���'�i��'Z��С��
�*�����<��'�>9���?�����DӼf�D�%>y�Vc[$Z2����͂1S8 a5G�,�M������?��sVU̓����h��a��UJ�2�`Պ[$7��O�d�<a�K�#��OB�O�h�3��
cs�U�pG

�AY%c2���O����0 ��D.�d�?���F�XJa��C�Є`o�v�"b,y���i��ꧬ?���'h��	 r����]��h��@�7m�O��
����5��2I���8�mՠEg��s��C�$7��>&�n�ҟ`�I埐�ӿ���?)T�\�w���"
#���D@O.L�&���r�|����O|ݓB�� ]��!���*��K��I"���'���'C���&$��OD�D���+�gyB@L�a�TH��X;)�06�/�DXSI�a$>!�I㟼���8��b�B+�&;.�â�æu�	�6ǲɌ}�'Pɧ5&
\4T�$��4L�0�11��D��L���<���?A����$\�'��@��W�_�D�i�%�]���2��L��?1O>A���?!DKWi�r-�G��vl���
�o�z-͓��D�O6���O���x$��9�����n�kD�qt&��	���˴�x��'�'���'J&$��'1��a#��Q)eV��-���>I��?����@�$r�&>�H1)P�r$����87$p�պ�MC�����O��$�O�A��?O��'��qZå�X�e�&Q���ʦ�i���'��ɃM���AK|�����1�켣r(O�[N�kG��:|l���>!/O���*�i����^���y��15U��|�˓fE�qT�i����?i�'3���=n6����5T��C*_0g`������OJ�� ���3o|�F�%~���d�iIЁY �'���'���OB�I���O�T80����=r|,�2$�=�l�1lDx��T�'a8�%�]v��B�A�0�,ȧ%u�j���Ot���$�$��'�՟��	�vn,�(S�
� �BH���@y
����$,�d�O����Oj�ɢ�G4u
�@ �H�8i�J��v*����̓B���	ɟt���0�<��G�da�+��v����3N�e=��'�"F�#}�G	V*Y���?��X�N-hdk3a�:<��H�#��.jC�	�|�D<q�F���0�܄L6^�r���<L��a"$H�y����-^7ڙ�qd�?� 9���U�yBxm+�nV�+{(�᎗(k�r�9gԱ\�N��f�)(��Yu�X�M*��jfhY���"BĆ�d�ha�c
����M�Ѥ�Pxh�g�/��I�0	ޣQ�P��hB�o��k�Щ4�ًr�B�e�ܚn�"ylk$�9¶A����!_AP����'�"�'I(�S���i ��+v���xA8bzB�!ٳ$Ԩ�A�>� k���d�'���#��;,B���RdF$<� �"RI�?�  !�W��b{��ٵ�D��PI����@�D�O��?1Kr�=	4Nt(B0F�[Y�m�ԇ�	�I��q膣BA@,�!�an����Fs�I�{ty�^�7!�!!IS#mĬ�	#ct�Qy�Oj�Ĺ|�G�<�?)���?y��X0O (����tL�ź��?�P5H �N<Pb�"�L�*��b>��>1�N���זH���(�V>" �j��	�9������Փ4Ƕy�)��H@��V�I��q��tP=킄|l��	������b��*S�ؠmvցz��*j�ȓ=�����?D��#��0w��-Gx!)�S�gX�����ԘY,:�f�]�^X��'7��R���kV��'�r�'-:��џ��I6E����a�$1H�����\
x�	�t��50�&�)�\[�s\|F��ptb�̄ uV|�*X�c��8V�-���'~:-P�	D�~�xeF�1p�'J J��?���$�<��JɆF��PcU�SK��y���]�<H\�kϲ܋�$Kw޴9��>~���'����NolZ #�%He�ͧS6|�Kq�˧iA�D��ȟH�	���@s�������|ʃ��ٚ�QLX��0�)P�I6ZW�hȇ�ɍs���b+��<Iuk�$�l�a)W�p��xa�mZ�\��P�'%38Gf@ �����<�%����ɔY� ��(՛B��u�(s�K �IX�'¾q"�Y�L�Z`�
�7����
�'�0L��� �D*��ʘ�3�Fܸ�'���������o�Ɵ���l�d��\ Π�d�/�DXRm�� �n���'Kr�'ŰsAjؙ}B �O��k��3���-RH��an��Eyң�[��B���������51�('<#�<�#���d�	ߟ0�	f�4��]�@��2��X5�|����?����s�t�!3������5q	"��m,�OPt$�i�NE<3�U0w�ܦkm�0p�4�7���$�O,ʧ.������?9�|���&��,���}֦�A��C�.FѨ�y*�������; |P�3�����c勨IMb!*����O H�����;2�4�djPXh/N�eza�'s��'�B��O�d����k}֐r�Z/�J��?O��d/�O����MJ�|�.0���ʝ��L��I �HO�ӌ&��8�l�}�:m���)��	�ƓrHICᡐ�{�`�J2x, T��gx`�#P�9�!pU��/(�ȓg20�Q��1vX4���h��Ϣh���4i��-�.�A�OBs�%��U̬A�󠂭6�r�1�,���}��UQF����&t���҆̏ua��ȓ��b����%YH�� �����1p�iU�8S�����	z�)��kF��Q��ȁC��= %�%�
���%�xe��ND�:���J�l��t�ȓ;Pn�Y��F2_�����*DK0e�ȓ7�v�������*s�E1���ȓO~F-A� I:���`"�˃Mt�ȓ��*fc#Qw� 2J@� ��aP�X:7E@7��X�4�C.u�L��7�T8#����#6=r��N+6�6P��VZ!y$ǐ�,�������(6���ȓV�Ν"ч� vQ�Q�H�D%z�����+A�+@����.VC�	�Rc���]��m�� �Nq^B�	Y&ة{7��<=����`�nRB�2i��(W M��B�r�	��=mNB�ɤ}ힸ2�B��!EA�V�E�,B��N��h뷤"*���"C�6s�(B�II� ��n�;a��e3` �:0C�I�-�����%�RE2揈d%
C��"W���A��;xE.��V��1&B�I� ��y𤝚�,����8�B�	#;^�R֤�N�&\�fUs�C�I�9�Rx�
΂=fi�*׫j�B�I	-�f�!����4N�9%�Z�2}�C�)� �MH�K�3E��m3�������W"O��dǞ+��K�5��|��"O$��Ä�<�0��FA�.j�)��"OT���=T�����ӃO�;"Om�����z�ԬSՂ�a���3"O��rb�l��;U�W5i��Q�"Ol����2.d ��
�+�ʨ��"Oq��0W*LQ��?|��6"O�p�k8J�*����=vk~�V"O�����V-�|��L�YT�܂�|RL�]\���ǓO�z�1�?|�&!x��R"��ɳK�j�a�!��>�8�E�l�T�'�R02�y���p�.0��]�-������ځD��	�s���:T�	0>��xkuK�$>F�#̥_	!��[?Pμ0�B�#9�����O��		�<�8�bEp�)ʧe�f�[3�E(I?�p�P�ï�R�ȓB��T'�.�rh��*�T�%�,(f�(�D���ɞ544���K�h�8!0E�pk����˜1$��e���2�� �D�'glqY�x���'(F�@п\�B%���$�P	�'�:�B�f�VQ��N�z��
�'�@x�B(�'�)�e�@A��'�@5)Ir8"�	U�I�EAx���'��i��B劑k!C�@ɘ���'����U���a\X�K��h�r]��':RHXe�Z�L�Dي�`�)H�p\J�'vv�B��6B��>��C�'ְm�wA�����¥�&�H�K�'y�L�@c�h��) ��
���l��'�������gt��
Q��a�Q�'�$�g�6C�@P#N�p;N���'6�ÖD�;+bL	0D��2p�h2�'E�D�"����=�(#y ��'�M���)Ȅ2�	ŗm���[	�'~J�0�˄+��8�Ѝ��^^���	�'�H�@S,�${`P���āM��T
	�')�Ij�@���
�j�58C�(��'芐� �.]�U���Ѓ-̜�`�'�����H��0�%�qf��@�'� �pG�_��b\:u�U4o&��
�'��t�$��!\	��Id�Z���k˓�(OJ`�%<F���Gj�OQ��"O�lh'���d�Y� 2kF��!�>ѷ�0����O38�0��BO�j�X�R'����'O��a��(~�zy��ܥrDfT�{r�J	B���dV
=έs���9+E���U�R�
_�|�cO�*��}���X?�@��HUK�xq�DU���PV,3�0T@8^��bD��Wz B��%�$(t�f��V�<=ÄP�'	�$Ba�6pdH4�`��6�^نȓP ~X��^� ����JB�\�����t~	��]a�5�S��yb�-��	W�O!����	(�y�"����eK��ս,��詠���Z���G�0$���$Ŗ�j��驳�Il�~	��R�<�C�׻Pi����GuN�	U*1� #��vo��ɉ�=��IGF2����䉢w�"���A�`��qJJ8G�����!!'�D��޳R�h%?�IS�u�E�S�O:|����)D��S'��	�qjQI[}a��떃�r�cw��vU4��J۟"~�C�؊O����ҡ�([Z�ȓ'���uF�=/$0�# �f��x�=�$��D�#\��g*֯��O�(K�"]�fH��jT��:��'��r�͙%��q'I���!��G��Nx9�RR��'�0��ċѐPGp4{ �I��d�_I>`��Aa#�".�鐺l��4��C�v�T�B�Ef�!�$J�i�ըׅ"���#+D�r{"�H�
G���\+ԥ�1B��s�� �@Z��Ҏ5���'	-��TJ�"O`Y�oH�F�E�0��pv���O�U�g(B�o���m�!`�?	PG�8�f�!�EO(��[��EZ�8[s#��D�R�%L܆B���Ƃ4i�M��G
2M�l*`�A����g_�V՞��Ǌ\=Z,~౰'�|�v��#֎6m�<Q���:4�O-i��f�F"�r&�b52�S	�' �`�aҨUx�ps�nߩ1�V�hj�z栌Y��k��c�K��yL��#l����h~L�T-ɒ�yg�	=_����Y $�:Qs�mN�V�6����O�Q��@�W\��i�ψO0���Q�<�ꔳ lՄW�
X[��'+&� P�ʺLހss�C*8	�1q�ʁ�Xe칒�۔m�<����3+�}�+�"Uf�R�M4U��)̂�O"�[��G
*(�R� �(*�1,�|:�E1n�r)�J�0RǮ����u�<�S*_*T��j��;�f�#ƇlI(�'�OQ@�Q Ƚ ���G.uӑ>�ݥ%�pqB�a��G�`=��^ f�2B�	-2-����*Y�(����;z�0��&K`�R�[!�%���rCG�|Zr�	�>[vȻdK�g�J��V�Ւ3�^����Z,����
X�m� �"�@��>O�x��J�@��P8��"��H��l�aX�$St	1�LseA-`���(�^VK��2"�B8��&ڢV��l�~jwf�F����QG��<��v�Kt�<�j8h�)��@иk$�X�MOH}RF�GƼZ'I�,�BM	1/���?a��?d�P��Qj�u� �E*N|���*1˜�z��+�c_�{��)�������B?�t�3���OK��b�x���$͊w�@�����2dDB����@&1OE@�������u�'�ҭzӄ�4N�����HNBa#�'p�xM�P螏(� ��d$4�p=��Q�Qyx8���;��1mH�Ko���'AF���D�G�j7��e�>�)�����x��S�t���Ȑh�'2�!��6C��1���D��ђ��7��l��l�!����<|T0�kZw�4���^��'���� iL��9ǅ�^k��0��'L�����BO�DI!hJ��SPnЇ�
l����\�����]��'��Q?)*3�S�1�6�hrmN?�P��\�,i���Xl�4�Fz�\!Xm�0�6���$ͧ"�X�xdG�V��B����@C�,��G�v�h��IDI|�8�N�z���" 1� IӦu�&��U��0v�1+�{Rm��IÆ5&��QS>�:���C�&ɉaŝ�a1�d��)��s*j)3Ba"�OGe
fBD]"��6�h%z���MC������io�!���TL��2EEG$o��Y���2(Z�a+��'�"x�3Ƃ�'�@�6K�d�L���� �J�s��n{E"t"5d\�hO��A�%��Ru���^�HH��O*-����	�P4��I�'4���@���j$���v\��V�E�rP 2�#A)K��A�<h��ab���vQ�I�d��ʇ��;f�����h���>�Ӥ�z�lX�gܹnd����Lz�j�#Ŗ%A�Ɯ��I�s��Œ#��%ېOT�B����_�H�P-;փLRX��ݾp�0� H�n~�Ј�e�)^£>	`�y���m�L�@f�O��Ј�-E��ys3a�{�D���'dl(��ŋ�I��ڗ/Z-?~Hj ��02:J%�S�W
51:��S䝒�~R"��<R�ϓbo�%�Ug9��$Vu��I� �&��f��f��<"S �d��I�Mc�E�r���[D�M�@J&�m��'�
������h/���+��`f��� j�
(��O����'R��d΢=gp1���Q��$�N?9�ط�ē��-�w�OJ9�㑚�y�,��K�Y� ��|�zA�� ��0?i
ґ"�]�Gg�$� ��uH�|�Ƽ0��GUy"��a`��Ɏ_����1���i�+���a�J��"I�P��a��L*R��\��DF�!YX%+�HLy�����
2�<9`�ۆ=�e�����!q�Ń#f�l��fI�H�џܢ�)�K�X��[�:p�I� d�����t} �Ң�.�8,)�X�$���A�C$W��m�P
@&X��5[T ���}p$�V<�vG�.&�j$��	IY><XG��.���Iu�^i�'$�s�h����
e�D�u�t�Ǧ�,l�̹�7��(
�~(� m~�k�*����ª%��`r�
۟4�(}�
�5v�\dF}�-E�0&�mʕO��?n�<����<��O�qA�iy�h��N�c��]4n,��2M�{vh�J&L,W���B�Β��p?�7���a��Ñ,�f�aqb�aܓHi�9�I>I���ħc�<!�!�ͤs�6����bx]��k	diږ��HF��Q�����I���n���͝�9~X���m,Y�r��ȓ@Wn��MZj	0�G�*�p�ȓtJN�����GLr]��K�f�����S�? D�!� �v�p�B%�P9*��ia�"O����&�M��P�̜r�mC�"Oz����A��ȗ���%�J�#"Oh���b݆7E8ıe�I�^m �h3"OX!j g�-g���æ��!@yph��"O�����
|qn�k�e��bl��Y"O\��aL��-�t���/L�kY�z�"O��ф��N�  �d���@����"O܄cǆ��,�p�L�M�Z�0""O �ڄA)�8���	�q�`8R"O����7��TR"�����S�"Or=��F@(�a9��Ϊa��|.!�\�3�bLA!Dr�B�f�H�!򄋛G�`���\Z��D�ߒ:h!�$�#F6��4.�(S�ޕ�P荼T{!�D�HR�����g����(�!�Ԣ3(�DX֯�'�!Q��_�!򤂑r#T��%eK�p�B�LR�!&!���?�d`�!OEΤu���H�V�!�Hv�4�Vm͕c�\��5	�=Xq!�	�<cCTN#P�����)Kk!�$կ
�4��1�Xx��2�ɧH�!�D�9S�]{�Q nK�0r���	!�$J#X7�A b�OC���Ɗ��!��:[\Dy�R(d8j�8kݪp�!�D�CkP:ƦU\]�E�]t!�D�IS>�p���G>t7	��Ib!�S�L�4�0,Ao����IϽE[!�d��en�u,5̀�GbР(<��z
�'���*���>|����q�_;�٫	�'oa�5Õ��Jm��Hʨ�s�'}�ݸ�E�:h7�|Sa�Y4O2Q�'q8I��Va8�y(aO 3�r�3�'��m(�䜷��gI $���@�'3v<��(M@<0��#P}��'ʾLh��-<<8�&�ʨ95�'�e���ץ�h����ތ<_J|I
�'xp����f�Ȇ���J)J`I	�'2l1�'`�)���f�J�f^t@	�'jn��A�7C�*a�u�8tuF���'@mH �8h� �R�l���;�'>�Q@'Dڹk���%�_�`��'�%�u��Te]�%WH��:
�'k���PS�\������9S�@�
�'^2%x����Q�Zu�IZM����
�'�&�K�-[�X� ��W��.Lz�ճ�'�����[~�|0�L
1G[ҥ�
�'zfY�e,؉u2���fꖏ+B��y
�'��Y��Ɵ< �C��1(��'-
1�Rj��\l�sH�79��'o���Ug#<�SFG�-'�
���'�I�Ծc{�ʦD��-��'B5��AɈKjm�r�ʳ�P�
�'�� WL�2TU�K=a�ɫ�'Cf� �`������?^F���'"HŒq�݀o�V}�����A�'lص�EL� j�,k���>D�`tP�'�\@B�
,yf��W� 5�>H(�']f9�s�[ l�D@��o�wOԠ��'�P	c��;y�t�7�K�K�91�'zh�i��ȻZPP�M�+~��aC�'G�u9�B�d�ĤBsϊKVek�'��8!��Yw)s��0�$���'�J�6G�3Xs�]Q զyK6(i��� r���]z�v�[�ɀ�;�% &"OJmXp�E$Hͳ�N�h# |9�"O��-�n�����~}^�)u"O��e���Ed�sg�ܘ`e��`"O����3]��Rp���Y<&�E"O�H�I���)�t @*&!D��@"O��:�$���9T2�"O�I{+��T�`�%حM5���"O&	�Íӌ�ع2㛵JQv)��"O�EC�K�%!٢m�`"�Fp6���"O�0��iĢ��
a�IW\p!��"O��@���n��2� �� �"O\�b4���L����=��ii�"OTy8�	�L��@Z�*q�V�hV!�-���	e�ަ:���Ӳg��dJ!��"rg�����H�lz��'"O8��D��e���[v��.R�,�t"O"�Q��Sc� XP��|I���"O�e�t,� wzm��@7DLlzv"O�9�W��u3�H!�.(76(H�"OP� @�׵V���BQ-�_$p c"OFY
��[�/2n�W���d�r�"Ov�4�ċ�`�Rѫ��TZ�v"O�����9�"U�f�C<BeP"Ob����ҝ>18��񪂗D#���"O������^�f9Q�A B�0��"O�1hB��|�\-��'�'��x�t"Ot�C̜zȠ!x��9pE��"OQ��� �����4m�a`�"O��:��n��do.=���"O  GF�V�v���r�h"OR�W)G3��g��dp"��"O^]i�كo~�2��Z���"O���㙐�D�Rd��gN�tɇ"Ot$2F@@�8q���1b�@@,c�"O��1��.bViZ�`�;��"O�xҡ"�L��3EM�5C��Mr"OܒA�U{�$��%/�2вT"O:��'�Y|�7`@�d�t��%"OvY�!̓#F�@5��E�#ӈ���"O��������tS��B� ��P"O\���6k\p8�Ā�!|����"O��iQ�З���ύT�ވ�d"O���O� :�5ɷ � ~��VW�<��II�4�����!�L��pe��V�<�!�58�xq��н":���U�<13.Ī%0	2#��/8<��""�@U�<Y���+�$x�UØ�<0��s&]�<Yt��Mb�a;�"�sN�p�r+B�<ɶ���i�ܽ  �E���0���O�<i���--h١��%}4��[N�<a�҈*�	`$���a�IM��(�<��FԤd���(A(�6D���'�c�<���n�.���%���$iU�]�<Aw�����+� �Ҍc�kW�<aV#�)z��pr�7ڨ��-�]�<��� &)2d�p�ыQ���� [�<QWl	�	]pT�f�N�)��]�#��m�<��ч��ȡ#؛���J$�N�<�͆���	C����{w	�P�<�̟T�n|{b��XZ�����]O�<��*��]?`\�A� ��$-���I�<��@�k/������*u�����D�<9�W�.ư1/5��]�/ۿn� B�)� �X"�4$WH���;�:��"OF�����ETyb�n�9��Y"O��{�
	E�P���ݿP:a�3"O�y3�3�pmV�t�2 c@"O���b�Ϻ ����Q/+�"OJ,I�B�6��	xPJ�%{��%��p���-5���2P��5��`A�'P!�$^d�z�lф3x�l�D�7i=!��Q y��퓔#I7#��`L�!�DU1cV�4P��~�*��D�!���Zu%��G�`�_%X�!�d�:�:���
I.a+��U�/E�!�dO��x�
�+���(�ꉺr!�$]"<1�s��$X�&)̋6R!�
�2x�b�~&�I����zM��D��xi�UP�� z*��ddG
�yBC`r�-+��Ѿo*,�[&�M��$�Op-ٵ��@-��{��3c� ��"O�d鵠җc"��a�щO�b�e"OJ��Vh
3m����-�~b@K�"O�|�R��k�V� )|�&��"O:�;w�ܰs�����J����@�"Ov<#b���L:�p�åR;?���qQ"O$ev5,�ڐX�gBL���"O\���i�gUZ��Q5z��e"O����N>K�>��EĎqm�ݙ"OLZ2"�^��KG�JND`+�"O
z��ЌQ���J��D^T��4"O�����39���`���s����"O�K��̇XG�P�vM�x���Z�"O�	ʂJ��5�Z�����ْ)r�"O� FƬF�B��$�H��er�"O�8�b ͆����U���x���a�"Oi�Ve �
f�F-Q����"O�+��&Ն0�w�>�R��2"O��EkߏHs�l9�)L���"O�ӵ�]�Aհ�p��$7lցA�"O: vm�p�9�`灀qiJ]s�"O�3Șfjm
�&��e�8�T"O��;v)�j�J��G$�-MZеj�"OvX��� W�6i(�텛vFpD ""O���Q/��b�t�{�6P@�8�5"OR+-ք=�Z�jC��f$Lt1�"O2��WjF�=T�{rM��c6*�q�"ORH9��Q
w�.%b�E��Pfm`�"O84�v'A7n1��2Ám-P!�f"O��C���$xT�s�j��>��"O����(|k��$$ǜA���["OP����1�A��P}0�z3��y��F5A3 P��P�A�B���O;�yBi�����g�]0��r��"�0=q���:I�)��W� �@zl9�y����bӮt�ņ�B�މ�G�Q�yr�Z�K�@rfg�=m������0<���D�5I&�
��X�"ASb�P�
H!�ݹiF�j�d��БJ�4�!�ĝU��`d"$�H�U�C�:�!�D�?��2���2�%9RBծ|�!��#A	��ܶb{db1�G�!��T� x���ߺ|
���!?�!��ڑ3�1)'��4��{P��?[�!�䀕^�8�ql#��(�`�Gf!�M�h2�u��D팕�ǀW
[/!�ͧy�����4W��q�M�`�!�� ��(��M5��I�nӐZH��A"O�q�	>?`�;�'F�V���"O�2�A˫`��� ��W+Zh9��"Oԩ7*P�}�0��G�|8$5�'c剖U���"
ǿW��[#$���8B�	�bEh䪐
E�q�� 2�C�I�-�"�ِc�ԁQ�:B�I<|8��! �Lu�x�2E�.64B�	�wM�q��Q�+:�`��"~B�I�$D:-^���ɡ� +8ܲC�Ɍ9��P`ao�5@/΁�!PDc�C�ɵZ����	W�f|-��g6D�|�7�� ���KfȈ_�l���4D��y0,��R�gm��Oe�x��o6D�\����T!����D�3Qc3D�����H58�be\��n��Ro#D��0P�I�X0D�+�/�i�T�B�`#D�`�#�P&ʝq"��)&.���5D�����N%d�K�B�=R8X���0D��s�m$�ԙ���U�C��@Zb!!D�th�D�#="x�0��V¦P���3D���.�(Ml܈ �i��>RV����$D� ���>P����F3Qs�+�F!D����e^�$�B�! 5pT�b=D��@��K�y9"�UmOO�LtZ�<D��AQ�ӑc�J�:�瑮^�4�*�9D�\��czY�h9aT t��M�w�6D��a�M��Z��U<����.D�th�,��<�� 6n���+D����o���\(����CWh}���5D��r�m��sV�3��°/�6��ci&D���Ǚ?�<�m*���0/D� w�0,;�u[��):-]�b�1D�X���܈1�|Y��)w8y3b'+D�xℏ�$�r�r�!��H,��(D���B�_���26�'�l���#D�Ȑ@�s(�ɨEd�<�T���5D��q�+�$[PQ{"���!�R�ѷD9D�|��eͮOt�a��E��ES�l9D��Q��Pw[�m"EO��X��!�w�8D��q&�WЌ�*�	Z��N�"Dm2D�[q돥rȌ�԰q���#�:D���q�ז;�H���M�-E�9�3.D���V��\�
Ai�ї=���P�/D��qM�8���`!A1j7���&�.D��K�iT��b�� B�-�����/D� ����9"԰�wĦg��ݢ��.D�0+fC,�*iʓ*�4�Tx@�,'D�$sr��
y�`���2�v���#D������RJڵە��+x��qZ'� D��ZRLK\x����T�Q�&}A%;D����n6������N��k�%:D���&��ADF�0a��qP�Q��=D�� a�@ 8�hP;d�V�Ż%�-D�����Ǻ>ŢQ���f�f�bC+'D���Fl��B�Z���k��#{<!�!D����6
,
Ŋ�&V�E�R��- D�PxP��^�&u�$
&�~Dq"�>D���v��J+ZU��KP!�J$؀d D�TC��.].\a�(��u{,�cS)2D��'t{P4�f��
)��h���+D�t�S����l������Ȑ��*D��;���|q���'�3R�<Y�=D���rc�3QX�:���w\��$:D�� r|Q@�\c�|+%�4���3�"OrA��@aI�8��*}BE�`"O2u�ƍ��t9(�i^�^9)�"O���e�j5�L�sN�p z"O|���a�
ES��i�M�dE�"Oi���/l��p�m�	`�lB�"O(SE�RQw��a��
"�A"Op=+K*jsl,�$-��6v �5"O�h��S�^���(\�E�U�/*�!����[���%>� �07���I�!�)h�q���K����5퓬"R!�A����� 3�x�JÌ�!�Ć�yq���I�H눜�'�#�!�H&đ W-���.�y�g�t�!�$п kr����,h��t�H*m!�D���Δh���B!JR{R��#"O>����GOl����P�D��e"Oȉ�	% �������/I�ց�"O*�ے�M/@���fIB�J��x�v"O�\P� �:(�p�E�'���A"Of�I��f'��h�Ŗ43i�!򄔋#6���܆Xt�"5!��#!�ٴ�uCV� �.Voӡ^q!���@=��شR�d(�8O�e!��:p�4��6�ѭy#zM���4rW!�ǋ"m�D��λ!xH�W�_
^K!�Ďo��x��!>��X(��ِG!�䏁x:h��X7�^��E�2!�D�f�&�0� �$�3A��z%!���1��� p�� /D��g%n!�?j�rc��pL��d�" a!�dޜ3q���e�L�%��e��cܙN!�#\���vש0�*q�ȝp4!� �Q2��B�C�w�HX�&��-�!�D�w�l�3
=��y�O��!�dPU!Ԉ��ğ>)��c#�ۋ?�!�DB-/��Xq�S%Y��F_�!��O&[	��h����q��y ��
R�!��y���0Ág� � "`W�9~!���Q�ᨤ'&=r@� ���kj!�d]�78�R��RQV�EA�\�zF!�I=��+Aj�&"�9��*;1!�d�9je����۪3(�+�&m!�X�s��� ��m������^�v�!�D�TN��9"�V>l�TY�2���7�!�$��v�1������LȂE�!��'p宄im��T�̀�qeE,�!��oN|t!�
W��j�ߧs�!���@9�u�'�6� �+�\
M�!��B�����O'F��@��a�!��dx�J�ԴU*d�U-ˠx}!�dʅV���G��p�y���45�!��(���ƤL1 �j���MT�KS!�˙h�Jq��m "�B�ΎRG!�$�!^n<94��e5����!1!��T��2�д<�aJ�A�KM!�d��TL�����#U��p˱��<3!�Դ^�*� 2A\MQ��ԥT�/!�$M&.ahq%�Y;�ȢX�C!�$P/H��C ��a�𔘑�I��!�dV�[8��$+�/F�A7���!�J
R� Ő9
xa���%�!��O�;�Qv��8�Py�E[l�!�D��:m�p!���*��pC�D�|�!�� �\��a�$s�iX��H�{�8��R"OD�@L,yȌ����B6<�~Ձ"Ox%�db�49�y�] @���W"O�0{f��Mv|� ��C" d�͹�"O��1�K#4��RSh1t��!�"O��鐇�Y�H��u��,#T�|2f"Ot!xD9N�����k$��5"OX��H�%�*܊D,�p>�@�g"O�ɚ�@��@��B�E$��"O�`�OƮ/�|�seMA�<0�""O㧖���C��8Y<ʤ��"O�x5���E��D�D�ҙg-~8 p"O���Է|R��;�J�\ *�"O쩉��
�b�DL7i@?=�%�`"O�X��H�gV��rj��:�I�"Ohd0�#��3�X�ț	z|�"OJ@'+�+>I�� �L $����"O�A6�!,�n�����5���I�"O>�@����M�J�(��)z�"O�!U�دB�*����8���ڭ�y� AxhJ8�`ĐK����g#��y�`�+!@�LsC�Z3�5��i	��yB.Y�O�bY��&�Z� Јaֵ�yRCqB�1�bO�.OEtL��m�:�y��/q�e!����}v����'e$𨥪D�EW����"�5t�A;�'ܘ�b�"n�pр2FȚf��b�'n�)�CNI�K��-�� �+j7Ly�
�'���H".�  �����(�h�h�	�'p�� ��F9N�ұxrK�_j\���'NPq��K�=�V�qRE�AE�D*�'f�4�l�<,A��,Z�:��'Aҝ3cOէ[��;�I03Z,��'g4Ma�g��{5�X5A<|N��C�'ڰ���5Q�����	C��j�'�����B�iFtLXp�@G޼
�']2!��'U�L�n�pTn'���'�����@�b(���ghƥhgp(9�'��c�I'8�B��ݛsH�u��'����C��rR��I�7���Z�'-���G�S�?�\ �Ӹ�B���'��tS 0)�؝�S�)���'��@��C���ݑ3��#@�h�'�:Ɋ�
��x�H�d���n�9��'
N� ��ŵI��cB�gA@-��'{m{�a�"�d��@޾jԂ�#�'���XDI)K�k�h�'u���
�%���q(��dA��
���'����_�(v��P�%_�* ��'4�{�+�+-
�g"���U�'�`$�OK#32���ɽ~6��I�'���k�;_1⡥�e� �	�'��\"v�*T$He���"p�ظ��'�P	��g՗)4�ء���k`��	�'�^d�@��O���P�@�^8�b�'��a��'�F�(h�(Z�WW�(H>��� �x�*�ka֍R�����'���IW�(����a=ސz�@b�C�ɮZ�t��7d�4۴�@��C"�C��N����fG��T��_
L�B��<��Xǫ��WU@���_
s �C��l���s7�V�d�c3C�-�C䉫]d �HB' kMip�W+טC�I{����u�%�
�T�۽$����?��S�? ��PR�)Q���bF\_�R1�&"ON�+`dٷLr�](��;E��L��"O�t;2)�	k̠]�e���b� �C"O��� ��(�v��4a�9P���g"O�P+PLä\	�V��=;�P�O��#�`�|� UkE�\!A�p4k%�0D�h���T#{���$�Y*6��cE-D��P�J�&ܑr��)��!��A-D��i��ģyK�����l^�t3�� D�T{UG��=ҵ��o۩\�0{7	*D�h�d(W�D�HժE���EN�5���)D�,{�H���䘔'F�~ahC�5D�T��H�c�8�*%-����3<O�"<��샋��|���ck0mg��x�<9��I�x�����8"�����r�<� �P�E*��I�H<�@Ԫ�h�<��<<�J:ƠS�>Yl�k6��o�<)L�I�D���

\�嫖k�<��(��|}(�*e�ܚ$��$Rg�<9 CKPb�
�Rm��1riy��'8�OQ>�g�͝ &�6��;^�Rl{��=D�����Y)��RS퇧6EN�9�e:D�4��`ޗ��ܹք����	�
%D�L��F��eBRKC��mAh=D�k�&��n%Zmk� �X�Y��<D�Ph�oǩE����9k�� `:D���֭	���ڐ.У�P|R�7D�D)Ҩ�%w�v	��:&���P�/+D�Re䃋3�j�9� � 6�T��5D��ŇӚ��Dy7e�@����%D� )H��;��)9�V�"!��Fc$D��
�eX�0N>iA#LV�VG�ڄ�"D�̈ƣ2j�Zb%�5"q��8�?D�02H`{��RLF/U��cCc=�Ib����H��;�G�"@`�a�W1O��B䉽!hz�+2N��|�(p`'����B�!Ey�$�3�`]�u�(�%O��B��q�N��rh�#��E84��"g��B�?-����o�]Ԟ�(W@��C��4�n��!.� ���@���2�f���&?�S�҄ Kb�He�ÓP[�ă� f�'M?mgΘ�7��3d��=�����l/�D:�	G�O`�t*�P�����k��p�	�'_�l{�oP8��̀�� �8��'F~U(����?.Ht���$ײ��'�ƕy���{���#�T�m�@z�'��@1�UH�ʥD��b� �+�'q��@�) 'T��R��+`od��'�hTE��#=�zU3S'�\�^=��'��ɠ �}Q�Ah����QƑp�'���Q���ĥ�q�(DD���'W���]��ީ�V�� P�:uC	�'���FZ=k�Rؘ�/��N��
�'��Kb��:��5�%��*p��[�'1�k�j�yTU��BL e���'�����%G�Iر�
���{���x�Yw<�p�I1_=Έ���yr!�� 	��B�+mp�[',3�yBl�9mv8c�C7�Z�im��y�A�I�����G^�b��	Ԇ�y����'�:�J���ZiL����?�y���K� a����V�Ԙ�C��y2�	�j���CT���S�D��y�Љ5"A�у]�I�0����y
� ���a�Qd�H��܀7%aj"O4�b��2wE����"> H��"O�p`��4 ��@&U�dj"Ol@
���;�B�7D�{�|�v"O�0�c��%TL9��;if
	�S"O�3�� �v� ��ˆtt1�"O���"kVi��x���#Xp��"Oȭ$gџC@!уC�Kd��"O�2G�4��ua�V**;Ik�"O���'�5�����2�-�`"O�I�Sk6	=>P�c����"O�P"a��V������̰��t��>LO���p�e�4�բd����`"O�4R�ޓ!>�A2t�\Hl�@�"O�u�b#O�|[�m+�� ��fd�!"O���"�+N�Ɂw.ԣw���t"O�8��ET�R���i}��Bc�F��y��I�B��e���a�̭�/��y��;(�C�Q^��jb����O�"~��jL�='T�SТN�ް�Q�H^�<!ᥘ0+A�0`�m�-C�%�u�	f���O��T�H.G��i��&C(�ā�'��@	�κO�H�ؒOQKX�T��'^�M���Q��ƅ�j	'o�qZ�'�Iq�ߖ��P�	Mx���'��"Q
m�.h��?q�@r
�'k i)U�FuטP����V\)O����|��i���F�	`oW�p!�d�6@��e1����(�l��Ά�!�$��N>�UrvJ�=	��E	�(�5!�D�"�eB`
)S۔�8#���K�!�Č�;��Q�p��>)��)qD� H�!�d�u���x�Y���ַU�ўT�?��O�V(A���.�h�@cޚ�!򄊗+�"��N�S�p�4$΂E!��̜!�t��W�P�Va�V�\%�!�d:p�ce� 9�(��WnX
�!��V�2!�t�BOW�X%�ܡQ!��H�JuPz֌�S��	b�(v�!�=���RFD�V�|H��E<�!�d��7�!��"�7Vcl���ԄI�OF�=��*���(BDR1�)3�)p"Oܱ #+P"-' H"���H|��"O�, �C�&^8��0�8�i+"O�5[�凳A�����7��Uڳ"O��"Ac̠&�LT9�C�?\��`;�"O��`�	�0Zꑻ���v���e�'zў"~2ө�5�LY��
׺)gtt���ϗ�y�(�9<�E1R'3�ڠ�����?������� �����J��5��!���bh.D�ˀ�J"?U�Y0�oٱP>�:T:D���m�L��D ֊DZ�LQ&5D� R��ՠz�N8)4(�L�P#!�'D�p9�M #h�/-S�ʧ%&D�����P/	~ͳg"8"@��ë"D��i�W�2�>%���?� �2�j"D���pH�0� �j#ʙ�5���	m>D�8P�Y@3 ���Ԯ��ܣ��<D�Z lU&!&�$�SdR�!2��C�;D�x�i ��*H�!#O@���Jg�9D�T"�xA-#��ڿs�(�a&2|O�c��S%g\|5��L<�t�H.D��(3��v�kE-P�Yuش�f�!ړ�0<����n��g	�^��}�6I�|�<� �mX1�)A��Y@Ѓă�6R"O�|�t�>!a�����'k�:Q�"O����ܔߖ����;��8[�"O4�A��[�!���a��3x�L;4"O�e�p�Ȏ�$� įؙ ����"Of`JP�\$n4]i�e_�i(x�v��%LO��0c�h��-��n̂d� �"O���-mH��9�m�>m�(�"O40%���E��LQ�*$x2��"Ovk!���l���:hb}�e"O8���;�(i�'P�	NtX�"O�%�SG��V�\<��2ͨ#$_�<�V(�9���`N.8��x�7JX�<��n�v�� ��,f���#%�T�<1��w��IAh� �pH�^x�<!0�O�W�<�h�OPB�-���p�<�!�F�6I�L�h`�Q�l�<�2G؂ �؜��;Ma ���f�<9��m$�������6	D��&hCc�<�g�5F��m:b�ʓn�����+�_�<���Aa(�R�����X�< ��Y���q�"ڋx�00��iY�<�C$_*d�n1s`�|y���ԃ�V�<����<ר�*Ʃ��|�(��2�]w�<�qf�'% z ¿1��i`"	w�<Q1�о8� �2�[fTu"Io�<�%�&���	R �?3��1#��B�<���Vw�a!2�I�a �2�m�D�<�`n˝kˌɉ���֩����C䉙B�d�p6lҭH�e�z�C�	C�֙� �n�Hł&��-e�C��z��	[��	Pdyv�[�B^fB䉶)�z�#��%�&�y`��#�HB�?�f�kD̚�q��kڒU�B�	�b�Z�*'��*�,S!`9&�C�	�Lt���ԇ˶鸰��MS��C�I����p�ܒtl؈Z$�� 7��C�I�_|$�Ǫ�m�p�S��dU�B�-r���BO���7!�?@��C�ɬE��$A�fސ��2��e���$d���s��gʭ����?9���)q� �O�� ���ȅJ�xRԨ޹-�>�����Z���*m�P@"��s��ȓ� �(?	�&�Aԯ��D����8xn�V�E�$��(a� G%%���*���esv��cA�>/V��6��ԥ�,�}`�
ɚSF���	u�'�~JR�d["�k�OϢ4���ߓ��'�Ȕ�V��,Gp��7�G�6�D�a�'ub<!K�{�j���ϴX`����'���S�<���BM�T�&��'N)����L� \��-֛N�N���'����Ə�	K����D�h�*�'vl�3�O/]�8�c@eR:��0c�'"(��E��s��x7
���0�'�@���"�;c����f�S(~ܼ�Y�'ح"Q��"��1E3z��-��'�d��f
^�z)^,��b]!r-~,k�'�(Z��5sQ:����\�i��d 
�'���@��7���91�	�LUJ	�'��q�	�o?@K �\6�Huq�'SrLӒ
X�.{ެ��[�u��C�'�nP���.WV��Hޥ2���J�'������m	ȰDa˓A�B����� ����
N!;����&`	5ʈ��"O*�SOG�Fl�
�@4h�a0"O8���R�6m��^�,X�"O4L8ǡG7�B +g	�j�����"OhT��X��Z�%�P!,��lK���=�S�	�j^f���݃S
��1�j� !��;r>Z���g�$V �iaW�Ѝ&�!�dM-�\p(�E��)�<R++-�!�·_bLI�4�O�A��M��鉿l�!�Q�q��#ClɎk��C��݂g3!�@�d��m��AOq� `����O��=���X��h�+Hd�d��h$Vv��|��)�SB�8WhF84ߤ��-Ȯ)��C�IW���#�Ɏ��F���J�	�'�F|p�¯Ft�qi��J���	�'��L2�␈��}{GL׻=�� �	�'�L��`��eLt𨍧^�Ȱ��'.�u�po�NSX�����[8���O>����)X5�8LJ��A4G������(N�}2��ؑ�c -$��X�U�Z�G>��(D��a�i�W"�K$�ܶ#<MI0�$D���J/Ǹ��.��x*&MJt�#D�\�F@[+9$�bD�+���V� D�[�ꕃ_��̸"�)���K4�=D�@��$�|wBuBV  ���L6D�lZueR�;�6့LΔt:���c5D�0��\�BC~M�gKY!b��PR$	'D�$�rb�$~k�i���ڼ1��lǀ#D�XitFK�.B*���K�Hۚ�xT�!D��j���&>�!0��X(iDL��?D����ۏ8�q�4BՇ>h"�6�8D��sm�3y"��b��ԥ(�$N<D��P��ƿ�̴qV�2�ڍ��:�$�O��O�"|Zc�#x��26BX�w�����p�<)��C�8$���!��u(bp�	i�<�i��&��������1P�o�<I6	ƊZ��Vo_�/��V��l�<�wO�������K4T��S�k�<y���L�`�&k��O���iS��g�<��Ԩ W��� �5�,L�1i�k�<q��%pe�4bU�Nu
��3��g�<YR��2\`(P��^.^4rT;d��x�<���&�8�'�, bi����<�!#�0il̪(a2%����y�<م�-�ք��(�&l�Q:��y�<I�"�3i��A��;a˚�����J�<����%piKr`�7ײ�;�FHy"�'��y�0O�����%U�6��eʨ!�v�z�"Or`ie��	�DLZB�	!)c0"O���p,��	h$C�c�x(�ۆ"O���0   �␁X&�����"O*dg�����)�� �h�����'d`-x .ɓ#��U�Wn̳E~�D��' F�b#�I�T����K#: ��{�'`�X3r�	�pn�ݠ��I�0����'��Q��`p�a F~Y�'��Qc���3a�jew�0�D�`�'���J�;���Q�#�"h�'���p�% ��$�Fm�> ����'2Q�%kB��8)�enW&
7�x�<)3&�g��p�̨����s�NP�<��C�^k�A�@U�'���K�
�E�<I��_�L�( I�w[����H�<9��ɕ)�tp3�W=�z���D�<� 8�%�T+u�t��D&ن��q"O�M�֩G~v0�g�ɁQ�V��t"Ot�C!Z�?U��"Bh�:sY��{B"O<��enU_��D��fĬwG&���"ORHÎV�5S�����" )�5�"OBِ�)��W`p�8v��;�`���"On\�P~l���OĿ?q��
�"OV��E"O�oΔю�!TtL[�"O<!��W�zf�p+�ߺ`QnĠs"O��s��߿=��PS�PMB��"OBː&,_cr9�j^�&'�q�g��J�O���AE��~}Ρ2���d���';��Y�M�qO6TA b����hc�'�� �B�#z�>Hc�I�~��E��'}R01�MQ�y�h��)�p�~���'$�ҵ܃C�&�ō�aB�hI�'�^8�cX8,q�A*��̋P̄��K>���)˞Ul�9Xb$�����A"��FO�{b�$!@��5��2���0�Ѯ&;!�d� ~�0���/*��pE(P%G�!�$�)� d�b�Cv:\bǓ$!�AW�Y�V�H�=2�b�F�	!�$bR�I2�`�(�V�7f�S�!�ď��L�K���6�Te@R>#�ўl�'t�P�7���vg`1ɇO],���sC)0D���f JAo,Eڦ���C�lI��,D�ܪ#o6a(l�(�C[!�v�{�'D��c�ԵKy
��D"^�.悙
�3D�$0����y�S/��D�Ъ�!0D����)����&�� ��-9@:D��{�g�?d*
�e�p@�i"f�$D�X�Eh^�S�F<X%F+-��Y�A$D�� ��T����3�	���P��"D���ы@0dY��`�[䡙 �+D������}�,���U�
����+D�P1R�J�HvYI�ˑ�9�~X�%D�(捖�(�A����)~��4e8D��cc�m�F�r����`u�7D��a&�[9d��M�"ƞ#��9KVJ �Ot�>�jx4��n�ꐥ�: 2bɇ��R�{W-_@Ҫ��DT�p�(���Yj��!U-�)gg�%��iȷ5񒘄�pW8����q�|�JdY�I�杆ȓox�02��k@�� mZ�`|��2� 8V̘���"���}6�U��	X�'�(A��E�'>!z���&�kL>��,2(�Pbhױu:�H�SA �5X*���kh�C��2�FP8�fQ�lU�8�ȓo�`�8�#sj8���:i%�}��/��Ȳ��L��t�e �8��@��Mv�l<T�5�l�9���ȓO�BX�����i�����Y��a�6L�f�κ}��1A7�O9/����E���BB�$?�a��!��2 ��ȓ1R
�x���>n���	"rbn�<q6d�1�()0�	�g�H���i�<yF/��>fıЩ���P�DL�<�̧bQ$�Ǐ�{��Q�1-\�<���(u�}#���1o~�p�PH^�<�Qo.o�B\���дoJ�8��o�<��b(>N��!�-0�����m�<95�+7r�ŨDJY#&\ �*�,�h�<�p.	'h�� �f�J��0�N�<���a|T�2��^{"\CU�F�<� T ��Ę#j�x��͝��tK�"O<��fI2p �0��*�2�� "O��� C�X��$ۨ���+�"Ob����T���C3����"O�)� ��6�Yv얳��$p�"OTq��A#{�*�jA��/	���[�"O��g�D!��x�	�	<�
�A"O�
�P+%�@	w��J�&Y�#"OziÕ�#e&V��ѭ�##�b��V"Oڴ�p�J�U��81#�C�4F $Ң"O\���
zh��E�ʤT,`�H�"O ۣ��7(���P��TwL0��"O�PA
�0Ԇ��@�o}JD"O�D)叀.%zP!��ݤy�� {D"Ojt�S.Y�H�R��@�9k�t�s"O�!�W(<P���+�$
�Bb"O��ɂɃ�l��
а8炝D"O"=���
QQ9qj�$U���D"O�\�Pg�!Wv�ٱ��k���"O�%2V��z�x�H0٠*O�l�$ T�8�ZRn܎\��U��'��i"��0�������S0H2�'�%����2zD��WC�*F����'�v\H���_!���fK#F��K>�����Y��21%Dn�P��,�2T!�R�֘�ۥ`ڢ:�x��69�!��
��h]0��mߺ7��QJUjZr�<Q���L�*�v�X�8pZS�Nl�<׊�;bfv�	U"S22�Bj���S�<	���5
�u��kA.t�8���ƕI�<��S��z�k/Vh.$)�D+�J�<�� J����
�a��|J��a�<�˥|k�wOz�6�{w�S�<i�L���|� �d��d���S�<�AC"n���"բZn  q�G�<�q�S*@�"��ƞJ���9�c[{�<���	�^����{*80#�Op�<�0�Ȓ��j}��PċF�mؕ�ȓ)&��c6⊒W�&TA��3FɆ��ʲ�����o&R@@Q0��ه�i���!w.�08��<����#>��ȓp?r�d LLf��v� J0�ȓc�X)3M�0s$�ɃAσ-p؄ȓ"��b��r.���*K������*?n��Q@C�B� m��#UE�Y��1�H��̅�l�sLR�rD�ȓy!�r��4MǦ��q��*�Q��f�ʀz��R�1���c"�ލx�%�ȓZ<T�R��s�\��SBL�`�ȓ_R�Z�v\Ju-V'���"OLt�`� �$z���s:,i�'��% $L�=6H��u�ݽ	� )�'m��b!�|�xI" :rm�'D~��6	ǣ�r`IuF9,Lb�'�N�`�	��(����!��XU��'� ik�F��%������u�f�9�'��ut�A.*��TEG%l~$���'[R�ad�I�΅��1�
��e�,�y�� %i�����DD�0��lcp�����'ў�Ow��ڷi��i2�Dʑ�Ii"6���'��!� *�`��A�J���9�'��訳n�2'.� �#BRb�`�
�'hl�T���I�����߲F[:1��'�0�k���'��2C������� v�m��2��D��$C�3	����"O�!�ڕ?�2�0�_|��E�"O�$�$* �:)��{�M��n٤q�"O����k�:R��MR�f��v���"O�b#E�0z(��Ñe5{�hcR"O�Y[AAY7FLnHaC"
����T"O�L��]�		�u[Qfˋa�d�"O����+�"z*p��(R��z�"O�5���im�挗4^�D�8�"O���Fւ~ZmC�aI uI�Q��"OR�:�%r�:��@"�+<*��s"O^�JV�M�/�Y1C�d4��"OLy{���*P�\�R!5͞%�!�$�~���`�$A��髳�`�!�D��`�rpʐ�S3�D�)6@N�z�!�$�g^��+�̏�B��x���~|��p��(���g*�
����"���b�`"O�R#Ν 	t� �������"O,�@��}�e�����1cp"O�H2���Z�عC��;�� �"O�;��	 #�,D�猊8�jT(""O�w��a[�/��O�v�#���F�'a��,�?�4|s�l���v!Æ�y"�]h�tE��x
 �ҵ,���y����z' �
���n�<�0�A�8�yJ@8p�8�d��Z�:P1���yҡI�a�I���A'Q�n,(f�T��y�� ���%��0@7��0���y��{8*�)��ŝ4�LuI����yB�k�@���߿1��y @��F��$�<1.O<�#	r����
�'�P��d�#�y��@�ܵA`��'��d`��M��y�J��
�6�[��X�D�Vȣ���y���v�bH;5�J	PZ�Ja�֨�yR�]3oC�!�	�ˋ�y2���1��!�#�

��q�#%�y"�X'Nl��V��z�<��F�+�y�j�$�zu��Dē-�A+Pn��yR����JV�Ķ-r��z���y�A֯GǬEjGȞ�u:$ �F����y�nP�K��5�0�	w�:�(���ybc��I[pE�9{�pa7�*�y� ��|�/;h19��y�&�>V-I�TG͋b�\�1E��y���(���ںW�D�P�[�y�W�0,t85N9+�1ՋZ�yR��iȘ�3�,���kT�A�y�=a��J�/ٕ1��Kt����y�,-r~���	ο/25�Q��y�ǝ$@�(14a�*��l`��"�y��J��V-�RJO�JP�8hBC���y"ll�4#;E1D�x�E�/�yB���]fА#w�ș6�ek�ƌ��y�h�wJM���\\���CCB�y ��9���Jb���@��6���y�!��Iu^XR���.(�Z����yb@GV�5�@h�j0�81��ɕ�yn�r��tj�@]�i>�c��T��y����K�6��kJao�XQ�`J��y"��.���'�\�"A�	�(�y�H$�>�q��*�>m{1)8�y�.��C����GZ�/�rP��l�!�y�*��@
��A/Z(\!0���y"�
	[t�+bH��3�C��y
� �Y��'�=",�u-J�s��`�"ODP�eXF
���JF$[���B"O.|�p,�+"[δzi�%��#�"O�#�o�T�����<3�,Ѷ"O��Q���i�f��D���h��E�!�d�r�
9�T���,����f�)�!�@8�:5��ڥi�T	:��W�!�Ċ�k�@|*�J�5��i"�ɵuh!�$Ԏ7ltth���x0�X�IQ!�D/N��`�@֦~'�8k��Jbj!�D�U=���q�ۣn���D�_V!�$K�Z<x�CGl���T� ��
L�!�� �6�K�Ċ4#�n!QA�9!�$�=Y,����ۡ
.�\ �iS4i~!�ȺqR�Q�
����ǎ-n!�*)½AE#ګ\
��ǆ�	[T!�$ �d�(c�����+�/��P�!�D��N�t5�"Q�����W�!��9,Ubq�┕r��a6h�;�!�[�e��e�!Ybmr�U5-�!���qS�G�!v549��e
6n�!��ʒ^9`��5L��a0�e�f���y+!򤛣$���-O�@ȳD!�!�D��q��� K����`�C �!�d�3<���+�a��;1̞I!�$�w`���w񨬹'A*/!��
ھ��B	�4w�29��o͙"
!򤂸v��lQ���%{�� ؐ`(!�䃡#m��m[�N^0�$��#W!�-(ȊTC��
9Bp�K�Е/$!�$Af!�I֎S"*D�@ ��!�$�3���92���k�(��J	�O!�$P���i�-[�=#�iA'!�dQ4�١Gڙ�(�j��1I�!��\ @��@��*u��`{U�ؐ�!��� ]�ex�+�����oL�!��¨VMf��
4}�
$�([�!�M2�L�	4	�=�
�I��S�!�\�5�b5zgGL�|�� Y7Yv!�C6	Sn�{�T���8��]�l��)�)����n�%�Vm`��S��Ո
�'Yޘ�ǣ�+H��F��{���B
�'&�`��`�+_��a:�)܄=��E�	�'Aj����U�\�
�w���:x ,��'�er���,w��f� dX>��'�	��l�P�d��4�S�\o(��
�'�8��ӆ�4L��[�!�9N!.1��'���8�)͌*렩 �*[�Uk>���'ͨ�ӡm�C�jE��U���i�'~pa��^!<�B�A`ʈ�F\���'Pf�z�)Ĝ�B)#�$R�Dl���'c��C��"ho�!����s�&	�'�v90��\43�����Ň;�$�
�'ʹݙN��j��(�V��=زQ	�'k�(�DM�G�-�4D�K�by��'�Ld@�@WfW���#��C�����'���D�T+�!���X-:,���'+1�C^���y���j1��'�ܐ�ϒV���S����r
�'3펍g�����	{a��'{�h!#㗅4�4���J�/0�b	�'�d �l�M2�%!_�T*e��'5d0�C�w]�u1�(sl��B�'�
���b����erS����� (��Ąÿ&X��#�8Ԫi��"O�RO��$���:���*%e�D"O�5)cH��[������lm45x�"O =�4���zX���)�tHp�ʢ"O�B&��2���b�'v3`ٻ$"O��`��4s0h��/J50�"}S�"OR���Э�f���V0Z�H(y�"O��y�aR:`".��I@��\$�r"O�0��ឆ:�$<�(N�����"O(բ/iU���E�z�J-Jw"O��@��4���J�ǝ�c]�uK0"Op9QE�'dR��"GQ*H[��"O���#b���@��;>U�I��"O���$Y�X�ં�מR<�Y�"O�Q�V�*���h5#�
K!���e"ON���C�
���!��K�n�x5"O&u�b�3o��؛� 3,4P("O���F��"A0h�@%݅FXTh�"O2Q7J	�Z|�2c��<�p`h�"O\�3D���(���Lxމ�5"O��g$W:>�LhR�fϢIf��"O���1F��{��Xq��@I��d;�"O&0��*N�L�˰	:75R�"O�����^�[|P�
6HI�V-&�	"O q��ӏ:誸���ϓC��	�"O�T���	x�I��F�h���"O����I�N(��P��;[�X�V"O�L��a��BJR�i��l�b��"O��r��/�@e`����,` E"O$��d��u��x��ǶA����"OX����-p� ��7iޅG����F"O��1�`3w�܄b�h$"�m�"O�1��^>�����ه/vD!0e"O.�+� C44LR�bD��1j��s"O�z�"I2%���HD��)Z��"OZ�ٳF�� ��ZuWHz�� "O�-���WGD0}�c�Q�4d i	�'��T�4�
?N<�XB�	ʬ�
�'z��/ժ/H��N8#��K
�'O�0��l��@d̢cC�S�ͨ�'���pe�]��y3%���nA�'ޢ�#ANBQ�x���wᮤ��'\�0��+��}����G�>rި�
�'3z5a���WcH|��c	
8�^�h�'�%!C�h����g�PX)
�'.�a(U�ȉ%�X��e�M.0��J�' ���@�
tV@{J�]��y�'w�rs`��Bi�͝?52|��'��b���4"$�%,�`��'�ڬ��OF�O�+�CӨ%�
%��'^JAY�N�3��u� ��NJU��'�A�ʑ���c�i��2�,P��'Eh���DM���� *����'@,���4��$R� 3�f{�'�NU��j��m�&␂��b���'�#�ފ[Nҡ���պ�P���'S������5EnB���ʀ}7lq��'��96 ����'�[�E����
�'�jY0f�@���:���9>�&�8
�'�H�
�fB�&��W���9��iR	�'�J��I�]b�,K��̳�:$)	�'����^��h�l@Jt�S�'K��Yt��0><�yJA��0���
�'R�Yy�l�U���F���7�B�k
��� ,x�4k��q������:K�*��"Ou����Hp�^�F��("O8I��(�0���4��1$`4��"O�} ���-��a�P#��p�Q1E"O�%��)�@��A��YW�Q�6"O�HX���b����AU
CQ.ac�"O��/P2[��GV9H�D=z�"O���b�9$j�,jȄ�3"O��i%PB2���� �H)(�"O��B�N���=�uJ#Zޠ\��"O�Eq����P�狂8����t"O���{��H˒#Z��S��p!�S�och�NH����P�6]!�X*l�Æ�� ,���	lՒ2�!�$C�/�Iȶa��bE�њ/�!�يq4����P�o��iC5o��7�!�䜸Pീ��K�s��[��<	u!���~C YJ��"�T���@�T!���P@^�� �ڮ&�0�
S@��!�����L�i�+��9p��)�!��M�g{��%���ph��O!�dHHt��3"�`�� ��Y!�Ɯ.h<�D���K�����q�!�D�'J%��I�F���DAsnE3�!�dȽ[xV���χY~��0��D��!�$6��1���<hP��wn �0�!� `)(��D
�H���0��ϡi�!�DQ�L���5�]!X��s��F�f�!�$��^���x��ǹp�\Q��_��!�]�+�:)�֗dD�D4� [7!�DV3�J��C�և5l��
�M0!�d��i`6�i�= \�����/!�"S�����- ^��C��#!��)V���H
 ��y1��.F !���s�v3s*��9�:��,
G�!�Ƽp��8�b�6R�p��+��1���D�&�8��B=R���(���y���,}~��y3�E"7�^<�3���yR��C�ڕ����|ܳÙ�y�fU�2�ə�{�J�0FA ��y��^Vnx��@&ޑg��q�� �yR�F3f�L�r�bR(�~-y%	��y�#�!V�D�d�G�,�PƤ�?�yiK�1���#qoūE<�G��y�.�d��Q�y>!i�c���y"�
�T��9Q,͑wuD}g���y�ɗ%��,#ec��r���E�9�yR��8f��(�F� @j\P�
���yb�ʣ'p�$쇠48[P�y�*U2p=X@%�'�8ɹ@�
�yb�ә!��x�Kǉm��)�@4�yb͍�d�Űف2�N5�gjJ��y�M�zg�!� ��0��Z$f���y¯סN�2 �P#�^�<�ÈW:�y�S�Pm���6)I��Z��y!�,h�nX�DK�9!���E�ŭ�y�m n�(h�瞄i�i�a%5�y2*�&m�ݘ�FL8v���`���ycC�9v$����-@D��n�(�ybi��d"-����,��xV+U��yb�^�dȱHP�)�H8�p&��y�S(M�R�@���p���ʂ�yr��5'!�)%V�f7���1�҈�y���Q��!Um��s��9ā���y
� �����)n%��v�O&rQ��"O2��$3ҵQ4m��#"O�j��X��ʜ⥦Ӗc��m�@"Oܱ����	%{���������f"O*!����82"�PU�����"OL8
��Ӣ�r���)����@"O�}����z��[e�R̈ac"Oxu�fĳHW�]1�i�-�f���"O�����5Ob�=AG���b�x�"O�t�FB��)A⑮!�H�P�"O�	X���X<J��aɒu;V"O8<�2�E"/���D/V�}���A"O��� �ԍA�Ҩ�� �������"OF"��¾Q�D��� Z�z�9d"O�U�Fl����P�Y�S"Of��MW��v�$j�d�ZX�2"O�]���YDj!A�'؝� �+�"OHi�΋�J)jhG�J�r�ȑ"OJ���@�_�N�����2���a�<��aT���y&.Թh"�t�Xb4B�I�E�T%[񏍡��Y2@eŕ)VFC��v-��֟>����+g�8C�Ɉ584�����13|ͩ�b��|V6C��76N�C�Ċg-Dr"I�m��C�I�`>��#F�){g���!A�\|C�	�%
J+�BF�NV�Rψ=�B�I�Gz=a��%o�����I�l2��'�ў�?��6���^�ܡ���O� z��)\OPb��9�,n��ek�*Q�i�4�e4�ɠ,(az��]�]R�Ԧ�:H�^�
��,��'�ўb>��m�(vTj�⑃jO��P�# D�|�F��;��Ģ�lQ�Oc�9�s>���*)ayR��_6���i��M¤虧�y⇛		=��3�1u�����J��'J��뉴\�l�Z��Λ4�*�$�-��B�	8Y�z`k��"bdN���$9�nC�.W}�tB�'�&6쵃c���\#?A��)H�$bMj��*~��b)��Pu!��	f�j�Q�\#D�� PM s���G��I�N�
�@�[?pb�J�����y�L҄Z8���L ;8D���������hOq�@D�sK��W��HdDB���8�'m��u{���䬕2:/r��5'�8B��B��2��i�.
�x�P0*.��C�Ɉ�Dʥ��E�:X�R�f��B�	/P�81�Fzt&���f	3��B��K�t���O	C�ҴХo���B�I�U�v�J��iS�|*�I�}m
C�	�jU�,ycHՏtV�09�)�	��B������uNכيx:�J�Af�aF$D���`��X���qb�#d\�S��>D��a�l�=n�X)K�OM�����p&:}��'�45��A*
<phʆ�<�@��6r�I,�r��jQ0dSn\ѓ��p�C��8,qx�V�[�<�Z/C���">1c#��D�S��DǄYY�S����6�D� �#�TP�����z	,�ȓ��)b���֔����� �ͅȓ_˺��ҢpT3 պn��ȅȓ���̭qMB�H���7�����-�:�SܧyT��
��N���F�S�F�ȓ�r0�D�ȼQ����#o����?1ӓg4�����A�|���(�>]��A�ȓbB@����R�ND�$XD4���S�? ������*�,�82,�-,V2�hP"Ox`b�,�Jq�e��ӣBA�Q�"OX�k���*x��j
�9.R�k��|��)����`���h)��a�)d�FC�	V�&x#��0>(�a� �C䉧vl����3�$�+�ˠl\�B�I�WV�$�Ҥ�6�"M�+I�5���V�ў"|�n�oK>�Cc��!G�j(�w"@x��FxbɮF��d��Ŷl�p�(���&ɘ'��{���\�"���c!⌣����hO2���� fb��v�Ӎ{Ő9C��5=!�� K˨�3&n�)��I:B�-|/!�$�͌(%�T�*��1�&
!����U�M�yF�����L-7N�o�Ο��?Q���A����6fX�5�(s�*S=ax!�$�B�P[�Dǖ;�Hs��;W�!��r`�!�r5�e@ Dm��D{ʟ�d���uWҐ��ˆ+@�iȀ"O�=���v�d��eaU�s":�2P�gx�8j�#]тu��n =�D�da%D��`E@BX©���A*#Vq!���S�'wayrI]���	 ���uh:�0?q(O�\�LS�@S0%��b��V�iI�ɡ�p>)q*\/����琔'���s�YA�>�D*�$]����O�tu5�7>f:Iʰ��T���#�'��,!�O��6긑pm� R�⩙�O����L<�'�ē/z�T��h�-����d��bS��Ɠ(�X{R,�7lt#���J(��g�$$�Xӓ�0�p��O�o�z�n9<O�"<�5��3"x��e!��_Y����gk�<�� 7o�d��̂!1�,Ca�Oc�<)F�E�
e�`�_�H\�"��u�<I���Rl�dRՉ]%@/��z��[n�<aҏ��r<r��ĤWz� x2�Vn�<�%§pbQቅ&f�x!P�Sn�<�gn�,6�|{��(�B����S�<����,5����:I�	%aPt�<�"ϑ�It��5�׹s�X�N]l��`�'�V,�q��^C�
7�W�_V���'� )Ɗ(Vt�i*�
L�Q���O���$��6���H��'m?�����/O~!�Ӧ� �����i׊�x��<+h!�$�g.	��K�s�5�"$�YJ!��)}��-#b�Q=���C��V!�d��S�mիCӺ���dR���If��(�ޝ鄡�	M%
\CbL&R��P��"O��h�F	�>��cC�W!���#R"O@���?t�lH�	D9I��$9��'���/6����)�+�IԝZO!�dY�G=����3�D�2&k�O�џ,E���.s�x0���A'O�H�
���y򮉊���*��ϽM�����	��yr�1|��������?b�Y�����y�%�a�l�P*IA�YcA����y"�B�B����rˌ3d�0 �@���'�ў����3��*c�{�!��]�N���0Of}���m�|j���l�䐔��^���Gz��ty�d�ay<�0��>� ��y���&R_6�2���~�X10�,���y�Έ.a ��AHܻH���Yc���y�ꖳEerȡ��+;2*���P��'Z�r��"l��&Ǚ$�,�k�'�La1&�H�G�JI���)#)�5����M��y�[?#=y�WV��P���>�&��p�Y_؞��=� &�XacȈxyb1�ץ�1�e@��'H��n8�4;�P
[�T��I�8�sf8��p<�ة)�V�YR��!1c�WiAQ�<�R� ���JI�rPy���Ԧ��<	ӓo�L���˂d
XS�#�qY@�Ɠ�����)l����ƃ=b����ʝ��&4[�Jպg#"k]�q�ȓM1�*
�Id4B��d�l��ȓ\:u�$!Y�2�����:}��<�ȓI�><�d/�%b�T�&�@B
H��	~����Ɖ��JrF
?5�B���2D�!򄅈s�����DL [Al�+�OΒ1q!���.H�~��ln��*�#чyj!�䘁�e�g��	l�eq���;1f���)����mޭ��  �'B�R���o0D���%+� ݛ㳕8�D� �/D���u�5T��^�Y� �C�-D����fՌt�u��m7F���&D��q2��:1�db@#B�h�<�0#(#D����2&���q�B�%,H`jBH?D�t�$��*N�"��ՅLt�Ą���;D��Y�D�'e�śÊ'���i$"/D��A���{pXl���:@b0�v�.D�\�!��,@j�1�u=/"�{tD+D���@��h�� �fE�!J�
�X��(D��Igo����؆�հ@���)��#D�t�R�f�h��D�T�R0t��) D���U�Ն�(�Sw_�X����+D�\9�� A�VkǃhD�<[ta)D����9� e+�/�!�M��J'D���7���-q�xCN�2<P�q$D��#f�9�(���o"���V�!D���r�	H�2�0Lڧ,
l[b=D���@V�W4r�@���_��9!!<D�)CM�s��aD�U>�QH-D�4��G�m�n8�:'�-��C�I.].���ߵ
�R5���ؒ��C�I_8-ڵE��#�0=�o�g�nB��8B�*):l�4h�[��C䉣6�U`��Rtd-���s�^C��0�D؉�N�����#�nC�ɕm)ʌ��[9�n����<�dC�Il��С�DEB��xr��e~B䉯ie@416�ٺ-���t�Ρ?�DB��)W�$�r@߅~�����ό�L-�C�F��|�'&
"Od��X�˩q!�C�	3g�>���i�仕��xv�C�'99L�Y�IM#7����/��C�%��5��x!�a�2��C��B�\�s&�2rE��Q����7MtC�I�e/"��@�ɐиB,��{�PC�ɜ���	W"��;P��6�AA΂B�	�{�XQbEX�
; �A�A(B�	�yob�B���,q�T`U�{1VB�I�N�J ���hi�"�?�
B�	+?C���B��6�Lů�:dq�B�ɛ
�XYP�)Cd>$jp����B�I�U����� Px)^���@�8�B�	`�x�h��R�r)�S��Fy�B�I$m��Yz6�Z.f$��p@$�`"�B�	
J9�mb�0�,p9T��R�Ν�d�56/����ѭb+.�R櫑�2���(A�!�$պ]���5���z��!o2!�d�(����5+�%H��8��/y!�� f�sf�K�N����GQ�=�軓"OD�
"O�\��1ȣ�6t���� "O,M#��C��&�Ch�����"O�=��K!^TXhSe*��b�\�c"O�4��(�07�$�@�'�i�0��"On�۔!^<�hQ��ϰ6��h@%"O飵��q�U�a�(B���� "Od<Y� T&	��T�c	!n��2�"O�]:�8e{�)y�L��0V"O��z��$b%�X���	(8��pi�"O0!���Sn��1*�&�h���"O�a�Ə��s���ڵ�9)�n��E"O<�s�U. v���E*U��i�#"O�U)NHцA`ň6U���"O�|�@*S=.F����a��"O�@�Vċ+@�ͫ�G2r��"O��g 2�к'�L�q�A)�'��!�`W3T�>-S !�?p���b�'� �,V��|�9v�G�r�N�k�'T���ȕ,�04R& ��"Fj�C�'���SfF [�`�j��X4�vi2�'4f4�SNO�Y�V�ti�
ީ�'�D��u��*,�����PqfZ�A�'�����P U��ii��`i�U��'/D�b����J��wj�6\rШ�
�'/8�31���9���'��%]0}�	�'b���2��,�@$P)Z�K�h���'�|���@;O�h��H�'s����
�'ǎM0�B�,������w�rd#�'�m!$&�>ɧh������5)6E���J|�P�@R"O6M1��JDBō)�X�۴����ĭ�VT� ��'��#�^�J^(�0���P|�S�P~�kv!��Q�P-�S` &+��� �Z�_���B��U�xL�CTH�Q��>iw*D{u�#�hO����W�p4@�:��>�|iS��1�)k1�ߊX�VC�I;r3�D�,(t��X��Z({��D-���r��FN��S�Oh�}h���"q�q��l�v�v���"O�$�D�\�C�&����P�Z�I_����,yv^=;�|�P9m�3-�ڤ�W�f���?�Ob��4e�uܾ18&�ܹk0�x���av�+4%�`�C�	�e&����^��dSA��*W��=�������@c���O`�Г���p�r�$2��' �|	C@LŜ�a�Dׯ��I��0�	�$,	�N~�")O?��dJM6*v���Ҫ��z�.�K�'�D�<)��#Ӿ�B��#.���c��z~2�F�EY������}8� 
 M�6"��,�4n̨m�n��P�=�O0\q�h 4|��dks#ܞh3<��\�SPh��Q�-$��ա��N�,�1��-GV �#P9D�p r	�$	j��ࠌ�u�H�cA6D�@r�Ш:��)� T�h`�,��� D�<�/\?�~���U9*4���k<D�$9�'X,9���,Ӹ(Hı��=D��X�-��r����kP�:C�E�R$:D�T;�H�!~	�1R��unv�#1d&D������B�<�X�LZ�"�T9�aF'D���%�����a�qØ�6�&Y)��3D�0�G(�7R�؁����`$|����2D�t�ªX��	r-1~ޔ�a&�%D��2�2^���6iL��c�"D� 9r�HT�xKş�Y��a�U!D�LC����˅h1N�v	�c?D��f�.��9� ���N!�ъ.D�,(�K�$]�a9����`%*A�8D�0��kU�6n>ɋE���BMP!%z�z���捧������� &@p1�<�Ȉ{bfӶo��� "O�;�	�"oY���6�\
��`�p1O�$��Hm��m���lݰ����A�F�
�p���ɼ;�؄z�W%ѲQg<k<���^�0ߨMX�m�7t���wji�P� p���2��I8/qO^S����/0�Q0Ri �ӻ�DyR�Ȃ��\��ĳ�VB��-��;a��!�ǡ=�x���a	;�&iQ����?�C'�gy��<*�������uI�3�˥�y��ܶS �HS�
mbµ�.�/9�iu H5w� �V�*/�r}ᒃ�Q��'_����eG��u�jR�2�����MA�@aT"LOPEhS��$K����½S��A�C�|�|�����2��hQ���6ԝ�wI���t�x�pW�?ʓ;<��I7��K* ie�!\���'�yU�K�_����s��p;�A���B�U�� �u+��|��Z*>��Y ��̘
ʈ("Ly����C�\3�̈��	�:@�Y� �_��h �4�� %��`���-@i>0$a��f5 �!�ޟx1J#I"K��wM��"��u-��I�W�5�1�74��!���"�ޕ*fH`�iߡ&.�3��L��iْ�Gr��!��S�F�Ԭ�@*�����O���)*���*6>�۶OU�q%��������y�/U-s"���5�I���"㡓�>��S膌3���Ғ$�
_�zԣ���~�$�L�N�,R�#<�� ۜ)i��W���� \e�I�V��А�@]&�P�X�XͪPE��h�|2�%��>�*q*�D˃tR����`�?c\X�)�I�4��I�Pb���jۢL�Խ�@�?���@�F��X�������B$���OX�Sf���&C��!"��Ez��.]�55�U(�gv��1Uo�/���k�T�`�\�}EZ��5!J�UDq�iՈv֙����/Y��[� �h�Z� AG��̢p����T�ĊGOΊ	��`
�U���3��E�azeЫH�r��!�[�I4`Z��B�/vb0R�lA3����,��*���'G!�0�'Fl�P�
��Q� ���_Ռ�rMB� �(4�b%�	�!�  �wb2Z�
��M�8"�*�1B)���ɐ""p����@�w)�ٔ�O�uZ�^2���I�eLl�:�"�T4�J �[�4s�)p/��hU��&
]�e@r�O���;(H��B"�ӈ?14�{&LD-�<��U�.|c��I�PC�	qRc�7V��S��d���#u$Y&4"q�A��x�'^�kįۣ����s���Q��Q�
�Xy��u��6H_�<��螖&�>��.��R�p�Ò@M���C�	�"kV@`�*{D���2
��U��#<���^�;FР���5�'qfF�h��D�O�UCQ�8)@���s�ŪA��%5Ƒ��W�nl��n�7X4�U�����O��"7���=N��"� >2��
�'E�
��Z
_'���M$[2]�	�'���
�=1�
��)î:��A	�'�ʔ���H<}�25�p�� .�z	�'�0y���L���o�'T}3�'�T�K!� 
5j�q��վ2r��'��hsd��u��B�,}�	���"D�PY�`��H�R]����N̩� -D��O�m?����+�<��Q��+D���0kJ"yQNp��]>B̜̙pi#D��Y�n��B��4a��; �Z�Z�?D�*rA��k�
4b��@�~GN�ؔI(D����I�,F�M� �ۋ[*>|�� *D��ۥ&J
,Y�%D�gz��!��<D��pb�ݞht�i�Bǟ�@��5�1N?D�ɑ	Ќ��@K�<P�1#l��㞜�<d�LBh����qYda���n�<Q�	���ЕAӂ>�m���أU�(�� �߉��>�cn�KrU�D�� 07�1F��gx�P�KG�30� !V\�,�p�@�3TU���*~��a1D��E���4R�8zA�W�,�b18�c*��W�/�vh���ȟ�@Eg��;'��z��Y�X�"O�M�tH"/�Yأ(7	��|yp#�N��)�OX��R`'�3}�J��dn�m*��M��itg����x�l��Ag)�G�F�9�$��g����"�BF�͈�M.�O�	sQ��>��MB�kL����' ����C�nK���<OV��b圼��i'MyM��CF"O@ҵ+ң9BldR#��/"�s��|*T.( �#V� _�?�R�.mU�����
E94���4D�� X��3��n,�\�G�T3��j�Ʉ*?�<L��R���#j�g�g��ɣ� iZ$���ԠK4�˚�!��A�1"4���<�
�#犉�uw��1d �E_���'��=��G�~UH4����:��8�����(-;��I�EG�i�J�,�Ā��M,%�B��0|iĜ��!�[���3�K;����9���LU��k��00�!�BK��T���k�.��B�ɘ@t"��df����W
j�b�1d��&#���'���D�,O���TD]�u�zu3���M��@�1"OԘ�AذP�����	1cav�#�i�:3F*�s>�|�DB#]��X7'��$�c��4��=����28���d!���ghƥ	ap�"��+�ܴ�ȓ6#�� P��}T��3��X4�L�ȓ}�lip&�u%����KI?✇�yq>�	�΁-k7��7������p�W��0�k���+��Մȓi��ۇ&#<�&i��Q�:6Ԅ�w6l�
�E��Abb�ŉK��ȓU����TG�l�Ҝ�2��L6D���v%Q�����w�N�fĉ�ȓ~T��NM��1�F�GfD�ȓW�v�b��9��a�`��<T\��ȓy^P��	�f҆��.
&S�Z	������Lw�������Y�ȓ>A�7
ĵ?�u�VO�>o��!�'��|�s��^HVFQ� ��'���V�*(/ ���NP��@�'D*` $=�
�!��>Bpr�k�'��4���ʧ
�@� �΀1j���'������%�.�˔aU$1�Fi��']ưc.@��a�[;ϒ���'�|���ĕrC@�&�ws���'�>�Q��k�ȴy�I�o&n%��'hb�p�f�s��㶡��3�dM�	�'{4	�/r9�$��K��x�v��	�'5Pa ��B/K�����O^-&J\���'�ti+���#;@��@�i�	ʎd��'�B1��BǢ1�hm*'��=[����'�L@�q ֋~��P����<s�X��#��2#j�����Lw�)�ȓ]��|)WEY�|�v8b��s�Z��ȓv������5a�@�&ռ|�葇ȓH�<��G��
s�1v�ӑ��݇ȓ��EELC�.��{6E zs���ȓC�:ݱVG΅R,Y�&CF6�P��m�`��O5>h���X�gY@)��\�L�z�#�>ҁ��f�7'$��ȓnU £E�3q�|����<&ąȓ#`�(����y�����䎴}:`�ȓ�B��Bʮ^&|�f�ݴ�,e�ȓ{�@�t�ّR��t�75m���UR���e"�3T�&Yps��zp|�ȓD�X�Dk��^Y���@�L���f��)BO>H^�)2�ɿe�ۆȓ���iSG�d�*a�3��?5j��ȓt��5C�薁jpܨ��O��6\p��&�6�k�u��T���b����oP�bІ�4F�0������ȓc5#���HE�-{R(£X#XE��VɾP��oC�[N|�����]��ȓv���C���" ��U��@ݡ\Zh���{ڠ��L�KNQ�Teݣ(V��ȓcdy@�k��a�΄�D"��LaH�ȓr�ZE�d��	FP�q3d� k�����S�? ��
�/s��XY��t>�t��"Ox�!t�6n "�̉*.�kb"Or��vŋ$~�ᖋ�>x�.0�"OBT��i��C%�Q�O�>�'ep��JS5�N�Ӡ�]w�	�'����Nʎf!��1Cb��JP $��')�Г�ʆ{�D��!AY��'���`@MY^�������;�B�:�'qR����Ɂ��P�$�g|4��'��݉�, �IF��r��!^	T�@�'	$\��_�6>Fz'
֍e�4��'� ��4⊪Eu���@-]�@Y�'�F����ۂ�QQk�=P�����'S��Rg��S������!?r@b�'�(��J(U����u��E�'��a�)�d;�8����n���'�L��$�M�R�4Y�s�Lv"QJ�'v���"�`�,�±�V�L�ZT)�'�����v��D���۶
p8���'q4���V6.�D1V
Ԏ m� 9	�'m�he�_�S�ll
��G x��x#�'��4�c��n09B'+A�p���'��Zc�	�-?�YY��$�8
�'�8��*rD(k�J�%lF�
�'R��BR�;48���7`�	�'�RUY���o��]x�l�-�*�y
�'��t���$4,2�q#*<�0�
�'�R�p�A��*k`��?3���'<�X:��Vh�dׯK�2�M�
�'�`���K<I?8a `x��1	�'!4�R!O/��xC��+}
N��'4��B��V��-��(��D{�'ƨ0vܲ ������O371@�@�'���eG7T}ɧh�����A�u�<d�+M2L�b��'p��B��Q�e�����L!�6Ԋ�O��G�e�Ǔ,�TB��������*G�~yن�	�|���o��k�8`A�%��
UCT������L<@+�|,\�b�� _5F�2��M`�'��J�C�ݸ����V�PTC��ݰ$����$W��!�D�Y�YX����zm�4(�}t�[�0!V���7K��)�'	Otq#+�f�d�h��4E�r���'����Ŝ�o�4�����j\t�+O�e�r$��\y�Y�%�/ON��UlAjG�@�!H@+��'#B\{e�	^�2Q�Cc㼘�@ꐼK,jq�� �'!�D�!bی�P¡^�Y��p��g�!�ў�r�Y4f'�X���ḩ3L�S#.ӹo� �R�F��tx�ȓP؜s�%C`��b`���j�O̱���±r�~)���<E�t�\I�!땆x��&�`�!򤗝~�T|s#�ŊAf
�3�Bޖ:{�	��� z7��,t�x�	l�}��	Q�A����Z��p?�6㆐V$�Q�"�N��Y��#@0x���㨑���x��C7��A�T�SR@)��S��y��G-&>�ԛc�B�j�����]��y"$D+w��a����p�Y�/��yr�L�v�{���
'��@���y+���L��%�kV��y��ˀc3�	*3�5��В ́��yԍa5���cޒ/�T	�Z�yB�	j��9���~�+�$е�y2>�@�)fŘ(vn�Ѓ���.�y���@;����f�.w�,�a�A���yR��!!��K�h0
��fm+�y��V�B�˕N�.j` �Ônˎ�yk�;D�&�Y�f��v��sd�y
� �T8�*���4|#$�&kj@h�"O`�T́D�ȱyP�y��x&"O��V+�v���� �[�g�x�U"O  `��OȘ�1��73W���P"O|�ї�Z)����[1��d�"O�m
�MѠg�(�䈐�~���Q�"O>I	�;�j�{Qƙ�4r�Uc�"OС&A�� B�� $K�.E���"Ot��%Sk+��3��%�$,��"O��Ǜd�~I�����+tݛ�"O�q��#R o�
�[!�H(_�}J1"O�ᒀ(�"ݼq�҈��S�옉R"O�r2��$����0����x�to�+&a���O����>�(���7HH�� ݆N�Hˑ� fk�C�I��& (���9ۼM����[��� !�B��]�H\w�" ��Ɏ���b�)�""DJ9����2W}(����P�5��l՟�yr ��aZZ<�拫J�*ё�Lŀs �0�E�g����O����ђ%~�ł
.\�f�<���/X�r,�tlY[?9���-^d�
vcx>� ��ʴ�Ϊ&�N%�qB7D������'w�ौ��9�TH�����@"Ǭ� h��G���d��t��A���B%��Ż��7)L0���ѡ�$Q��ެ�g�8t����R�~b��h .͊zz�{GH���;�,D�weB����I�IĂ��4IJ��t<!婒�|`L��
5�lA%)+eH��&�)B^	wf(�6��2CI�Z��$A��E�1a|2&� 4\�Dbؒ5�A��$���4�i����Yk�`�'�����O��#���'qx���W�0=c�%��(��ąȓt�ʄ���9j��ܲ���N�ZH*�덹o8����]�y�"ӻYg����a�u�s�a��#��A �M�n�@dQu�*4��z�"��M���[�i7Y�d!� �]�7/��{�I�<a7d���"ͣ�򤎍h�p$�҆֍m�4ձ��KP�y�Ɩ�n�:Ɂ��S}��! ���aT�[;�si��?	��G�����8C�K�NUj�6X�׭ړM1O4P����O ~�FښOO���  E�j�a�H�E�<AQ�P�E4<�qC,讀�%]'
��=Ѳ�&�gy��4���#֨�+Zz��v�-�y�剒>�:@��ٶ#Oz�@FKղ�yR��p
<c�_��A��J*�yB#�0+�P
0#�z��EC��yB�ڬ/ֱcT��O\���W��yB�OQ�� ���@����u���yBH32��	��\+��K�[�y�є@��U���# �������y�
H4� -�IÄ$m�|�����y$�M�X�ԩ��GFy�P矉�y� ӊ0�.5��!\�Xh�QSI@��y�#�C�d\�G�_P56��R��:�y��9:��ej3	_YV�{UÕ��y2��X4�s�(ѰY�|��tO��y©M
Si:E�/��|�g �9�y��T�V��u�/���1��т�y���E{�"�a��xhCg���y"��]%���G sN��J6C�y�'x�F�qu�	j꜀���"�y��Bvh򂇟�k�Ċ�IÕ�y�힂Kv���bw(*HS�#!d��!��{ːr���L�����^9|�"h �!L�x�!�цIMjY�ģ��\�t T7iXe���4L>���d�C�"y�f;cN��M4<��y�&F:`@���Yt}�AO4x��IC��c�կ�y��Na����DE��*��ѹ��_:��+����b�^8B��"j2�LѺ䢰���B��qg^_�<����0��2��K �d��5JP1>D,]#Ӟ>9�������	����4dY�v�j<�6l�?>HC�	���F�I�;[��8Feڒ+�eB@`˳h�����E;�O� �m`��D5d1��2B�Ĭ>��M#�'3��b�ů;��Y39O�i!�D��)�}��8�(�JU"Ot0�!$Y�<=h8:qd�<n���cӒ|R�S=j���3sB��@?u"��Y�p�ΝI���;�Z0�<D��X���.p��ѐ�A
T�遊���:w�<i0�'����	���AC��a��\��_�4�8C�ɯ]A�B Kش3�z@H�k0T��E��#��ec�'�O�XS���y�h���Q�dQ���'=j����U&\S4)�K8�$�T�5u���#��Lq���t�JA��@�p��q�u!I�-�z)�=����D� �J"�'=� lbT.�?
�ƴ����83��ŅȓLtP�"�]�$�P��q�֮KTٰ��/g�ѦO(���Y���Z5$ƊU��!�r�&�
$+D���6�ܿ/�AU��(�ʔ�u�k�$��'AE6�h��D��@��E��YR��;�&E�(�{2�ؼBjV@�'�!�e�)�8��&V���\[	�'���b�'I��A���O0�	�')��#�) D��J��Y#	"����'�ƌ��GK |%��aD�&��{
�'4\��#�����d�r6��	�'vn�Q��ŗ!Jlڣ/`�.���'�^���Y�@�rT�Ue�<�a�'?��"j��
�
|����_H�M��'�p�hvś6 4�E�_�J)+�'8�0�`HbNV�J���_Zj���'��@8f�0C�:pZ�`��R=��')�zcM�2�*��1�ވz\���'��a��w�I��ND�i�� ��'[XHQ)Y�C�2Q��X�`�x�[�'��%��!�tH�m��N�a] �`�'U��9s���i��4]����'�pE(�c׮�"�a&���t��'y�݉���l�`f��)$���
�'pt9��ԓHu��Bu$��
��H`�'�Rh��́)�34� . T$��'��!@&�U�i�r�[����w�^ܡ�'m� ��L���s�X�U��(��'$�1�d�T�>/Xx�	��&�
���'U(C��0]�Ε�ӌ˩HJD�H
�'s��1�G/fy��#�kɒt���1
�'��s�	�F� ��*�o+����'dn��F�(3D� "�aب^�p#�')r)�s�
Ԗ�bSNҖ���)�'6Z��0.eg��������'R�)�v-�ckJ��D�E��!��'��ͪ�R�/���aaȷJ�j���'��D�v�2pL���胛�с
�'�J=���۳�H0��@��
�'�����Q$4J� T�v{bY��'7^���$-[%��x!�m��)�'��1��D�R�6Й� W;12��Z�'5DA22K�0AI��q�hǧ5�)�	�'2�@���9��=�UkǶ?�d���'��E�3�ĽEQ��)V�}r� ��'p����)͂$9>x��[t����'�v��Q��A/,�ǅD&���;�'y �b�$K�%��ޘ�	�'��CW���d�"ݪ���|�Ќ��'�N�v'��ab�K��c�$�`�'�R���&֊�X�1�C�_��xQ�'�H�Sc�>��y��D_Ȓ��'C�i���J�4H�`[D7x\��'��銧�)g, �r�ڀ.�İ��'���R�Q&lu$"c�҇'�4���� �qx�o�R�h�h��4$�D2"O�X׀ˠ	8���1�����"O�9i&��q����G��iA@l�2"O
} �������SdN�i�~�zw"O��@Q蒘D��A&��Lw:驐L��0�1$�'Uдs6��F��eR!�3�.܂	�'����G!�
�0���+�����'�T�qm��#���sqF�6�R�B�'z���䬞
' .����:8��ݰ�'$N��fz���E�D�6�^ղ�'��J&/K�ݪu�J�c(1
�'_�
�N���d����%�������y"��1�l�x�/�6O`�@{A�.��	,m����梚���S������_d9�x� ��~}��(� $�qg�3��S�	#}rA� �N�;�Ȇ$
�TL��̟�W��ɔ83�nL&��zN	,C쪸����!�t�F�''���:Ԏ*�̀�0|*g�Y�=�rlA�7#�y%	S:r7�OD��6jR&�0|�J�u����M��n��!���t��ۆe��m�S(��0|�!��sI��à�� �Jٰ�c�Y?AEޘt�E��m~���X����Q� շ!Ęm�
�*ň�3AʛuRy�4���)�'0bT�Z̈́؂HA�'F���y3f�)e�N��T}�;�iJ�>0��'|��C���9>�Q3�ʹ+�$�'M������z��H�r�2��cO�O=��i��ˌ!�a�րQ�gT|���O(���A#Ϊ�O>yC��.l ���PC��}���R`�a�����84�c��>-8��'�`�j@B�&w|�ʞ�@6@�/V+%6hz��O��I2��H�O B��ʟ v��L��>���?�?ig�P��?A@ϓ��0|"v��~�BI���K.��{H�bƸ���ğ���
{y�O>e�wɍ+X$��g�(�(`/6D�l���5d�:t�ag	���j� 5D�8kB��&cy���QS=z�S"�(D�����>�^՘�#p�HT�$D�����U5�"4����o4��#D���j�2�8q��hR@r�����=D�|�F�0h�r$i�*�_��<cc�=D�P�#b�>/{h��TO�_f,���<D����ʸ9��H*=zP��7D��BD.�7%�I"$�4E@2X�j6D����톶!�zp�Ai�;}J���)3D����1�őB� X��0D��3t �!�%��e��K��� M�!�	[|��� A@�V�X9f%�*d�!��>�d���B������C�!�V�:�3.	�w��+�b��@�!�_#9��m����&Z�ع�̃�VT!�K-X��b�@&U̴0b%M6!�$
��0�K�I^�9��E���!�d��n��-���)5ɈEkO� �!�dܷb�$�Uf��5�֬�v I6�!򤑇_/u�a��7Z��qr�R(j�!�ב0&&�2�'ڑ&�����9z�!�C�4nP�A 	?I�|��#�0gz!�d3s�<(H�\�K~µ�p��h!��6aYԱ����J�;p@�V�!�L%��4j�%�P�|鱴H]�l�!�d�34��4*%ҸkU�T���?b�!���.$6 �BD�]`Ҩ�7�G� �!�DϽ�V�K2̍ bNY�!�!��M(M?�0��؊#[�d�S�͜/�!��i JsWBB�oV���F���|�!�$���H��Ǆ!vb��A� o�!��J�fA����!�Qa�YIBJK0�!�ą�,�@�CdN�bp偰h�#�!��ڶd��J�+��ݡ�d�,?�!�d�O:U�f��3d�����TD�!�� H�X��W�uW�qi	�FH� "O�ܹu�����C	U,Ur��"O�}���_$aQY�(6D�B��"O�(�&��G�B��u�gz�}"�"O���G7eH1�hʯB�`(IV"O��Y���'�R@HP0[�p��"O.,��e
�w�p\լ��rʲ�"O���$B5.��u��kG,z�j:c"OH��ì�dӲ8R�7|����"O�U��
A5��19t)D���"O@�+�bV��M��1)��t�b"O����$T�F�k�NYA�" �"O��G$Ka�pА-��_��`{�"O6��eJ�&&NH�DL��}P�"O0�qʉ#[8E����0;�t���"O��K��0Uc���Q��s�"OH� c�I���5�p�������"O,lKDE|����Bn�!��Q��yKͫU�<� ����Z��S���y�m�4@�i�i@����Ҥ��y��*>O��kS��$T�u�q	�y�%^�s.�)g���M)��#��ybMM ��+�Ȋn} �� P!�y����~p"�gԑh��=C$���y�1s�1�¥�lQְscbߨ�yR�E�DT:���_v��#+�
�y�G�	`����j�vmpdM4�y�P �FN,g�l9Kѻ?>j�'�n��@k���R�*�41��z�'�`����l��j�k@/@G�	�	�'���
��P;@�R�c�3���c	�'TB�"-�I�b�;���'>�+	�'sN5�a�B)Mg�X���Em�:���'��E��J��g�N������1�'�W�yo6��5gE�z���
�'�F�%@ء�Ni�t�[�o-f��
�'dd�1B�I���&��`��MA�'E �+��@�cf�$P�I5\��E�'�d5�rM�,��_�_�r��
�'�����L�
�4��?(�P���'2�x
��Ii���ЯP�����'T Uæ*��>�H�xsa�-;J����'���h��`��A�e�l}�
�'��0�G�D�w�ְ�2���YZ�=C
�'�Z��Tpݰ���g(M�2B�I0�<�H�a��nt��7̚C��C䉋}^�YA���C�^dȓÙ�W�C�Ɍ����l�U�R����ZX֢B�ɔDr6�SP��|~eRe�Y�+zB�� R��a�N�%�`�8�(�\B��4|�ؔ��<�Bi���U4B�I+�(ـc���&�	b$|u�C�&d����99h"�hS/R�j��C��+pn���!#
U� �ө�t�nB�	�>j^0y'�L��1�W�1C��C�I�"H�%�)@�2n��Fj��m�C�	���J4A�����Y�鏬!��B�	�6'\�Qb/� /��� �#NP�B�I�IL0܃P�:2ֈS��]ǮB�G� ���P�^��#�B�I-��Pf"�8_h\E�@iܛ@�~B�	�TZ��S��
�~)�2��$#�lB�	,�@!qf��S���)��[E>B�ɕS���Y5IA�f�֕�Ѝ��D�zC�)� ���`b�67s P�ւцw���"O��w�M�Vq"\aq��}YnP�#"O�i�֩G��4E�!�ʧ.�y�'"O�}�1��=8�X�aR�)n�Yg"O~�b�AۗtA&������]��Y�"Oȥ�����P�� j�/̧k�|8��"O��qנ��e
+X�5yb"O��KׁÜJ(��уפ5O��F"O~UHE�/W�8�r:m?J�"0"O��h�럲��{�F�|!���A"O:y���Y�v�S�,ɄA�9"d"O�y"��яJI� ��B�1��-ã"OB���$W��Q1Vgݰ0�ґ��"O꜈��6{L]��Q� �|� �"O^�1F��qX�+�o�/UT��۵"O�y[�!H8:	�p*��285��a�"O�AZ�A*>-�(�Aۚ�th�v"O(k��A�Aؼ�c����Q�H(0�"O�9��nR�l ��� Wl��ec1"O�|IT�
��ҁ*��սP���R"O<i�!�=T�Q��}�E+"O��P���%/9��@Z����"Oj�����#��A�O�J�p�Ӡ"O�jO='^q�/��*�n57"O�P2 ɞ�NM�怅�t�dAe"O	Y�g���sf���\�-z�"O�xr�:`���H���"O�pxN�7d�:�+$���.z��2W"O�50m�6L�e�gHFO�4�"O���o�F=�a{ Gmb��؅"OX�2��E�\m�}+�D��E�g"O�0$�K=x-�4D]�C��Icq"O���DĲS�����ř|�d�J4"O��Í�=]��D��b�rċ�"OJ��(	7^&��AcDU ���"O2���97����ְl,���"O�h`c��#��p���'���s�"OzMh ��J#���^ O��J�"O���t9<���K �D�X�;"Oj!��i�̜�(�2m����<D��Z��׾X��9Csn�, �Xa��':D�Ȃ�͵rH�yr�ة,>Ix1 9D�P�掍4̪a�7=�zX�rB:D��"�b�`@Q%C�v�p(yQ�*D��Sb%�<G�2�K��F�,��gb4D�4����+i������ӄQ.D�;�1D��#u�>���i02L�<H��#D�D�f�ʈk�[�v����=D��K���]�NPR�1�찳K9D���'��7D�fGVa���qE7D������=��U���Ha���g�2D�L��Ȉ�,��Eŉ�L���kR�0D�h���7S�(� f
otl��+D�LC��8�8�(��G�h0�5c-D�`����~2�h��Jff��KcN7D��n�!_��-�P��w�Y$�2D�TSP�!_��r�E.)+�0cF5D����B?M�����2!)t�x$�2D�d(A`P� <�m��A�:M,H�r�0D�8`�+�|� &��1��* !D��������
�f�,;���Q�)D���4mI�08�J���w ْ4F2D�x��oӊ@U�]1a��7����$�1D�Pe��-N�)X�^6<�Lx�D):D�� Pc +X�x� �K"�>@��"O�dGo��*�8H�'�E���KP"O�Y8���	�h�b���.xh��9�"O��	GDA)6���Q�'X-А"O.$)F��So���"�CZ���"O.@�R+VSf<e�Q5uo�A�"O��h�iI,�b���b�Hd���G"Oz���&VF���C�)c$�}�1"O.�#�)��A�(��C��C�^��"O�X���x)��5`J�q�%"O��p`�Z,Z��䁔}иq�"O�ı��CH0|ir![�-q�|��"O�q�cC�
��l1t%�]�)�2"O�,��Gةg�,��'Dϥp\$Q۷"O��ڂ�ֿ#bxt�� ��!v�QY�"OzmᠫZ&D���"*����r�"O�5�HK;�*�"U�U=�0T"OL�'"��>��U�Α�NQ1�"O�a�r/�2�X�L�<|��a�e"OdL{3nR!�Zl9�ᓸ|� <"B"O�RV✞Z�*�F#E؂� �"O:�z�hԙ:r��3DiK�\I9�"O�Q�?�U��
%v��9v"O�T�$ꋐu&FM���H��(��"O0���$D63���P��v���"O6ȑ�i�.0f����
�N�Zt"O<�
�!C�w���AQB�� ���u"O`Pq�cؽ)���' ڍ>w����"O�A{�$ߣR�H9��H)ڐ"O�i�c �"w�iY�W�Vy��1"O���	M�U�p��T�	,g����w"Or�@��F0J��3�jY�p�"O�8�dG�K��!�IǦJ�"A1�"O�q��D@�Se玛=�����"O�\3   ��   �  q  �  �  �*  F6  �A  �L  iX  3d  ho  �z  ��  ��  w�  ��  ݤ  !�  y�  �  &�  h�  ��  �  p�  ��  j�  ��  w�  ��  A�  � �
 S / � �% �/ b6 G= LF �M �S %Z i` Wa  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�?O�=E�t��A�t,1��;Sb.�{c�;�y� �_$*�#�]�K� ��e ���y2��#/��Ļ`��'@0��OT5а<����A6�^]7灦m�H�Y2�'m�!�$��6�yA4L	*���Э�y��Od�GzJ|
r ��+6� T&Ǯ#�挡GnOs�<Q��^�V�ґ��Ó�w�HȉuL�1u�qO��
�S�g�$��x�૒�
_"�=��J.@_��d��jD�e�䩐/L�6t���W����t؟)6f%0 �"�B93�J�##�$D�T ���9i�rea�8�,�pR(D�D�a�[G~L����6.���&�$�hO�ӡ�v@��C�K@��E勺!��B��eS&s#Hۦ%BMS�cH<e�B��5�����r~h,(�kF��8C�	�����TIәG#�����c���� �i�aR��:<�b�fC¯�� �`"۰=�7��<U��Kƿ}���a���Py2K��,�b�cǅR(:3��O���'ўb>��S��!���1ĄM<P�C�./D�$�ǈ�.�@�� �K�,��,D�� �Б0#+W",3�T��U��"OTmP"*K-j;LU:�#
<B�q"�QVH<9!H�?�")�"��fx�͘�%F�<�0/հ���u���Q���D�<a@/�O<�h3���%L|0pRg�A�<Sꘟ(C���	�7|�E�7�R�<���ؼ1�&D�3�׍�业0�4D� r�;XC�j�Jٮv��	Gj5D���g�� u{p��"�I?$�\���4D�`�u�&.+ �1&���{���
�4D����#ۉ9Jl���D�^��cu?D�8��Ζ�R�-0 JY�r�@"D��v�ܵ&�vs��&7�V`�4"D���$�ε(L��ފm������ D�H�p,^0Iw�u�!H�^���FC3D����m�[tZ�3#E�u�<�c�0D��37�N �r8�Wh�� n2W�0D��QE������	P&Y���E/D�d3���,T������7�����9D��9�ښB`@��@n�'Դ��%3D��0qDu!��V)Pj!#H>D��#P	)��ႆE
��p,?D�����81
D�Y��ɍ`)��CJ;D��Õ�ؤL:��9�6D9l-!!,D���,-A˚� ��e6�w�6D��(�o��݉&�Մr����ă(D��f�ͼ'T��ql�����@�8D���ƉԘJ(́�b�"Rʹ����7D��%oVTn�����3��-#2c4D��b�(Ώ-|�0��W�^�ЭIe�3D���U��`��ꅋ��"3�%�vc1D�<��RPf��g�ƋB�m�%�0D� ��MK�j�.}1�Ŕ�f�Y��4D�d;��X�l
��A��{�l5D�:��̀S�vͪ�bʝ@R��V�=D�d	�*�q98%!4�F�
˰��7�;D� r��5���P����Dl��6D���۬U�R����� �|k��6D���(A'�h��T�t����23D��t�'u���0�߃ :���-+D���g�XM
� ��]*;%d��C*D��(�G
 ^�FX�2&\�\n��+D���c���9�,�i�gY��Ɉd�(D�`��(��a� V�bg�Y�V/"D���4g�'ap�)�㟛K���RGG;D�ܠ1��z���e�S�9� !G�7D�(:��R4��O�4��s8D� B�ܖks���4f��[̦�*%�4D�HB"�8Y�Tu��b��o���V�.D�����(���"l�D����.D�dYbhˏM��` �͉hK����-D�$PV�@�V*db�/�^Yd\rI1D�ʡ�"6ҹ;R��!�z�R�3D����l�Aul�#dDm,��21
0D���Ug�T�������>��-D����B�,$�4�a�ܶ>{�0�k+D�H*W!�-� 8��M!O�r4��
*D��3t�γ)�v�[�&ϰ�Fx�e�<D�TY��^3V��a���xd"%F'D�a
��^#XU�FG�ٲs��8D�|"F�Ǆpp�a{C捎+��t�4�1D���2�T���c,���ܳ��3D��2��V��x�;ϢA�w�1D��$ϊ10�T�Ҧ#�l�p%2T�/D�� �Ӥ�#�L�{���\�<���"OPe���}� ��]���+�"O���O��~IRF�/wD��A"O�������y�ޤB"���T����"O$9��Έ9��@�KN�k��:��'r�'���'�r�'D2�'f��'���B�Nom����&Ђ*Q^1�%�'��'�b�'N��'{B�'�2�'qj�[�C�#J���!Q1~�r ���'��'#b�'m"�'���'��'	��5#P(���,� 2]8aP�',b�'���'r��'c��'W��'"f, �^�������S��zw�'b�'v��'��'m��'���'CZͰ�.�]T�C���T\(+D�'�"�'O�'#2�'	"�'��'����.�26��)��(RW���u�'�r�'"�'0R�'���']��'��u�"@��VY,�yg�� ���)��'B�'�B�'���'O�'���'v%���%H\j��M�-������'6�'2�'8�'Z��'���'p����dϞ\�2X���e�2$���'��'o"�'���'{"�'��'�(y�P[�(
��4#�$���'Qb�'EB�'�B�'m��'�R�'_�}�CKW�}%&1b�iY�r�<P��'���'���'���'3��'�r�'��a{r�VnÄ�'��,X<��U�'8��'	��'���'}��l�����O��r�=:ޅ�uB�!���kA�~y�'��)�3?镱i�y���;Lμq!�
�����#�¢��D�ܦ��?��<��aT����F��O���i��zt~����?�$��M�O�瓿��N?�B%\�����J0��mj��*�	�h�'�>-;���+`����G�` ��B� ɣ�M�'KP���O76=�|��R���ˊ4�FC�8-�d�!���O�j��ק�O����W�i��$��i�d�R�!�TR&JɸW&��w��x��e���=�'�?	t oA�%
�|�x`��#S�Ĝ���-���Ŧ����#�Is��|1���9imZ$��ӷ&n�?��T�|���p����?36���`�!.�"�	u���ӟ����N�b>����'�P�I�|���Dg�4��C�
��HЖ'c�I�"~Γ=-�\�ŮƧ �.k@IВ5e@P�}��e����˦��?�'��@f�2n�"i3��ny����?����?� ��M�O���z�8|m��4`�(jƞ �� �`ܒO���|���?����?���Y ��	՗^�B�z�Α=�8�k+O�o�,1��	ڟp�	m�s��PcI�;�X�
��P��H�E�'|�7mQ�Şq�� ���A����f��`IR�"�HV�R5#��iFn *��ȯ�t%�Xw�O|��'�*ـ�ǫ6�(Ѩρ�R�̣D�'���'���5Y�${AX��3ڴ8�$U��'$� �0�I��}�(A���հga J���?�O>�'����E+۴�?���Ň<��(@P�#\�
&K�3_)����4�y�`@�U�dirv����]ǟ�S"Y�Y��}�HAv��?(��V������ԟ,�I՟0��̟��Iu�'B�������2�t��뉠#��,��?q�Z�����:%��;�M�M>)Pə�6�JE�a��r�)��O��?)(O�YJ�Is�4���	h�攀�n�x#��eݞ܋�/�#nD	�J��䓣?�����������## �>���s�,�P�K�M�̴�.����� �ޜUJK	7���	�O��������]�a������3PĪ��ʞ�Q��ޟ<��C����I���KSO}>%�O�B���vl"���}�`��-�
������&�<IF���0q�'�	��yk���0[���!�{S����-4�h*�4Qr��2�i�=�:�[���",�4�P&!(�?���T����Db}��'�������b�VeٓOJ*B�"�9�'�"�o�f����b�Tm�'�����N�*s�ܮ v��Ŭ�0i?�<Q���?����?���?	,����i@�:�z�e��ń���ڦ=S�CƟ�I�&?�I�M�;x�M���+�(1 +��"�ใ��'���|J~zգ4�M�'6��HG�%�]PtGX�d?�h��'�tLXb�Pǟ�If�|2]���I˟��Dϰdʦ�)�"��j��9���֟���ҟ��	Uyb*p�1�i�O���O�4�n���8ї��6���.�I���d�O8�,�V�ơz����s㋸[Bd���<?��'���|�'n���'�����?�a�	,o�ӓ�ΔD��{�����?i���?���?�����O$KBCQ6
#�i⢍�8�$�a�.�O�En�2'��'��7�9�i�Aa���=|+r����e�\�&}�\�ߴR���iB�m)��i���e�\1���Os����T>H�����t�(Mp'bEL�IKy�'���'��'B�\JZ�Z ���B��Sfދ7��9�MS#����?i���?YM~�! �[��Hx���L�P�ƬJ0�J.����O�b>�	��#nZdq7�R(fp�y &�<�2��[Dy���(o�D���oX�'m剺-����GL�.g={[p�1�����쟄�	ݟ��kyR�d���0B��O:8�ϓ(3x��d� 8������O<4mm��JN����MS��'����ܰ&}��A����/��!���{�t�s�i:�	8.��)��Om�A$?��=� ��xE��[,�q�l�p=<����O����O����Ot���O����O�`$k�6({�t����,Q�F&�r���O���O+x�8T��2O����O�O$5AB�,gL�]����`1VU@V�ӦWE�Y���o�PEl��?�s����%͓{���ӄ�/���S�ʉ|L�B3�ָ��aُ<I��0J��iUU���џh��ޟ��˒2ɱw$�	V�J���F�ܟ0��Yy~�t�xw	�O����O��'I/�%�B�L?R.ڠ
+�;�e�'/Z�+:�&��O�O�ө]���w �8Q4��1щ���,�ڕ�H�b��C�Ly�O}F�	E{�': 1�ƘaN|�S�#���҂�'}��'�����O�剐�Mð+I�;�$���E��4Uce�R	o< �+O`�nZi����	�M�r�
&��MRfJ�b4܀Hq�Q�f��i�ـ2�i����D�&+�OdK�<!t��9nZ�]�KR嶬`�c��<�.OZ���Or��O���O"˧vDE���#'�>�j6FOh��5Iյifd�h��'���'��O���v���'gv�QҹP�4`H��B�7���)�)�
V���nZ�<���,[�Z��GN�\Ω����<��ior��D�:����$�OR�C,l�U�$Hf��EǕc�V��5�'���'G[���ܴ*|��?A�Y ��oDv�%�%�e�2i���>���'��Ш�H<0X���u�,���Oz`��lůC��X¥h1��D/A��֝"�?���ƒ�$h`���[HC�n��?���?����?��m	ڕ�.�9�?���?y'�g����#�[�<ǧ���?��i'�$i�'���'�bR�p$'W�G��i&�Cl�2���$;��U�'��<1�4j'��n�����Ki�����@���'py��iv��/}�h0��VI��(Y0J["�J��'k&7��O�d�O��D�O6�D�O�����A@��ձ+�T!r�kϓP���pP]����.���O��l��?�ş8�2eB�>5d�q��~&�c!jHW��)�I��M�u�i�^6���`˧����(�b���៷r�8훂{,-�U�~��h-O򵨵֕�?�0���=�M�-O���r��oߺ�b�Je�	���O<�d�O����O�I�<���i�b�Qr�'��<�6eEKzL1�B3a䚙'�P6�#�	���$�̦���M3Q	6W���#F�9�����2G�b��4��$�
�XX��'@����F�n�A�LX�&�"'ȵ�'�C�g�"���O��d�O����O���O<H*�!�#���+ZK�Iq0���P��`��5{��$�O��d���{Fo�����D&�H�T/�8���@��Xm<��"3a�7
� q�e֟t��4�?�öi���Z��i4�n���`��O�Y�i8��
�4�8������}��\���'��D�'<�7m�<����?���?�٢C�fIq�����Ơ�>�f���O�˓T��"�%E�"�'L�^>���'��/�
TBw��l�5?�R��!޴oR��|ʟ�y+U��_��A1��O:�(��ю��<�@)F�^�n�D@:���e��ם>�ēRO�P��]�w��h�%�� w���0��'E��'{����OC���R��ֶ4�8h����t0q��/�j=��OF��Ǧ��?!�Q�TsشH)\pj	��b��s��'$�����'���f�J_�֖���$�];�D�XyZs+�����\����7���(��ly��' b�'���'&�W>C�ަd�0�q�	�37��)��� �M;6K�?)��?iN~�~&��wE�R�!*���)2T�c�ʑYV�'��O1�n}z�+x�r�ɰ&t�ؠd�T\h�d'K�g^�I�|F�X�'s�`'���'�"�'�mI�
tBLdI� �\�~�)��'��':�\��ش	G ����?1�,�0Ū���x���"�ꇩk4�����>����?9I>ѱ���)K/�\iR "R �<y���Ku`*�M%W����(��d�O�p	/�����9�-ߡ�bZ�h�O|���O|��Oj�}�;)*�m�Q�F�trkЏP
����<m�V�Nj��'�R6.�i�]�"��nƅ&��aP4:sKj���I�4�	vnT�mM~ZwP2S۟$��/Đ4T�ɸC.�z�`�y4�(�d�<9��?q��?���?I��ϦY�Ty����4[�\J5���������C�R�0�	�X&?�	�)��%�J�v��%�R�Gb��)O(���O�O�O�a��C�����Ȩ*�x��b(�+~<�GU���ɋ#Q�Ҡ^G�	cy���
��Uc���1&�l�r�J�<1�'�2�'�O���%�M3fH��?y$R�`���Ye %��H��?)!�i9�O\�'d��'���B�l�S� 4� t���/n�]@�i��I;�(h@�O��&?	���pu�鐃O��2�E�;�~�	ǟ@�I��	���M��d����ԱC1�I�B,��q�<ш���?a��
��v�B�5�	�M�H>!4H-u�2sˆ	!P,�H��@B��'Q���sӎ��(5��6�z�$���A�h!�e��3 ���B���;C���\��+�~�Py��'R��'��4YULuj�C��Tt�C�w��'�	�M�e��,�?����?�)��;�C�6a0�@�W�c���1v���;�O��m�(�?�N<�O��LE�� G�vI�v$J�A�����ML�Q��m��i>-8'�'RJ%�h��ś!|9�$���B�&�ן|��Ɵ��	�b>	�'G
7�^<��q�%�(<���P ]��E{���O���ͦ!�?�tS���޴D,Z�
�a��0p$���T������'{�f�V������ۣC�]t��ANxy
� *��s��7x6�JD/�)f�ʃ9O|��?����?���?!�����P:k.�8ӊZ�H9͊Eg��j\��nڦ.5XA��០�Ia�s�������S�R�&�mڡ��!l��C��	ԛ��OVO1�*(q��w�L�I�UK���6�J���iA�]�Vn��	�l	�t(�'>�q'�l�'�r�'g
,�BD��k���z��-on����'^��'��R�h۴2Pt���?A�x�8I��.Fg�(�`/��e��8��d�>���?�H>A���tn(�"�B�3'�.�XF�J~rjgl�4�3�i�1���Y�'���	6GR��u.C._�"�hf㓧d��'�2�'/��S�p���̾O�X� ԋӍrW�I��CV՟��4\�Ht�'��6�7�i��3ĕ�w��)�1�N�i���d�r�����h�Ir=nW~�i�%g4����"]	�O�:E4dt)#:4laI>1-O�I�O����O���OH @Ц�N�"��#dÃ9�0+c�<�r�i����'aB�'��ynV$5�}(�D��]c����P[�4�	۟�$�b>�bed
+d}x�fn�6a�hǭ-�Xn�s~�M��
�\�������Ϗ,ނ�S��M"T����
 �'?r�'�"����P��z�4o��Xϓ�H=��gN;\��]�$�
�]�Dϓ({���'��'����?���?ir��&�SCշ�����0xن�`ش�y"�'����X�9O�i��>\`�EZ-��{��F�d���:O��D�O��$�OX��Od�?!AHF�x�m��E#J$1�w�u����ğ,��4p����'��79�d���p��-I#X8n��ߚH���O����O�	�6��6M9?����)b�j �F]�Ll���$/
h��`&�������'m��'�Yp�K�.)~5ыU'�t�j��'��Q�(�ߴ)�=��?�����iӈ&ĵ�G�£����@�7��	'��D�O��$=��?Q��ϖbg����k������ӥ��t��#K�E��ԋ�O?�L>���@7hزXc�Eo�0E�"^7�?I��?����?�|z.O�nZF��r�.܅w`��Hǽk�j%xI��X���M����>IӰi��yd@1g��Q
D�d�4��ŋq��nZ�<+�ln�N~b`g� ��SP�i#R,��W%D�
�d}�7�D�W��$�<����?��?���?�)��`�ܑKX�qDӾDD�x���`�`c�`��꟠��y��')j6=�X��,�81|������9�8�pE��O���9�4�����OFTQ`od���I�7�z%�ÉN�:�	q�]�L%��I�W�8���OX�O��|��'aQ"©V>#��	���A���y���?���?�(OHPoZ�XV�ǟP��1}(����9mC�U��i��?�S���	ɟ�&���� 
|���N7��)2�9?!�K(�~AI�4��Ou�����?���eW\���#��!��8�+�$�?���?I��?	����O\[��w����e6��̘���O�\mZxg��Fԛ��4���(�H��
�!3Q�i�E6Or���O����=wQz6m.?�c@i�z�&
p��5!�&@R�Z7j�/W��%�̖��T�'�R�'���'J� 2��9D�~9��=~�xL+P���ߴ�r�C���?����'�?Ti̇G��-
p!MUf������Iş\m���S�S(s�J܃cN5).��YS)/Jc�AH��D-8���\���k���O��N>q(O����,ǆ[��u�t/Z�[ݒ�����O����O����O�i�<�U�i�FlK��'Q����	�}�����ΘX�� �'��6=�I���Gݦ�C�4*Z�&��%���ցe�̜b`"I�d`��i/���$Ipp��O�q���>.G�!�h��;�␠������O����O����O���%��ך��#͈[Ŏ�$$�xj��	ݟ��		�M�6'�|��T���|"�3 �U��ŋ�I�!���֐O�O��o��M�'��M�ߴ����?9@�
�NV!s� x� ��
Fl&H�0c��?��) ��<�'�?i���?vLڮ�F27�E# �Lݩ�I�?q����$ަ*�IKy��'Y��|1�WD��|�. xR��)5d�0��	��M�i�O���u���ю�,��9cU�P�>dd�Y��@6��C�"?�'c)��d���tG�p�v̞;F�҅1���ĸ��?���?	�Ş���æ�z�%˒}	@�a�ʄ$7vJ����O:�8�'�6�$��'����O���IF5@�-:�/I;Y1�����O`�d�!;�6m8?�QFy����dy�N�%N�� �"p�ɘ5�L�y�T�d��П���۟|�I�D�OD��	�e��p�:���k�*SX4� b�n(8 ��Op���O���v�dZ���#���j��ӂ�V(��!ǚ=��ϟP$�b>"��Uڦ�̓��. {|H:��O�H��J(`ᲢG��`'�P�'���'��MY�͚�Y|d��gZa��d���'�r�'PRY���ܴ1f������?!�1E64�5 ����a��g_@�F�
����>�$�ih��/񤎦3��8�Ag���J�/��E�Opx����K�)�"�'����?�"��OV�CS� Z���� �[�F8�;6��O����O���O��}B�P�Ll.��`��m8E�$P7J�#�?���i3�	��'���{�(���.1d<ag��oH�Y��ʕ�5�����to��MÕ���M�O,x��
��*!� �Б�(S�<Xa��M�vNEkw+�Ĩ<�'�?����?���?aRg����5)4E��K|�\S4M�?��$�Ʀ�������	Ɵ&?����0�U���<9���@�L(��O&���Ov�O1���C��
��!�Yy7Z��)G�{�:6_`y�O2��������rτy`%FE&��XRL�A���$�O2���O��4�0�q�6)6t�R,Qr �0�ߚ,�:��K'o�o`����O����O��Ё'�f�@*G�l��d1�FH'%�l��Ӥ�ԟ �D�"M�)�<Y�'��K�-e��O.N��!��<Y��?9��?����?9��d�׆4J��aB�ݩP����@G� ���'O��qӂ�� 4�������i'�@RqhȃW�&A�+NCm|�Z�#$�I�8�'�T-1��i��I$������� ��(�����gJ���\
�O�p�Iy"�']��'���*��q�̟1YP:�Rw�@{�b�'��� �M{���?����?a*�,�a¥��w\n��4��2��e�����O��>�)��%�v���
]>b`#��[>�{�j
�6��d�/O�	�+�?!�m7���"R���� �F"�hٱw�:^#����OP���O����<�!�i崈���S�����Bx�h���n�	��M���>i�� ��t�#�S
tP���F�I��,O���-oӮ�:RR�'e��b�+O��  �%�1��(Ӈ@�EbB5O��?����?����?9���)�4Q�50p���?� �#_:3s�ln�B����Iß��	B�ß�Q���;��݋_q ݻ�,����.Û�?����4$��"L��9O88W�ۜ'�
3t_d"M�4O��ɃH��?�E;��<���?�V!�tH����^���a���?I��?��������A+S柸�	���QN\/9-�L�#�Q������|����IϟL�?Q���k (|В!ڡF@<���F~�%ùC�謻���ub�O����u+��/�,�S �xE]��׊>jZ��������؟��IF�O(�D�A(ɂS��::��Q$C�3>�Ҁ{����S�<�1�i�O�.*24A�gg
 �����D�O����O���hӀ��ڟ ���!3��@F�[0�u�sj�9�KT/�	� �%���'ir�':��'n2�'2��N�ͦ C�ݴeL��@��<��i���?9���?�O~Γ:d8@�d�����!�ы*�T���P���Io��|��?�i
;Nh�9�Z\�rD�QO\�1�^h"�$V���DF=j�� R�Z���O��7��xn�|��@-�<C�������?���?��|�/O�`n�4���ɋGip`fb���ƨ����_w���'�M��B!�>Q�i�x7M��-��+A;�)Pp�H<kɨ�@�L/QŌ�o��<!��5z��0/�^��'o���w4�1���+;a���gH�z�'���'�B�''�'r��I��J��gmj��	 &%���*�O����O oZ�cB�ӟ��4��) �T��-3�ڬ���/c���<����?��I��9�ٴ�y��'R@D+$��>l�HI�͈= ��� '�-~��I���'�	���ڟ��	2<*x�B\f��ݪ3�<���-�O*�d�<��i%����'�2�'��S�4������D&�@��X�Q�F���IßD�?�O�ҹ��̍)�`�����[��-��aʷ"B� �`�
bX��S�	@�+�s�	 &6��p���~���Gd�T���ܟt��֟��)�PyB�`�pD�b���0���
���UcfP���G2�$�OEl�M��	�4S��t:��ej��sz��#�C�ԟ��I�V� @m�<i�OT��Eڟt˓/�P�D�l$Y�C�ʪB9��̓��d�O$�d�O ���O��$�|"� F�{���ui]�4!S��	@�6cB�A���'�R����'!�7=���Ti
]\$�9��dt�YF��O��b>�c��@���a�$y`��Ȩ*4��à��&�@�� �OP�K>�(O��D�O���tp)�TO�!S�((2����{�'���'��	!�MK���)�?����?��V+i�4����ޞ��jGA_���'f.��?����B��)��SF���0���as�	�'���"BY����9��Ų�~B�'��M��uZy�	K3�D���'��'�2�'@�>1��2b3��Q��!� ��@�?`� �	��M�ЮZ�����?�;Q��Ur3�H�R>�hZ�-�S� ���?)�'ݛF"��0��v����6E+�t�Ҩ��k��i�F�y�kFxT��'���'���'�r�'6��' ��6+=x�PQ���� �
-�1T���4K}�`��?����䧣?ɤ���B�ܝe:A0�	��v�Ր�^�����<�H<�|����7&ْ��ˋU���r���>��c���r��c�GDf�O��`��T���_;}p��BE垞�0����?����?I��|*)O�qlZ�h���%B�P�rC�"~ԛg��:0rY����M��R˱>���yR�i*"Px�lM�N���v��#�Rї��!)������J�G	�t�Sy����y�ukl�r����Ka�T�2o}���	�����ɟ��՟��"Hߍ/�h�pc'���XӧԷ�?���?���i��O:҉f���d�<i�[����q��n�]0c�޹���?I���?��V�M�'�ܧ�� �5��O�7~����<>ܬ�ӭ#�~�|�_��Iݟ`�����@���ce� ˈ8q*ּa���ퟜ��Ky��`�.]Jà�O\���O��'o���uS)^H �0���	�"X�'7��i����v�|'��'z��l�@
�>dc����x�H��	ئS
�l��m�J~�O�X�ɇM�'2���	M����R�T�kc�'���'�2���O���M��TH��Jsi�
���B��Ա���?��i\�O0��'���UhF�b��
���p��*(Z7͉Ȧ��`�A馡��?9 ��p�F���F~�I�r�$4 �#X~�F�+�f�%�y�Y��	ޟ����8����h�OH�q��O��"5@�/$���@y�������O���O������UҦ睿qb�`ZEi��E�j��g&2kN��4,��&F1��	�&�.7�z��hqL��|ނ�*�	O�F(t`a�x�'&H/b�n�b��oy�O�d�&E����,�,���YC.�]r�'�Zv�f_��@�4��ŀ,O���ό>��|�q��W��l�n1���?��]����4W��x��_.����U�Hue ��d�a��ݛS�S9V̓�����<V^��J�$��mAF!72��9(����!��0+w�r��3V�\��Ȏ.~�����qcu�J՟��7�M��w:�ѹ#�=�`[R�T��p��'��'v�я=��V������x��sSz-��$�2��Lx�Q�	f5pM>Y-O^�?ѥ��P�^��P'^����#�B~rbtӨ���N�Or��O��?q )Uh�ْ5MP�"N��򦁳����O��� ���R�BH�3r�W*J���
�lC�O��!�fӊЗ'��W@�Y?�M>!(ORyjtלx`��pG�P�X M���O��D�O����O��<�Ծi%��
��'
zݒ%��P�@%	�*}Z��S��'��7�*����D�O��d�OH<�B+�2z/�i#ɍ�#Ŭmz'#��$6�{���	�M�d�p�՟v˓�*�;/����Å[;M��B�iQ�z�����?����?9���?A����O�,ـ�$�._�q���	~���Ȃ�'H2�'Hl7-	�.X��O�oQ�M��d�J��(�4��(7.�\�'��	��ӰSA�)oZ~�n�4*)��X#bE?64�5����\���]N?�K>�)O����O
���O�4j��H m��SQE	G&j��B��O����<���i��0@%�'�B�'�哵q�X�y@B
�g~*�
�"�B������X�	X�)���H�;��d'��R��ׂ�?h�T��U�M�^�擝���4�ďf�%�Ν:ib]�f� g����O��D�O���	�<��i�����Q<@��(���X��ւA��'�Z7M:�	����O,}r&��5m�x�2E�>$9X��a��O���M7LW�6m9?)vMS?T���yy�GC@�~����)��A����y"Y����֟����p�I��O݌�Z7��3�V����@�z�4�ʔ�aӦY�r��O�$�O����dC��U�@ ����!S�� ��h�.)�	�&�b>�wEĦ�͓t�S�C�z�Z�)V���̓4>(a�W륟,%��'J��'���`�I�a�@R#@Ԟ]��1�1�'���'6b]��"شN������?���o�h�P�?)]�09��D�,�"�>��?!L>��hՈwE
% "���v�ƌSSG�<�����y;6�*�M�v]�(��2Q����O>ٛ�12��a���(�>̹&��O�D�O���OB�}��X�@q+aa1���O��̚3i��?9��i��$���'r��u����݂��1�nO7)�ƙ�g�A�mT&�	+�M;�i��7-D�5,�6�c����)|:,���O��}Z�g��.vH��	Z)o��ՙ�#�g�iy�O���'���'�b7\0i��&��Rb�� �I��M#%KA<�?���?)K~���R@��"��>|u���f�דnZ&�p1T��۴/盖m+��I�4���+0�������iٱA߶� �M���ɳc?�!��'u$��'n�y�A��G=@)�n�xP`�'r��'�r���$T�p�޴a�e��dJe�%,8�燑T�8�X��%���D�Iy��'�ºin\$�cj�x�N]�4/H$X�p�`
W�͛&���j`�����^|�������0���')Q�z!:����~����џP��矐�������B �	ڍdc�>�:�Ӧ���?����?��i�V�7U�$��4���а�W�ݴ��!`��*A�`�KH>a��?ͧS��4������HA�<JAI�6y0j�ʒ��t�`�	X�I{y�'�b�'�BIJWM�HcR�ֲhP�����^���'K�	��M{"C�+�?Q���?�-���[���%��ՋG�lc�d2����OF���O>�O�S�B�4��-Ђ 9���%�5�d�)�NӉ)=��mڎ��4�XH��'�'�\��*�'c�h! �@�U�T�'���'w"�O#剳�M+�A�0�>$��MA�&�Ч�F�j���++O�-oZ�"��I��yW�]7����hTS��}
�͟���3u�r�lZA~Zw����7؟�˓@0N����k�z�i�k�7r������OH���O��$�O��d�|���[;.�\�ӥ�2`	<!+A�\�-ǛƆ�3v��Iʟl$?����M�;A+lU��b��'����w+S�0�x���?iJ>�|��$�M���� P���L�ZC|���+�f�h�e<O�t�7$��~��|�R�l�I̟\8ХO*	�^}	��՛��ę��U֟��Iğ���NyBOk�R�Ԋ�O|���OH6@N2=��)7(Q��apc$�I���D��۴"݉'�f$v�J
}5b����&/�X�ObĘ HF=Q)���I=�?���O4��΍w{�d�5n�B�.�����?����?���h���W}�fu�4 ����x����'h��_Ŧ���2?���i��O�.[;'U��uk]�pa&�Qr�3~���O���O,�C�u�N�gX���L�?����(G�
����ű[l�dꢩ�{�Ipy�O���'���'���Ƹ�A�5c��f�
�n��p��ɝ�M���<A��?�I~��h8���X�rF@���/ǩU5���\����쟀&�b>
Т��U�<p��GD�A���F+'��n{~+��D����������I)\6V}s�	�o������$}^���O�d�O��4�˓G�&­/L�!��cs$��F܇xR�̓�jE�/B/b�����(O��$e�<�lZ ��S��D��iB D ��I!(����'q���aC�?��}���V�(�hȾ%if({Q�LT����?i��?q��?���Oǎ�R��ԓ��o��w�N��Q�'���'��7-�4>��O�oZm�I�)��Q�#F��Ȭ�R⛊ߒE�J<�i�j6��:y��Kb�H��D���߅(Clc�!� ��,�h��N�n)���'�e%�$�����'���'!����A>u�Py��C�0h4�'��Y��޴e�na*���?!���I<G9��J)Q&:iZя�7g[��7���O�7��C�韢���l-�zS���b�e�X�8T��+�"9L��ݑ ��x���r�b@l��d`��P��> ����f�9>o�A�I͟�������)�hy��oӺXpNY�L���%�ټ ���h.��O����O��o�W��c��I�S��K�uN�Zң�] �{&�NBy�)B�&�� X�'A�$8�Poy"�L1�����(-"�x� ����yR^���I������|�	�|�O������8L�|�Q�P̩G�s�����	�O(���O�����P��睭)��0"%�G�EPp-�V��_Z���	S�Ş}D�aݴ�y�`_���q�T��l٢�@��y2XXLq���-s�']�ܟ����}q��)$� L� y�#�$�t�Iџ4���'�7-X<�t�d�O,���m�� ăfZJ��6�B�9��t�OZ�0���E���4/�(N��Xa�iBq(��Q����ƛ�Zx�I~�ѥ�OPx��)�To�u׼Ha4
��x����?���?Q��h�N�DA9 �p�`1�)C:���O�e���_ڦ�(�lG����I �M��w�bUС G𲀹�(Ǫr�B�B�':��i�p6-
�3Lx79?A��B�Z b�)�&��d�@fG��Ђ�6}f�jJ>�*O���O
���Of�d�OƸ�s/a�X�"RBƅu�XB�ϥ<A׿i�)��')��'��O*B��0q%�� �K� ?y(5B�i��s���?�����S�'�&�ې�T�F���(�N�a"M4D÷�M�V\��m�%!��1�Ĳ<Q���@�(sd�J�J4�0H�6�?���?����?�'�����͐�e��$�3F�i�y�%�PV��&c��D��4��'�듼?9��?�0��< � ljmSmFM�5kA.��]�۴���֬%qH�O�O�N�h@B� !O�AX�L��a��y�'B�'�'W��I]!h6�jWd�	�P�l����O����Ӧ�Jb�m>q�	��M;N>APdקb��A@3�d�X{�b�Np%�\�IП�	ǯ3/(6�>?QP$�'$�H�p2�I�bF\�sb��>�j�	���O�DaL>*O�$�OR���Ob��Q:����P\T�O�O"�d�<qW�i:�92�'/��'���9�F�x�mSD�X�h;��c��	+�M#�i=O��P(X)��ɡ ��5���!�j	 E�Չ8�~�%?�'p��
��)p���1#6G{|i�
�w(�*��?����?��S�'���ΦY�5�G��0�rPk�:$����F���u��'��fi�Z⟜C�O��l}�vq�ĸh'�m�����U�����4"ϛ���^��V�� y��D?h/���~�"mV�[�8E����:^��A�O�<�-Of���O6�D�O����O�˧ 
8�t�i����b��2v=hH��ij�k �'V�''�OWr�g���.Hx<�P�5ަ܊wK��u��o'�MK�x���P�t�V4O�Ѻ5� iѲ���ˀN����?O�	p���?Id�0��<�'�?��æ^���v� �⬃��?a���?�������c�������I���Yd��&I��A������j¦�Y��N��>�M���i4HO
�AfU�&J� �t��3+S]����AB�^,!u���B$��!}�C៤����*%k��Z��0�H����	��\�IΟ|G���'��x���7
�����_�1��H��'��6M��u���d�O�mg�Ӽ[�u��1CI_~���o��<�B�iƊ6͒צY	3n�ڦ��'���7���?��_��%8��ȑ M���"����'H�i>�����\��͟@�ɩZ�R����1�X4J�D�;0(��'��6-�U$����Ol��9�9O�L1��L�z�f�� #Pu9ҧ�T}2�'I�O1�j#�� &h�g�%�^���Ή%;�Lm��/��xt�ʓ'��<r�a�O��	I>a-O<���E�'�&p[}�-��o��?����?����?�'��$�צ�@�)����&)�n�CS�� l�$I'lUߟ���4��'�<��?A���M�6�=v��NƻO�`}���Q��W�A�'�Bt����?�����w@�9��T2X^	p�ܺXj���'	R�'r�'lB�'t�U���A<v[.q���(:�z8[��O���O��oZ�#�)�'>6-:�d��}e
�@�j��"s:)�螐5.1Oz��<I�Ǹ�M�ODIhVF�rE�wJ��|�V���ƀ D*i��x���O ��?���?a��	���V����Ѻd��rj`0���?�(OB�lګKT�9��ğp��y��gד%*9�G��Sc�T!v�����^@}r�'��O�S)'MX�7&�������ԕ)��r����bcR=��~y�O厙���B��'����&/Sm����h; ���w�'@�'���O���7�M���CF0�7K�2�K%��1<K@,��?)7�i��O���'����Ւ ] 9�B�x�`U/KQ�4�'��H�5�iY�I-%?�-�C�OV՗'��c�@K=0�]Dj� ���)�'	�I��I���I�d�	z��'ϞH��05�T��­�f��
3=b6�6>�����O��d/���O��nz����S�Td�$ytƝ680�}��֘�MK��iMO1��1�6Noӈ�	�6���h� 7�P��ڝJ`��I�FՐqz3�'���%�x���D�'+� t"L���4$�(\SJ�@%�'?��'*�W��I�4]�4r���?I�'��b$U�Y�%"`��j1��")�<9��?9K<AA	�n��9��
��V��1%E
`~r��52����B
9`�O:����9)���!���A�^y�캤��,`�"�'�'�R�sމI�(E��̔��T�E�� A��Wڟ��۴Vf��
(O�)oZi�Ӽ+Q�6/v��Ꮘ/4�$\zc��<�`�is��qӈ����u�T�5�P\*$#�(aKǩ�����6c"�tҰf�"����$�O��D�O��$�On��\��9�ϗ�K��<�A��C�\�}�����B���'����'ހ�Pp&��NIh��6���Qe�>yT�i=t7�c�)��;�L$y��Uc���0?Ϯ�R`�װg���c~�\9���O2}!H>!-O�9��!G� S��a�hL�p�g��O����O���O�i�<I��i�>�:5�'܊�:C�[*wȮ��@���Qr�q���'��78�	�������ߴlD��C\L>&Uxw�A�M&H�w�d_jȚW�i�Ɍo����Oq�r�nFY<����I�"^b���ˌ�����O���O��D�OP��#�S�L�<�� 㔆3�D�����7$$�	�L�	��M�2��D~Ig�*�O�<��׃?i��3$��d�Sw /�$�O��4�P*�`�b�8O̼@�o�� 
���ٱv�Щ����f����h��ry�O���'���Q�zM☃�n���}�V9}J��'��	=�M3U�<����?�-��mp2��x����*GCJ��☟ :�O��$�OZ�O�Ӑ<Tq�`�ؖLn,���<?�ɣG G|�Yo�~�O&����}�za��ć  �h�F+ǁ#vh����?i��?���|�`+X>{�@��,O~5n�   hb�FgA�'��X��%!���D�"x����X�ݴ���?I[���Ix��c�ķ�����A��3�
�	Ο���*�˦a̓�?�sF�j=d�	�:��DʃqIx-)'� H8,a���Ea�$�<���?q��?I��?�*���)c �#J�B�*�şA�B�j̦a( �V����� %?��ɒ�Mϻ�V���P�v�� ߹��������Od��'�i��M�x�8g���4V�%�c����ވh���a��>�r�O���?������OZ="���K�	z�����?I#�ݒ�?.O(�n��wFjU�'G�"#)R `�`&O�j�R�'F"Ru�'���<A��?�M<�AӍp�RD���o؎]��Ɲ�<q��y�$��㯛�'h��+O���O��?q��OڌӥjV�����JF�����O���O���O����9kF2����L+�mHgG+��M�m/!���D�Ԧm����	
�M����4����9j���"wL�q�xm��P���$�覵��4Z��&CCϛV4OD�ė2�٫�'o����w��U����[4��8�2���<����?����?A��?	oξ|j�զ�e� Fb]����\ɦM��#�m\A������O("�'�f�i��0צ��ɳ7�+NX�����O�@�i>����?e2#���p��a�Q	�A����LV��*1ley"A9Du4q�I�y��'t�	2����Bl�1[��)�iT�|���dDۦ�IPH[ǟ��,�P�rmR�h�p`D��˚ៜݴ��'lB��?!�Ӽs��?i�)�l�P�0�
!C2N�\�
�4���)�4���O��O�����T1�F:����ZL��a�[�a�re3@��)��hȄ�|����7�Q;�6��3���Fd�	!��^�u����dɗr�(��͞�V�|�t���u�ɦ�@����$D��(0t6��!����hè�R��>���& �70Y(v�*kl�pH�*:XnH�����xd�H�Es&|
b�@�Isf�!�Ӊrݠ`�u�Ī>Jvt9u��d\b-���Q[v�J��E�e*�U�uN��r�ȱ�h�eӆ�]��M����J0v��	Ny��'��Ğ�=��+�+"�6��$C��0L��<�r�(O��O�'��'� H=� ��6|�Z�B2�ΊF�Q�1�i� 5XZ�I���)�O��O"�ĈD�B0�J3.��cg4�*�K}�卉B�b���O��d�OL���Op��H�g�!Aˉ�)�!X!�U  L�D@wF�<��?�����?���6�ұKb�� �r��3��>~t&����1��5�'�R�'N�'y�	��QR�)�:Мs�M�w���D���o��P�H��b��ӟL�	,�����b�jy�@	��l
��`��0P�@�Iܟ��IFy�J]M�p많?q�AK�U�zh�iA6(�V5�v��S㛦�'��'���'.�CG�dȱMJ���P��L���3%Np8���'-�Y�`�R�؜����O���v)Q��
1zd��k�Fl����G�̟��ɣ^!H�?��O��H�f��>,�R�n�WD,Mc۴��G�gzf�n��\�����������zl�ѧ�w�� ��J�Qw�i=��'�J%�� �� {�>��e��|���B:��6��*�l��������S��$�<����<[d��Qmۂp`ZE�\1{'����Oj�?��&2�qH���_� �����L��H�4�?1���?��O�M#��Xy�'��$�,Xt��cU6H@"�z �d�O-�u!��O����O`�j! ��9볧��v������Ҧi�	�V[��K�O�ʓ�?1N>��|D���L:a�~ �C\�lQ~]�'^2���|"�'r�'�削N��� �D]l�RTZ�5���x���
���<a����?i��h��:� 2bE��:��̶z���7j�'�䓎?���?).OJe����|$Ɔ,Q��eR�L��?-.S�dU�͔'3B�|��'2���# ��� 9@�����!96MnĢO>��?����?�)O~`Z0G�N���'s����/Ɨ,@�sAY��DzdMp���D&���O��dI1	l,� Q�N%��Xjw�XR�2A���i�"���O�ʓH.ܬ�6W?I���d��8�,!Bう<'������C��I<���?�CT���'���GG\�0��B��4I�e�P;��X�@��`7�M��S?�	�?ш�OP��7���c�鋍!B<���i���㟼�ɞ�ħ�����Ϙ}������&fvdB'�|��iA�o�ܦ�Iǟ@�I�?-�K<ͧ~Ƅ���,Z����V	6*.Έ�a�i{2�'�R�|ʟ�d�O�(��R!dJ�u�6�~�Y�1#ʦ��I��p��!e�d�YI<ͧ�?Q�'2ޔgd�$E����fY^���4�?�N>!�S?�Iȟ���؟�ǂ�(o<C��H�������6�M+��K�)b�x�O�b�|b �9l�����
��0H�����O���<)���ɰ<����/�X,����!�b� 6�:d�t���xb�'�R�|r\�֝����h�ᙾ��5��]�>�7�Ol�OL��y2�'�p���ӟ$���+�8m�p�Q�נU�(�G�i,��'c�O��D�<񰮍ƦMQ �8i��A���&�@e��� ��O�˓�?yT+����)�Ot ���%O�#��/� mz�����E�?9���D�PL�'����b�AA0���?�0��4�?�+O����#$X��'�?����1M�8��Q�G�_߰`��ǚ@t�%�d��uy2f1�O�լT�,̞���Pqc����i��	"1� �4V`�S��@�Ӱ��$�-C�D��Oʶ,�1!�j��vX����ڟ��M|�J~n�0�2��c�/ H�����)[\7��3v~Z�D�O���O���<�O�25s͘�	�R,���ͮ�؝��Ou����E�5Z�1O?�3&O$jLxkd�)��S����M���?��f�`�-O�Sc���>Eƌhs�L� �<�[�	�.NG��<��B̩1��O "�'$��> �('��4L��y��!��I4�7-�O�+�	u�i>)��Z�iݡ�D���9�̰l�4E�Lg}��_�`f|b�',�Iٟ0��e۠��so��aHz�3�$�?�	�'4B�'E�O����OJ�rA�ޑ �*�Q!���u�t��C 
G����D�O���?��E����*��e� Ȓ	� Hw@Pb�G��M�)O��$������%TT�7m�����2��ֶ�����lX�'mrS�����
��O�B��5�x�Q���DP���6�Y`��6�2���\�I�b>���@m$�Dś$z�ȐnR�u��݃��Z�v�']�^��0��M��ħ�?����B�32����M)g�bXw��S}��'��ɀ�����P�Sqz�hp-�!�5ĩPv� �WA�&X��HEg�M�T?��I�?���Of�w�+��k��J1�%�D�i��I(N
��	.��'��禙��R�X%�R���^��\��Bcӎ%�k�ަ���럸���?m�K<ͧo�ٛFΗ�G�2HY�8�Hsoג�MKm���?����:�9O��D�%5�2����NY��n�.4�<l˟����L1��� ���<����~b/��
s� ���ä\����Ũ�	�M+O��$=.�?���ܟ�ɚ
��$a-O�.s��r �2����4�?icE�A�Isy��'�	�֘-;Bd�q��-rv�Ҧ��+7���%i����D�O����Oʓe,T¦�B�rˤ�dl� ,��1%���by"�'3����П�S�`ͫoh��K�ȓWi�$�@�ĘYo�������	��t�	䟈�'9n�0�v>� �@���ݧfg�2�I�� ����i����@�'���'�"�(�y-�s��G��8��AfC^@` ��?���?	+OT�w �`���'���*9�y��
�l��� Q�iӀ�D�<��?	�F�-Γ��i��e`ǯEv8�S�[1a�;�4�?�����A
���O�B�'��$��U0B��_u�����$�)�t)�O��$�O:�I4j��D8�$�?��WK���xm����o�Zճ��y�h�,c�y��i`��'���O�Z�ӺCb�C7S�����w%؅j����}�	���SS�k��%�,�}:��C	h}�Y2C�QeU��J�(ƦQ`�O��M����?���gY�\�'%J�R ,K
s�fa��	�\�6��Іt�|q�>O�O��?]�ɶ,�� ��O��3�f��գN�F�(ݴ�?���?ya)�(j���uy��'����|����ύ8$2�m�RIT�$���gy)Q=��4���D�O���B�J��)j>�8�� H��-nȟ�$퇩��d�<a����D�Ok�I��L��`�5#m�p;�װQp�	�O�D�	؟��I,�	ܟ��'���&��0������ɽ57�
�O�1iʾ����O�˓�?���?)��Nw���Ǣ>d0���E� ,ZT�Ipy��'C��'�剠?4�ʚOct���
�~��%�����'#���4���O�ʓ�?����?����m��dM?=Bbԋ��  ���Q��O��M���?����?+O
��C�P��~���i3đn�څ�4��
� �z2�����y�'�']~ő�}2��I^���ؖp����M����?�*O�}�`�d�$�'F��O�&u&꘎E^�: �Fx�@ :��>����?�� �����9Of���=iBP�$FF0{���Z�R7�<yT@��_����'`�'�t��>��/l�e �j�1;�4P�g�)lrEnZ�����6_M��	���9O��>�y�o*H�� 8�>I�Ɖk�����¦��	��t�	�?X�O�˓z��()H��
E	?Lu����І�M�uĄ�<���?!���O"�)��O�Lq� m�R3�3f�b6M�O����Of@S�̆L}�U�H�II?�ӥX[e���;��$Z�B��6��<���S��'��'Ě$t�h��Kk�(Xi�Ф`�����.Uh�`%�����`%�֘=1����U ���\��T���y��<)���?i����DP�!)�%E�6%�����%}�I�`�	z�	�d���&OP��b۞L#h��Y^A A,�6
N�D�<Q��?�I~���M�D���ќP|dD��#�'*Ɖ'l"�|�'m���U"j�>S�pA��IT��Ȑ��Cn���?i���?y+O.���@�ӕ::\hb.pv4�3eV f��!i�4�?�J>I���?�����<!H�|*t��|.^� '�4<��Y���u��$�O�ʓh������'��t��0��S����ny�!�h�DO����O��C�6O��O��6�"�S� FK�L)�r� X��6�<��! �c��F˯~r����񚟴�� S;tYa�S�a�0�S�y�\�D�O���:O4�O��>��'���.s�3(N
�X��vӔPX�
Ŧ1��ӟ����?���}�'
Hm(���$B�5s.�� R��V7MI :���.��-���������	\�6D��Ѯ1\h�c"�M���?������3�d�O��I rA.��$9�$��!�ɏU<�6(������?��Iߟ���"d,��0~�<�U,T5o�͟�ɀ��'�ē�?�������`ۥ_�Arb�'c��%���C}�Nй>��\�x������	sy�NڀDr-��T�^��bCj��
�ҩa�K7��៴&�����8�0.T	K� iau�H�n�aA��Z�t��	Wy��'/B�']��MI��O��ըaƚn2��3̉	0L�%���M��Ɵ�ɛu ��Ɍ�r|�P+�6@�; AT� �&j�O���O��$�<��gH��O^*X�$��ψI �M�G:Ɂ�%n�f��;���Od�I^���"}R��ZRB����WLȡ져�ڴ�?I����dO -/� %>���?�X':,�C��0�W`��V��b��I�Q���I]�~�F❰V<r k"��E�640dAHԦ��'0.xC��aӬD�O:��O�q:`ZXU  �J�gG�>�F�� �i�I�����?�g�Ix����-����]3$�P6�q���k���$�O�����x%���Ipb�����V �E�:i�l�PشM�:e���Ϙ'*2� f�d0`�e�n����'�/jE�7-�O����O�hPW�y�I���I�`�qj�`}D���D6(�F��W�F�@�<���?��B�q9�ŕ�{3�z$�4o
�l�0�irl��C��O���O��<���~��S��n@bm׺P��	�'u@�C�y��'S��'���;r�P ���E��p�f®U&p������ē�?)���?i+Ox���O�ik�@�*(!H	9�Ŋ&Uɴ��'ݿr71O����ON���<Q�D� ��I"]�P�c
�:L�Ե�b��*v��&[���	Ry2�'a��'��|J�O�ș�X�2��e	��w�����i���'|��'R�I�@Ӱ�j������F��`�B�B�2��) ؈����i\rY���՟t�I�j��I��T�Qh���#[rZ<���@=g��-l�����Gy���4p�'�?Y����� ����W(h�&��g��8�I��_�D��Ο���'g���u��'��	�-�`uS&"Y�bjx�
T폸8R��R�0`���MK���?Y��bU]���6A�Pܐ�
@96K�=!ǭ� Mi�6m�OT���7 ����O����O�Мq��֮�#�/�j�����4W�֥26�i�B�'#��O>@���䋫�<+�C�i	$%��J�o���lڥK���Id�W�O[��)QŘu�:����d�L�$�B�L�l��]�YMh2U��yaz2�0������=�FԨa9���D�4�&��J�&@=[#�?&QzM �8�,��B�ո#n�)�S&�.�HX�H�:xtݛ��52y*�@��.:�� P��)��ҧD�����	���.;9�21��*kf\IZ�h��<Ҁ�'��&G����pI��ś'`����&q��$H*0���MB9��'���'Ȃu��'��9�� K�����z%��(+�����u�����/R,cb��.&�G~B�R+J���`pe܆A�F������P�p�̱fb�\wJH	,jn9��c4�g���	��|�e�2�h�J^8FpL�HUG�j�'�џ0Cg�Ό�4�&�[$bR}9�2D��3Z�Œ#"��H0LQr�Co�Z�On�z�<�(�\�t�Iq�t%�	T����Q,F.d�Q��	�0GG�|C�'�R�'�p���C,D�$a�C�6d���T>X�W�T�$�q$W S2��.�+ �!����g��$sb"׋��'���{�Wpvx�zw�I5
�XDy��E��?����O�h�bW3&�`i6�ڀ6����'���ʜ�}�}���QN4����L��0>Yv�xbLڅ��"!
�8I�,j$���y� ͥ"����?Y/�̡ )�OV���On� ���{d�����ǡx�Pȥ�T
>����DDW�Ĳ���̘ٟʧ��?���M�HX��wclY�E��Ӗ��2�WrazFi�a3����OR)�D��^*�����M�E{�+U3M�����O��S��P�h<�q�7�^�S �J�+���C�	1 [0��ӷp!:��f���o*�#<�)z��:ݒ��?N�,<�^S��?�C�,G��=z���?���?�����O�����ƒ(+
+O�V��i�ҟl��]�Ѻ�k�hS
 ��	0l�ʔ�F�5���C�ܛ]���B; �(@m�
�P9�V��?�=1b��X� ��Coh�ؤ�b	~?)4�V֟��	U�'R�	�G��B���;R��@AUkW�dY�C�	q�z��sO���P89���O6�=���?ݖ'�l��Dglӂ��u+���C$̉�Qz.1r��O����O����,���$�O�S*f�1ȳ��9j5�YG��������{��rA:�O`����YH�7�
%�}��BOl]��Y+*X��|r�M��?i��G�����/_9Z4�q�gT2WW��ȓ%���pd��j�$��x-��U>� k�-ڢW1�,"e J�8�� ��|�֌@6B7��O6��|z�mm\�TjϚ!�t2�h��w]�]����?�[��X��蘧�
<L��d�-j��1֍O�0�Q��q.&��	���JĂ\� �y�W��*X2$Fy�C��?!��	��UZh��i�aȩХk�!�S�#t�d3�Qh2�0h�	0�a|bn8�$�<e�I�G��[ ��'�zL��a( mZß��	M�D� 2�'�!�8G�4�� @��
@��#�ҥL1��'1O�3�H3ܡ�������	��x��D'��O?��M5?c���DH�(A�Ds5LG%��H�3�O�b�"~�ɦA��L;�
F�-�H��3fք�rB�I��\2�@Q@Xx��UCT�v�T"<q$�)J�'͋O��S�HH�����̎��?I�Yf(�
�����?���?�� ,��O�C�+b�y�
��� �f��[i��0b��}b.I���<J�� �0�¼��b���~�\���>Y@O�e� �ϓ9\j؅���M?�w@ ៈ��(/�ٺ��=��CK=�2B�I�j"tz��/
��HV͓�d�P��ᓋ|d�ڴHs��`��R�l�pP�B��o�L(���?	��?�w#���?a��������M7F)��!�����M_R�t}���НP�`��	�u����'�@�P��"�Ė�-����Ҷ��	���I뀷X	l��G�b�dٻ�#-D�*�j	!�ˋ�[��	���� q�!�D��	�0(��eLs j}X׃H"v��\M��0G�ih��'�7$8�IXEB�*Y�Q�a��_�*�C��]Ɵ��ßX��)&d�\��N>�O���rć��[���
����Ė�G��u	�")�'|�|A����ޱǬC0^l	��	�"���1�g�? �{�ˍj(&]8`B���vIV"Of!�"*V=m�a��f��f�xu�'lvO\�Ƥ^�Mݬ<@  ��2��5O* �sI�����ؕOv� �'���'̬�@�}H�pb�b˒'�"ES�-R
wh��T>#<��#ΨU��'`�r՘�+|<<{����O>�	�������ʻx0�aV�C�R�"��"�)��4�� �Y�"��5O�"4	��'D��&��X�y`��=�9w�:�_���U���[�(ß|�=��u�ڙbn�O$�d�/y�‌�OB�d�O6��Eɺ;�Ӽ+�l� i�4�D��#S}b�ZgG�s?q�#�}x��dgW�ⱁ���y�
x:󌫟4)�	!�Oh0Y� �:{��Ef�0��j��O�1���' �{���<�^��$Y�&?0*g��%�yr�"7�8;��v�`�S֍L���#=E����94c:7͞�8�n��2�T
�z֋�cKpѸ��?����?9��	�?A���4 ���?��L�2���.C�z(� +e� E�����I�Hl��	��h�	�3���b��W8&�hh��ɇ]���Oy�6�\�@�FyX�Mڻki�h�""O`I�lkq@��Vl~���"On�2V�A��9�0,D&2����0O���>���kf���'`�S>M��N8�T;��$ ���i�ތP�8�������e/2]��@�S��T�$楳s��\)˃e��(O$`D��7�>=�uFK�n���bF�^�H�<�5��TD���J�_Z��q+Q�wF���&��y�
��'U>���"OhFZ�K1%C;�0>�%�x��@��~� ���Y&6�x���yR���7��O��$�|Bя�,�?����?�(��U�l�#e۾F�fD
Uhםi�|Xx�������(@]�Ы�)+��Iq�B�O>V�{C=�S��?i&��H���A,/���� BÈf@���ؘ�����H!�[�&�I�4%��@Ȣ�yr�څ+��lR�E4G V1�.݊�O(XDzʟ�j����%#�iX����&�SFM�O���@�rx��6L�O���O,�d�޺��Ӽs����!&��WFW�s��j�JQg?1�ϊgx�����sqNeIFV0Ā�&����'�O.��pG��n�R��2�֖!,aڗ�Obd���'��{b��x���
��Q�q���y���UsR��Ֆ?��@@ � ,��"=E��Bӱ}N7�J�~C��r¢M�eu���)����D�O`���O�i6��Od�j>�ɒ��Q�t\��ӸH�y �?mMZ5�"c=H�	J�P^x�t�aD�
h(�K�F�!
�2iq�-�}�x|��ß$)���S�^Ox�`���O������p�D˫�ƴ!�e҇r6�=9���C�a��+��k��0��cW#.!��&�8����%=�<�z��V�M�d�e}2]������M���?�/��Pq"��T@�� ��L�ZtA�O�\R����O
�����|��8�|zE0iZ��sB�gM�yQ��z�'xbZ��iӏ�����U����F��Q�\� ��O��}�ש@<N�
�$��cD�N�l�<	�A����K�2(l�Taӎ�d���L<��<\h�r�iT* �))j�<��!�'����'�"_>��@%�ן�������$��|��\�@!�[��	�P�i�����u�S����@�<�j}!B�؍n�h8�"\<E��,:�S��?!	�+��y:1$M�5�XQ� ��"��0�������"N�	
�H���	�.*�c+_��ybd�6(w|��D�Z�<�,�+�a�O�qEzʟ�U#�EF5�8�gC�${I���O���Jb�MP �O��D�O��d��[�Ӽ�PM�8^Y�Y���R�l�u�W��|?�@H�fx�:�ۃ �
*C'K�
����U���`�<�O4��#�l;�]��-�8ڠ���O�u�a�'b�{� G:`�V����G��d�Vɒ��y�꛷
�9#���fū%O��U@"=E���%��7�2*^`��c�&,&p��R� ,^���O��O�x�E�O��D|>��+�O��ֳO��)A��=��9�-X�F�|�@�����Y��H�5MT��E�w��D@�|bE߱�?!�|����ҧ@U4���[�d݄�S�?  ma���6��!j�	])j��#"O���ʞ�r<��ɓl/v蛆6O��>�"#�6�����O�����AXP�q���
��Y�BA�m���'7lV�}���'*M {}���ԏ<����9���A��9~��M!c��.G�)Eyr���V��"�R�D� �a1�):��<9̈́�(fgπ4�x�T�C;	ģ<�@����Ie��&�����+���٨�� ���?!' ��I�TP��Oz�؈�h�n�,PK<�nS�GO�$�����;�@��Ȟl�'��y���Vb��A&'��q����cA�y�Ť=]H�:�瓲騁�0���yb=w2�	EkJȊ��M�y�Hܕ0����'Q'm|�q�,�y
s)T��i��?���ТZ��yb�ݹ+��dX�͂^�"�P#�R��yb�A�q��Aö�Pu�M��"^�y2$�W��iw�X< �S���.�y"a��,;����8;�����[-�y2�"'N�Ո�/�,1" �[q�ڮ�yĨ�&t��&	�w����`GC	�y����Dx�M�v�D�j^��y�͚9�%���t,���$	��yRm�y�ĩ�.�j��Q���y��&��}�V+V�x(��Pr+���yN�?�N1����$k�yQK��y�@]3C��̃D��0�z�2Q`�-�yr̟+r.0��
��rU#q���y�I�;���1���5 {��0�J��y���9s�d��A[�-�85C@k�#�y2�N�*+R(� iľQA��鷋��yB�"h�NȣF��Q�����H�*�y��і,/\,1�o�4P�Z]Zf@�$�y�
�´��h@�J=�E�`��#�y�傻$�Fh��fn�:\�06�y���AI
$�0�X�iŔQ��(.�yr�ڭ{:��fc��\z<4��F���y�)V$khڽ��ΥXc�l��ˉ�y�`Y�_*�	��'�|���X���3�y���w'jX&
�%S*E�lH�yb�V�@/X���Ù�瀀�7R��y�gނ$2B)c�*����)�BB3�yRϖ 5���.�j��G �Ti\yz�'�x0T�nN��M� O(M��x�ӂ jF1O?��'U�ʅ˕wU�E�̆9�!��!(�&�#0����$�3�R�D����U�t\���<lO���@�a锸�b(U�W� )2�'N��$`ɲf!��Q��R"k۟Q�n���P0�yҥ
�}��$�̗��S����(O���V��y� #}d�٨4,��ha�"l�j���$Yk�<���¦�Z�ـ�@�2�	;�&N�>Lʱ�Ԛ	�ɧ��2a�>wE���´w�\�r���y2_�L�x���hEhp�u��|��hx	Q��=�'L
(=�P��,T3h?�A	d��m(<Q�4F�DK2D�v�l``mԒr����ȓN/��˕�@W��9�do�x�P��?�qE�U�)$<|9��L).�$��pR$�(�/[�|�p��r�N�ȓu48k��Nq�<AOA�}���ȓ'��6�O	�J̐1���E���ȓ�$�2MJ==x*��S��~�`�ȓ���H�K
%�&���ËF#N�ȓ~��ٰ��!]�`�@ڌN.��ȓ0Z�]{��T0FIBE
�9�ȓ/2�)�H"-`2��d$��ȓ1=�ܓ�j������Wb[3K2���S�? ��:OO*}|:��4(^���5"OX�hp C|�i�d WmP���p"O��(�	�m� ��d���XL�tp"OH�Cb�öiv�4�wa�nf� BE"O$0{#���б�n[�!N�T�g"O���d@�Eʎ�)S Y�s/�+ "O2 �,[/D�Fi�a^B����V"O����ي@zb0��m<-"@\i�"O���G��'�2q�m�#92�u"OY f���n��������� "O`����@&�@�'��/��H�"O M���-��53�	O=�6�r"O��C�i��-���'_�{<�"OzE1��>fN��p摷Z�K4"O�-AԨR<t�P�$F!�>�"O���GH�DT�q1��%\��"Ot3�7"N���,Z`�}	b"O�4���B�u�r����d�f=�F�'�b��$���:#t��J�̆\����CVz!�#=�ڡQ�K�0��t+�._�'��Tkg���Ga�����FID�����ŲP/!�֗|�j�{&`˾�X�"�Ћ(��O� :�E?O�Ƞ`����Q�V�R"j6�q$O�A�(�^53���ztˆ/E�<PB�I�C�6��1虳�sƊR�@���䘱�b���m��(��8�3�0j�B�,D��{��ͶT�LU+R&ʕX�~e��<D�Ы�呌_H�	s��ɣA�j!�-%D�P��'V�4� ����!3:@I{%�!D�d %�f��t���A6G�9k�H!D��J�PZw�$z�hU�IJ��y 3D�$�E���wY�YI$MG7v*��`"�6D�(�r)QR�* 	�I�=.^da��>	S	Y��p>��(˗/�f�"G���� �3�c�\��Y�18��I�D;�#T���{4�H��ȕe/PC�I7#����r�D
y�
<�kź=Vc��X��Q�]��hw��y�Ot�IaL�b��D `�U�����'Hi��V�*�{ע�!�"\�İ6�ܩhA��_yr0�g}¬�%1�숋%�?jW֍�bF<�y�� �r0pp��0�`lC�:� �##G'���֖p�yroC�0��-B�Aڎk�8����T6�0=�$e��@PIA"�;�R�S��ׇHu�yABIJ{X|�2L>��x F�Var��,X�� �"�����!�&���bejN� 7\b?"G��'T�U�dF�+(0(3D0D����@�Ox&�[&EH�yh:��P/��T\�o�%҄����Lu��?�'�ů�G@�ѩAN���BN:$�����L�/��a���t@2lbw�*+�E�Vđ9F)�`J,�6�����	'T���*#'y�aQ=Gl���ʩ������Yx�]��D_N�� �c�/4�@8��09�h�x�jU7P_
��Y#�������i����I�85������}�y�Q��;L��X�|3
���Nʼ�~�Î:��UȜ$6��i��V�?�|�U�
�I�` �C 	C�R/��'��ܫՁ�M�@`2Cb̧�F���í)��}�� �&R��y%g�XQ:ݘV��7|�"-{�'lh����d���g��"M�s��r���J~lZ�&�9+�ta�S��?i�N�F+$��Bb�M����6k��c�JBI�p#��̈́y ��j��$�&\��yr�Aڕ4Ķ�H��T52����ھ�a6�F�����O�|�dJ�p�\ta�!�N�A�G�	�i�c�G����U:t��@���>�,08��Q��.�ѓ�� �pb��ӗ��-@Bp�����C��(��rӉOM�`�&�8�S�78R���'F�{���Qj>��Dx�D�d� �gYZ��Z����ݴ>ᓯO*|�'c�2�z-+�T�x! ��2"O�B$�I���H�æS-!<�rRM��u����{�:�ƫ�gUaxB��.!*]P!�Rii�J%J����>9�B�Y�H�A�-�	:��)��-��h�*y�a
�}bC㉳C�E��h� �B�Q�M�x�#=����<�eb0�7�3� 
@;�P�T�KD��M]��C�"Or@�V	��4��qR5I@ uJe�iT*�򇋊V��A�O?7̓;!�"5�B�6eePHB��H3W�abj�sJ�cW��6��1$�4m�`�䆳>��� !��hC><O�Eq�A�{< ČLG~-�a���	�4��'���Xt���h�6���%	Vbz���E`�sFHONh<��G���ft���"FmZ��`��B?A��
�950hע]%{u�ʧ�W*4���؉�ԉk��I�Ń5�ܺ#.�3�y"`��rMK�LXS�;��~�fx*�,��M�᎛Fg@4�З?5R�c�<=6|�c�C�`Ѫ�Ì�L�Ԝ����, D��UoڧI�<x`Ƃ���Ԓ�o� . R��ś7��h���Q9{6�(%O0t���ˍ�Z���՟=�V�K��I
mغ@���ޏ<�d����׾:��6SlA+�jņ�Tep������B���PxB�F�?�	��!K������κ�M�E���;bŌ�t��Z��ҭ��d"
�����0�Ñ&��EH�^����'�WC�<����:N�0�'P�T�A�k�9(zZ���lY�(��x�L*~F��OKrD�q��&��Z��M�V�̹m�<i槛�v��ه�I)-*��Q燍)l��X��
�rVN�	W��K��R�u=�5%!ed��s��]8��AÉ R�~}����ql���Ѧ'ғV�d��B���t@uh�v�|�j�K:��A��fN&��pkd�Y0CI�(�d��Px2ķuL��B��!6�0��ș�?Y���N�a�-�
݀��7 ԗ5̈�@��A̧u��j4&��eX��{e��D&�@�
�'odh�bÁ��z@	Ç:�L�(�N�k���3��<ؠ2��T���i@?H�x�CI�<3�R����6a݄�¡�3#�O����H ��p3�.��V��~��zbm�Qq�q1�&��k�9�oيgV���D@�l�%J�@���pa��U�@2!�O]8�I��ꛞVÇ��x!�䓋Cp0�`g�_�@��b��R(if!�F���Z�g�8p�g_�>d!�$�CF��צ�[n2ŉ��םV�dŋye������<���M�2&�k�H�*(���I�����Ҏ��<	��C>�N��㩙�5�r�s2�Lx�<A�I�G��� j�-#�|CtM�u��k����$��Ĉ��H���*kl�3�l܃�*��"Op:�� '},�@d돗[Τ�z�
F�gu� 2R�|R� �ꕃ0�ڼR��R�����D2D�h�l���z��U���"q$�O����ή3�H��d��z�L���Q�a���R���v�{�-�^��7Oܴ���J�:D8gX4DG�`Y�"O�'�я[�T1 ƲL1~dч�ɍ(� $Z�O'�'q�-`�ዾ�J�b���UF���ȓA2�����f���S#L~]�H��y�(y��V�X���*�N���ȓl{`��3�F$b<|��6>�RH�����KBk}E�Q����H�i��V�l���|�Es��@�K�h��@#�(���A �;w�*%a�\�ȓ<8�%ɒ-�_�L�0�B�>Х��'1���!f+��*en� AM�Y�ȓTF���#�3!�T#��ÛO�����	�4,�V��2�p	�l� �l���/8�EJ�l�`���B�e�t�*���!/�D;�̽"B'Ѳei�؄ȓ���E�R�Dn��9�9��߾��C�z Y�\�}�\u�ȓ�^]1�M�F���0�Ř\�i�ȓ!+�)юg��m;�!��.���X�V��1n���a�/�R`��f�h���*�`n��������Մ�tXA��.���@��@'��G_L���jLQ���C
�5��B��D���8�کs�!��L$ESa���<]��U�MA%���Ll�D���d��݆ȓcJ0b��
'�;�@\�ޜ��S�? ��1	?#�Zd�b۠o�t�I�"ODM3@�͵Sˀ����ήf��B�"O�݀� pYBPa��X�?о�"Ov�v��={Hp����-9ݰͱ�"O
]�v� �B�-��I2h�
p��"O(:��
�pyub�#C�h8�S"O��*�`��"��0F��~�|Lrd"O,��c��=J����z嚡1�"O����@C�(9�x�(u"Od)i͞�-�XCě=��8�%"O�yuL��>%��%ƙ���"OA��f�1l� �`'ā��:'"O�%�wb��(�0�C�S�oz��6"O�a��� Hp��r�I�' ��"O��(��ܾZޖ����W�]&�tʑ"O��J�.�<k`�	�dQ�f����#"O,�0w��*�T0+!nC�O�T8�"O���%iԉx�!�1/�73��"O�E��
�5|:�qmS�D��l��"O�A	4��-`U`(sk;U�� t"OnU`d�Zpy��[_Q�-2�"O��IU�:'�B�kgI¥";t��`"O��#ј.&(C�%΃'6rU!"OB���̯[�~	Z��X,5 �}��"Oh�,V�]�DQmɛ4@[#"O� �"�J1K����Sh �<�""O|����5/r�8A1,�B��"Om8��Wi�����LT\���"O��� FS�(�2��3��� �"O�$1׭N�)�QR�?:�H�"O�)8׌ѥkS�H#e�82�~�˳"Ob����7��i�ܟ�nA0"O���1		�=Z��+˪���J1"OTLp����Y��҇GH��3�"O������k����]:��8"O*�j��V�B�܅�v��%v��᫦"O①cM�l���Ж�Z�W5�5K�"O
�� ҅z�)8`�ڗ'&�	S"O�xE��:\�H��'H���Q"Or����r�f%C���C�N�	�"O|\ t�8D|��m��R��Lv"O��
&)D�b�x���)j�l!� "O�iQpMȼ�K���&����@�y�
H[��.�%$^�� NǑ�y҈d�@(�� �������bP��ynʷ{MFi0���<��@`���y��4	'1j5 B+Ѕ��M�ybn���<��$	�54��҄(^��yb�,R t˦�̇!��a�ɚ�yҊ�F���� ����(���y�A��z��{PBF8Ne�	��yR�Y3M��a�r��${��#bf���y2nN�R�����䍻D��48A�Q��yR�O�A0�d��E�3<c�P�qb�.�y�d�
~������V7�6�R�ć�y�B�e���;d�J��Ԩґ�ю�y"e�t2�(sl��?����P!΄�yBlN�:����$[7��̢����yҏ��4Rf��� �E���y�ψ17�t�@fm/*�B�SAʀ�y��H4-��MY��]�"'��cЎ��y�ˁ/y4�}�0O�	���W��7�y2�i��4rc������L��y��M?�, iuj�4J�Z=K�N@:�y
� v�ᰪD�(F� c�ߣ+����"O�<S�"ͮ2��HM�U�*�"O�LٓbS;}Ä]*%�BZv)Zg"O�Q釫T�N�F��j��L�"O������%tvu�%��)v���"O�l1�C��;�콘��J�:�5 "O�H�΂��KI#e����DԺ�y�ą%�>�إ(�&Ɍ�8�l+�yҁ
�{����e��V�P��HǴ�yFX�1��U�hتdVd3���y2�� 6��%��#֥j

��F�A��y�d9�!!�N�fPʙ�c��y�.A�4��H�ꕬXE�d+�LM��y2GҔuހ����N�\�Eֳ�y� U^N�Ir���G�4��@O��yr�NWc��kT*G`=�'�H�<��-�,r�����.O���hJj�<�t,ǿђ &&ģZRZM��kM~�<Q硊m��4JoI���Q#�\b�<��V� ���d+N������KT�<7��g���h��Hy\�0�h�R�<A씢]^�ի�1m���t�R�<�"�B�`(DY�	Y�R&��(4hAU�<)�k �#��1����
�vE4"Iy�<���]��XC���w#\-��$t�<a����g�vh� �6
�bmJ%��m�<Q�B��0ĮJ�`a�p���_8�XFz��w���'�`Ȕ��K?�yBa�i�@ � � gv9!�Ǐ��y�*�\ؤ�Ѡ�z>�9�D��y�	�=m�A���Yr�@�rd��y"��S����A��}��\��ƙ0�y@��Y<�-j�AJ�$��E��]��y¤�tr|D#D�9� �C��� �y���e^�[�/N� ���	��y�.d�:�R�J�U��9�BS �y"MV�On�)�)�K4�&��3�y2Тv��Lo:B�I��%�y��ƮD�Xꇎ�8�h`$�A��y��TjJ� 5�$ |�Z�KU��yB@�"��BҨY��X�jW�y����^@���:lJt(#�	(�y� 	'C},����t0��sɜ1�y���=��e Ug[��H ���y�&���y�⬑X�V���ǐ��y�&�M���| $�s�!5�y"�H�vL��s�\+%eA��
���<����
���վh�����[�L!�B�UÀ]P��wzP��Y1<�!���`:���iN�%v��F�l-!��M67�ȅ��ƒX���W�т$G!�8|��,��(ճ�lt���!�������eɚ<;����pc��a�!��$5�m�g�
3q�DQ�"��.�!�ߨv�j�y�B^�c�2��A�!�^�,~�@u �=WM�̸ X���EE{���'��H(�C��5�h4)�'S�
D��	�'o�����L�{JD����?L���	�'`C�F�Q��]I��;IɮD�	�'u4��e�=�T�t�أ2��H��'�(T)DBקm�$ܸ�*��&���!Ó�hO�e�eJ��$㜰5��4}Hn��T"O�����ׄf-�i�Y�g��%�Z�Yw�)�'�حQ �u� <�0���A��5��S�? f� X�YT�٨�Þ4x�����"O�<�D�|9��w���U�p�A"OT� �HE*A|,��*
-��9�"O�$���p��J�0R��"O���T�4�����)D%,0��@"O���u!
�N�ڕ�4)ϯ^�B,�F��F{���BD�LdK��+w�BxRa�
�!���J<�)��Ŝ�%.�!�?T��3*""�Nd�gd	�L���/�O��ɢA���yӠ˸{�`��@(�+��C��-d��:�D�7&`��d�1rP�C�.@T��O�4X|e�p��8_�BB䉡Z�Ӵ��.˸4٤i��[(�C�	m���z�a��-��Pk�*SC�Ib�B0�&A­��!�S@�P�&�'la}2KI&�j�ٷi��HZ�Y&�y"o�*2(i+5o��N��(�i��y�O�q5Jya�b܄D�,)`����yA3����+hq&d�V��=�y���n#�R�'�ehV��0Ι��yb�l���⁒�[��a$[��y�K��� 篆�]�l���L��y��R	9k�Iٶg�%�@gŲ�y�N������m��w�@�8�y"۲[ ���^�a˸�ڑ���yRޞa6��a_�$��$�������?��'E����H�(��ez���Tct�s�'N�D�*�\������7p���'\.�3t�Z3��d�$�V>C]:P��'� �Ė�S��횳j�7�q	�'Z�{�g-���#�!>����'���S��m<���"������'̀|�!
�;
��Ȁ��1۸<�'���rs���X8�lW0�(��O�х�	 QK�}�fn_�I�6Q
�D݀ar���$�^y2�Y2b���C�̾A��xA ��=�y�A[f�@�d��7��8�����hO�����H��L��b��mS�Y����!��\�mp2�@��'l��x���a b �V�����@V�֖~���swo�2s탒G"D��z�߼Id�sd`5 >�$��<1��?�O<Q3�f��e��e��P +��q�G"O�i$�l�&	rT
�;~"�qc"ORq� ��Z��!�)%c".���"OȵK�-�0;Y�x���-!��4"O�A!�ӻRj��r�]5y�Z�@�"O*l��(�g��!d��:v�^M�2"Ol*�MK$�})�]L���1"Oh��5�K�q�L�J���S��Q�"O*���� 3�2�!�l���*XkG"OH��@)�JYBq��R�!j0�J�"O�u�,18k��1�CT'<hP�9�"O���Q�ʍB����̊772@��"OF��6jS�b�Blb�d�W|��"O��2�1�tt.�K�24QE"O��Ѧ'ë J�Ԫ�E�R(	)�"O���Bڀ%Nl�v��34��b�"O\�S�g��j�B�ar�'P (��"O�� �$� xCO�XV4��"O�$˷D���5�d��M\��Q"O�r��$
�ʭ�M�  >���"O��0rφ78�����=W1rT�"O��C�+O�[,��6���) ���"OҌ�+[�v%�����M�k���:1"O� ��#u�cV��jc/�U+~�a�"O��r���
en^�B/�+W#4�r�"OV�
��S� �6P�RNU�j�ԥ{"O^)�Ə:f]�]�'�^?�|S�"O,�yb/s9 �#gO�|?⼩�"O"AYc*� vq��F�`;0��"O��P �G�^itlҷ��3],��a3"OB$��.Ȋe��&B�t��
�"O�y�s��RԖ�Za^I�y*!"O:L)���>Ȝ�P��չ4�ى�"O��i���w�� ɠ �#W�̐�"O�X�k�*>��a%�ϐ�Aj�"O���m��>�ެ��d�s�x�!"O0�S%l��6k\MѠ�F��4���"O�Ų�D�P@ر��
�Rǀ��"O����[���q�#鏣Ƙɬ�yҊ�<��1����1>���8�L�yRb��$���'�9@\�b���.�y��'h����$/3(�P�%N��y���!38�t���*��,aIZ��y�%�l,b ��&�F9�����y2���� �����t�تeE�y��V�cv�z��_��q ��;�yr�R"�Wod��Ã�y"l�!dȋѫkܹ	B��?�y�.�&�V�����U�fhZp( �y�@R5L���U!ÔH9l˷���y���\v(�!EQ
Iv�y�#Q�y��Z�q����AF�M�P�ೢճ�y2���%.
���lЛJ����-��yү��w�J���6�"yIKP�y�#�%'��ũ��8f4i�֪�1�yb D�pSB@�'Q1��P۔��yB�^*e�T��1{��s�� �y"BK�1.�� �h� zNX!�����yR�R�a�6���L<s�Sc�J��y�)ڌ<;^H�cC��_b��cC�� �yB`��v�n����O�1S�J�7�yB$D�2Y[6IK\�MZ�L5�y��k~�ոꑵo��������y2�(!D�)��άg�ڙSd`ȹ�yr��(W��Ţ��Z
}�4ŀ�y"�޹R��YS��&	vx ��H��yR�D�cV�rm��z,A" �y��:S��)�I;/���;�c��y2)J�0����T�$<��W�a�ȓ3��0 ��c2�9����"Z̄ȓ�j<���A�[X�u0�NC����c�}��K��v�`lx�g�O�=��Y��݂dW�>�����.@0lg�M�ȓF��J�@�f4$(�2+Ҩ~��A�ȓG�ٹ�&X�Bx���M"$D�ȓ<�Z�`�]�2�Pfn��g9B��ȓ�� (�ެ\�G��� ��[��;4��:�6Q7�J�X� ���B��ds%`պ%Πr$'��^��q��O�D�j�g� yE�h
��ѝ(��̆ȓE�B��1�_�FoN4�Ŀ���ȓpu�ݳ�삌4� B��#L���ȓk�d9t�I�vord؁�A�956]�ȓ�6aS�a����kUdʞ9`H�ȓx�lȒ��t�,ћ 4/�|A�ȓ�l��B#NZHT����0 �ȓ.	�# H"D�bci�,1G����S�? ܭ�D�D;o-N��6��[\�"O~�"4%�8V��0�vn.ZDP�xb"OZQ��f۹��b��y*F!��"OT庳�G�3�v����;"� V"O��y��V��1Ŭʡg�����"O��e�˿���SK��m���!�"O.]��
<�ܚ'�O\U�ZG"O�T��NHʠɥB� 8d:w"OH�ʗ
�~X��`@��'I�FT90"O0,s��'g�,�E��>�h�h"O�]�d�[�Q>�,�I�"�<�"O2ٰq�ȑ0��y5/��|�vP�v"Oh�w!���Z3DI(m�xz"O:�x%@�?�l�0��;v,#"O숃A���+w��;�cQ�\?�t�B"O I�+W�)O\!��'�\A�t�"O��t�&m�29s��1�P "O~ac�M)BH"!��c^ص3r"O�t���8d�M�b��c*O�``�F�<��
�*N:[��'����Zj.��FA�^o�C�'R���FO�'<h̭˃͘EB�u*	�'S�
�a�d��YP�f��5�j���'�&����f;L� �,^�B|��'�p��#�90R���RnP��	�'�3�%1 ��e��#W���A	�'�R�Sp#�03�)8�a��j���'��r%H��)sP"��6|eS�'�~X�@�q\VA�b!J;.��Թ�'����D�U50R���+&x����'�H��(��H���ԫF^��"�'K���t@�\��B���F�T�i�'V�JC����� @!D8Ԝ�	�'��t�@��%anI�aI�>E��t��'�*�C�B߉�^EҐ�Q�B���'D^����L��E��1����'���!�g�*Q��p8��+�'��Iw��[��q�b[���Yc�'��xA���1g`��wc���
�'�
�����!h�{l�l	8P
�'�t�B�h�:)j d��kB����'�xM�cO��6*4b�
�hT����'ג8P�(qMx���7d/<�@	�'�@ �����x��Ȍ�����'�:D3���I�¼#��-7�hx�
�'�2�Jw�@���s(M6*����
�'߲A��m� <2󄌑4��uQ
�'���k��=qr�]TDJ0�~�ȓ]��!AL�+CU��BE�D�̄ȓ`a�s+Ѫ-�L����K�F�����?g0܉&�K�Bj��a(��K�1�ȓgFbp�V�f�0)vċ�
��\��H�
���i#f3�س��c��ȓ!�\����pȅ�� ��S�xt�ȓ
������L@��w�Fe����B+t�+��@dT@�4"C�c�`P�ȓl�,�{��	�8q4%�T�E��i��~殸C�A��0w6 ��H�"2��ȓ'T�dpU�ߝT<$�D.��/�jh���V��SQ�K޴LJ'��p���1�5{�dV9Ji@L�AI�'Y��ȓd4|L�Lݍ䰙h2CV)7B��ȓF�h�ѯǏ$�H�Y�Ιk*����9AC��[��) @��/`O����S�? |��`�*rO��Q���	����"O��11o�:`#:T*�E"m�~<iW"O�)�gtS���p�T���K�"O"��A�����L�Aъ~d���"O@۶'�l�,�ɆIX��"O���3h�������L95�Vm�D"O��
 ��p'�sAKF�j{�i��"OR��x�T��i��p�F�Y%"Ox *����}�]�F�Fn��I�r"OFU�-���Z�é5y2�'"OL���
$rb�Ac.�� zf"O]�#HɃe�"��Wcj�#��gA!�$dKFh�@Pp3z<���)t+!�D��A.z���|$���F7!!�dрH��"�@V�
�����I��O
!�D�Yؘq��˽x}N��A�T�ў܆ᓑr�D�p�U����R *S���6"OB�3Q��
[��%1��V�"9�x;�"OH��+� ��@��7T$ �"O<�� ��<�+�a��^���"O�\y0'��R���ӹ¹Q�"O�m�����j��1 �Ɠ�2[H�ؠ"O(�Q!l*!M ��Ć�#+o�Lՙ|2�|��'g�O�a P�i��)��#�HC��;�	�xE��')b\#�nQ>󱋁�$y�E 
�'qX88A�Ǽr|��Ƃ3Fmp�'{����m��p@��#���>ݜ�'��t��h��a,��x���<1��,C
�'r�7���}���a��W�0*�@
�'��A`A�>j>ժ�
�1$cxI����:Oj9��۞&�j�V�!'+��!�\��D{��Iݻf�QrTj��JXYXr!V>@c!�� f=��	$ �j=�j�߄gK!�=;�F=�VH��\�1H���D!�ĉ�{VP1���N�l�k����{$!�X xRM9&@?^�$�Q �K�n!�D����/=x|����L7��г�'�<�r�AϷ?8{��<�����'�axR%	$X�eТcH��ఄ���y�ds���v,L�C/�X�a����y�*%ap��U��?����L�yJ�1�lTa��Z�iO@���ڣ�yr�ߗ?�hш���e���ˑ��y���m
F��P
�����B�ِ�y�+Z�?�X���KWE]��I�hO����&ގ�)�g^%�ڥ�BƟ
�!�DR�H����*�;���BuD�?�!�䆁L�eB���p�b˴�!򤊈@LF\��NM<�t2���(�!���bt%�+�쵠�Ŋ4J�!�$��~S
ٓ-=x��Śr�Ōv!�I;R�"u#�-�,D9$F�:uvў����)8�6���S�L���pG�?#=�C�I�-<ۅAכ�D|��+f6vC䉼x|�0�&���>`{n\�A��C�I�W|��4Q�0r�ݓ���fpC��]�(�`S
Mx����י)�4C䉽f	`�CҀђ*�L�:�˸a�4C�A	�a�1.��0A��hq�B�ɇ&E�틷�Әq���d^�]'�B�I+D"�p[��J�)��x��Y$2�B�I&x��%CW�7/�\�J�a�o:�B�	�,u+"��J���Y�s��B�ɷ	K� ��
&o��j�kG"O� J�2�+��H򘻖K�^)�B�'�ў"~�eE����s��k0p5�tŏ*�hO�����'z��qaw�q��Զ�y2V+�u���Ճ���� ʿ�yB�'�TL�U�	�v)bl�!�y��˗������큁�Q��y�/G�]���1�A{�t�@Ț��yB���"&X�z&����<�y"�R��4H�� ]����%�y�h�b: ���o��2��<�y���!��I��A� �ͨE�y��F�)�LEc�����-��(̲�yb����]�w!
��\k�-�yb�0i��)��X�n+!�E�y)CPv|٣���ewD� (�y�II�i���h�[r�!���yR,
�ڐ%�pɂ^��<y0n�)�y"O��2��٧��Q��<��b�4�y�͔=�p]��?Z8&�H@���y�C�ļUh���)M�����B���y¦�t��HF�L�I�V�E��y��y2.��d;7>�hm���y��H:f �@� 9^8��¢Ȟ�y�űx�`�sХV�4�~]*R�F��yүY:�+R�"�Z`�f����yRN�!d����_&HY.qȦ#�!�yR���+�P�4a�4�����@��y�,T�TT��ȇ�w����c���yR!@`m�`9"Lã	4"���R	�':��&�S?j`�x('O����p�'/���D�L"RrX�G҉\��!	�'1�yGNٜT^�Œ�&��\|s�'=�����O���2�`�yC�ũ�'j0<3�� ]�b%ꉮqK4ĳ�'�`(��}�AK��A�c�ؽ�'s��Ac�E3cJS�%�l�R���	a̓e?��kT:d� %I�k�?dʤ�'�a~B�Z���-K�����g����y��b��Ȩ��I�,.���!N6�y��Z�a��)�qሹHw�(�5�]��y���w4`�q�$�L� 蔀G�y�EЦoY�Rq䊳@O4e���M�y/g����Iu�9�����yb�ǼS|��߭A��h���y�ĉ"9�٩��Ո~b�AB3��y�*L�R��`f�� ��y2�����OJ���0��yB�ɜ_ލಡ�n@��3u���yb��)�VD3ňøJ�tU�D�<у��i|����5FmJ�g�L�<i���J3�hӑf
9�0h�B.G�<ɑk6x7�t
�$+u����fB�<�g��~��d/ީ��%H��A�<��S��TK�ME(!��&(�~�<ٗCX5�¨&کU�t���Q�<G���+?�����@;:�Y���V�<�Q
��:Tr����rQ��I�n�V�<��V��i�]	�b��4�{�<��fB?���ѬL��3���[�<	����t�Гl�c�Z�j ��W�<qJ��{��hu��'�0u�g��O�<�@�,F�qp�%F�*�%��IDL�<�������	7�͡�H|�<YCbL)��-�E�4���a�aC]�<� :�23S���#����@��"OF�ϖw/
, ��D	����"O<�Ȧ Vg�&���	nh�{�"O,\���B(M���)���6��4"O�QD&I%tB.X�G
2{L:��"OFhS#hH���h�'A.6&$L+w"O¤@E�.G\M��W�J� "Of-c�NZ@�lK�Nӈ<�!T"O<)�C
���M��fG�@�0���"OXԡ�J 7)���Ԫ�n��q��"OP��@h��V��h
�{�$�k�"O�eċ}��Q�(W?a1V;�"O���t�l����E��� �J�*u"O��(���|\~���e��xKW"O��j�"�	v~pX�EB������R� E{��	�%UB�Rl�~߮�°��c;!�Q�3$"��!Ȩr��
�1u!�䂲m�v�2!�[$?�`�!�IH�O!�W9A�*��a�$d��9�E�V�!�D՗���D�+P�qRba�!��3r�t��85PhD���E�!�䊍�h�E�W�U��m]�d.!�O����I7^,�@��9!�$���5;@��
H�Y
�JݲV�!�יM������I�l�������k�!��3*�{VრDA��h	X�;�!��7,���G!:5�(�j�%d!�$Vg0(���ά]�@��"cP�I\!�d�"�<0�����Z���M�n�!�[ .U�a�W�"o�������Z�!�ՂZ��p8F���$O���R+Y�P�!�d0(���3G^?��AP�	 1L�!�@>B��`���!?�r�`�/O�!��^;l_��"�Ϲe����Ѧ��2�!��! ���q+�v�h���K0!���;p��|�o����PX�&12!�$�ڈ����/����ڵ~!�d°TG<����T	o��5Y�NۊwK!�EY���䪔2H�~p��b!���	xH,t�a�Ȍ=z�]CBmؐh!�$Q��(Q���(pB}�-�H�!����)����}Y ]p�랭_�!��S(?�̐s'�XT�q'j�}�!�P=aK�Ak1�%5lXA���@7!�d�Tf]֩L1 H6hpUh��91!�dđ}�`�@w�@1Af6�(��¹%%!�S7Gk��
����DW`9*rg�9e!�$@�^�.��bS�ES�`�e]?.�}��']�F��FYt Mu"�+@�M��!�M8�Hz��J)�~��!`J��!��1T�p%Bbgڣ<+Jm�3!��Ia!�ĴT�H� �e��m#q�"O,�!�d�.$�Q���U���T���Pz!�ć��V�c֤٦C�Vb�Z�gk!��;_h��R�Ǻg�xUyì\�ef!��.����6Y�K}2�Iu±R-!�$�Ud�	�Ab{��w��!�D�/&��"�D˺j�Ą���r�!�  [D�Bdb��y����t��S�!��hN�y�W��0������&o!��%O�\HES;K(X��"�)Ai!�d
d�� �˂�iD�H�'��v!�d�3&΅��ș�!�2;�eҕ4�Io��(� 8QJ^���b�*R[��	��� �(���IV�B� �&��R�zd"O�Y��F�7����e\.���C��'1Oxx#R���C�A���T����e"Of8K�hV�S&�N'�R��"O�59��	<ԅ��B{i#r"O��0Ģf�8����
!:5�}1�|��'ZazrP�4����\�8��b�T)�y� �:��}�N�a�0I5����y2N��9	&�J�CA�SZ��%L���y����ʧ��K)��I�.�y҄�=�F�P��G)L՘��8�y���1�����(��KRZ��HE��y� Κ+pP��X-} "�6j�&���0>�FD�G�b%���G�bL��f�u�<i3ƓX���ՊL]"�"r�}�<�D�۷k	B ��b�@�Y�A%Mcy��'�T P%ɓJ�d�"ȱ{��b�'�PݫS��K���!D�
3X]�
�'� �I��4o�\H1���7��K
�'����F�QY�R��s+�X ��J
�'|��s�^$�������e�	�'�*8jd]��l�(6�V�z<й	�'�P*`L\
5\t"uc�8~�B$�
�'t��`LC8vn����+F�	�'��<#�ٙ�\��������R�'�쵘��ǾY��� u��?
��4�
�'ˢTI��2Am��s#�& "N�"
�'
� O�T=����8v�6E)�'Ͱ��7j�+@������s^��H�'Q �Qc:�(=��"b���'�h�u��)����d[�ޘ9�b�'��hC����_�bPcv�<��)�	�'&�u� �K�x=��!^ig��K	�'J|ux���B�����ċ�Z����'K*e����=[�hC�)��	�����'���*�aݎ����'�#}�J��'$��i���
V�3,D�z��l����1O�$�w���!O�C�Q�P���k&�|b�'�az��W"�Α$M8��'�y�˰<��%��lM�>�@�%K�>�yb������qP�+����7�]9�?����� T�`T���/�p��W?,���ȓ;Ƽ�2Ơ֊5V6��e�\9w� �ȓ�T52�?�R��'��8��(��	�<�K��_� ��Q����Ҥ��Z�<)�G��1�x���*�(&����m�<��U�x�ا ߻�HYʤe�<�����+�4A8�	/ O<�+У�jy"�)�'AQ@���G��=�w�^1E�l��D�$7�0���?\�����n!�$C�;�v�a��ӢWަ�#�N� c�'�r�'<�0��K��>L�+��R��
�'�z��0FR2 �F�cХE�N+�8�
�'���Q��5Q2����M�Jnf�!
�'>hJ�74Z�񁵇߆ID� ���hO?�)CK�TDX5I�  �f%b��Ls�<�ǥÕs6@I�ük5
�Y'n�r�<Y$�Q��CtBA���	t������tx�h���<�0Z�[ �	�1/�ԣ��x�<�փ�4U\qw�M����X�<i�b_9X� 9{0/Q����⧉R�<q�0���V�٣	��`��S�<Ȏ)�����P�8^�D�@�Sg�<a���K  ��U�*Xm1��x�<� �i��Α� vde�!GW.]���"O�x#^| :�²��a�"ON527���m.ց��Dӽ;~�s"O���ĭʛ^\B��i\%$8tO�UQU�͂��ƨ�+�R���J�O�B�	�t@��͋2��p�D`E��nB�IG�t��v��{n�L
AL��C��B�	%v����F�&5c�7⟜{Y�B�	�s	�8
��Х=�	XRiӈ@lC�ɨ#�hA+�eS�/	�L9�N�?n
JC�Ʉ(}h$	�Enr���a+��B�v�O �O��D<§��hc	%v��!CHla�!��|��x��,ΰ.��d�X͆ȓNba���z]�����.�E��4 1��X�H��9bFN�"B^�%����V������ϓ/D�Q��̜vT�M���5D��Zq��%:!��Q@fޣp)��ڡM1D�� K)h�`KBARXr%
�L.�$?�d$�'eF�d ���C�-B@��'5q�C�4z�օ[��'n4�Ӧ��?,,�B��w���C(H�֍�FC����B�%_l��&.W	hX����5dƊB��<o�Iʄ�U;6:���Ь|�B�I�@(�]���N#(� �.
<mFB�	#J�x1��
��$b��y+B�	��
(r��Y)p���w@҈pwj�=Q	�o�n��̜k��9ׂJ�\�6���r3����!o"H�Z��^G�t1�ȓn�VjA�X��V�p ��>��ȓkRݡ A
�Uހ3�Nb�8��ȓP���2D@ ��,�+ ����1n���ˉk>d��5'>STx���It~�.r�^P��
T?iqT�igb��hO���$��\ ���
Z:.���i�l܊Y�!��@�o6���Î �����-��D��D��d\p�&��d�j�ju�^¤B�ɚ]�p;��R-<�H*�J8�vB䉪�Ȁ9f��4�HH��iƓ_�C�	,Wht���D	X�A�P�<y�=�ç:;L�j�LN�1�s얟#/\���cP�}{a!]�bH�a���z%`5��V0��,=`��!D��~����[z���Ăi��ҥ�L�%���ȓJ|�X�MU<$�����F�%fm�ȓ^0b��®FJ|�:�ɑ"j�H��3@|1�@�}}��J��9vH���ʟ��G�V)��ϟt�"$�D�ĀB� }&��'�>�		"���c�Љa�� ��M�B�8S�E��ղ`��QˢǔqF�C�I�b�|��ȈG/�x	R��C�	� f~����5b���J���/-�C�I�c*B���d	�����k]�@�C䉄p�H��%#Ď]�A2�B㉗�@uzDG�� P��`@.i�؅�9��p�a�Ӹ,UH�J$�_�%r�ȓ߼�r��!;���q����	+D�<�ŁJ1�Rp���G�9ώ`bm>D��	v'�I�ё%e���P�zj/D�ī����g���sf��:א�A#�,D�xɗ(^D A��Q����ǎ?D�Lb�e��	���&�/c�#��"�D�<�,O"|J�d���*���d�,��M�3��~�<q6�va��C����܍-ΞB䉌Q`��J�y�Fy�+�28�~B�)� V��3g��-����!c4j�8@�"O�<�s��!7������=8�|ܢ "O6 $��&Jfʝ�!��;�$�'B:O��!��L�{���A�/֊Jn.�h"O@�x��B�f�~l �Ð5KPd(�"O� �gs7� z�@ŕO6���`"ȎxS��u�p0aG�0�ʆ"O�a����m4��$!�he�%�&"OF��(�{��| ��-)Xz8��"O��w�@��aI-Od�<��O$X[v�5jEz� g,������� :D�����'�����/�s���!O4D��+�EPI��*RI־U�t����<y��������������خ9�Tb�`R��Oz��	Y�hd�k�f��	c�${!�04'!�DZ�1w���EX��%3�*�!s!�䐾U�T���l"l���¢F=�!��'['�eb�k��4���W�!�d��P���iK��� ��a�!�$�>Ծ���Ë"|�f�2��	_��(�B\�Q���AN=q�4��P�)e����i�,�x��T�	ĸyC�1�!�D�RtP��	?!��H�.�V%!�Č�j�Ղ���h��!.�6!���K%�]����N�+�!�A5A��8j�(K)�1�Q"A�_�!�X�ke�5����*{ 4�jcV�!�d���X�#p��0
����Ɉ9.�ċ�x���$<�'e\`����ӑ
�x{V)�*s:`��>sv�+P U'�l���f�XƬ��ȓR�${�`Dd�X��ZD��ȓ�����ɈG@���ԡ\'O� ���I~+^�G��q���m�:��ܠ�y���<P-v�b1.�q_��x�,���y"X� ��q��g��e|�CFA�+�hO����L�eN�9�El�-/S�}�"�&N�!򄉝���ze�U8v�C��8L!�8��9�πg�}�1a۔}I!� %1�9t,��f�����˚QC�{��Ė �L��$�����T,�6!������Wl��47�١���@&!򤜲K]Rx�׎�W&|18�ʇ1
!�$�ڒTo	=>��P� �J���c�'\耘�ɍ(3�!����8�u��'x��7�I�s�^x�4i85~�h#�'�h	z�M^S�$ �'�^�5~~�i�$ qM*���Mۮ�"�E�!�Y=���whK�0۞9"@��|�!�$2!,z��%mǖw�Lr2I"R�!�d[�J��|�G�X�,�X�rV��5�!�D�P���;��,};�e3eI2�!�$v�H06n��&!hD9ײR��{���J2�Ń!�ymvMB�#\M���m�'���Ȣ���N�9��td�����:D���	�&��42l�c �`	��9D���`�Xr5p�*F	v#\��`"=D��*�eM�%��3���.���hį<D�Xa2ŉ)� $� Y�g$}� D������3}�"\�ڼ	7���L=�����\�ܩ�h{�>0F��vۤ����x�d�`��#Ő�I��	80����yr��aT�h ��1I���q���,�y�.AU 
Ɠ�=��zd����y�-�n��`�&/�ج!,ҥ�y
� ��B֐Z:�X�����pQ�"OrL˓J��Yx`B���B�֥���O��?�'f��[�C��fk�J�&x�ె�	R�'ʐ8#�LC�0SZ�{�m�V��=�L>�����0u�@`�f(�9���X���o~!��G���
���{>9@h�.ou!�d�g�%��m 1.�D�`%��7g!�d�*yF�,���ĵ8�~����I�!�C,)��uy7&E%C�(D;���H3ў���c������1����eV�fubD����=�yV����7�J[Wh�sk�(�y��@cg����CMx)`�"�=�y2�Z�%'�� �	4"��P��*�y��ǉ=3���t��7Fԑ�d�^��y��.l��� �1��Z�nM�y"H�o^���d�������d��>��O�QA�Zv��<�"�KjA�f"O
���g�1.���1�"ԝX�9�2�|�)�)�1��ifb6Z�`�9l��B�I5 RhAáP�A.�-�P���܅�I��$H�v�KP�X��E��:��C�ɱ;R�P��.��E,�(R��C�	<A|ք� J�N:r�I�m��`4C�	)G�D���$f�	�f�Ӷ(ޜB�	�Y1�\;'��M:Z��P�Ga�B�	,C�.5�!�&&���@EJʆf�8C䉹"^n���*wl�aȔo��*����R���X&�R�Tl�*WY��sC1D�����W�B�P�懝o��Da�k4D�|P�)��M@h���`C^8�:�3D�db��
v~�$���q1L%���0D�h �ǭ�V���윪d�=�p�0D���B�"�(fGZ&��i�0D��Fn��pX8a��Q�vq�aJ2D�8A .��u,���
�K;qZ�B2D�tj���:O%�DPA炌x)��b0D��a��Ȧ~�I���[�:��:|O�b���6d@-H:�� bH��4�\���7D�ȑ!��5�T��Pb�*��sDc1D�� c�pQ�@P��ϳ=��D
�;D�Ԛ���M�|ٰ��_�����8D��g�F�pʸ�@�+f!���'W�C䉲�6����H ���Y�K��L�`C�I�.�N�� ݤ	̐��ٝ�2C��T����D��0&Jv�ZG��.C�	6�I�#@� D3��V:�C�ɔ5����m��$�����ӽ+��B�Iu\���b��Q:�QDPj�C�	�Z?��y`j�0)����N���B�6���	C�CԾ�[�&��'�B�I4�@��!l	8�a1�'���NC��>xP8�;g�K��H�����d��K���8�!E9X���$�C�>!�ȓE��L�д	e���F*�v}�ȓ7c�����$PR�r�K�+\-�Յȓ��0��J�=	����g���ȓFT��1�C�`��X)�/?r�Nф�nE�&�Ö[uҬ��OU�c,���ȓ}u�a�2����� ud�6Oy�p�I�`��^�)�'L�BaʔdK�Qj(�c��g.���'t�%�E͂�_�,�{����	"h��'���i#���V�P���W&�!J�'�
]���\(�ZI��KȫG�h�0�'-�9��3f�
�3nH�9��� n�:�	�n%  iDo�Z*��`�'y�� oE�iIL�����t��g�O"��#�)�DPA��ػ<�:Iz&g�RT�ߓۘ'|$���1y�)���3�niJ�'�\
�]�BPa��B��.G����'l��
�
�,m�,ގ2PHܹ	�'�ԙ2DKʒ �����j�;� �'�
��"W��RT�Z�+��Q��� �'E�: ��̑�bU���I(���蟴�?E��
H����=���� �b�}����S�N��T�����ĒO��y�*OBD�w��Tq!��T��V��t"O��b�_���I��T9~��c�"O^u��oF7a9�#$��5��P��"ObQ0��3L��D���F$�D �"OHq�5��vQ�s�ܺ2���2�'�ў"~�%�0��q2���5&I�I6�y��u��(�ᗱ��M�� 7�y`�8U]fm����r<�h��"O/�y" I+p_&��k��kg�B#�;�y��!�p��7G���Sj2�y��"0�Upǆ1Q�ܚ�e���y2oϣnhy��`U�$p(�*��?���S7r�@��ފY�+��_�,0; k-D������.hY�.O�x`�l��`9D�(	r�K9����̇������5D�`�FB�N���,	��r$:S7D���A�$&_@p��n����%���0D��X��E
QDv2��Ӵ!��A#Rf-�O\�=���3m?+�2eJD��6a�5�� dNa�$��.�r��t�'ɦ)�ȓFڴ|AR���y^�E�A T�F��ȓ{�.�ӓ��<t���ږ��:&�b��ȓ9i�l���E 0���2i���ȓ"�h��@`�J暭����,O-8q��VѨj�@@���-�1'C&n�p��^���g��!;�9Z2�B�_�`��JN`�17m��	ϴ@RDO������乖nJ�Z�
X1p,J�J$��?
�h`�p5 �	<H� ��0e��5T���.6�hre�J�n���}��B�k >:0�p����0�`�ȓ` ���� ;���Ye�T�Jn����CQ�!�eT�H�)�5��9|�a�ȓ�X�34�ݒ~�*��g�j���%�<Щ����] (��Dg��@%���&A��2(���u�םM`�B�I<f�xr�ӥ|�u��	�B���H� FE5�R]⃣�=YHC�	�8�&�R �!=C8��ǃ%[��C�ɫ��d���R'A�$)��B'-�C�	>�`��S�фdm��	��Rl�?��Ɏ)K�#!�N���1���"��'ma|e�6`�x�ڇd�.3qV�k7���y2M�D�05�B���~�-�Q'D��y�ھ_iLቱ��C
�h*0	?�y�r�N�9q�Yf�  �h���y�M�,]�Z�f��(�2,������yRo�2[jXq���%j���n�3��O�"~�qgF��� �C�4�V�[!L
o�<Q�Q?'.I��,�V�H��B�k�<iE X3��8����3���e@�i�<�v�ȇd_��c��_�v�
!Ɂ	�d�<���bh�`S���P��8�Gd�<� XL�4��Tg��|���P#"O��Y��\�"Q�����`��-"�6�S��@��D�ȇHѶB���Q���'s!��̴=�\A��R-�����4	o!�$�T,H��!���"�~T����8C!�(%P�2B{�$`�j'^!�䝕7/���nH�%p�98�)�f�!���V]h� �F��$
�
0`�!�ˤ�TD�u��/Y�$��ӥ %g/!�T9���sP��5��sZ,�!�@�`��e!U"Z��n��`j�|!���&>�x%��N<C)�Dq���4 !�D�S)� �m�'Q\�:!&��!��B�2�0@�An���s%'X��y"�'�"��`��i��u&�H2l̨X�pТ�a?D��2B�GI�0��(��BՃ=D�(�#FF��H:���Bi:��?D��b�	�l/��	ġ��%z�=Ȕ�>D������0l�P`��C�)�5S֏0D���Tc٩1�Z4�HB�%����T�*D���%�L��~1K�)�*����E*D��2�O-n�r�:1mԿ�F�P6$'D����a0wb�;t��� �aa��?D�ԁ$��4XN��@ß �����h(D�,ȓ�Cx�ms�!Vz��1�&D��Q��H>Y.Z��Ж({�Y��&D�l;' (�ni�ꛓp&ʕ"m?D�\ȧ@�y���z�$���<D��s�?\ ܪ�Ù���X!�'D�З�Lk�A8c)��@^�Ð�9D��S�L� ��L�rGO��&�!���v)Ѥ��Ha0�h�>)�!�D�.��ēR̠A��9�ߏ`�!�����9ٕؽ8!�}@�R�\�!�$J�_��5[rK( f�� Gݿ[B!�S�+n�}I͏�Ԩ�ц�<V�!��$&LPb��ӝn��8)o֎0<!�$F��eKF��(ܨ$U0B!�DD",�L���%���H�K�.!�[!6w�D��/�
"EA�I�q�!�$�~<����$
5�J4AW&��p�!�D�ZM���b�+l��9j���H�!򄃺K]��х�D `�.y����:�!����w�lt��m[�}����/��7�!�Ĉ��ؠ�tc�%�f�zC���!�$Ȭje�u�Fhφc�B�Xs.-E!���>/�Z���"������?!�D  b�
��o�*3�!�bω �!򤈤g�:���&åk�$%Ҧ�F��!��D(0��dk�D& n�xX���}z!��д-�4E0�/���v����)^�!��^-af�ק0!��4ia��	!�o0�`PG�"0�L�a�NU- !��ߖDI�(��%r���2o�{�!�DB�PM��q�)M�/τ(A�k�9`�!��"+g<����'N"��S�!�$��E F�"��J;4&MҧJOl�!��3I�z���.���8Q�sg!�g��2!H�%	��iB#��p!�D��:1��^�F��ш�$Ub!�Ę�.9&����N�8��O#WF!�#ܚ�%�$�j�3Ӡ��X�!�Tk+��i0���x��XFM�{�!�ܥ��l���r�sW+ZA!�� ��z���nF�IZ	?�A��"O�$��h>O�%�ͷq#��ɳ"O�Q��иZ*�x�O��p��*'"O���ޗ��ꀯ��Z򞵹W"O���ǒ�cȬ�� ܡ0�V5x�"O�h �7�^i`/�&!��QT"O*q2��ǲ{J:�k�$kƈ�"O��։Ɨ)����ڴ~A6$�s"O�Ix����5�`a��煾{Z���w"OZ����D�@��4�Є�5,F�J3"Oxȋ��K�^7|�c�㐱{�* �3"O�rH���K"˦|rNA"O�8��D�Vj f�;-� �P�"Ov��AB� J�Am���~|b"O@�q��<tS&�P��^�a�� 3"O��0����r�� ��O:��B�"O��{'�js�PH�D]���b�"O���1��-*�K��-8M���T"O4�QL�F�d�CF.I�u<h���"Or�0�i��H� r��:g5`��"O���dO�^Q��RҢ��:-ibP"OlXde�_�j	r�� a� ��Q"O��2�ǵ�JI8EiԈD����C"Ot����?�R�R���:���۳"O�����U�X ����+�8��"O&uS��B�2��� �]Yb"O��2�,[�k�ڄ��c��;��[�"Oh�
�ZP���F�ؼ!��P9�"O��ZV ��.J�Mj4(XB �T�d"O�P��׽gۄ�a&�� z]h�"O�m���m��Mc�b�2L�1��"O6���(�2!Ꚕ0�/�[��} �"O���G�˙vAvā"Ύ'AQ0�:�"O���'��x(�Q���(Sጁ:P"O:qy@#�85!(�ps̜�:9�hc"O��Ӣ�<5��P�N�kW��q�"O����_8[���٣JU�Y��8B"OB����U� ��I�f ��"Ov��/�jW�4n/�ͨq"O p���T� ��uo�*i�(�$"O$�x��O95�D�1�CQ!6�D��c"Oh0��D�eu`�H�/#
���8E"O�M�Cf���1�N�K� �c�"O�U�Ơ����	:{�H"O��S5��Z�a�ֱ]���"O�ɲ����P��i��"�= {����"Ot}�EeV����� K�+�d��"OH�z��3Lo�8���?����%"Op���	[���(��h�1D'p�`0"O�N ]�^�rNzx01P�6D�� ��SBj����9�ڥ9c6D�����[�qWj0�WbO�vز�A2D��
��	L�����gs�)��4D�t����nEֽ���[Z���j!e2D�ad/� ;� 92�W[�x=��'2D�P@"��G��l����Gv~��$`5D�x����x&����e� sL˟N�!�Č%7���#�!��t��&�E�.|!�̘k~�*$.�.�u#�6!�ذ�L9(0NN���cb �7!��Ӣ;Ū9Q�d�Y�eN�u!�$� �Ll���&(c�Ӱ㞠W!��%Z�Q��ʕ?��q"�~D!�d�k�����T�c�D�Pt��~$!�� �q0�FT��5���}ۼ�؀"O�!EB�KVt��p�_�L�|\1�"O�T�ѪϱZR�X�Eɡcմ��w"O�KEFB�$��M�5�2W]��	�"O�Et�4l0 ��1&9THC%"OZ����aH�#�:7�U��"O��� ܢ"Kĭ��*ǐA��"O����"�-��p�a�M��8LX�"O�ui��G4VG> ���_< ����"O���m
!`�����EȕW�ɀQ"OҰ�(ȴy���6&E�f��y�"Oֱb�MMHR0Յ�(g�e�!"O̬Q�NA��-��FI�� UZ�"OƜh�C��mS��߅Cg�Ix�"OF���Bp�H��M_PbD,�%"OF�q��!��d���׃/b����"Op!(҇\�B-@|�x�ڶ�e�!�d	���5��B|ځK�G�|�!�D�>��a(T#6y�@A��ʐ-�!�.��������3@�~ !�D�/����Ȕ�� �
{!�d�
f�ɢM����%�O$#!���E�Ai��C�+���`"�z�!�4������M�*ab�G�
h!�4d��A�_vR2��!�K�q22Hz��F��+�!��� ���C���z����
A�!�ɼLH���C(�� K\�=�!��9y �
�8��r��L�R�!���8�
\�F�s���v!����R���O� �SV`ǔF�!�d��vZ�ѐgGϻ9��=�T�P�@!��"t�����Ό/��x!i�)5+!�[� +���%t��jR'�3'!�D��Nx�'@�YvRY���4u$!�M�}�	R��Y%_�>�F'M!�D�r�<@7��9Q�FyS�_l!�D�
z\��S�CZ�k��8�v�]�*c!�-l�Lc�(�M��QYq�2Zf!�D�61H�� �1�������,O!�0v�����Nk@hzd.P�|?!��t������3\���M��}3!��0x'p��C��G(*��R��k*!�DH4[�򹛄��b
d��mʋ!�D!
����P��<4��1�@�Ʌ^�!��Y0inxQ���hr����!�$�!hY3�dB�$����Gn��c!��,
����*� 5A��˛TH!�D��� �)�2�hZ���21!�=eyZ}�p�H����`��?S!����ra��@b
�h�҇2!򤞴o���.�'0��LjD#ߥR�!�Y�ZxZM�G�P���*d��?�!�$U�t�`y���ݿ!!r�j�(�V�!�$��<a���%	�%�܀�Dӫ_�!�dS�[rYcE��<B�R��2,�!�RL2.t���"��yg�\'no!�D�1@�$�«R�QD6��Ee��1!򄘠[�񩄮E� $���BE
-!�C.SF@A�'ĝe��Y�D�A�!��˧
�̥��:����#M�'W!��[_�����s�p�&��5b!��
��8�R-�>4�W(uu!�d�<h�*� �z͛ŅѶ`K!�� �e��)V�eaf����\��c�"Oء(A�F�<mj��d�Q.*�fӄ"O��1M\$����tɶ]�r%8�"O~	ɗ@�sYjW�&�<ݲ")E}R�i�a}�ԟq�]�UcS&�%f�M ʸ'����%?�sFA�j�(\��g�2(�gD/D��r�_V��B�ʡ=,�D8h+���J�c�@79�UQ�$ ^�P�"O��Sd�U$5΂Q���Ϫ�|� "O�5�A���C!
�I�7&�h�� �'!�DG����ËE�G�6��f�E�tO!���6��hJ���i��n8!�Y0V�6�+��� ;S
],!�DE�l������?�ZSI�!�D�20��9w+��0Tk����k!�&H��x��U�!��}"dŎ�Y�!�D�|/�����v�Ԥ9r�!u!�Č1fV��f�b�8�31#r!�$�./(]A�> Ak�虡 X!��]M�~��Ή1<���ʲvS!�R/)r�[L�&E��c��5z !��[��pX��b{���w�R�@!�DJ�+D`�򧞢[��ŀ��S!��&��Y��g�V/PH��O<!�ڃT̤��2C���B�B0���b!�L�-F���������qH�/�!�ڮFM����8�.i�W�V/v�!�Us���q�I/'P>hQ�S�Zs!�D	�D���w��>���8�,ֻ}!�D��f�V�	�2S��y��6G���̇+�6�)G�?�Ĺ�w� �y�Ǆ�u�ХK��ȉFO6=�V�ʣ�y2���Iw~�B�/�8z��u���0>Q�'Pp�	�!`��-V�M�uU=O��B�I?1��=耪Fnd��B���;BȢ=Y�'M%B�{c���K����bC�B�ȓC�.T)��Qv���\�s@�Ԅȓ`C05�w ��G��D(��=O����(����J��!���$&�:XQ���ȓ|�����LZ<����1�t��y����0�F:����d�ƮU�0��a$ ��^!<��p�J,i" ��Wv `v��1X_H�1a���l3����U���5鑲 �6YAa�����ɇ�;����o[[��!�,G+1H���:k�(��C��;E
"J`%���q����!x���)�e�5�̆ȓ��M�UFY/�vԩ��� F����hO�>5��F�a�f1��߹~�	q�8ړU�ў��X�e�oШ)�4�գ�`܌�'$a}��ƮOTl��DU=}b���w�U��y�,Z�VOzh��%x?$�0�@
�y���9���ہN��o6��2j�
��'h�{��$�z!Pd쌋;�T�Q��Q��yRឭ;�8�!q�;�.�qqI�_�9�O~-�08@�֍N�� �'��I���	и� Cܺ����F��{�M��4�p �bdEVʌ;g�ˠ'0n�FyB�|�pGK�VpZ(@�8o�.���L�t�<�#%ƕ)�P�"1�Űt��31J�n�<AU��5-0�И���ky��B���Q��hO�'S��IrC	J�����(FzV܄ȓ�|y��/u*P �;Yf*�Ez"f�8����uW(N�����HU�yBp�)�y
� R��%���<A��#/d��ik���՟���O`�ק��M��H�K�t��/���vLH~��4 ���ĕ�)I(�&b��D�ᛇ ��ik��h���'��'
.x8Nϵ`�TH��S�wp�Y	�'.��)	����j�jG.U�	�'���A�o�Z:@��bZdI �')�O�s� 6Ռ�S�Lu3��Z$�f�'��x�G�$h�����6�Q􉓪�yB�)�'a�T]��81�>쉤��M�AΓ�p>��J}���N�'���8��_-
t&�'�1O�qr�ʫJ�h�3Gξx��98�'w������@}�"��t�����'�f������ᡏ՝<��(��{��IJ�U�Tc��SE5F����0�1�O47-I�T� 1Q5�`�`��`��6N���=QJ~�e����C4��T�E(��M�<�6͔$K�8�ꅚ	V�\
Ӣ�Ǧ�s���s���k�m�?�ps�\�~�F@{f�'-�I5��@��[�#:l�A��/NV�B�	,�k���9c�@��E��G�Σ=�L<Q��t�������ǊZ�KcԒ�y��G�	�%�@,��Nn�#�h/�y"���be�4K	�*�|������y��)W>p��I�
��MH�$̮�yr�![�pږɚ.r�X�GB�yR�+f�2�!eaW�jDD��m��yBiQDX��[�����k�?�?1����/�@�#Qg#�(kˎ;,b�a��or
��4��{Ͼd���\�v����?��(-H:t�"�Iz�)%�K�<�rN�����f
J��T9��G�<�UD�4�����,ں�2\��B�I8`��i���U�Ap �E/·B��B�I�ptZ�i���3P�6��VO�)yޜ��D �$G*�>�c�U9�*`ۂ��'��|��׾$ʰ�E�N;12-�v�C��y�B,����p/ߧ#d���F��p=�}��F�x��#���QV�	��Щ�O��=�O���!�F�F�lЁ��#F
F�*�'�l]�ӀS���aR�@˺}P�'�(# �5k��t����9G��B
�'��0M���8�#��S:}<j�s�'��������$!֤O4o
�� �I�����D��<`��I���%���R�ͅ?$�B�I�74L���O�8
8Z�I�X�m`���6ғl�"9w�;v"�黄�W(Q�`�ȓ/��,�r�6b�ț�MX�2ֈ��ȓ0>�A{�F�!b|��m�����ȓ-1�\�Oy���BF
=p˂Ԅ�w"4d��ƐDrB���M�6-bZ=�ȓt�m��]�:�*��Z�1r���	g�T��츤`�� @�jӃ8��ȓyFt��d������G�u��&��y �G�8�$K#C:���L�� ��ꁑ#���4�]���l�_��O#=�I|��*҂(,Is��6)4�I5�w�<��B6{GZ���/�|۰�Kv?1�'��'?���ɚ�Wt��R��fl#K�'�!�B�L�0 �!`�O�0����ɶ�(�'��6�O���O
(��J
?.#�	���aV���"O�ĂP�S�+��a����D?OJ����:���.@cXf���Pv�!�՞XP 1�r4<@Z��ny!�$��S��`K��P�,#�h˒CIK!�� <̠a�T�J���bX�XD�\h"Oơx�(�lgF�s�@"h�Ia"O�<����s�X- �bѲO񢬙�"Oj����J�L��A�@)cb�K�"O���b��#����1� B�"Oҽ���p:u(���S�X��"O�i�5��>J�8�X�LR�Ԛ ��"OL\�u�B/IDδ��Y'~��S�"Ot��N1d�)@4������"OR�� P�T�U��M~�i�"O�8��:N\���j:C����"O�� D�'�2�g�����b"O�)9�듘-��<���݆���pV"O��H��5}n�r�Z-g��{ "OR���ȢY�L����Y�5�S"OJ��ch#6x�iw��:-�|L��"O.��-��*bG"˰}�scXp�<)��֛Wc>lj�FO-�i� �Ho�<�5hӨ �U!U��r���lB�<!1,_�hM �5�J���� ]�<�wMTk��*"�F:H�h���PF�<��̞C*TZD��[�A@�ʘC�<1���e���� M�J, �)�|�<��4��|����55�,P�w�<A�Q�FT�p�W4��cC��N�<�D�	8�hp��I�]B�k��I�<�U[�1G֭� J��.'L`sEhIF�<yAMd����{����t�Y�<y�ÛG�]��j��l��F�<q��� �31=����l��+\��sT�٪T�.L�\���&��ḣ�)5N����ԵL�T��$�L��ȓ/�l0z�ʎ(-" c���T�7D�42�İ^�r�ɴ(��H�p�
�g D�����U2�҈���l'�5�@)D�L�
W!�����I�rqx#�s�(�'M͂=W.��T��0� q���6���oU�L���P�\2A��P������2-
T�`�ݞd�����+Mhٱ"LT�D]")�5�U�ȓ6w��
��B�	e|��t� O�Ą�<�9�ć*TE�<2 F��]��P�ȓO�L�ZQ�RwBb�#R�.P ؇ȓ2y��x�G &�1R�@��ȓ5{�CU�N3;ט<do��KJ<��ȓg��tcΉMلC�m�cR���aڰɡA��o�H�zѬJ:D�p܇ȓ;V�'�ƛG�hL:d�A:v-F8��G�`	��D�<MO8B��<���E��0Z�#I���q4M1���7��A�ށY�,�Ү� GT��ȓ	��aꐍG*aP�٨#`!jT-�ȓ^��Q� '����"�W%S���XȤD���3��@qU+��=��ć� �&��F暯f:��/_2'`��T^`���3�V%(ÏG);jP�ȓ~	hQ��%S��Ah�K�)�,��S�����Y!Q�����UqP���2�X�"���Si�7�Ε�ȓ4P�js��.@"��d���\Pt��ȓz�x��ղ{���5��ui�%�ȓ&��8���VO��pwGY9�ޑ��6G���բar �W ��V,l��ȓqښ4["���0�֪�2z Q��"͂e�g�Q=D�I�G��3p��ͅ�S�? ��X�C����!z���3`"O<�@���"=��Бf�/0��l!�"Oʉ+�`�<���A얍D4n-AQ"ORphŦ��v(���#S&2,3�"Ol��(@_̒�p#*&p���"OI���b�B�숼i�i�"O�������I��k��/6*�	U"O�#@or��l�N�̓D"O��93Ɲ�\ap�K	�r�P�)�"O��X�ڗ>�}��� D���I�"O��č [��'J��D��C�"O2رCǹY�vL�siP!z�,y�w"OI�a�%AIH���b�Dj�"O��wH��U���P1��I=��kG"Ol"�J�>4ٜ���A�����E"O\)�Ԧ��
�ش��eײ�E��"Ox�"dj�%_�<i�^�.�i�"O����X���S�i	F%#6"O��`�"~h �%Ӑ!�j��#"O~�(,&w����ffۅj�RH1"O��H�,����ӕ+�b�Td�"O
A;�i��:<���0q�\d)�"O���� �}�p��R>��c"O���:����E��0�h�P�"O\e� ��B&ȡ��M�K�V�"OȐQwj��|(<E;���R"I�"O�D�k�'zX�u^����υ<D�t)�A�M�]���&8���y�G"D�t�!f�f�>�+w�1�rm�.2D�T��2\��`ʗ!r�"	B�1D� sC�Ђ��EzA�0{���k(D��x�-�U�<�U�P�9��{�'D�lA�Z�~8X���"|�`���8D��+T���O��8���x��%1�9D��#�	�&������jM�w�:D��� AهWK�Q3�k��O�tM$k;D�L��L�ws@�ꑁ�)+�J-ˁ�6D�,��Ɉ
�.�2��N��Ȼ�/5D�`G�.��H�j��pl���7D��[�S=�M�Í�8�69�dE3D����셤W��I�	��֨��.D��7cT/k2-�2*>3?D�C�/D��
����p��ōlB"���+9D���R$.VjP8B�^[z�hu�9�Od�1�U=�yB
�H�c�K h��L��C�y�-�	��lT=W�&]��q,�"<�E�?�`������R���sl��R��8�)�d�ޅ9��JQ؟��A�Q���D��~��f�U�"��"��[B���iL�#��L��Iĭ^ 0�����%Ϲ�:M�@k3D�pk�逖ae�������bw(M���O
x)�Y��9���qO� �cI�|"ħV�v�\�G�FHX82���a����$�� 5�� �g�z�tpC���*��8C�cԴw�����'�ɺ}B�ӏ��O�P� �A}��̱5ދ2�t��V��/7�2������/M\�'i�V��8E�I�gፕ:I�,�*ĸʆ���;c�ti����@��/�8y��cF�F�sD���.�T?�˟�<��nO���$c0�,Ч?��E�j]#U:�B�Ƀ=Ղ�N�q�š礌VC���P,K� @w �}G�PDx������	:h���D�B)^؈�S��."'�����?���
9n��6���.9J$)�(lbiC��J� %!�$�3I ���ۤdKڬ	u�= ���G�d��gA���OJ�1{g��7�5K�ϳeߌ��
�'�$!{fHζ;�P)�w��+L�D�)"h��f��t�3�y%��S��?�S�
8����-�	{�Tzv� >�x�S.�Y���� @ FL��򭄔`��1��-;?��e�+��kH>E�� �4@&׈?\5Bl��b�P�9r�'}��i�@	X��t�P�؟a�M1���&�" %�H!�+�'%�.���%�P��D`hEÓ�9X@�C�		Jvd��J�aUp��բ�*���0!�G�����HS.}�~&��"H�>Y��*΃�!:�d�Bh6���2�<	����g>�Mץ}��p�I��=�di����#�J�ӑ��s�4�D�ĉr���G���m #$��"��q_*�k��Ҡ>�����䘜G@N�ȓ>n�X�Y�%!��68�ȥO�=r�"�*<`hԩ��-�'A����[��$��-�{Z\��ȓ.(8�B(X�m�Ԑ��D�Am5�"�B�#����9��|B( �'���C�����>���,,�Px2 	�	03�ɬC0���eP��B�� 	�6���*�'p�b�+ϕ$�Lpb�εS~�
Ǔ=S�4b���9�JY�'�Й��$���qAW<M`1s
�'����q�X�#?*�p��A�B�ZP)	������(�t#d����S�����ړ���&u���÷p%����3�BY�pKǦ�h��g�\�Z�&
j�v JB�JҔ�RUD-��I��(AsR�P�3����6=�!ȃ�u��� �}f�'�4LS���0� Ȁ�B&&6q �^>�;`㒊h�09y��OE�4��'M�|�\�;dB���e��	<~C ]CJ֊oR��P��Y�}L���wD50�l��fe	
͒E�g�<}K2}+cZ?�`�<O�@�fջ�刦	M|��e˽a���G!vZR!G�υYET1x&�]�QW�[��t��d��Ue�q25e�dP�l�XA^%�=!�34$"�*�#(C�� 2��@8���`�]��C�H�Yd��V�M��j�k �4��F�k�j�4O�O.M��@��p=ч��E��w��02h� Ʌ�i��T�bn�$a2럼Q�^��#H�Z�D!f&m�����<����)C^�"t�M;e��3'�6D�l+��څ#b�`ѡɓGH��J4�ӴQ��Ax�&�$� Y�٨@�(i�hZ�!c�S#&�@nz��gI��L��]bB�F�B�1�ģ�`P(
��#D卡7J18��8S����`?@Q�8j��ՁF�ΕU���		��4��c�
;�h��I�L�<rN�,h\*<��	�1��5PRD�]٬x��F����GcDn,�H��H�.9Rf�[?y0N��a�	&�|��0�� �i��t����T'
�2�Ov�����	�"�Y�H�!X�����	K�Dmn�6e �4�x��
`CG�(�z�.�}�<YPJ�&@/<L��]*h�a�e�� �THRDBB<����!bW��
$D)4D�Op�G>�����S: cS�P�4�؍��O��$�G�A���U�J+ ���ĄN�ؐq4)
�F��tb=LB䙄omA𩐆	�Bc�(�-[?D�ȥs%�M?z ��$<O̱K�.�K5j$�U(ŃT֦��
>sG.)�f%q��ʥ/��L�T�k��nY:	)�J1LO���#$SX�HZԁ��i�4�|�!_�e�@vf�;I$��ՏE�@���M gl���ȕ!T�x�a��q�DMo?!�䆚O�`� @$�?!Ј���6�z����V�Nf�[�m��$��ps��J�p� `T>!�ր���ڡN������]�.�Y�-�ph<1���j�,��AD�3�ZY��;d�l���B*$D�qӨ�*)D�#�J�i�"��!�D���'GTD�p�3� �C�8�`ӓG�qc��x,��C@ƙHҬ�8�&l[�L�8T��dd�!�Z���ʂ�g�v���	�����F�P�r�c`G��VfqO�9�����2Hʴ��fV�|2x��㞂�M{E�IغS�d*�<�6�I��qT(Q�<L,V�(5��N�m��Eс�T`�f�z�
R�Co��vN�=F	���'}��Ȗc��D=��!��-���	�'q�]@�%���R���%���0X��?�qn�!h�\��j����z8$�F�M�ؙc5�A�^�������ywV��`��7�Pi�j�'�����%߇�y�iz>*�P]�0X�����y#�&a6���s�l��9��2�yR��oE�ŭM:\1ƈ��`�>���ַ4�t� c��Cx���Т��4 lA2k9d�ޔ�' ;�O���� 7T�TeG�T۬)��ݦO���a%�ܰHW!�0L�d�N·wv��c�R�{'����*��]�� 3W�;�S	o�(�(D�`��[�Lp�B�	�"��	���f_$����E��6�D�>nD\#pJ&:<�)��1s aF�1Ne��l��k/��g�-O��	'�I!ܴ=�3o��I8Q����T�F�xL��0r�7n樆��vs�qi��(
�� ��
l� �Q�sA@>�~����{
���s� PИ�B�^����qk@�#\�i����MH<9 )*����)�/?z���u̓>}򜉀�5�l�����S*qB�\�j���e��X��K<	"����Zt���qUnҴL�`����Ə|�t%"��U�"c�"~��)�*۞�Ƀ�ݽ��6g���0<�­H�9���pY� N�'��Hr #Aߚ���)D��@� �reN�2%~=��8?�T�\�fO0�"|*�U=�Û&��u�Aq�<)pn��L��BНS�\�2 �oܓw�h�	�%H��I�%����冒|�����T��a��O�v)9S��}�B��ȓ8�������	�R�2��_��ԅȓV ��)դݡ[`\��6M��"D�����&�B�-�r*�C�a��l�b��ȓ3�z���.p�0t�B�j���ȓc�64��GF*ct^Q�F��6�<x�ȓ<�<P.Q'!RH��"�qXQ���l���$E�b��%4���<�ͅ�C�|���D(ee2�O�@IC䉨i��A�GN݈o44�3�OzN(B䉨oP@�
���)3��
�1<nB�	� ���=���%oU�7B�I�P�΀�4aS� -�1����w�B䉶b���PwE�/U�����rg�C�	,d�$eˮ0�s���&��C�;1��"��4"�<E�!o��C�.�t{�.�*M���!䍞N�rC䉗)�����.��ACgꈈ$�NC�	>U�dPp��U�e y�`"�+fB�	1m=\��ǯ��ftn�uAT<{�B�I>�XuP���+ ظ���+P?(1&C��HA$yB�]{v%�� '|JC�ɛ�,ˠ��)�*��Џ��c�4B�	n"^I`D��"r��3̊�/�VB䉥xʦ�#(5��Tr��K��VB䉆�����'CP��֦�i��C�u����d�ո~�>��D"P��dB��p�h)�����١�"HB��������mDڥà#	�4j�C�Ɂ��̃b�FYVD��bF�f;pC�9�8�s/ׇ`|�a�ß�'��C�	?�p��3b�q3!�.]��C��&��PrE�� ?٦�����2D��cC��9r�@�a.V�yј���`6D����I�.�؂�dR�W�	"5D��k���4}��T��%�`��G5D�{c�ֈoY�t+BM��^���`
1D�(J lΙ8%B���R#y��x�w#/D��8�*ʢ<u����\�@D{�.D�4��S
�Ѐ%(S�H ��E-D�dS�,������c��,��$K7D��fg\�p��qIC*��]Q��)'D���׏T���Ѣ���C3��[tI6D��Y�M��F=0��P��Es��)D���Sƛd��5��R!)�0zeA&D�4�a[F�z����D1�jTз1D��#���6I��	B7�ue1D�|��@=S&�U��e��0�Q/9D��yF�V0u��!��I�Xa�|�ƣ6D�\��+S=?��d󒍀XBJ�+K.D��K���8>.Np8�mS/b�@���/D������+�s�1k����0D��z�(v)�%�P�Χe@����$(D��3E�";1�!�7L�Q8�1�'D�� �X���͋.�YRG�;I�.�	p"O��@B/uhTU�� _��F"O"0J��\"�����/��]���'"O���H�K0z��,�.��t�"O�� I��bd4���"ov���"OФ1�7]��p��O�4_~�T"O��"gA=f��l�Į��F1d|��"O0��#�~��*׉���3`㞓O�!�,2=��Ҡ�@�c��I2!,̌'�!��%�@����8�E�����!�d�w<�"�cG�lc2峳/��(!���-`f�<�w�}�a#+�����z	�'�艓bFQ5A�\��ԯ.2�QR�'�����n�%��OAjx��'����k�7~�z��
�^���'�"�Y�e�(.%� ��2�T�1�'���L��I2ic d_Pg�m	�';��	'c��+v�D�ZWY\:�'�T�#I�����4��*E8�T��'U(EB+LþI1�-۵i0��1�'��a!UAB�8B�dI��B}�V�x�'��Q��+Lc��Y��h{D4��'�0`�5%"`"`�t.ݔqRH�H
�'���R�\�4�H�˶���rL�'%(�C�(�O�I[��͎��M��'� �7)N��`(��Nʉq�4���'�8y�"%.�&�#�A�sP49�'/,8ʦ�OeV��+�	=5���'��i���:Q��*��)�I��'u��`�ɻ����ɖ]���'��q�Hǩ;�h�q MR�l(�'j�9Zŭ�rr\��a��C�Й�'�pʅO�V�9vB�(��	�'sL$ѕ����JiR#���:t��'�<Y �W��ܡ""cզs��y�' e����{��áD��Gz�ِ�'�Ȋ��Z�J��▆԰0p�8�'u�E��B�^����5'���(
�'nbI�r�֔0�TY` �ֿ	����	�'i��q%K�u~Y��̙;ۤٱ	�'�Ģ%.b�E��F6,p�	�'�!�WE��;X���?]Ld��	�'\�(D��K�e����($�rd��'�,�#����mi�N��B#���	�'�� �N�j%�����/t�|�	�'��M�'@�}�v�I�%5<��	p�'!R�pB͚,0z���͂�0��x�
�',S�Ċ
^C���@�,�
�?�(T k�t�����l� *��L�8��$D�L���T*f��Y���z6\	�#%�+�v��r�)�h�^Y��Y)�!i�
�4� ���"OX�с���d���^1]���`$�_�Հ	F�I���@��~IĈnފH!ee Q&^=�SeC��y¯�3�zQ3�O;Vp�@�F�<!#l�4i�SU'5m�y�e��*�v�P�AK�����_#��=��l@��:�((ά�%�A�*F��P�@�>i��,$��k�èpjb<�R�8~����� �Ivy
$h���T���X��	�+4�ʴ��M�F�j�P�Վ�!�R-�TL��c��[��i: ��c� y���ć2N��5�f?A���Oh��%�%;��R�,#RI�8+1"O���+�u����W5b*fd�&�'�j9W��\�fes���VX����Ҩ 9��Af�Y04�f��>|O�k���0�ٱCCҕ�����є���93�W�j^�I�	�'��P�+X6CQL`��D�JU@5��������&ֲh����~� ��9 �\S�Q�aB��0�T�b1"O�5�5 Ԯ�J�!����J���A���]F�� LD>N|����R	��A)��i�h�
��#@9A����bJ�0?��d>F�9dh��PrR�X��a~b�Ч���|��i�e h�G��yj9���uf�~�)�|j�Xb�Y�D���w�=T��(�`�U�I=��!*IIr���wrJYsVO��9îq��;��B䉘=�M��	��b<�+?z�`��Q��%��$�|�0��~&�X��I���5�쀹;�bԊrg'��R���G��a��B9\�|k#șbJB�X�$�SI$���	,$�Dy�Ïв=�Z��T�9��>A���'�R�T�����2'B�(P�$�(�ȓ&�ڹ06	'n.�S҈<C�O�H�$ ~� ��d:�~^�P94NK;%��K���\�A�ȓ�qc��'k��������҉i`� 5��I�%5f�3���|R��U��1�ťܳ�0�!� %�PxrlH+f���h��E
T-�� 1H�ON��2�_�s^V�P��'�9�i�>z�ı(����ͻ!�'y��K��Ļ#��й(O�t��EA�a�m(��͘9�*(�O��؁�e�F��!<0z������X�@*X�sC��lzӧ�Oj�����x/���.Y'_��,*˓-�V�s�2��I�/j|*����x����Zn0�벖|��Xk:c?O��1$���<Nn��Pe��t �C�>��J� 8�Xj�0��i_�1��O����M�U�7�z�Ӆ��l������G:�lڤA�-rZ��reHs��[��>A%ʒ/�p�>�O���a�xnL�I^)ȤX
Ot�� �(@����E���+g��b��{�$�bt
J-�0?	�I�/}J���ʓuN���E��y8��eH��,C�%����:'جl7��l��9�t�q	!D�p�K�$O�}b��A F���x�;}�$[�E�Ms��
w>���IS�t�A)��(�jy��e7D� qT�P�����[�aF���`U+$��O�H���@�Ӹ��;��-����dq�� QJΑW�~�q�Q�Q��mdވ��EԂ"ެe����$�m�F�ڸ'�2|3��	Z�0�� �&K�%}b8��7GU�g7���dI��d��*��S�iit0 ��	|x5�Pi��� ��\ȃ��G��Ȫ0�J�J��E%�Ih:A� �,��5Kn4]�`,����-�"��d��11� ��b�A�lp(�U���3R�e�"���y���'4bQ0J�y��x����Hc�>i�GCx���(@HE� �OT����3�~m`�N����JbNY�)F��apO���%�Т@ԔccM�pQT̈�<^�5�a$��4��dEz���ۅmѡ�8��L� ����׊P�UN�%IX�dat,<O�D���&OR�pq�'�<�[U&�$��詤���8q�`��E�Qo�e�P��Mf~U�3�'��0�h;]B.���Y�FI���I>�Egْ@E���m���:酬>��(r�Gi�J�i��0|���1��2yh��ǂ�`�<�m�4<�D��C�{7h0�s�P�k�vQ���O�̃�C�&�@U��e&~�'gw�<:�w3PE��dպ2�rl
&�h��A�'���qBֱp�Q��_4Tj�J����'f� ��t�b��a������u��g�d] f�h����	~DQFe\q�azb��:�8�"^���5f�ף��F��Q�*('ys���.r8�$��N$\O��	�(T
~����փ1/R1I1��A����,O,�!��,eT�$��M��M�P��g.���HE�<�a)�PI0��w�&��� �q�1O$��F.@�s��R��vfD���$Gp�	x%#�z�<q3� �Z<�pEC"h��ÒS76�:-�=���;�gy�ǎ�\�6�ֆ<MS�L������y�ܞxql���BͱN��Jv.D��y��M�-�d��kQ:.�P+S)�yRfZ�DS8��FOQe�
���3�=D�4c5FQ�%)�S MY�0J"��F.�<�g�A4d��8��'�(�����՚BaƂ(^�0�<^�P1꓃fЂ��j);���$
�5��P��xH<�`�Z)H�b,!P��5h+ft�ǫ�^�'�d��M�%Z:�0����&4��s�j	�g�Z`
AI�y
� n� U��l"�sG �o®�#�i�$�*R��w�� �O?7��\Ż���./���X�a��c!�_�F��K @�+Kn +����`����He*C��H�
��dH?v�jB1n.Ԁ��F!SCa}"�ӌG��$�@'�w�"Ѱ#��7V
n-����'%l�k�'Ǩ��3.O9��TQ5���
Lmx�����)���#�i��$�D�Bg���:�L�z����=��ȓtt��3��̒� �Q�D̈́	���b(� qhB\�S�O+�i����C�����%�t�Q��'~X���S��|��3�=D����^N�V�
)\dʧ���!�dT�A���)%�A+S H�J_orv!�ȓ6h4��Y9��-P���$u�^� �"OHE*�˗#�t��!���\��"O������k���R�"G	�RxZp"OXYA�l߰w4͋���O_��"Ouؗ+� :��}rc惜E�D��"Ox��t E8TtTH�L�����E"O�񅅇rL��r'E=1p�*�"O��a�_\�d�.і<L��ؒ"O�x��}^��!ɟ�^�0h�M;D���ժ�3���%؍`���A��9D�7�� L�4
3��h�
s�6D���E�ŵr[���;%��ۂ�2D��;�ý"K�}
Cj� 28��:D���kd��������:�a7�$D��2�A�vFQI��X�d�x��#D��x1c�NUD��S��;z |��F�>D�P�>��I�� �@J~�R!�.D���� V�T�U��S�,�|�T	(D��Q3�E�Gb�q%NQ�T�d��-(D���u�Ƅ3�4!g�R.5s�L96g*D��!��!8�Ѡ�(.� Cb�7D�\2�ĵ1��� �B��۾6�P�<�Gj�	��YRr�I�%l*�B䉟`a������
"���vb�R�HB�I�G�
ͪ������m�n�B��:n{�,��ƪH����YB�	O�0�Rs�əj��Qf�)�"B�.@�V��s̒?./�uQ���^pHB�	}�~���:����B��1j�C��aHj�YC�G�SW�p�kK�eݬC�I ���C�lZ���	���,B�	?Tr�j������X��w����+A�0mP�l�r�n���޼Sl#>9������P��{�xu(�H�y�<	�K#-�P�#N+�<����m�<Pχ?y,p !j\�X�D�s���r�<1�h�z����`#�#q�%Q�OZp�<�v#]%d7���#�P$`�d�C�<AS�ߺO��}ذO �e� l�$&�|�<�
y<� �w�>���3�I�A�<A�(�|�t�ţ^	.�P�k��u�<!vÙ:�r�z��Ti�0���Kt�<�u�M�č��o�
Ȗ4;�K�<�T�P�S�\]�ak�7G�H�B� �H≪o��1�)�S�u����O�']s��7��2|���-~�<��|J>�$�P�k.���/�i�bB�K�
ᠡ����0|��a�
B��]P��	rڐhAgŜH��(����)���
���?�'����Ъ�if�,�dE^7�i���(?Q��<o�9�
ç=[��.ئ��b.Z�@��t�q�~y��9h  �+­�Y���7���S'��4}����ׄZ��};��'.H��^[}�{��÷^>y'>qj���3L��8�bўadz5-['&��9�dm�	�~�K�(i�a�n
�2��@�-^@�"���C��6ऄ#�J���A�'�����<m�ℛ�
)��qUiV�Ӏ���'��Q@��+J� 9��π ����8i� x�k�.{8�:��'J
���-��O�D�Z��i?E����#<@ZP�C' �l�5�I�9%!��[>,޸=� �R�F��0��]	!�B�*2<�YW��Sxθ��ʔ�!�$O�r��5х�S�,�I3��V�!�d�(!n1��ǡz8��E��9z�!�D�}3����&"�m���w|!���c����bb�3p]�e�33!��^�N��a1��<P��]�b!�d�/͸���M� TT�ږn�&�!��eU�퓁`�,����-��J�!�>��(��=39츀�eM�/�!��дo��mar/B�8B�ӧAd!�dU/N�QRc�0;q��b��*!��>Ö*�	Qmh���옊I�!�D��LzĔ��V�@mHm�U.��!�di���H�1�d�E��5i8n ��'(n�C+ �R���%^��1�'��Ųr Z	q����^�(�ȓL��I�,ݪf�����M�$�����h�,A����iX�/d6ȅ�!j�ј�`�7E�QS!�	˔D��U�4Q����p�d��F@vn*�ȓ@-2���#�pS�K՘A���h��a�"��7+0r C�J������ȓcv��sĆ���4�ڑ?��x�ȓVU�AJ�l��,�*�ւL_����ȓtƴ8ȇD�15R���hD�?H��m���yb��NS��ct����|��cd�T`���%<M䵣�Ñ:3�nL��=@R�����n>�K +_�O3\t�ȓ<`q ԥ@�
��"�I2&�ȓ.W�i3䪏�7O��� ��3�"��� ��`�A�v��$�d�R���ȓ�
����_�c��	ע�:�J��w�r�5�
H��)���4"����ȓ��� d*�k��I���3b9�m��^)�9ڣ#�7d��j�$31��H�ȓ ���kgƓ�$����H1;���G����/��9������%�X��k�L	�+�r�����y�ꀄ�_���)t��2G�4p�E���J*(�����%��J�?��P���`�FM���<5�%O�G��V�ҫ5�ṫȓRxy"��Y��]`A�פa��L��N:�r��K�k�
Th���F��<�ȓ��#�*��*�6�� �ߡ
����T[0m����x�FIʡ��fP&��ȓ_�Y��O�z P0�j@��Ćȓe�Ԑz����x0����1%�ن�D|��xiȂ����l�>8E���B���Ђʋ=EMPa���T9vZ����;(�і�ɳM hh�5�s���ȓeX�8Rq�ՆU��(��͜av���ȓ8M�Z�AR��5��a߾[e ��& ����U������-���|����w%$,��P8��̲S5r���<v41�   &niq 뙬']jd��b�n)B��Gp������e$�-��Z�<LJR�_S�~��3��(r���ȓA`,H��Ɵ�lRV�� 5��܅�v�����G˰p(���AÜ9��P��I��SOK�i*^@�@ۏ.�1��`h��t� ~O�YZ���
N����S�? r��ᏤLC
5x�-�	� Ze"O �b�	�=ΠI���5~ P�"Oj��NR��X�s%�`�V�	"O ���W9��5t#�*y�J	p�"O*M���X���U�G0 ��"O��8����kj�pv'��Z��� �"Ol��ㄑ1U 	��� CXLP�"O����m��Q�c/�0S"O ����O�� ��̽���PW"O|��%EB�Mش ��?�hX"O��3rg��?~�Q��%�f-c�"O���6n�ȕ:�6^��l1�"O���5�,@�t�b�\�$Pp�"O@��n� ��U��.̊x�T�c"O4�1�JQ�QqƤk�` *B�x�"O hx���Sɼ5t!t,�� �"On����G ��ѤHTg"O�<)���yY@0H���'/Xi* "O�qc��˙$m����i�{��A�d"Oa'�Ѽz^�� ibaF�BF!��¢N�%�b��	��=J�a�r�!�D�Ow2��@l��Uj��#�*�3�!򤖔Y���r"`�T��Y��8���Dć:��P"��ݛX�J�����y��_��!u���jda���y�jװ-��$1� 4m�bV��yr�\�
6��pB�L�&Ф��e���y��Y>�|�T��s��d��C�y�A_#M}z-`#C��G:�2�F�y�2!�z8i����(�q���y�%V�,뀨�5L-*�$���y�ݩt����4a2pq2��5�y�G d���XaE�q����Ɇ!�y�+R꜈P�	�>xب0d���y+U1R6  ��8θ#����y��N{�|���@�>a�%m�y�S�7��D����%:�]�ՊZ��y�h�a�BҖa��Z���!�lG��y��%8ez��#a�2PU�5:��]��y��2X8@P�!7���(��yre=BF�L����2)��g*�)�y��&Oԕi��"%���Ñ�Z��yb�Ķ$��j��YR�� ��	�y�h�15J�K����"��HO�y��JO�T�	���
��=qBI��y��h�D8�0�U+@���h��yR��7
BB|�4��81�ab��	�y�h_�W�� ����"=tb4)���y��1	���ua�29Y6�!���9�y�D#��׬��-���8�@E�y��Ii�P�SÈ�T����j���y2%�"~U��*,D��̙f�V�y�oؠW�����d��)V�jlC��y2��zꚰa�#�&�����Ά��yBꕚ(5hd���T ����yB�Y�l�,(��ȦY���͡�y���mn
��
"L ��jT��y2#!t�8�  I��~{"��E��7�y��K���q� zS�@�M��y�.�jG6�[d;?C��c�T4�yR/�s�惌5��@���y�G[�eQ�Ɇ&A�z�d��VB���y�K�.L�*rf�vTD�R����y�
�'� �.�
%-��X��[��y
� B,H��sX�#A[�Tި��"O�8����T��qy%e�<p�I#�"O�� D��/��A(2��;b�>�J�"O.��������zмa�"O�9"& */Z�Cf��/�6,�"O�1�T,h����M��5�@�#W"O� (�%<��3lB�$���%"O��z�k�}[���!K��*�I�"O��Ӧη��� ���?ia�8��"O)�R�{!�8�C�Eg<� 1"O�ċ�h�tTx�ț��$a �"O�-����;w��Ò��=��@ig"Oh�x���@(օ��.�zE��"OL,)��SQ�ٱA 	j�\�1"Ot�"Ê?wPt�@�}im��"O4�*D�;n/B͊�-OdOdhrr"O����2�����0�2�k�"O�蒋�9��0cBp�� X�"O�<�H�9r����bk�-Z�m�0"O�I�T�0´�x	5&�y�"OD�3R��Nf��2낤j#R`�"O�)���***>��
�x��@"O�s�jC�J�T��03ܨH�"OP�)H&LD�i�$%LH����"Ob�qb"X�1�X������"O\Lq ���CQbH*d�l�[�"O�<hg	�	Ra��&��v��P"Or8��ڶ<���[c�S��))�"O>T��.��Z�(�����~{b���"O�!wLق�8:CDί7�,S""OR��.�>gJx�K�)�l�����"O��a�D��Q��ˢkݓ	�lMJf"O�A"k@��䩡�ADT*c�2D�(z7��E}�C���sP9!�1D��a��4�ese.��^���R�-D���w��\Ƀ�T8>�U���*D�8aQN�A���E�E:�� PU	)D�؊��Ǵ2ƦY�%B���)���(D�#�@�M.����"(�<ɱ`%D�t	�nú]�V ���[j0�cj$D��)t�(��5�7!۱�e���!D�j��G5�"��i���Z�?D�x3FcX=iC尷�9|��B�;D�$mJ�rݰ0JA@-�� ��M6D�js�G�@*e���D�H6D���iP�9B(U�@�[�~�b�C�E6D�xQ�ÂF/~�2%lعD�T��2D�p8ㄖ�-��}��/W�����/5D�<R늾{���J���$ d�P8փ3D�,��X#&�JE�IJ��,LC�+2D��x��U�/>�S":8����0D����M3B�����e��!D��Q�΋Dc\E���a��:D��b3i?�VM!��ݰ~� �ѕ�8D��Z��ɳn�D���\�E�1`$D�����L���� Z$!�a��D$D���Q�D18a�U�B�S�}�V���$D��ѓ�Թ�Jh�2"]}�,� ��,D�pBD`�i�zx�W�UuW!86�*D�(8��1d&� jva��Dn��:��-D�d�sk�=wZ� R2��&�X�J6�5D������#�XB��6v�H���	5D�4{�!��W�<�nת8�&���k3D����m
dARc�W��4�""�/D�� �,���R�  �I
�3��"O����h@��q�� I6"O�y���K�X�$EB�¬5�n4"�"O��ꒁ�<��U�5���d���"O�{��Fj�0b���*z�e�"OX-���R�A5:-���۝VR�%(�"O��Kǣ8���u�B��S"O!�e��GU3JC
�us"O�;�(�_�t��(�
RD1D"O޹�4    ��     �    	  �*  �5  PA  }I  T  �]  6d  |j  �p  w  \}  ��  �  /�  s�  ��  �  ^�  ��  �  4�  t�  �  ��  #�  -�  [�  ��  ��  ��  � %
 g � �  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�	l}BK�Ej����&��-�uAA����y2`�8�x�ؕ� �q�E��yR��6$,���*��@
��*�yr�NF^�Xx�L�	�:��B��䓘M;���i�Es��ؖ��&��Kg� �!���H`J���`B�<�dG�8l�O���\�Y��a %с"�����KM�!�;]�lڃO�6r7��
��ʯ��@��;�XC�iP�xٴ���A�ޔ�ȓ%K�M�u��	rG��S0KK9��an�!�x��7>���YC啾(���%���=�{b�S��:)�j 	�%���y���"�����(�'�t%��lA�y2a� FB���4'ϟ���kЈ[�y�_3R �S�G'�.��$� ?�yRh�j�
�Ƀ,��v#Z��S����=q�y�$�&P���Zni��"��y���3?��*�D֩l�¸��HՋ��Op��#��b�mDnϖp���+$`DW�<�$iB5MAiB�biܸ�u�O?I����9O��M��W�?w�sH�&}/JB�I= ܒ� �LD*s��+Ǉ�Zq�C�ɵ]�䝻�.�=P�]�c�:+�B�)� �ݫ2�ʰ.7tH�Ӌ�v���"O`qB2�ܲr²0��ō_\���N�Q?y��Z�]JꬩH�մ�3&�=D�<H�D߱Z�����Ҋq��`����XE{���^.J�t�ѱKϫ1_�A�RgrI��'��i��6H����Y/C佫�'K��(�J�]��90a���U��'/��qa��
	>%���� ���;�'8��c�Q��
$d�쳏��R�O�D��E�+����ҫG�0����'"�`���(F�����W��\;�'�faZd!�1� p	aP20��'Q��S��'{���J0m�z�Z��'�(\p#�; f��zV���#1 �':\`y��I`�I��Y!%� ��'C�5����'�*�c��	��'�P%�S����r���F;mz1��'�8�Ҵ�P�5�d��g+�/�DL����v�K�DD=P9�@��N��,��-�q���u���x�͝�D\n��?Iٴ�O�6x6Ah��T<�Ы���s$P�ȓ:�" �W�	K�M�V�wN�܃�Ot�9u�g����(���]%z�Z��e��
��$���-���vζǦW;M��oZ�E���&v��rc K!j,�$�#����O��|�O3zš2E�9�tK�*)/@�k�'�flg�,h�����&�t��'��}�p���_[d�Ae��3�R`��'����� ��UY�O
"�!@�}�'ٖq���
 wJF�%h�'�a��B��r��ظ'�%q��H�'{N�hg'&P@�c��W�Op��B��HO��i�OߖRԺ�����a*����"OV�H �}���ie���`$~	�|"�)��0�>%�'%	H!�C����C�	�T Up�GG0\��)w�H*�C�I�������,5Z���1��"m@����������G:�����CΜ<�e P-o�!�&?���Z�ƈ�.�5���f�Q��D����O���c����l������y���[��Z���!@���(�y�a�/� ���R9����yR��&(���� 4�241ē�y��� -!0"6�<^��Ayp����yZx9����U�F�5��/0@Q�	�'t��C��9��r�R�#el���'��P ��a[L�h�ឹ(O�`��'�
TB�Cu}T`	s�X0s���'x.i�t�!8��w���D�
�'�.Ԫ�˙�T.@���M)}�n9	�'Y4dq�kޅb$�P�T}h@	�'eA��c�
.��4��$�mbI"	�'
i����;�����aϳm�J8�'-ў"~"B������
�1k����U�<�`���0�����N1{aB}8��M�<iRd ,��	h��'i���@�"Bn�<	d�[�e�<1�ժ�";�� Q��G_�<��.8qh#��0D�Y"��^�<�4IR�N�z "Wn+:���!EZ�<�qh�3�	�6OU�AR�.�lyb�)�'9��y3b�%��+u�ӠpZ����%�*��O)/B�����l���ȓx&����hl \�����X��ȓPYt�Y�慟Q%��;𫌓"����S�? $Mf��[f�SÎ49j��V�'*ў����i�t	1�EZ�@���3D�D3P���}j蹻+]�CHŬ#?A�)�'4��<u�H�V������ӿs�*Ԇ�6�ص �A�*}�=�F��"#� y�'~d��gĶFu��!	q#Na��r��]�ә���'$�[V����Yj�C�ɓ*���8Bk�6,�9��,��wwd#<����?�ad	!����`МS�R�bTH6�O��Q޴x)�@����$1������J)w4pQ���)��<��m��9�^`h��J�>����|8�H��I�cZ
�S7`�%��(�`�H�x!�B��;H�f�۰KA$& �kP��'�ў�?�j$��1��`��J@F�N���8D�4�� �')g���s	_�)�,A;`-:��y���[B�׭W�_�([RK]	I���D%�	�)��}�2)9 ���_C���d��(O?a�s�P@|(ى�F��i�M�P�p�<�p�Qni:l�拶�~4�-Dj�D4�O�8���,i�Z9� >.����f�Dj%�\�@�H5�P��h#j��>D��m^@,6�1gB/p���î=D��a��� �`�$Y�7�����<D�T�����LZPc�#X�r��kk9D�D�6��+B�@.;4��q�7D�X+�p�}1�(ң@��L��1D����˜>"<ĥ���O�&j�
/D��`�G"].� �o��/���1��9D�|�A�IL�%	�+�]�*A�!D�P�%� G ��j�����9f/>D�����̢U3��1����C%��;D�8�Ŧ̏(��I����=��d@$D�\CR-J�a�f��H6а8BL,D��Y@≥3d
�{Sd<=ֵ�/)D��I�L�Ҏm"��.V�R(D�J�	��/^�Q>����&<D���hV�J��M1F�\.���1�%D���O��RKX�zd� 0S� j�'.D�������FI���7ⓣ;��hh@�*D���/�P�TФ�R�]Pp��#�-D�H��a �%���D�g��K4)'D��y%�[R� ��@5L�"!���%D�T��� &Fʹ[���!?�a�9D��%�J*����D>9��k%$D������'LJ$h�KYTUXge"D����e^:bPnM���~$! c%D��	��͹KL�Ӧ���8X�$D�bkVQ�3�F�tY�)ď>D�ܐ����
���LO�d�ޝ!�.<D�p��Q<i왘�Iȷ!-���V�4D��K�hؘ*����#[�Փ�C>D�P8��̸_��e�UlW8�vͫS�/D� c�ύ%d �-T�}��)c7�'D�Ā𮅖uX�ɱ�'Ѐ:m2���$D�����I�4�d�g��}Vl$��6D��QFZ�hQ��Y4m�/�p���3D��aC��>'@��lD�J�Bu��)2D���d�BI��%FeW��0�K/D�����Y��FO:O�Ј��-D��z�9zΥ2 �H�$���M D�$0��_�H�P�h���9�`����>D���Ո
�N.�=���� } 2��7D��ת�� ٔA�Ѯ���T���1D�$��?�lU�<8�6@�I0D�� ȼ��f�?��h9d�=攣F"O&Q�'�
 :ƽ3GN:A���X#"O��@�A�UA��4�� �*� �"OzG��p���,P1Jތ�Y�"O�pa6�$͑ HO�K�x	���'�r�'�b�'m��'���'�b�'�Z1q�'�j���Z��92�4�!��'l��'Kr�'#�'��'���'�"��!�I!�N�y�"U�7�'{�'���'���'�b�'�B�';*ɂ�[3�n �Y�����������x�I����I۟p�I��8�I�$���A�2r�p0%3WքjSGY���Iǟl������P����`�I�@��
�|8:D�'
�bwv�8%�蟼��ϟ���ݟ<��꟔�I�`���P�!$B�H��h:7.S�B�vD�!l�ş������	՟@�I�$����l�Iǟ�J��]�&�����-ѹu��	Rè�ǟ���������d��ϟ��I�� �	şЀHQ�p&6��iG����Q������Iҟ(�	؟��ڟ��������idL=u�� pt,@''Bl�U%Hş��IşX��ןH����x��ƟD��ǟ��A��&sQ��pdhT4��P������������Iğ\�I蟖�����ǟh���Ajp��B䌫1 �|����
�p�������	៸�����	�$�Iȟ��I<i��lzq@@�%�L,�B�D7:��h�	��0�	�`�I�����ß��ڴ�?���LU�&<qd)�"͹�r�I�X�L��Jy���O��o!n�(�w@B~��� �(�,�`Q���*?�W�i��O�9O���Y#;]^8*���~��A��X	��D�OXb�O�r���4�����OR�p"�C�BUT\㟘z{�(��y�'z�	N�O�T��J'd,�11�P�r�,у��}�	C��;�S��M�;e��A[��L�
g>��'��� FP���?�'0�)�/f�±l��<G,�-�����B�8� �KQ)��<��'�.�$;�hO�i�O8"mC�*P�s��:)�b��:O4ʓ��/כf�Z��'�|,g!�|���b�_�H	���C`}b�'��3O�G���$�T�=p�l0�(N�@����'w@%E�luɋ�Ĭ �p��'����y�PS#�D�/���C[�@�'���9O�\��ɪ�
U!`��1a\�@�5O�oZ�cQ�\���4������\Y�u1�)mz����3O�d�Oj��^CN7*?əO���)F2L� ��3�lH���P��-�H>�,O1�1O����	���@��G*�(`�����Qٴ,��Y(O��D$��#��Z񡆸P�8���J�V�	ٮO����O��O1�����$Q�Y�X����� �6���l��M�t�U��<�ԣ�1�8�dV��䓳�˿ �thU�H6`�-�ًS���D�O>���O&�4�<˓pM�v��V\��r/�Բ�h6A�,��bG@?A7�i��OH��'��^�2��|�ވk��BJ�b(b
��j���l�}~���%T�H4�ӱ7��O�G��t���L�=v.dJv�ĥ�y��'���'4B�'���ɛ����X���;d�JQC4+*g�����OP��䦅IV�~>5�	�MO>-y���+$�Bm��)S䕃HaP%�(����S�SL�$m�Q~�9s]dj4�S�&)� ����!���<+�
��K����4�t�$�O��\ ��UQ$ E�;���=)٪���O�Z��F`�T���'���O��$��B��Zĩ˪sR�=H���1�y��'����?���O�"A�$<I���8_b�26Dʀ"�H���2IH�+tQ����-{A��W�	���{Ǉ['D*���(8����$����)�tyªh���HUcO�QD\8[�F̸�~i15!S&4����OFoo��7��I֟{�C(Z9�pE�ߢx��ٺ�M������ ��n�Z~Zwc��`5�O����'�4�`��x��7�տ����'���t�IɟT�	�d�In����H�����z���1�K��Z�6�R�O\�d�Oh�#�9O��oz�Uб+�'��a�A��T�G@���I_�)�=c=2�l��<A腩|f)9t%+M�(�6d�<)�g�KV��Ċ�����4�`�D�f�B��%CX!����I]� ��$�O����O�˓,�aQ5~*�'\�	(�e��dڼI�$I��¡	��O
��'/��'K�'W@�X�
�?28����a�:�@�Od�D���|uH�#���?��O�tH"�E)D6I��(ڃU��z%C�O���O��d�Oܢ}Z��-8Ŋ����Ȍ
�o�3c��u��|��$�<Q%B�'�6�>�i�!�3��["~k�$��:���it�P��П��	K}��oZa~Zw���yc�O�8�#w�N�RP<e��O��n9�@�i�I[yR�'��'1��'�R�k�0d�]�PʖK5@i�)8.O��nZ5�����$�Il��`��i�;�ԥ�%�d�54i���$�O��� ��)@aՖ\p�'�U�-Z5*B���
�c���9(�2"K�� &��'c�ciƾw��`^[�>TC�b��fA��tg��J"`<�p��9x��p;U!�yJe�
㟴y�O����O>��]�(*����u�PH؛9W�y���`o�\��!���J~B�{�? &L����+�^	9Oˆ}*M�t>O
��$�7|��ɢ㔺۰U�3�Ǝ���d�OV����K6�5Z�i��'Q*�QF�m��j�%�'��0�4�|��'G�Oq�xF�iT�	�J�@����,L��� ��y�V�AN|��D=�D�<Y�b��`�>Y{r�P%F�����V��O��o�-y�������l��c�� Dz}#E��'^�yZD�]���r}B�'Pb�|ʟR� ��#�t�*O*�R	�6�)��D
��z�`Ĕ��tRQ?�K>	5�tm(�e��&�Fe��NQ*���ϟ��	֟��)��^yR�|ӄ9��ʋ_px�9'�T�+�Bl 5J�b�����O��l�I��T�����f'�hk]�(Y~,���˟4�	���m�c~��
E�6�����h���g`���:V@�(��d�<a���?���?����?�-��A"�Ѝ{��3@�כ
���9G�ͦy�u�П��I��,�OD��'	�6=��d�^�S����&��P���3��Oh����4�Iz%n��<��`�	�jy����L<4�j�+F�<�`l�ZC����+�����OL�� �1 Pi՛~,�Mj�)C4|����O��d�O�ʓxJ�V��������8��ʝT��Ա7��*�,I"dNO�Fl��şT�	Y� L��t���D�J�zs��&e�J�0��� G�%{�P��|�WH�OD�:��,=:�����X,8� �^�
X�ȓF8D��"J�u���s�+���,n���ƴ~p�I��Mӊ�w/ֽ"�	�*2���$�&rÝ'["�'I��cM�nZW~Zw�p��e�O��}p�Y ��T%�N���H0��U�I}yr�'��'�"�'2�g�q�Ub	�dʼ,"q�� D��I��MӢ�X��?���?I~�t�� �h݆{���b�R�-��m"!Z������|%�b>J#D�/?v�(o��CI�Hr@_8+�6��RC$?���yW4�䇈������,��FRZ�8����60�����O���On�4���:����M���K>sʫ�J*��Q�E�R�
����M{�bl�>���?��SY�`
��$a��ó�A6msJh���&�Ms�O��)�I�����$�w��z6��7|d��7��(f�QӞ'b��'���'��'B�O�Rc�1��1�O�y�>|2&��12�'��,k�ĩ��2�`���ߦ%'�4"PmG%yV�p�E�
XpZ��"��(�	�쐔�
ަMϓ�?aD`���Hj�D���=`��'~& �1��O��J>�)O��d�Of���O�s��ϧR�*&���Kh�İ'��Op�ĩ<�q�i�dC��'L��'r�S�(b�!���C0u�$�J��b�������B�)��?U4z �@AZ�S�5{$���L��#P)�qX*O��?��A ���	��t.Y)֬+���OJ�D�O�4��!�M�O�˓-a�V�Z� �%P�h��|H�K���!�ĠAR�tݴ���?�CZ���	<	b�`H���2N8챪�D�N+�x��˟��s�����?ɐ���`�z�����$P�|�ظ��`٢F�b��%`�4y���<����?Q���?��?�(��Y�/�A�4��wL�[�"�ahĦ��G�R柠��柘��r��y��#�p8Q��ZE�[��!@R�'&ɧ�O �@Y��i�� ]?֍�a/�h�D3��E���D݈�f���'/�'��i>q�I�w`�-`��X�.�dA�AT�vu�Iԟ$����L�'�6-> ��?�c�-$�𳥫P�#{�qr��ŧ��'����?�����so^p#�e�&]��	�N6|Py�',����@O�A���:�������D�)�T��1$͛�N���p��I��U���JeM������
g�h0�Ϟ�Z¬0A�B�'d���O{��=:*�Ftq�\3� ��ߓ
�y�ɒ�9��Z���tY�H��腱rbV8{�&���f_���!0X=>5w��`qε	4�X�p�g].O��}�u�ynhÐ�	�?�����i�/+���0c�;5�Y̈��L�m->ȃ�̏�PX02� ,�di5��3,aZ�eۻJ�ī��!�M��H��h;�S��'B�|Zc}�X�mJT���ʳC��­O&�JF" ���OL���O��FhN�j���;��}�/C1ͺ�Z�)Ю��	Vy��'�'c��'�
�6*C,5�<xЧD�<S�Y�7��=Y��X�l�	Ο���cy2f,x���ӡ#�l ��/��D��%{�7ͷ<������?���M��pk�'NY�D��|6�n9���[�O����O��d�<Ѧɇ6�����\�� �7D��
��ڕ����G��M�����?��M����{�,�a�聁T�[�  ��H#�M+���?�-OhSA_p��'A��O2���%�Bٲ����(�\:��%���O�D��$����'6��B'K	�p�����r�oZyy�TJ7��O���O���i}Zc,�DX�LK(Z�>ME'�(J��b�4�?��Q-�"���L7�X!���(�)TKۛf�M�+{\6M�Ob���O��iVK}B[�|a�)B
 j��pB�"o��)1���0�M��Kِ��'*���  0"��#uA�0a}�U;�_/��l���������s���!��d�<���~��'8�����K'� ��È��'K0��y��'��'�D<��eD	U2AJ��196�I�+dӺ�ă>[���'����H%��8� �1���"`�|���^�O���ӅP�L:5��Ɵ(�'�2�',�\�l�4���:���_~,P�"E�Hu�]:�O2��?�M>	���?1�
̾L�<�����^�zȢ�N�@qvH�L>!��?�����""��ͧ&�X�E�w4��)�FH�7.hmZJy��'a�	ʟ��Iן�2I�E2��T����l+؞!K�	�R}��'!b�'1�Id��K|"����o��|�a�Y�1"�@�+��g���'1�S� ��g��'#�S�P�p�
�0Ym<�
R��	��,�۴�?�����$�L�Xu'>��I�?�X3&���-��Q��=1E��2�~6�<����?���?�O~���ED��7"�B��[�`>B���ʕ�m�'����ou�	�O��OP�b�hLK�F3�*�1�ަd БmZ͟���şl�I1���<�/��v�҇�����    6�������M�4B��?���?�����.O������S��5O9�h�4O˽S�K�OP�1�)�'q||EX��qȰ�V�ƈ��i���' B&R�Q�)*I���T!�VژL2�NK�p/Y/$�u[���F짉?i�'�$�C�AB$'���BH@�݂�4�?������\����2����/ר�𴂡�F�1W�M%���.�I�<�'��K�l��TB�� {�Za�w�]I�-��\�|��� �?1���~2��zV����A2,Y�CF��M[� �`~r�'E"�'��	�b�C�O��}��GWU��LrgX;H�J�O��D�On���<�����)�Oh]����\8��#�8o���B��J}��'/BR����0}�x@�Oo���3+F]Aw�?���W�{!b7M-�	ȟ��'2"�H<�'Y�g����E)Mir$p*��u������'�����0�I�Op���芗Ǉ�hT����\<E��i�&�i��͟,�	��t��@��X��X(��%P�oGm̪%�FΗ�7�<�eK�7	��fm�~�����盟L�ղ�G�49�<g��@�`�X��?q��'�O��M�P��d��Aze��O�m��e�JQx��ߝ�Ms��?i��zY�x�'�F[E(@�,��!�U���� µ��p��2O��d�<9��$�'�XYFBW%,�e��D�D�4���~����O���]����'��I���?S�Q2̈́c���g���1�o�����'��������O����O�Q�c�;В0�ABB�fԆ�XA��i�I�c<J�3�O~��?�/O|�����Se��llX�Ç�� I�82�Z�0�f�~��'���'�"T��-�-cm�}�ָӥ+�3�PQ2k܌����<�����O����OdX`�n�m�d!��M�*(�PIش�ΑP���O��$�OJ�D�Oj�0>�i�D4�������i�8��+4�L���i��Iǟ�'�r�'�e��y���s�^Ր ,{3RI�u,ԇP�l6�Or�d�O���<AV�ܽm����֘l/FY;���
�3�n�-lR6��OR˓�?i���?��PX�eAz����@�����~�lZ��H��Vy℀' U�맩?���jE@�5y<H��t�h��3'���	���ݟ`CAr�8��zy�П4�!�$	�\6-�@�2���y5�i��9d��+�4�?i��?q����i��H��`��o�eD�,�Ks� �D�OtL2�8O�X?�	�'js4aw��!Tf�'&�<ej|oZ?#�lq"ܴ�?���?��'2��I^y£�4Aa�v�������&��E�L7m� ��d�Of���O��B���UJ����8 u��+$�87��O��D�O�ӗ��g}�^����M?i ���P�!(�m��T��`U���	uyR%�l?�O��'�RKB#D��E��"�0@�����a��7��O��r}_����jy��5���eG�]�l$]p�ə������+^��<)���?!���޹%���`�[�P��T�� ��Z}�P�,��yy��'>��'����Xd%�9)�ȃ�j����������'��'9BR�`y������GF;Fg��۱�D�p dE�4�M3/O�D�<9��?)�4$�eΓr��Ԉ�N��\����qئ=xֺip��'R�'��I>8Z�!K���������dĭw&�}+�b��z�q�iq�_��	̟��	�:�8�I@��4a�U@-�>S�b�
էd��l����}y���0,��?I����WAƸr�%[q�өZ x��Ӕ*��ʟ��I͟��E����Oc�ӟ�!� O�z�иD�̯h����ѱi��<0|E�4�?i��?q��t��i�ib�ƅt �e#���>QZ4lg��$�O�9$1O��Oj�>����T66�����D�MC6�[v�ⲑ`����M���?1���u]��'�NѪcCE��Y�&!àSD��v�e���B=O,�D�<�����'g�)+�뜻d$&��^L�Q n����O�����K���'$�	���[�N�4':����H�^PrYm�h�z���)����?y�S)|� ON\!l�@^s�h��W�i���9���$�OTʓ�?��M~�"��G)&���)j���'�8�ə']�������p�'1@=qu���A(�@v 2D#�PѶf��W�
���D�OX˓�?���?"�V+aXn���==纽�c߯e����?����?���?�,O:���+��|jg.5"�40�q�5�� A
ҦI�'n2]�L��Ɵ���+?��S�? ��z��W��b�:�HQ/��!�S���IßP�Iiy��X����?q���KELMcCKL�� b�!;�f�'?�I������|xW-(?	�'�4�`���O�IrV�Y� A��I�4�?i�����Q�|��=��-6�OL���2��}q��JBЪ�B�FVX��'��'��yRQ>��Kr��1N���G���#����"�զE�'-I��f���$�O����p�ԧug�Sl���%F�<`Y0�`�Ȯ�M����?I&@��<���?q���O2�����bw��Jf��$��!�4[[��g�i���'w��O������ ��Q��nFPdV�`�Umڟ?L��I����'���d3���æUN,VbA�:HmZӟP��ş��c7���<Q���~�&��)�)�g�پ�*<�����M�����A�|U�?	�Iҟ�ɦ)j�X ��E�[dm�2CR"��ٴ�?i�)F�_��yy��'0���֘3-�,u�4�N�aZ�)2Ec�N7�O<�W;OT���O��d�O*�d�<���T?|%6���\�w�� P�a�3k0��`R���'�2Q���������mK��
��OK,|�s�
`u�{�h����<��ܟH��Fy"!͑X�B擵W`���Q�$��X���ܙk���?������?�����2ѺaZ�N��0�YH��I�$�(@XpW����՟��By�cV������K�O�.� �^X8*d�b+Ц��A�	П�I>YNF�	D��C�y%�8�hG�	�������5�F�'<"Q�ؘc���ħ�?q��q%�9����=S�4��JC�䣄�x��'����6a"�|Rٟ|��d	��t��dA_�("X��i��	�5�`�[ٴ%��S����S���1c�����4�,2�-P9���'uߝP��|��	ր8���Di\�,
n,x���02�Ƣ.8I.7M�O����O(�)e�	؟�AdGR:�D�愒'vдM�sO���MS��<�L>A��t�'�LT[F� �"�P-�qO�R�D$��Nm����O���[*��>���~�"G�Ou��j`��9��maB�Ǐ�M�N>iw�K�OF��'s�I��_&����γ	4������+t-���')�p��&�	ҟ�'���P�:�I�	�Z
n�)�ğ<E�4�-�P�Γ��$�O����O��^���'%�X ����?F�$��3��1<�'���'?�'���'b���T�J�x@(�X�-Z'S��P��E\�p�2T���ß���Py��X����e�� @r�߽A��K�配5���?y��䓩?q�i�����WJ����S
o�H��0��<�H� P�`�	ԟ��	DybJ<���2���a>>�Ry �g$>�Ԍ��N
��)�	n��ԟ,���^#*���[�����fF�)w�$ن�͘i����'��_���6�����'�?��'�0��4@��k�~�'�˧?�b-�b�xB�'~2#ҧ�y2�|՟B�;�!������r&�,w�p���i�	�e"ԣ�4q
��ǟ��S����7��Ё�V'r\,ġs%W

���';
�y2�|R�i�<y���dO�?L?.i�P-5����;H�7��O8���O<�	�}��ڟ�ɓ�X��F��"�\������?�M3ք��<1M>A*�H˓�?�SbM9t���92*�p �2@ɕ�X�F�'F"�'.H�۔%>�4���'
B3�*�������Z���Aߴ��'Y���D�O6�D��XI�!��ͤll<�;�D�X��9o��q��=���|"����6��irC(
�|`{�a�1rf�''�R���Iޟ���ʟ��I�GB��8�M1Q�D�T�� ����˟��IUy��'?�'"��O���	�-�!VIF��lh�T�i���:�OZ���O��D�<ISA׶9��IS�B�������^�&Y����)j���'���'W����O���: E٥ F�Ȭ*q�	�m��꓁?���?����?Q&KA����O$ �5]7V��<A��OP*D�x��Ȧ%�I_�	� �'�t}�N<���K�"8B�� "*�v 
��`P�.M���h��D��6aj�Y�Ka'pɳ���,n�!�^*h��q!��z��g9b浪���6Z�� Pm�1�f�\�d����Dٛj,Z����,v:��'+�������'400��M!XI��+R���8��=D"�%�,�`)��l�Pp��F+La�!kӌʯ$Ԕ��0.�<$L�
��wHt<�a*�5�0�+��2.�(��G`g�R���Oz���Ov<�;h��3ˇ8�\�ܢT��c~�{�A����K�'�&q���\D�'��fZB��Ι%l��a�,��x�,��#PB988(��I��p��$
�uܧM��k�I��E�)L�5y5ƑV�LQ�����L#	��Oў�f�G&R}��zU��+� �QUC9D�La��%n��l�q���h\��P�;?!a�)2)O�U�ML(���X���9�z�4�?[��i�Fj�O����O�dLȺ���?1�O��)���H�]������@FW���È]SRt���]i��P�'����ӻQ����u���C�Z!���;��=cFoM�i�}H��'��=�3�ʾ5�� ��HW <�FQ�R��?���hO�⟄iǭ�� (�"�ϋ0k����6D�<B�n�&kΉ��&��{� ��e4�I3���<� % f����D���B���"r4|��hߟ����KN����p̧j�$<��P�L�����O� ��wλ�0)RW�=O�ଠg�'����W�P��|U�P������P#��\�c�JP��!5OzK�'BW���h%�����`�)H��0h�?�	h���p"��%si$�򕬈�!����=�(�ݴ���Ie�^�P`HQP�W������D�whj�o˟D�	|�ħ& BF&ڢ�끅ٝs��y�G�(i��'HY ��]�w~1O�3?a�O�#K���G��>h������y��N�)�>��sHV�T2��� :!)�堰-�s�$�tq��'G��'��e����+9��q��=2،6��O����$eb�v탩�U����	�ax�+�-Iɶ/X7|H`�PG9(���ǲi��'FRcΓU�t�B�'XR�'%�w��y�DЯ66���^�^����3n1��Ti�\E���|�Dӫ�][V�L�e����w`�%:%ړO5�T�-����"T� ҋ��	3��v�!RJ�����?���h���S�gy��',f���X�%L���Bf�&7���!O&a	�N�+�1P�@�1��A�7��ڍ�4����<��	=N"�e�`��9�f�C�G7�kEE�?���?���N#���Oh��h>�)�h^���)���
�
�h gT�)�u�1$׆rR@4ٳoWx�8��UAaI˓�F�aa��� ��YQ4`܋t���C��Mx�PY4��f	�Y��	A���,�p$
�W�����O����O���?��BK9�� I��?m�`Uq��U!�yR$�f�"Dq�oٿ�JLJхǍ̘':���hO�i��?�¹�Ql��p�r�� -�!��"!ц|R���33�JA�R��9E�!�d��J�2|�%�<�f�$;�!�dڅM*Dq�]��-;�aI�!��sX���wbZ��$��2n�'&!�$N�ZV�v�ۀ��a����0^	!�Ă��^0��9�f 2��͉%!�$A/nԾe��+хO�d����)#�!�dO(S+�y�G� !�|����#}!�dj*��aw�N��lD��FE�!��R@��2�B <����ׅ޿Td!򄎄"[��
bm��줰��9(I!��&`�N@�+��a��ݻtM��g!�Ĝ'����
1#��e���k^!�D��V��t�\�|�X,c��
s�!�Ğ�`5� ���F������S�!�ė�@x�<�f���婦�q�!��=9'�Q*6#�'T�*̑TM��(�!�D�A�E@`��R��̀bFøH�!�D��P��HDـ��,)�Ʉ:w!�$)5&��TGڎ�������<k!�W����w�4#��@�u/W�u�!���>߸�@�%���SQ��!�ޙ#咅 ��R?3tT�j2n�6Z�!��a6�Z1 *
\P��Ǘc�!򄝃~��Y:��9`%*�ff�!��dU�uq��Ө/DM�d�3D:!�D�<X5j�,[�L��<�&E��&!�ʤ[_p�ٷeM�<���uj ��{��'��9�B{"�W��5z�n88��C�		wly#6B�+{����t�ܫ^,b�� �b�7K��?��ӱf�<�&e�ySf����"�Of�����)-�0���	߯+
��ˇ���:�l��
q�<���O��h�
3����'�<�uj(�`���,�u���O��8������y�N_�|������n�����V|o�Dʓ��a��}B����x�s�G+N�z��L��MS��/^���j��G�����'�ށ�'��Q�a���bK~�h���=~�����'w����Mj�V��wnW�<���O�Q%���ϸ��X��ϙU��c؟��C�j�� ?֤i���c��)��'��1�(X>"`����aS�8�X ABh��M ���0DK���	2d���\��iOӆ`��Fy����B���B��h�RQ#�GH��O�	��u��}��	��mY����L��{�dϝ�ia�a��&�1��(n��{Dh�6�68��S�? ��	c��|M0�a�7c0${�K˼ ������$C�fr�R�2��K��|2S���v�r��4�Hb�WgF!�dK!
5*nE2v]�@rh��P�Q�Vi�'�p��@�RaV%a�-`��%1����ܙ����v+�:�ީpF�'�D���F�:�Ɖː��F.��8�+^ּ�ɳ�܂�?)d�
�g���e�K�|{�,�������Fy�eͣڢ��VB�	��ن
U��OP�7�ۺ��DSQ��� Y�7�t��ג%��a��#C0#4���ƕ7j�p,[F��Y�2!�= X�P�[�D�$A��#�1"bj�۳�%M���I C�N�=a����y�0�O!&�����6�>�0Bb�6kNT��4N	G�<i��A Qe:��G5 ��C�
�&�Q��)�$Q%��O�a�w�^5�y���7S6`�C����uo��=^��-/&����d�%ѡC�p��x3[� )D%�.]� �1$�ֻY��yg9ғd��4�r`B,z�
�$B�bF~b(���ؑj� &��@$�M���üL�h�f���5�@�-Җ^�<����Vq*�I#`@|�iyr᝛ٜ �'���F۳Ko�E��X�x��,O�O�%�r��)_�^�H�IYa3�M�'�
���ĩfڼ s �l��᳧ h�H�h�ū<A�?���C	xea+O��Y6�_4��1Y*F�"U�'$
#�d�&DPv�|PD��o��Sb�&S�P��}RL��/p�Qf�F�'�������6U2���$�:qB����>/N���)�f�`Ջ�H�(}���Q�J�HX�u�W�,��=%<d���'�(���=_��\��hڈZ�:��)O|<�v��)�j��Df�
�"mC�O1��ыg@1~3��4.)I�
��8O���-�"�h���"0����=��Ҷ �F�ݧO�$&?!�5�x�-�<6tSQD[g�l}6���y���
t�
�8a,�4*圼ZU�Q��M[��N!S��D�B���+*4h�}J~ӈ�^Q�ːe��T8R�IW��`؞l0�W�wi*p �'dH�pBEar�q�*��!G��aܓ%qʑE��O`���
݊ �"ٴ��6_4�`S����tXT-����h��8r&*#99U(Z�z�y4b�a��q��V�����Y.{��֎Jq)b�`Aa *
�d�N��"͟��CB`K��I�_���W/%�hĨ�DYC�ɟ%�>*�� `��Z�IV�����S�r\`a
n
�%d�Y���Υ;|4�� ��ho:p�g _�/�a|҉Cx�|���E�Sf^;�T���C JU��ad�.�	�j��#|�'D"M�7�C�NL �93�ɴy�04J� �wnƳ)s``j �X�i}&u�ׁ@�,O�ԹĪ�%��ȪV;U��Q �[�,:Yf���*U���"���!e�� �`�P%�
)N�T)����:6�r��O���PD%�)zC�<��X�փW��@��A��xK�=V�p��v��93��I&(�OE���֮��'b����'�f9�D@�w�	s�Ol
Q����fuȜZÓP'Y*m�-vS�yD��v(�FMuָ�E
���`I%�\˟p�Uo�����%���̴BE�?�&��Q+#��k����)2v�9��hH��'e�t�Z�F�3wP�=ha�I�?�4�D֮qgt�A�,�	�bU�p�l(��(�Ơ@�ҿP�V��Ö�0.���v��#E��s�i1�aF�^N`c�@^tN=�4�'vԨu��#_x�Qiة1Tq��M�f⾰��R�x�!�"M�Za,��� U���P3�,&'��FBB��
��G� >0��
c̓f��]r�֑BmvM86o�9��	����8V�ݎIG��1�5!cD�H�21	bK��=����bK���}I���j[�2��I��#�`6�y�=�v�E#�DxZ�Z�h�I���n~��5� ��3Q�!�`Ծ�O60cg�NO%膣P7b�iQ�eS!s�F����A�.�
t!
דP��y�A��͖xz!�4��	�'^�<Q��d�G؞֘g�r]Iv���3�J�3F�W�v�,B��?'>r���\�}\��`��A� ٹ@�0O�p'c��{��`�%}B�0S�#eے� �*�o��p)�J	�0<ْ���H|0�[H!����d0�4��F����P�č8M��'��ѩܩ[��թ�,f�� ��$Q�/��hh���)80l�7��y��I?4�pa� g '@s^$�m�3M͖"<9�M5M%��J�IS��aUh֫C��U�P��tIa}��;ޙ
��T�O�6q!��Z��I��덉�Ld�˓D�󮄂S0t�K窌0��Up4�« "!𤔢��&X��r�`�`��.�:4�A�!����hM�S���ՍH�f��"!��X�2�� ��p���a ����a $��d�H���Rb ��x$�#�lʭ6�M���'R�@�C�NbM��h����H�R`��D�3�����mB���r"�����7HZ��;%�T(�ވy�
H���#<� j)�ЅF�
!N��#�=Ag�U����O�h����y�J� �z>������.�T��s���A���㫑�'8
m��EE��͙U��Y�B�Oۚ�Z�oy<	ŉ1CQ,H�2D!]��-�|>!EyR�2�,I�6L�%�?��DU5:`��y�D��x	���Doax��d�|�I4�f��y餢
=pz�dQ����n'�%�bdk��쑣o[v?9u'Y6c3�Y��n?O :�d_/(��ba#�;o�:5���9��V
7^VthF�� �����O�����&Y��`��xu�=:p�Xh<�2�5~T��Re�I6�ေ.��hs�P�C\.��	.Xk����$�V]?ͻX�t$@Ѩė�(�@�1���D}�FW"T��P��9���Ǝa�0��įm�|C	���a\�l*�S��s!@U�Y��E���[7B��T��V!�� ̓[��t!�"?�i��I%)�l�5��x�DI7ESs��2��Ƃ}��x�P���x�AR�&x��Q�H�6��ĪR�i��ɿ�~R��44I�3��kRN���Sy3�J1(��sh�%ڂ�ZC����$�/��ə��)6���m	8{�|M��%_4�0�`��K�XQ���3�Ǵ=��e���iζ<Qp��6 ���s�N.W�^q�ՠ٬q�#>�M�=n@�?7튎u�D���掭8,Ru;g��	j>�/O�J��1 �6���k��j��g�D�$s��m�w����8s�G+y��$Ȇ:�:�{Z�~���w?x���E�3%Ja���}[��C�@�%�r�C��m��0����D��ISדŒ�3�IC=;":P�g$�2"���'�Du�%Ć�)��H2>�8h�cCL.��P@h��ɛ�o�B������ ��dk6��a~J)k�(`ޖ*��\#�jH6�6Y� �I�yr�/��c`�i��cƦJwP]E��JY=���R�Ơ>I�����I�(O�� �Z<����V�ր~ɪ����O�����X,?���RB��1v����^+L)����<�za��@�h����H��PF�'!�&�������A��0!�+a2&�����'��B!ª��q�'��L�u���1���N�r�X��a�#8'Za#WeYXhE(�5\OV9�!ۛRh ��T0B�(�Rwo��0��d� ��
D�{�n�mZM�ڐ���ahv��ѣڿR����I�^U������H4��M�6,�lQ!�DY:(!,����?�	�P��@⫙�?a�dJ��?�yQ���#�D$H0�r�J�{Pυ+�O�r�.Zy�`�J�h�?ZdN��󘟸�hR�NĒ�·�:SH({D��[ v� ��'m|I�7��R}���b��>	�G1|TIEHY�>���*e ې0|�x�W����'�I�����ɵs�|�CHB q�h�sm߃R�X\�'A�\Q�z��X���Fdbx
gN��PR�E��4T�џ0 �C3R��	=-�PLr�'��M��CGK�,F��y�$�-LOހ�!hr<]�n��|�J�� F֏HV��	wh�0bZx��⪄�O�d��ɽ0�!��W�i.�Skq�O�0����� ����5��V�� �q@�R��(#��X�,��!(O��z�GE�d�@iyք$O�.lJ ��'�TJR��'�(��R%��:vn^�VL;�.��~�0T0�z:rfN��~�JS��'�L9�&�Ɵ��ĳ�D}��6�BT%��>Yu!���V�б��-L�ܠ�ŀ{q��*q�*�D�!Ov��Q�@5z�����A�[���!1O|%�[���f/W�/�p�yB�^N��L��ҵ��=#f'��g>���%��[���9#eS]��Wa!?�wNچb:��D�TN"���T�)��UX�w�qOb�h�,�<2��pAh�	�>qr�ݗ2�`!�	o�RۆH��y��Q�]e�ܹ�F	�PZ��A֣��G�
7��{��))ODJӠ�Ο����w�b�@��# �����i	�fUB`��'�,����X3A�, �	ɬc�b�[�'G�x�e!�ɧ���$�#{�8e�~"���F2K!�v�"�y�,��$v*�U�Z��!�D)	�������+oT����C�b�!�$�9)8P�١A�W¼P��:t�!��-C��(���Z!�tS��X�Z�!�D"U�����Y5�\ �TC>�!�0w�����[�IAdY�G�3�!�=A&�+� k��1WFDz�!�I[����p,�~S���Ѣի0T!��կ`X��%��i m*��"A9!��Z�%Ѥǆ>R[���`�M.[3!��E�^����끊�`���ΐ=:!�n����%��O��㳈�mh!��NN0 K���/��x(�HD8*a!���X�swL �W��`˦���l&!�� 
`��Ov��(��"b0�K$"Of�8�`�))� �C��6K�DY��"Oh(óT�o��h�G�$rM���"Of]*!�	9�`�5�N�w_fd"O�Q���׳�7*�IG4��"O�d:��"vP�!U�â ���0"O�̋�&	�9��i�c�V%�ތ��"O�q�Dl�7[��K��șg���b"O\��2��o�.8�S�J���@Z�"O�9����>�P$��$�J%4�C�"O�a+@0�u�V��U��Ms7"Op53So�1O̶-$��N\�s"O��mI�E���x�	�Ġ1�"O<U�w��0�Ĩ�����TѸɂ&"O.�+��LGH�0/x��ARB"O@���jP�Mk� �c��q9����"O���κEnXa �KQ�l$>�1"OhPpS��g�e��M?5�L��"O ܱ&�B
���ku��,�G"Oѓ��
i��I3��rˢ""O֠(�gP"���ɑCb�\�Y�"O���� �,?��As�KV�BAz�"O�\�$� <V4���H~�4��"O��I�IZZ��ps�ψ���"O��CK['|s e����@}f�"O�""+Ƭpl�Jw��rh)�6"O`ɋ2F&�<u bK�^p���u"Od%b��<�4���DU���T"O:t�i��Q|zdbS�K�lDb���"O���� �[j�غ�fÇkR
dy%"O����(+~�X�M�O�!��"Oh����,�"��K 0���D"O�]��dӲ_��`���^~���u"O|�r7��HS�(""��9y����"O�����O�RmI��	Ef���1"OJ����^��^a�� �kG��j�"O��`�É�x" �w��?=f�;B"O��:1@��XmR�Y*+;�hY`"O�A�b��C��eH���17%�]`�"O���RLI�6%)r.C$�4��g"O� s�o/d�1��,I�z�d"O\ `�Ý��Ԋ��̄Gظ(@"O
}B�及qs��jGk^�:H��"O`��M�*�
�S��L05." y "O�	Su��M���6,ĝS,(�آ"O8��`�ZF*�+#q:�pA"O����o�!V���BW���D^ �"OT���.�
����H��s"OLQ`7��.}���3���11���3"O�T� nȹC�pU��`��(�Ԣ�"O pS'cūv�~��ufJ�TRw"OH�A�'c��
pF��dFt�"O�ai��=�c�3s��7�6D���7����p��iN�>�j�� 
4D�4�f���Iނ0��瞬X�qA�&D��J@�x�5S%ަZ�f=K@%D�I�b�P����2��i�
�Гf=D�ls� 9���*	B��	�B@;D�0�DKD�\�0���0p�$D�ze�J�7f� v���`�>D��3&�W�bT5Z�¶-9D`;D�0�F��{6��C`@&-b���9D�b��ޫ�����E��1VU�7�7D�� r�
 ��i{�E��BqU7D�� ��Q��Y�Ѝ��`�O!���5"O�\��F�}�R�@&ϗ�^9D"O���5�_�
i�ԭ�/����"O8Uqn��ֹ`�H����"O���e��)�� �@�/�>4�"O`�S*�a�d�RT��($¤1+"O�x�$F�}w�Y�)�h ���@"O�9zK��\����批�@7"O*4�Zi렉�r��G?
H�*Uf�<!qOĭ^�V)'�ދ@V�i���Pe�<��N��)�)�)04�e�H|�<�$hT�;��qA��(lZ�#�/w�<����Oq~�i� :�`�Տ�]�<1B��u�ڙIv́7Y|"D�Y�<I g��_������4p���A���L�<�o�}n�裒إ	:��%CL�<��dJ>r6���B��:`v��b#�s�<��L�	6��i� �^�h����6�r�<)�m�(Ӷ�U�<=vJU�"q�<֧/J7HUX��[��UΛn�<٣i���6�fF*l*� Q�i�<A�r�R�y��Y!:�4� ҥ�J�<1�+@ "�(�G��*���MKI�<AԊ��5Rq/԰VB�r�j�<!f)�`��:�閯 b���b�c�<� �6YOhܢtȑ�Y�2���n�[�<Q��_�etF�:Ø(O���4�G~�<��ǅ}�L+tC��0��g-Ty�<��hJvpJQ@��@�Uul�Iх�w�<AD�J�kiFp��k�9g�"d��g�O�<q��*=`��hR��4��B�G�J�<ɔE�e���C����="b��G�<��-�&!�~ �)�V;> �i�@�<�E�-I40YPC䔆k�8�'�b�<Y�oR���I���`K�����W�<�&�̐I,,����G�B�#��y�<)B�>�mBaGU�x?*���Ju�<	���4�8)%��)�SW/9D���p��=D�X�!Bf[^�h\���;D��x��+��*g�\&*����5=D��s��E,`	2ms��Dx�����
7D�� �ӢHIJ��ჽ�l�8��5D���DB9<���hB�x;V)+'2D�0���֨k��t��-R+L�jU���0D�$#A�LX?�hJ�-�r�@؁I*D��X���3q�����It�aӲ�'D�hR�.�r�K�hR2?-Ƚ�R�)D�h��=,�饥.��u���%D�$3��=&m�����&*^Ez�!#D����#=c�b,!DIO=`�2����?D����\�|,�wF��}��4�<D��#c�kfja�3�*勀N;D������u����TH��`����:D�(P��r�fERQL�����3D����D�xN��$Ē��#�2D��IVb�r����,��g����A@%D����ۼ�Hh��̢b��s�"$D��7	S#��-��?�@�C�=D��QU�G�d*P;�'Jb��8X1�>LOT����iI�b�x}YF�L�S�|��2D����� �8�.$#�G�80�á`2D�X��ެa�����C��t� ��4D��r�*8a�:�ZD!� M&�)!�K5D�Pٴ��4k�J�k�	"r�3D�� �I�u�y���k�cѥsĶ�u�'ў"~���,R����ܓor�{��S3�y"�.xS��x�/?Q���F��y�*D��
���9Gtbg��3�y򬄬J*\�ӠM7C�� 	�FQ�y�fU5}ʸ	@�l
C�ȵ�\���<I��d����J�L��H�D��H
,!��
��E�b�ы09T!��HַD!�dJ��]������S3!��
J��|���7s�| ��h!�dHiD�������#����Bf�z�!�D��y/z�RVa�l���0'C�5�!�dR���)��hZ(6�Ĉ�AOM�o�!��;D@§��i�m��́+v�!�D�&Y@X�0g["&��Q��^x!���	 �B��qMn�,� ��'8�!�dD�J��������f��+A��|P!�H�"<�a���9+	&8�ˆ!nD!�$Z�N5p=1���{,]���T�!��<D�@`P�n�DL��K̾tt!�$�K�չ�*AVQ``KӬ !��L����aNc�0���땽G�!�T�����h��7�j�?C�!�$x�&��U*��rR
Y82�!7�!��A?�����7c6$h��j@w�!�ʀS]��#�@�*R.�;�Ԃ�!�ϧ4� 0�ǶS�yqeB�$f�!��<N�p}��˘Ov5+a ёy�!�d�Re!M%`�Q2�<j	� 	�'��	Rw!�/]�|��R �D��[�'㘝���D5]aV����[:<���!�'.�5�%M!w����,ȅEK:	�'���0Qb�>8��x��N
AF
(�'�8��@8B�$(!qo��<�<�	�'-�!{���!\�����<j��Di�'�,$�d�=MwNa���"cl�A�'����U�ǶtXz,��FY�W��P(�'���(LpX^��*�1`'@�)�'D��A����<"�-��B�4b�^ar�'�L#(9��H[E)K)��@��'\U Cn�&1p��+� <%ԚH��'�ў"~�qIC�|�,|*q��8��pa%�i�<���ڂ G��qQ"ŵX�t ��@e�<A����Y�$S- H��W�G �hO?�I/���BǠZ�-W�i(㦏�Z�6B����ZT�/�D5�!P�9!�B��9k���B��EZ؈�jϋ�C�Iu����!��'$�ݺS�͜��B�	�ĜZ��ʎj��7�ˠFטB��,nq���P�	���(�W�@6�B�	�5��i2 �	M���s���iFB�ɬa�DjQ&D@d����Zcj6B�I9:�>����1/�p��V��B䉧�rM�c�+�4衣�?q�B䉤,��l�0��I�x��ρ
Z��C�	�y��(��
�N�VPz��ԁe4�C�	(o���@�]
#a:�cQ�W�^�C�I"U�8yɡn��<15J��u�c��D{����#3��!�l�1��7�R��y�̹\F�!�J�0;vĂ��y�\>I�%���'3��b�B)�y2Ok�����I,�l���Z��y"���v?4��$��uvt��';�y�L�డãF�3"L�D�pE��y
� f�
 `A�$��cd"���RPA@"O��lʓ��µ��O�
�p3"O*t���4;���!��H'G� � �"O�(���G�܁�F�)�`\9�"O
9���5ze
@XvfݰNy��"O����$��ya&��K� �7"O|��PÈ�e涅��%; j�I��"O���$���s����Ձ\�N���"O���3녢��YA�AY�>~�)!"Ozp�b)�`�I�!�A1|�5"O�|{5>HZ�K&!!��P�"Ot\A3�ɮN`���	��ɢ"O�;�T=mU�D�>�⹲`"O�����K�|�$ˑ�H��6"O��3"
~�FiZ�
!�ٰ�"OTm�$��d^��)ȡ"��	9"O�X�c�5V��0B@"F�����"O���%^�)B�=*f��9}:�i�"O�9A��|k�PQ�D�^h�$A3"O�LRn��Q:,��Ä;:����"O����Q�<@�E�s������y����G�.��%ϐ|L����2�y�Lݭ)���Hߎj�	�Dk�<�y���$\u�t���ΧZ#�1���U0�yR�.6�LAJ0jU��3�N�3�y��6}*>�p��X� �\�h� S9�yb���#x��J�'DD��A��%�y`X� b�y�0���#�.� �yҁKX*�Ȫ���&�V�.�y��ĔEGڼ�BB�#2��P��!�yN�h�E�b!��(de�ZAZ���Q��m�G�Q�G6Lp���qՅȓG���z���Є�ˏ/��؄ȓ6rb��'�ܤ\Clc��H$Q
��ȓ9�	��k��E˓���L�$���:X聰L�/� �ᇀ�<����n�v-QC-4���m�D��d�ȓ0l�=�ԍ��]�� ��ԖL<�͆�Q�x��lw�FM���I��ȓy���P�� 72��� ��h���yg&�qd�j���Hu��VIt��te��I�BC�a�^(:A��&{�Ԍ�ȓ��qSJ5Q��<k�OM$Q:ن�J�>lJ�LS�BV��2�kϨ_�x�ȓ�2�A
$�|��j�#N�d��rh=��5A�\<
w�ڛa��h��|�i鵇��0����+�`�Խ��϶Ya䞽l�NQs aF2%�e�ȓiZ�G�Q�5�����J_(�ȓ[�q���!I�M����R4�ȓqqd00�^���ā�!�����"O�3@�&7�8�z�`R�D�D,1"O��ӂE�r�.�� U<^��8%"Ot��d�H1]L΁�F��k�t�"OT,Õ)6u�����O��u�Р��"O6��-��^�����JS!�J��hЈ���2�D�h��&,H!�$ʭ]��ࠬ�#'��s��[�pB!�]+'4�@�<%�I��`�Q!�& �� ��bY9/ĈE� S�-G!��! �Te�����d�G��@!�-.��� ���\��BKC�!�M"��2�	j���h�M7n�!��
<LhZ!�d�'�&@�1�G�]�!�� �ŀ����$���ߩ!�,ݐb"O�`�sn�.���x�";jg\�	g"O��9��ٝz��P�ga��]�ɡ"OR:7-�� ��N�W��dp�"O@�+s�
�4����a�6��"O0��i@�r���r��P3w�4x�"O��H�(�G�0U��ޗ.8��"Ob}�6*�PM8����@O�8@�v"O���c@�
���(�C�,��]�V"O����CWU��@�qbμd�VT��"O
i2�f�aL3恓(z��qB�"OΐKCBiXf4
T#ѿ2g��"O�R�Aβa�ȳ��1P�~�"Oj��Ag	"�M2B�݊�HeJ�"Oj�Rƪ"!��!Ri#C�
�)�"O~�p�Δ��>T:��W5PԦ��4"O���3��y�Ի�E��Z�pua"OVu#6�V2��K�[��t"O�@��B?N�h��CA��T�,��"O��Љ[N���t���Rt�A�"O}b��ʝ#�����@��/�����"O�XI	śi�n�;�!�-x�6m2�"Op	��Ø
P�a�O�L1��"O��kD�ǯ>?^�ĮԮ"�8� �"OEP�C�M�2IR�Hؾw�TMH�"O:T8񬌆n'�|��&��vp���r"O`����;+���1H�0_s@�2&"O.YYS�ϖ^h���&Ҷ ~��[W"O�irn�/�@1'X"88��"O��DI�q���%d)�b�"O�@SS�R3�R$0A�z� ��"O��`�C&��ۅ,���PY@"O�E*5�̘fZ�0	6��.l��
�"O������a���hT7:����t"O\QJ� �H��1�&*8�+�"OPTJ��t�a��	�"1\��"O�	ТJ(;b�)�b�u0�t	p"O~��k	q�@�w"I�_Θ�Q"OZ�[&�O>M��31b�5 @"O8S�c� �����hH9R�"O�|��x�\�2/�hK����"O��7��TQ�0Yp͕-A9d� �"O��4h��F%X ��ȹm� ���"O���G7>�W���Q��Hy"O��{@h�4��<C�	\��"ON�Z�a]���3�Q�^�R"O�I��HL>�����D_&4봈��"O�ɰtC�-~$��#M�؜9C`"O^��%�\�NT{�LA	C�d�@a"O�H��Z�c}�i�L� <�
�IQ"OH,����T&��P�q�� "OTY�'�A6)G�Za�˙z�N�!e"Oz����b�K��ert�C�"O ͹Pj�=Ol��(�(߮	W��"OH�� �g�`��$ż[���)3"O$���I)I�D���\�F�DZ"O��A���Q�	��aWc���!"Oh�XՌ��t1b�b�����A'"O�P@ ��1|�l��O�a��@�"O�4jӾ�z|;oP4x��"Ov�puH��o΀c�.^�}r$��R"O���,�?�0e��)r6�(W"O�e��J�(+�Q!��P���"O���#�ؕ	d8pbeN�K@���v"O� 19�Q�M[c�[;(b�"O֐�4��(��L��G	:��"O��Yą^�ua��s�˞�p��`Zr"ORY�����*X�c��"On����[���b�	��U2 "Ohi�/��,ct,�s���B��*�"O�P�N{�8��֠^)1&T8��"OZջ%lLL�#��(oB0�D"O����NԜ)=�th����.	����"O&)���]JN�4D�Z�p���"Oh]2�G�����Q��3R��0 �"O�-�����dΈy��\�i� �"O���c�C�JV���g�P8b��-	G"ONx���E�)Z�-��.ɚ��c"O4���%Y�\)+��߰w�҅��"O<�{?�T{Nֆl/��A�"Or��R'?Jx����/T���"ON40� �k�L:犛�L�Y��"O:P�� cN$�0$��x�"O�2���Ԩd��_�H�"O����οc5�]yעF5]�R��""O�� D�T���EzPh"��se"Ot�����[�*q 3��<B�Z�"O���B��uc�iӤ�Įu&�I� "Oh�Ѐa�Ġ!�"�K�
x1�w"Ox<k��Y)~��MrP.A�I���a"O�0�@�.�������0�Pu"O�-��
6ocQZ���wy��%"Of�kqKDNh`�Qe(o�:� P"O֕���=��E��#�ZH��"O�l�7jF8�Q!lG`���v"O.���G�[���k�j��T{g"O�u��*ômK�g
�!r��8�"O���J�Cgx�*v��3���I$"O<ܸf&F��s���4k����"O��`!(��f�����Nj�a��"O�X�"C@�t����m��B��5��"O�\�'�"��@ 7��a�Z���"O�jsi)itq��*�	)\�}�0"O��bU.ڥf�
%(3�ϏPTy��"O���{YT�5
��28��F"O0E��!L�0�����.)�E�"O��R2�+HI�舛%?�� 4"O���F,�t L��'à Y�8�s"O�yc��-#���>>��"�"Ob=pR�S<unn��%̆
TҘ��"O�]1��Q�+�m[�+D�Ja�!u"OPyԆG�7�Y�Ċ�<L��l�"O
�9��@5�6`��*�B����"O*L)ԨO��µ��"�.J4�pt"O ��S�S�b��<��	�+3"��"On�q���(P��c�H�Әݸ"O��b'/��H���$梙J�"O��ff������&������"OT�����8�G%ܲ^�����"OJ���D#�U+d�#N�@�ѣ"OXd���Ğx�l��(�����("O�	�$��6���%�N��<:�"OP(uN،��V�,"��x"O�ܠ�@��*�޴�B��8?`ܩD"OЄc�C͗H�
ԙԀR(����"OX��"ךF&�x��R9�V1hg"O�|�����+2�Ԣ�J�+a�0�RP"O>�bg�Pw�M���I��-25"O� ���!B;���2�)`���C"O�t��Ý0is�Bm�0}#8P"O�����C����۳��S>��j�"O�p� ]/+���`�$d)X��$"O��Z:?�UÂE�-B8��b"O܀Id N�aS)0�m�-b	F���"OPH�j��g���B훒mL�PJ�"O���%�h�� K�l�wH�d"t"O|( ��*L$D�Ǌ�1@ �"O~� u�F�P�!I��*z�zai%"O<%V@V*%V1����G&��"Ol���'Δ4BX�h�9_3��)�"OT�%J��viv�0�e+x��"O0���.H8+b��C��a�qJ�"O6D�F�!K����P�ʗu�x"ON��C�A�	���Hj�"�"O4���U(q�p����|�F�C"O ���g���1Q�@�bh�9R"OJE�稍�F�@��ЗS(�y05"O��H��>v�<�Sk��|�S@"O�șP"5�D�tl��
F�J�"O�4�e#�!{d��Cl�=�(��"O�����ڏ��s�'�n3�"O�t���I(��@�r��;��	Ku"O�9�� �l,hbF@�< Ϊe"O@�k�(�#��������*��X3"O���4�
�Bh�e��9�0��e"Or9��
#\F]��\<�R"Ole�#đ:���:����<�P\��"O@EIs�9E�h�h��H+�jU��"O���`L�S�:�N��QbG"Of�PȈ�n۪!h�DˮUs�:@"O�,Y�lU A����D2v�	"O6Y��֫rMZ�W뙶)�)D"O(���,]�9u
]��*_#O��[�"O�
�����q��f�?��LR "O�A�AH���D(���G�R�:�"O�b���\Yj�A�~�Q"OB	0ں}���◠�R`,U�2"O,�H2
͋�̨*�/D:N4ҥp�"O�`�U���Q�G�JCh��"O�lXw@ŗns U��a��J/�T�"O�����
o��i*qOm$�s"O�Y�� T�0�Q �=��`�"OKF�&%�
 �DĎ�F=!�$Y��� ��[�Rٞ�fi�*!����(��a�c��QG��(!��+n�P\�S��"{���F�!\�!򤋙I���;��J:DKY�����_c!�$�Iw���	T�<IB]����*O�!�D�dE��d�%,L@�c�'�!�dқa0�U�1kܴn���6�%!�D�uά{Ч+
�.��T�S�	!�wܱ1$٬uy*�@�'{�!�Mz�X���)�*irxٳoE4�!�D��.4�B�jM�p�fH��M�3A�!�d�"G�x�۠�	�etl����\�;�!�2=�Y��5
SD3��+ �!��s�nm�e��~_�t	�H�xV!�d�+:,�Ū��!B��u�s>!�DH�]F�x�'T,n�ԩ���'[�!�DJ�h�2�8����f�ў^r!�F�,���qL����١d!�$�����B�� 6����!�� �����sr�`Óq�4�#"O<l�B�8%{��x��߷2i�T�!"O��S@	 ^@�C���:aw@ȘS"O��_�
�Xs�DH\��@�"OPZa���f��p��PC�"OvyeES\�ȸ`.A5`9�)��"O��")3T���N�:7���j�"Ol��"՟p��Q�\�tm�$"O(����_8p���BBK��og��"O��ӆ� B�|�W��b*���F"O��b���!��]�r�����x�Q�p���9;�ř !�d^&(��V5m��B�I
f����]/{�����0C��B�	� G�	��l�+!QEԗ~�xB�I*T(ji������(�ӉB>B���RA!�ܿJ���ag	Kx B�	hl�P)�НxA��A��R�.��C��!�(�2�B!)~`�˧��d=�C�I(k)|�x�f�:Ic���w�L/��C�\��1Ҧ�T�We~�3��&0;�C�	,*r꼱sʆ�1L�k1��:H_�B�I�"��H@dQ8�$��1dA"`B�C�	�lL�<V
Y�yG��7���|EzC䉛sV� �v-�:x@�+�o�G*B䉰C�"M��	��bv�ic��/j�(B䉊5�iʖ$
e�������l/B�I<3V*5��2+�\�b���T<B�I��X���'� ���B�1��B�ɺpOڽ2A��#c~hp�߽T8�B䉳1;�ĉ7(L���吃eÀP��C��u��\��-�2l�
�h���t���O����V��V|Y0b%F$J�9�Hݳ�!�$�SƺH�g�)M�pѲ�_8V^!�č�i�h�c��0b��d#��)iZ!�dnM�ɒ�A�}�\I��JS+�Py��@t�P�b��+w�ʕ�D�M�yrG�5T�b�Kw��v�ؘ�T.���yrɌ�c90���K��#">��B��y�!��ZE
h@� ͫLA�d�6�T���.�OȸDo�m�f�ħ^�w�X
G"O�Q��π�p�F�l��Z�"OF���n]d̔-b��wȎ��w"O�5
�O�WbNp�B��:6�0��2"O�9�p=���Y�ѷ:іT�"O6�[w�-�*����J�'p��d"Ox��ܨH�\����R���3"O�+�Y�e\��{6% >d�Ό�"O�Ѓ6�+W�l��գS=i��p"O�|[ӈ�'rM��6����%�B
�y	o|��Q�DG_�MP� ��y����~�d
^:H,�t���	��y
�P�\�������@r'�9�y�ٴ8�
t�f/�@*�`��X �y�O�W��m�1h�2�n����ʸ�yR@��l�R�"��	 a��O�9�y҈�|N�LK¦_w�8( ��^	�y2L��,SF��U�3p�R���T�yr�:�>��v�658�x�W���y�C� �F��Ԋؼ-',�����3�y2"M- �y	��_�&��$�g���y��.��0�@&7��Mc�g۲�yR(�m�ڜ�GΚ6 �YBT/�y�y�\�p%��$/�.1ȩ�yb!8]| ,�4�@��ROF!�y
� p�ar�gjy)�jӵ��]"O&�@rj��f�|0���O�{E����"O�ఀ�U!D9�@ƌηޒ�G"OޕC1�GY�Mc�L1-�С[�"O: hci_C($c%�ܡg���"OpM��lY\�||ٴ䜫�$���"O0u#Ӧ��`�h���%Q�C�����"O�e�6ą%H)�嘒D��f��Ԑc"O�T��^�q�-��H�`�#"O�aA��ƈx�����P?"�m��"O1���M (BM!�cE,�v���"O�*� ��F՚� ���0"O�`J��H�b��QPa�;	��V"O�5�DJH:]xEj�%����P�e"O�
%B.b�*6*�8}2!
�"O0]	F��=����R[D8e	�"O Qʵj�.��	v�( `x�B"O^��NI�&)��@C��:m��%�&"OH]��N�H&p����p��D�"O6���'i)<�9��M�2�<dxc"OV�B4��#�"�R�ݒ$�6}i�"ONq�7�[&~@�U�ς� ����"O�����$#4��i�ЭJ!"O�=3*��EBeԃ�1A�"O@�S%m͒D��I�AR��MA0"O\��鉓#�R��@;b>���c"O,�1�B�D�0y�E-��~](d�c"O2����6 �!��.^�-^���C"O���#��N5�UP���yJ�!��"O����#�#�����i�O9�R�"O�aA�E:-E����I%��s�"O�9�f��)'���ۘ<NU6"Oб���׈�ެ8Q-��=���"O"�5��!LR4��fr.�"O`�0�~zZ�i�e�%bT,e��"OXJ�aۭE|�B�Oa;�T)�"Oj����"��BKZ�3�T{W"O����	xY���"D�M"��۶"Ot%��6uɠ�[#��"g^���"O40a���%��)*5!�3k "O~��VD�7_��`AB�T�\���"O `�V��m:]c����T֡�D"O�i�H�+�9��2/�
|��"O ����K�P=F=��n�H)ٶ"Od�ٰ+�3D�	.��Y��"O\���M�!�Ԍ�J�>>&�� "OR9T`��E�F �a-H�oL�(��"Oj	C�� A58�� ͎�uP�"O�y@�@�5Q�I��+��F�TH�0"Oh�&�W�9��`��#��*hjR�!�d�$]Ҥ1v�)Z>xݑ3���!�Hr�d�Y���4�U�Ɔ�!�!�đ�?��!J�"Iqe!���J�V���&�1�	Ц|!�d������2I,$2eF��!�$�e��L3���o%Ty:���r�!�$W�!�PU�h�<�1J�%Yw!�D 0pv��Q�H}��( �ƲRJ!�7u���q̋��*��0�!��@�U���d�HI���.9%!���LIƄU�-���%�9�!���:,�����C�$O!��<����OT�<�2�X ���!��O*$
8dHe*=�lA�oє_�!�� hTpA�]o��4n���0�"O���!��'eI�؉R�K�b���W"O8Q�T�J�&���U;3�b���"O
�u`_�\����r,E;8Θ�B�"O �"7��D3��ȃ)��8%R�"O<��Pd^�^"�D���	i�>�ۑ"O�EK�D�,�l!�,�J��V"O��w-ʤ����u,[�M � "O��Q�G��_(fJ��_<ZltxA"O ��lY�e�l �Á�(NP���V"O��+A�=h���#��T�]Ѥh"O�i���bF41���U qZF"O:�+���x/(h�箉 *A�b"O�mc��0��%(�.#M�H-��"Ol<���ME`@��ץj��8�"O���&�Q�B/L�N|@��$ȗ%�!��V�d	�NA�%�T-��cN�z�!�F��P���H��
��#�z�!��A�>% $I�|m���R"���!�$?���J��@�A��y !�$C��LɛEj �`��t:ǥ^�-�!�䇋&�p��d��^���I���u�!�$N+
G�d���*���"cdQ G�!򤁌6s�i���}.��5�!�$����+���eR�� ̻b�!�d6~��=Q�C^j����b�*�!��K1Z� �+!�{z��n�5�!�D�=
���{��'Ks�t*��P?iz!�DA��F� 5	�)U� !�79!���,��/:c��<PO:1�!�P�)��� X7-�V�@��?�!�N�dY*G6q�\`k[S�!��3Q���g	�3t�����\�!�ݻdsV�j�IK-ii�d� T��!�Q7�$�	K�K��I���)�!�dL�V?��c��Ǡ~Gj݁CFñ�!��n�<pA�K�63�i��O�:��O��=��B�xG��9Q�$=\	>�{�"O�Ր��CĖ�j�aQ/��"O֤��f�0]z�)�`�:k�h�u"O��Is�^�8������P�l��iq�"O��V�Rv�� p�@.Ȱ��A"O�U��T�U��Aܰv4��""O8l��#J5s������o��M�E�|b�)��,aD�{�����y)����K�(C�I �pQ!�իX��Mz��V�[ $C䉯:Dmd��Pc��C���k)�C�	�2̅��A�juSeF��#ҢC��aj>�@�ܔB��ڵ��F�C���<�H�F��);�+A�PC�I��¡Y���
�;��;!pC�	 6(���n�d>����bѐjq6C��*��(#�`^��|���J�,%6C�I���d�3�F'��ȐGH�K�"C�IV\\j�@�K$���p5Y�B�	4"�jX#�C�KF�	�� � gA�B�I E���*����셛6�B�	GV]B�K��y.�`����-mhC�9��Yk��Ƹ&��l��O�[�TC�ɆX+�Б��>^��GG�? NC䉡[���+�1w<d����4�lB�'F��e�烒�4΍3��D�.�JB�ɢY>�!ʢJͽ �*�իo�$B�	�6���*�@�$��͋7�S�^n�C�)� �Ɇ��a���Q1� �мP��w��Ң��<-Ҁ�j�Y�z���0Qc9D��8�������d G�L�d(6D��)֯Z?? ���DN�
<�{V�8D��Ҋ��b��x`D��/c2����!8D�$+�D�=��zV��t_8 ��)!D����j�� 9d�Q2�x�?D�,@���'&�Ty�)Гx�4Z�f�<I���S]%ΕH%���D�|��+��h�,C��:x醕iT�����9G잫�fB�ɥO�`�x�8G(�-�v/�,w�B�_>��z$k��Tz�9H��΀(�B��	+�|Ё]�F����ˏ�
C�	5mRD}���,h��N��(�B�I�Vy`�#�BD�Y{���nۍ6�ʓ�0?��'���F�8%cωYX�1��V�<�0e�Y�4t��DH�z5��^�<�/F.p�
DB"nÀ����Ho�<qa��*?���W���rK-JP��g�<92(3/��UI5g̲#�~���_y�<�$���6��
�I:"����R�L���̓*���e�P�.�l��NH֠y��B�U�aC�JB�2�
�42���Wu��	C*��j��p	��m�Ň��PJc�4P��%:W��m���ȓL�D��c�����hϭ7�Z���!� �@�� .�P�)S� V�ȓV��[Aȩ�rP�"�׫{��4��8M��P�GI.U~�D���&�ִ&�DD{��4�ȯK����F�'�n������y��G;SM~@[��Ï>��#�C<�y�f97$1��U� �����ې�y��զ%����d���1Sg���y�J�K�\Y�Ӎ��[��U[�'C��yHCQp�ʕ� Y�4��E��ybHFLZ�k�O�B�&�#��0�y2�&x����"U�db��I����y�Oޖ2�p��J82�l9k$ψ�yB�F1$�8  sM�%UF�%�P#���yr�N O_�q�ʂE�P��ܿ�y"�Bu&LQ�MM/7�8�K�c��y"Δ\�aQ�o\�'���:�c�yң�-6@,�G�7rR���� �y�-TL�P�+夋
K.�,u�L��yr�K�a��<Y��՝?����jL��y��\�xv>t��go���|��ȓ E�ɴ��8V�Z�ZRF�vU�|��#��P�Z��q�aڒnf���ȓ'f��PĊ^�PA�̦8��u��(
�����0P���@k�:8Mr��ȓB�B,�&�TQn�;���x����ȓu:L���K�cw	�%*X��ȓT����Պ�,	e��r`"� �6Ʌȓby���6�
�v�z���@J���ȓjw���`ɪuy�����:ކE�� �l�Ѓ�N �A�	Z�#����O����a��F��I�+�1v��q��.А�Z �_#�p� M2_�r`��"A��`��_�"��(�$6�P�ȓe(}�RCĝ}�~��F`��Q�І�u�(�i�!��-Bc�Tm �ȓoZ�ثV � Hz|�&)��7Y�5�ȓ�ʗ�7� ���ա\a���ȓf���ru	U�#���sf��ć�S�? �$yR�ܹLI�xD��?x��s�"ObQ��C�1UI~x
�HԎs����"O���W��S�-�Ub�!NX��"Ob�"�`���)�/�p=�@S"OЈ	v͘�8� �
�mA~�xA�"Oz�2)K 	�nQ`b��AV�i�"Ov�Z�5��H�'�'M�*���"O��h�N͠I��˰%��"/a�@"O���v��1���Pf+WZ	"w"Ol0�s�u� h3ń�����"O���gE��0y��dS�z���"Or�!"��Kܾ��P�Q�^�6y P"Oq�f�F�U�̨j���3��p��"O��J�l�]�v���?�`-1�Q�����?�*8�2��0/l��y�E�)�PC�� \�ZT{���I]\񓱩� T�C�I�1�\ R�)�v�(��Aʏ�-��B�I�Ԑ��O�#R���!Uw�B��N@�D��e��0`�ߚg�B�I#6tN�C�MY�\F ��e�(j`�C�	+a
�hӅ��P��VlB��C��4C��i�E2H$�i��M2 �C�	6w��9Y��.[���� _�RC�	�`_��C�& Z�J�C�ыr�0C�I�.�� ��͎�e�4���0�NC䉭uк	0�OS4A���BQ7N��B�I
U
�h��N�Ov����6qB�	�<�chM�)L���� RjDB�	\5����j��p��U#��γd�>B�!�\Eʔ��64�lQ�#�ͅi�NC��O�q����&%f�pr^<|k�B�ɂNz�9ӥC�`���'I�9#��B�ɇ48�㤅�x�)����|�RB�I�p֜��%e� y��R��03/2B䉯C	 ���A��U~L`ac�ϤKK�B䉾^�t���
�&+�JȒ���@p"O�;���ZN�Q�K0:�2,�"Oj�����?1g��b�F<�q"O��4�yiۧI9% ((��P!�y�u6����g��������yR��/)zP�{��̑edֈ�sK��y2Aݚ(7�| ��P5�|4Z0#���y��@�es�� 0hJ�<6��)	��yr��<6��᱓��w�CdX��y�.�l��,yFH�}%�LB���y�j���.�a'�A�r��"����yR(��fC��q-%o4�Yi ��y��.��A�'�]�w��!�
�y��

|,��A`ʹ|���Zu�J���0>��̝o_��3w��4O��rv&�B�<��_3+������&⦰j���@�<�%d�8L�ذ� �Ӕ|T`��R�<�@j@�F�4�A��ȼ#v��L�<YE�L�<b*l��I�]�\)���I�<�b��6q	��Dߘt[�,@��FH�<�C��x�J�bAb�=/	���i�<	�F��	�p�[�NғG.�0��b�<�uI�b��=`���5��  /�Y�<��#!!���D�,���p�UO�<���:nh�|鳀ïI��� �!FN�<Y����d]��1�N	�J��Yp!�RI�<��3=�乘�E�)^byS)�G�<)F��uxJQ�N͉8���S�Lz�<�MɮJ�i��(IE��Ls��^w�<� ��"ç�)m������
.I,�� �"O����l��]�z�ڳ�D�a�"O��x�dG-l���'�; ���"O�U�$"L�??�l!��O�TS3"O��cClFhbr̟g�U1"O>��58�3a�R
R��!ZE�'�!�V�}���Պ&!o\���m��t�!�$^�D�v�36�>04��+i!�D���x���c�t��7��p?!��X�*C�/��ӊ=P�NBT[!�D90pu�e癄�+��+����v��dXQ�L	?:����=r\��?�ӓ�n$I����K���(&�~�4��p���zw
�2��p�K�8�J�ȓ�pK �Q � rJޛ}�P9��`<V���'vm,�+P�ذ �*5�ȓ�$��L�:�ؽke�P����ȓ.����hU'o��ĒCG͓yv~��ȓd&����HN����) �V���B�\�u-�I��Q�ԋŉ5����+O�˓�0=��@�73�l��' X�?5�5"׋	D�<q@,\&G.��)w�@"�4"�Xg�<��*G:p�ˑD_���Y1�^{�<qW����9f�}�^�J�t�<�1�!/��8"�^b`j�
�p�<A���>7�S��|�Ą9�.�q�<q�	[v}!�(�2	 ��ƒm�<�R����T^���+�`�<Y�	@
P�D�Ӏ�NT�R#AT�<�Q▵n-U�
�p�"W'�S�<)E� �{뮵�u�B�R���_O�<Y��V�W�n�J��\ |m����I�<�I]x.RM�'HF�<�V`qB ��<��Ɩ�،���d"lR%�R{�<�1�9�f��B/6MH8��v/�t�<���� *�L�A�߻[
x!�!�W�<�2�T,R80�p��>f`H�7e\�<���%qPᛤb�#I�fU)�QU�<!��_ya����-&�l1"�l�<�ы�zx��/�J���@��c�<��9D�@�(����21vy�P��^�<��	��2��e�-vv����Z�<�Ă��)�Ô�H������Z�<	�A�8d/���d'��>�]a�Y�<��E�D��E��*M�YӢ�p�<����&C��wI_�>^�d�"�n�<���J�&J�`B�� P��aJk�<��m\�垨)`N�&2��봆�o�<1DmY�n��q�'�	c�00S�]l�<�Dc(lO ���%�	u��ˤn�N�<����A0�-ˠĒ�A\T��m�J�<���J��jQ��k&2p�(��J�<�BOݐ p��JE�T#BSb�2e�M�< D	�3���`�ĕU-�̻���H�<�GO�?��$+���p�{��FF�<���$V���%�q���kFkn�<���V��`;GӅ2@����Hr�<ɲ�D�Qd���;>� �����y�<鴍�=�<a��@3?�"���͈s�<��X=q�����O�+v��9�4��p�<	5��e�^刦&�+~5␨�CMj�<���&5n�M;�����H��Of�<!�1&'f���E��[s� ��Am�<	��	tzm�C�rZ��Pt�<� �+�G�-|
beH7 "�f,�D"O�%Rs�x�Z��@5(%:��"O������@�����`�aj�[�"O`��f�o�R�b�)!�|��"Ox��c�W�l��d!QcO?F>IH�"O���u��g;���s��� �L�@�"O� y!J�)�x��eg<'�ܕ@"Oؑp��Т���P��(}��D@�"O�� ���QS&�)Cd��b��X��"O�uC0@=U�xT�q"�0f���"Ox�.t���;y���u�F>!��F�L#���'�ѹ�B�7!�D�cP ё7�@�q�㈹*!�dx(���څ-� ̐�B
]w!�V�oȹ�׊ο�!	S&�0l�!�DĖB
x������Y�A��!�d�	;%2��"��z���0��̅3�!�$Z�%�uR��E-�P+��ٓ&|!���v����'	�)Ġ�T�I9�!�Dׇn�ެб�"<�f1����E!���%e���O���a *�D!���G���"�Հ(�l��O	&!�DυR�F���ST��؂�ޮ:!�$T?_|� J�ce�u /��.�!�D�Њ���Ä7TU�V�t{f�S�'���y4���pM~i�$��$g  8�'
�"@�-!&�I�Ç�e��8��'>\��)ߐ# X��uk�d��'u"� &ޒWb�!�ǀ9 ����'%��E��)P���HݢS�q�A*O��A��#l��b�'�#T�U�'���0QW5y�Ի��J3j~�H
�'�"��V̀9'B�Zt�8�~%
�'زhc��4��a�`D[�
�~ Q�'�f�i���|x~l���46�6�8	�'�\��E|���NI�z�>�B�'��Q+�/X^�z=�uD�x�8 s�'����'d_�i��ȴZ�Ji��'����&��A`Z�h�CI	�\! �'}p�2uĒDfF�pf�Ӄx����'g$�2oQ�SR����n ��
�'����ոh`)�!�9_w��A�'Q$�+SLߡ4��/*���'��H:`#	�or�z���z�F�P�'%8��'F+TP\�����d�Zu�	�'�ʍP�f��a�Btad��	N�Ԩ�'����R�A��>�zr��7С�'�T��n=~Rh��T�1��r�'�^�K�QF���(�<����'�6P����XNLuR1��3��5��'�3��nJ ѳ��V"(��	B�'�aKF��܋�k?h��'�v	���'Bnt` �5.v��
�'� ��g� @��Y��V�0vdh��'0V���E����x�ߕ/�ƅ)�'�� �bʖ.u��8���(\5��'���ɲᖣV���qNW�Z	�	�'�l��t�X_��Jr �Oy@��	�'߈h�e�B7B����RK��JQ���
�'�:P�3f ���$���9���
�'�2 Y0���h$��e�9{����'�&�a6�6�B��Ŏ�I����'&N-�%��*�ؘ�r�]/@��!��'�r`)��-m�l0�C�:ttA���� ���ƨ�~�Lx;6e��� %� "O��SSnH�;�����D%?Pp�؃"O �ѕ <#�~��V:��V"OJ���h9�NA��k�=7�<i�"O><�3��T(U�;%/�Y��"OP��FB*@�`tS��
B>�� "O�� b�5�6y���J����"OAZ�Ȏ6�l���iE/DV�`҂"O��!b/Xb5yf�4~[B�c&"O�=y�������
eJI40J�2"O��zE.�w���ےK�P,��"O��ڥ�04�B9�w��#Q�`Zu"O~�2�n�B�ʨC$K�9>�\{4"O�h��aϪ ީ@��� T�x�"O���T�/Q�q���R�Ol�MZ�"O``bB��6�A3Ll"dQ"O�P��ʂ<9�!�IU0>S��c�"O
���Ӻ9�|Zr�X �~�`�"O�E�e$r(�:g��F�0��6D�:�+�iv	)dJ��B��6.!D���wIƖc�����d�z���t�:D�����ۍ:�	ڃ�WOX	��D7D���4�Z{x�;E!�O"P�H%E(D�H��_58�T$�P�T������0D��:�U=}EX9��Ҡa�P�X�&0D�da@�Z�j�P��9e�* [��.D��
�c�������ڲa�5:�!(D�|2��-Ig�}�@gZ�k]���$D���o�M.�@�� ]�\F̌�!D���b˴~.�c5	�1mB����?D���&��9w��i��P4z�Ze<D��ᔁ_+2�ɆS�N@�QH%D��k�@_��2��bJ!�F��`�0D�J��-?���$ B���&2D�8�F�,.��`��+):h�7!.D�(��e�쐠�H�'�&�+D�,���Œ0<�iie�����ط�4D���G�a�܄�ҩ��&�Y���(D�|� �"s�l`Q��_��^���%D���FN�L�|50��Z͂�0�$D��+��Z!n��!��b^�Arv��w�&D�l�����.d���0�@'�X��a�&D������/W=����O08N8�6F0D��+�IƵn��5��Y���4�sL/D��)��+�eC�����8aF(D���*$o�^%rCU�g��P�q�)D�Ī��M�$9�t"P���QJ)��:D��r��0&PR�&։I�0-��5D����,R�I��(��h\M$!��2D���6m3.S@�4��^�hb&D�lhG�S�|�cRM@�"K��@�9D��ȕ$!(b5kF�0��x��<D�L+Ǡ��xl� ���-g�F,�l9D�|�B*T*_��h+	���"3D�H�4���-�!j1j��!qp1��,/D���Ǣ������w�ژy4m��/0D�`��CҙO�t�ǩL�7��<��O,D�x�-�d�ZCݖ7���r5E%D���7��`����#O�G������-D�$ڥ�̀I�hr��R�S��Y�c�!D����aV�� �ڶK�co�1��?D�Lc��ZP�r	B���b,�E8w�(D�4��oʱ2�NBţ�eӸ	�C�'D�P*5'GkU� �A�ڪc���$D�� (�)�'T)wT2D�DmѼ�RP"Oh�@EGGAF>��"�����Bu"O� Z��
�N]��
7`@�t��̫E"O����]>rށď
;@t��Y�"OdpÃƁJ���ɏ�	@�ۥ"OL�"`Y� ������0b:�"O��#T��>a���_�_�쀨B"O����A�&v�U`gr���"O����I%+}��� �.V  b�"O�a�S�^-~�|��Ǡ[%��YD"OF�p`Ƒ�����Oї0#�D�"O }�J���ak������a$"OƠ b�ԝn�v9#�گ2]��*P"O�qQPH+B�.	�
��#�4��f"OH��s--b����P�xi!�"O��JՃE�"��0�5
;E�Ly{P"O�Jw͒.�$�Pd-Q1�F�[w"O   ��1B<��ʀ�/�@ѱ"O���䁶Ӻ����M�4p����"O
4a��ȓ|�
x���Bi�(1"O`)e��m� Z��\QP���"O�(p�H�i+��P���/B>�!�"O�5��
��p�*dQ�e��U'<���"O�QB�ǘ�r�� 䤟
M���"O@�3�Rnü�";�P9��"OL!�Q�Gbbͳ�0�^(��"OJ�����"ؕ@��ȕ{~���G"O�m�Ƙ2]�a��
��,�0Ыw"OȌ�dgֵV�M�i�:z���P"O`��N]*-��� ���-���`"O����"ۊ�������[�T�ç"O��3d�'��	�(.�,9^!��I��P8Ptƙ�b9�p4��,�!��LY�|�C�ĖeE&P37�O��!�.u2�I�f�]4 >��q��4 �!��!�(��D� 7�p�j��3�!� �!�I�5�_�}�xLR�h��C�!�DNhA(��5fڻl��4I��U �!�D�;\߮��� i�z�"�Ȅ�p�!�$D�C��mvJ�r��p��B��!�D������b�����"��C�	��c�d�����#pC�I�A�����
����<zC�I�&���'�R�
� �M<IƪC䉝}\<k�(�8g������|K6B�	�M���
fa�.��[��I1[(B��*�xؒ��ѷ\�d�qc���D�B�~�(L�g! ��I�0!��[�:����U�1�0��MH!�.�d�( �˯0f��*t� 'Le!�N�{
T!f�6G�(('ˊ6O!�dέ`J�a��#�|a�֋R �!��ۺt���q7G �y%T�&��
2�!�	/|2���eC�/_�K�IQ
6�!�D�+:�IҠ=>�Ĩ2�I?^�!�DĘw
I8�l��1�y�s 2e!�D�&w|�,�aƵ��YP��GW!��<=�Z�5G-��H�M�><!�I�{��b���w��!s�Yj2!�ҥV�dyA���!b^ظ�/o�!�d߽O���R� h�0L�� �09n!�$�4��y�gfX}�Ν� o˸l!�@;t���01�K�޼@X��!�D�/.L�EP4
̓T8�CAe��a�!�� f�(�C��s�2!�R+0A1�"O�d*eK%Bh�����)����"OX!��l\�s�Z�K��'d����"O����/t@'���;�^Ū�"O�X8'Hn�����mE��̋"O�L�D�K�"6���ͲI���A"O�E8&)#B��@7\��պ�"O����F��h�T��:{���a"O�{�LW���\K���7kذ<�P"O����̔T�Ь����,wZX�"O�t�b�P�@d�J�nՐWb�PA"O��Fe��0|e��
$[V�Jr"O�}H4�nSXf�^a;��J�"O>�y��P�_��Ұ�F)O�>=�4"O.�q¨������ȅ�E�,Y�%"O�-1h��y�"�ȉ{�Xm�"OlmP�W��L�ǆ�e��!���O���d�!i&�E)"+�R�=��GϹh?��!�S���K~R�V�^�Na`�ď/��Z��̠�yrm�:r��Xƒ�|{�)y�	���'�O�UiG&ӫh�*��VHY�=�����'O6��' ���bP�� w�[-mA���'5^!R�ƀ�ne�%%1J<�Y�6���'�ޕ��ˑvn��HЁ��5�'.��q�+�h:�����9y�0�	�'���+v�Śy%�S7��� r!��'B��e���(��섴t���c��D1OJ�ɷ�{�l8��	��V{�\`�"O������[(pR��W4k`Q���	}x�p���tb������3P+,D�\;g��-��� !��# �jQp"�<A���ӕA��,-f@s�E����$��F{������zr~:�@ºO���'���y2�Z�$�>�Go�D����@�.�yrN�&��6E�=(Q��A�lC��yBD�5[c�T�Va�$dtZP�Z��yR*Ѷ&�HD�E/���l�J�@X�y�۩c�� �6�V�(1(E��y� ��\)f�@���
&j��#�b�=�OƢ=�O@��J�><�4�Ӧ����fd�'DM��f�/
J��bI�{DT�h
ד��'je��H�� �I�H3$��	�'l.5@�(�!!R��CM�"`pŋ�y��a���O���@���y��0C�'x��	�'/�����܉%����B�w7r����DJ��p<�$��l:�/% ���VC�<ʀ�>l�����_ Xpb���{�<	�G�m�@�
�m�W^]z��P�<a�M�#]*�H�.�.~�^ec��PV�<��F2�J3�B.`{�`�Ty2�'�T�o��d���N�YHv
���$��1��XR'Fϛ^���
v�R��Py�H�TQ��L �H��@���8�y��	9���Bq�Z;H�hɓ& 1�yR�J�RyH���TShTm��c��y���:	�����x\i�%���y��6{�m�(�s���
�CO#��d2�O��ʺ��(�-��?T��P"O��ٔ�uH^9���F����0"O&4�׏�,>�\�{�H�_�<���'������edv)h�n����KsIz����ɽk�v!S$�!"NM�P�Q��h��/�S�i5�d˃�<�;����D�Vp)0�A/PL!��9@�.Q�Qe��d��!	D�_�O���� �-:�O�$2�$915�ԃ�4݋f"Oj��4&Q:b�*���X<Z2"O���6 ϛИa�ף��'IBYP�'q�O^X3!�*L��y� ��&nP,�JGf�<�w˖�q�1Z�H��<�tR�&�^�<�2��
Z ��:��I�q��}SG�W�<�pdV�V��,�AĒ�B���r�i�R̓��=1��G?9�b�Z�M
W�ԝ�%��g��Ĕ't��`/���H�C�nY&D:�9�'k���C�6F�R����̩q�DMs���"��iQ3+0Ĉ!I�$G�PbW�ˈy!��(����肨|���a#%N�/�1O��'�I=иOƚ�ٗ*�F��1��)ȯDx� �'S�q���/	�k�n�T��'���!�Z��O���� 	(����D�(#^�a�GE�jv�|R�iKL�n�>q	�h��D���z���p�����y��'
n��q�P�*��	Vk�"G��������ȟ��[ �]	:	�!ZBM_�hB��d"O|����*��-����'��K$�'�ў"~JE��=O4�g�V�r˴�{�+��yR�,�Xyb�ˇ:{�a������yBF�[?���#�:פ��E���yҫ��wy�,f��bM�u��#	��y�LO	����@	V�`�=�#�G�y�`�f����'N�Y'��O��y�A�Y�E�V���r�¾�y�㓤>�(D�@�R�=�" ǟ�yR�C4u��ؘ�n�D��Y�q�U���'�ўb>M��%B�V2-̞�>�ڶe+,O��<��E0Y̘�F�)Z��e�`^�<!4"�-��P����{.D���Z�<�K�芙��_�0lQ����\/!�d_�G���Y#�l ��㔖R�!��7R��P�����t�BQc���!��^�KB�B9#¾,h ͑3�Oj|�B	/4~T���P�}onx2v"O�aP�dŷb&����5 g(�@"O��ñk\��z��Qߜ<b6��f�=�S�i��{8��5��*6�q��G	xc!��'�氐QhO�	� (b'G�9sўą�Ɂo���#�I�[։H�͠o:�B��p1\�HF�ɇ]�f1f���`�B�L�<�@֪Ĉ'���v�J�a�|B䉋4�(�d,�A��s�*Әy�nB�&�\�Ků��*\��6i�8~,O��xJ��c�pI+��&:T�@��$�����gEy[���c(�$Y|�x�/"�	���O�\���U�%���1`�%*���
�'#DX���\LG����&D�P�
�'�l��p��W�| ���2���	�'��y(�е/�xT���ɯ
)��	�'U��3�ā�Q�L��MJ"rV�8˓�'A2�L9uK:�ä�Y�hkz,#�C�	&�!���4r����B)��h�i�ף]��ID�'��SV�'�2T0���".�mA3@#Ps�����U?�P��l(.��F�WeVr�B�G�<A��4a\j���Xa@`�(�X�'�1O��'n���R2���>}����c�z���}�2�K���bU�P�@��?���F{��O���v��$��[7	�<X	��'D{��
<d����,�|�'�@�KE�(Hh��4�э
�y�$�1O�t����T>M�eB<�y�N���{����85��䂥�1O��S��y
� �H�B��'ը�yCKW�+]F-{a"O�a�疧]���S��i=�Qҥ"O��BPB��(�zlz�e+����OƔ��f��)H1�\�tf���'du�<��(ߋr�v@a�'R�3����U��{�<AtH¸f���+O�}H<D�k�N�<Ѵ�݈j��I(�柪)�Hud�A�<�e�թ�8
�l�l��U(d��U�<�1�Y/t�B!"l�Q�8	�B}�<	�E͔��`H�,�,41@�a�<�"�k|%�5��$݀5C3F�]�<	3!��UVʽY��$G\<����WZ�<YQ#ߝ#���y�,^�4���W�<�G�@�d�вB�#X�ݠ��_�<�u!�3l
��@䒟%�`���[X�<�f
 vb^S �Ʋ4�����QN�<y�)�A�ݒ�.�''R%+���s�<�C���!����Ɲ"9Ȧ]��)�d�<Y�<iz�)6�>NJ�
�M�w�<��h�r��S�P�70�ђ�_y�<1� ��]xzI� ��d���L�~�<)�m�>��AFc�J@����|�<�2�G���SaΘ �^�Ôl�w�<)����C@���EŇ�p'.(���u�<GF]>���3��-q p�B"�[o�<��$,�	�1-��3df�z7)�m�<!G���V����cD���4 �m�<a�b�S���К3�� p��^�<��� F���[f�
�N�����\�<!�;f���C&`Д"b�+��	~�<Q�F��<��pTf��0����@�<���-4�� �h�@�
5@�eGH�<9��.o��h�B��\ȱ��D�<�g&^��\ݱqI�6f�����*k�<��JQ�&~��!�m�X�x���HK�<�L�H]���X��35��P�<�(�? ���G@�o2pr�͟c�<�d`,V���@�`_;`4�A%�E�<1����eh�GMP*J˲���I�{�<�s��
���+���d��@	�z�<qRjHP�S�*��)2���$Z_�<!ä���X���&V��	k��NF�<1���@��ળ �B�2A����A�<�&�=Z�Ju�V�)u��� AXA�<�G� T��yb ��]i���!@�y�<���a�� .��pL@u�<�*S�M��$�#I'&��|9��n�<�2��2\-��Bpm�x��p0]i�<�*�14�S��T�\��y���b�<�Uh_�H��m�Bh�X"^xod��DYDï �����/E�\Z�fXe4�
�ヮ�:-�#�3D���/D�Xd(ՉǄڄ=؍���.D�T�#�S��� p����� �-D��!�_m��׋�+'�:i�� (D���M8}��@q��3��q31�)D��9�F�0<�j�(g��:يQ#*D������Uƌad٤Sx��n+D��p��H6����d.$� �2o#D���R�
8p!��
rc�a>F�� >D��RJ� EE���'=�,��=D��C�f"5j��T	�J�8���O'D���V�@�=�\�� �C�O���+7D��I �A!�C���`�z$
/D�4��7{�\c��#ιaa�(D�� �����A	;^���N�%g{*���"Odd��U�XB����P
��ڀ"O�e)0��j�GiӈaI�"O��C��P6�T ���ݷ(�.�`�"O$ �r�Ҽ5�E1u+Yh���"O���L�(t0j��hH�8�%"O4���Ń0�i�P��Ps"OT-#e�J�RdѴ�)�\�Xc"O|��uM�G��Ԁ�oN<Qx0H)�"O6���΃�xX*��
�T{�D�W"O&d�b���ܬ��mC�dPȰ��"O�5�A�*��d��a��*~8r�"O>��i̤sAl�����5"O�L�s*��*�X�r3k�E�x�"O�I�o-cO���h@\<���&"O<�@3$�d�4ܙe�Q(o%���"Ou[����ұ�I��I�X�"O̹���)�b�2"蜷���"O�-b���Df���E��i��Db�"w���XD�KX�(��'ڂP�R0yu$�*UJ�*6o1LO��B�ի'V��'��A��m�#TH�)��ݩ{;�K�'�
�J��P�!�`� N��bH>��C�M��Z`,Ԉ���� c�rl��;�I�1K�>0�"OV��cl�x;Z�1sH^+8��=�!�<��ȩ�S���,�F�g��Z�YR��+���U����E��c��J-��Q�s)�|��H`��J^����<�z0��i/�O ��F��9C�x��eT�&�^����'A�d�b�U;!�J���=O���]�)��5�Ë �J���{�"O��y���a����D�P�&����|��U�>��SK�%�?�AN
9t��}IWa�~�z���`(D�\���D<��Q���ւ�!�Fy�Z�áj�<vL������u֪!�0��^5�m)fIUf�hB�	�U8lF��i�s��K&�a� E�bsnD�6��q��*�E8q���	��2]Q#��<LO���T�,��p�'�ԍi��7+���'�B�)�Ҵ3�'�"+E�Ո&/r��tk (S2���{�H��(�@ز�S/x�N�p�o��a����ŦG>C�I

�B�B���>q9���!l�K��B�ɱ0��`���4S��Y��H��@T�B䉊���Bm4h��E��*��B䉜Nx�� �R�h����$�;+S.C� �ڌS��TrT���(A�k�B䉐0�4�ɢLθ'�(�1@e�"jSB�I���T�bI�P�,�q`�M���C��6��c!�ۛ?}�X���G��C���hsi\<�|X�#���C�I-O�0Rǉ��G`X��[�~`�C�	7~`04aQ-	-I�����ɖ0|C�	6V�J�1�$Mm��4����B����}q%A�]�6Ԛ��O�B��^�8�c��u�q�CI6F8C�	�n��S7�P��.��d#��C��(�,txtC� .q>�c��?k�:B�ɤ<VؘB�bCTR�`�DV�.B䉷&�<d�F&��{��k��_�B�	��Č���&U ,82�%P�B�.`���c`i�9E��,"FM^8C�I$>Zx*���[��x��mڤ^��B䉝Pcđ2KS�\�."���'s��B�	�G�2��P�T;/�X��u�\���B�I�,��t�5	�&��X��[��hB��3���s��Q#k��i1�-�a�T��dE3����N��cG��d^&�2�	��ā��I�N�m@�'���a��Ɣ�TG/ߥL)��D��1��hT��<Y"��?)� L�I�h�%CB�%�-�7�ԡ��O�PxB�A@X��se
܇bq������~�L�*P�0��Df?yp���d�R�*ׁ8�S��V%j�K�9p2�J&���C�Ɋ/�0+�F� X���q�$I/( ���!4���4�� AjY! �?	��)BE��P�*	�a{��AW Go��IFj�R5 (o9�����V�x�@`Q ��1Y�4��Ll?�U� `��J��)O��nՀ�`d�S��bSj���F(���/����A��� ܴ:�L�;��_<�F XW���$��e�3�$��B[UIjx�c��O�֬1�j�O�Ai5$�49�"���,���+�틩"9������-�*R)���B�d������
�!�$�|�P��%��,Ҍ�5��Đ�@P�(A�&��b��Z>�� 0��'�HI�bƵf�x��d�Z�8��[�6�b�	&y��9P�K;up�Tum9HޢPq�/��~��ҩh��]�F��c���&ϑE�I�O�[�N)��"ړ
r�����G� aV��'����L�U[+j3l���>p�"�	���\���1`1v�D�M�v^6��f�ƥt�#W
B��8[�%�X�@�� �}�q�ع6"������`D!§�y�	D�N�
��P���YrF���DK�$�ړ�,<O���i�2��%K�7'Yj��'�^��3̧�x�d��0=��Փgi��e�B��W	��B�0]Zq������4<��'f�������J�du؇ȓW�1kB��"�t��(�X��!��`�����OЬ���
�o$��ȓ9��=���\f|jyaD�/yY���tZ
��� �3W�\��Ų
�8-��/���JG6X�t0
s	�.;ö��ȓ2|D�YrDH�I��	�/�$M�`��	�u| �6��`g� �t� �
>n�y6g7D�H�ኳ`�hp6�M(���թ&�$��L+Ƭ����ȟbH[�ݟ|� e{��D���j�"OX�R��^+K�h|2��؅{���U+W{꽺t�O,س� �6���dR�	aG ����S��'���dP�Q)8� "i�8\c��լ�W�(d���A#P�����J��y��I�"�~uKa��E�X��ɟON�ȕK��P�8�֠R埠)���d(-sa.LzD��1D��;��2y�j��6)�.|��d�<����%Z�J8��Ί6��<�l>�',*�3pͨ$(D Y3�Y�x�v��ȓ/$�	p��`��!Q/^�o��0�PbS���6
ɑ��ύa�3����8F ˰]�j�0sgсP4����ci6�f߳(�Lw�A�$q��CJi�ӂ�K&u��RqBQ�����I&N��\@o0���jB�0�Q�-ᔉ����A�&[SE�
 %�%��%�G�=wej/}�A�6�B\�<�Z�St�lP�e�r�8�6	���@(�
�YXpy�k�m�!R��Qw�"|�0��x34 b"�P -�Z��>�yB�R��b��s�11(|�E+;25 +ǋ97�5C#�V�^n���*�������r<x��a�@]̍��*Ĭ\B�}��YNpa��ύG�`4��/]�| �$y䪆3J7��$���u�Wb��p=���r�&E��Xe~�"fmf�'�,iQ�`ݠL~�p�ǘ�%��y+�钗 � A�j�f��2��*La�2�"O�����ڈ[�l�2��J�$�s�'~���p��%.�ȭ�$/"9~�����Z������B�U-.��Ł+���*O���#U�Ti�a�4��T���K�6\�hA��\�a�O�n��0W�O�j��&Q������+Gd����'`�Ҵ�A� �0Ԁ�֫SF��7��h<~h�gF�Fx�ze�T� Tl��I�5������I`=6�ł�">A���FҢ�h���-$�
�p�a��J'iݤWV��W��!)������Q�<1�m��<	�Ä�x�(���u?a��*����@�L����G�v�O5Y1�M�UB:8����\�'�lec���%ܐ��G��>eMV�'H�4R��O d�� .���3�Ɂ
�����[�ޱ���:J���C$�[������9��Rk#+&iЏY/�����
�A���s�L7Rx�!A1�ӝaX��ڵ��!`���3/I
��I�m��) ��18���F�L�_!�� �L��$��!���k�gB��Y�V�Dv\qOQ>�:͉*T�\�K�����0H)D�\���@g9(�S�ʴ|pĐC��$D��Q��Xib�!����#��<Ɂ�%D�4Z��˔r��ivM�O;�@�'#D�x3�$�{����K4��t�T%D�����߷j�h��q��;T��iӄ D��I�O�"#׮�)�G��Kr�y��-D�����%�jŹRL�t��c�,D�� !��"t�\�p#�E��}�s6D���u
9��p�E�A���9D�L93
�r�LM���j̘HY�9D���"ӎt������	2	`#8D�d�$�ЫH^����J�6i�6���i6D���a�ր��5凼g��7D�0�F�#0fH��*2�py�/��/J!�DB����@����$6�A��-�	H!���N �$�)�QڒX4�X!!�I -��)xg�r#B%rĪ���!�D���[V+��#��� �Ȑ%=�!�ĉ!xk�܊"I��h������G��!���_j���u傆6-�ґ#��1�!�$��2޶%Xd*>N�9��>�!�DL�^�h!�3&�G�U�s#���!�䕍�D�AF�ڷS�fX³��mi!����(K��c��U�iqCf$"�!��ˢr��pV�9_z�EH�G�!�$\�d!b}!�����ge�~`	�'E�	#oÿn�0)�#�;T��E{�' ��d�vEhC�ȌVM^Y��'Z�FΎ�b0�1�a�A�0�:�*�'��!3�/m�@m;�-~9�'B�iΘ�q�~�ek��%)HE��'~�u���0,�D���"<R�'��A�`Z ��-S$ʇ�P|K�'�Dq2
�.}�l+���"
�Q
�'�tq��@�D��)C�bU���(�'[��"C]�}�Xh��#W��`�'����@�5�`8REKC�"��'���둢^8=���%�D2/��I�'�xa����$�4"���84���y�'/R��b)��e���5�&HX�'(��{T��W��B3ؓ/ਠ��'M��#�O���
��,�P(��'��p�Jʡ&J�}0�m�:	\ �;�'K��kA�ŶX{��f�z
�'|ll�G�D�\Z24�v�l���'���
UJ���d��s�b�P��'z��s��q��$c�\#_����
�'d@]�0ɍ�t]��a�|:��	�'�\���>,@8��F�?@nX�	�'f���i�P��$�p�X>j�	�'�����e����D��P�py:�'��m7�[�T�R�IɒS�tI��'�#���G���BoN�����'�,�`o��At~�:��
@���'�X���闢R1��+P��>F���b�'��,{�OTO�P��'4:�R��'}�m�e.*Q�Q3�kR�,��}
�'� �����
>Rt��f���&]���	�'3��!��%��@�������	�'��ݸ�,ۇ��u��Ȍ��	�'91���P*|ZؕF��P��p	�'7�-�$fʽnZHӤ�������	��� 0\���J�z݀ �#��
)�@�і"O�R4��.Z�}��O��t��"O�D�G#_s���a,§ �z@i�"O5{c� �0IBǌ�1��:b"O��a��3"0�#��ʸ*��"O�eswʣ_l��5jN4|�>t�T"O&2� I+���S�J؆;� �p�"O�zDb�hB�@3��7�2�c"O� �i����A��IW�xF���"O�2�� ;��
2�D6t@�r"O�����@Lx%Ӡ,�uvJL��"OL8i��M''v�]�q�ՈaR\���"O��S�(� ��+GIN�a�"O���t���l�Pe��1gO�"O�mG�@I���r���b��Y�C"O����i�����+F%��lx$y;1"O��z��أ/�	xB�D�ޘ���"O�Ȱ5)�m�̅ ��>l$,��"Oz��R���Q��ѱ��)<B,��"O��p�27"l�����=N(y�"O�u`w�Ⱦe\P��LDvV���5"O���b/0��	�ɌP1�̐B"Op���Y$�zL�7G�#�<=�eǻ)�Mrq�TX���0��~�����#,��Q���+LO��mQ�T� qb�'l�8��c��fi�ș�L�4q�0@
�'+� ��@ڃf{f`-�HIؓ�����BQ��L�5-�ʊ��<z�S�mT���\����.w!�Z�АC��W�J�`��ڎx)lx���86��I�h=���O&��ōc�R����[b��(O��PB���G]<��$��zP��S�O��&��E�NG����͡ ���0l�~Z�k�EJ���y�˃rD�u�6��2&���rb_�IU��JGC��H�!��F�4�3�˭Yj)xA�LA�'[`5(���JM$�I���#K6�2���7|y����,~T�C�	�2FN (��h0��T���yäU��6ʓBO\%��L��Aql�EM��c���7�� sq�74�h;#��
9�4Ys�B4l�F؁�]�2�d��C�S4$-�E���5PTհ��vo��ڣ�� n����$ܻ5�n��#့�~�L
�KY�a����"�d�*g'�&�y�A8p��m�D
���p�&❅θ'_�hю§~�?@(	��$ ��E(&�V��!5D��b%�μ}��h�c����*X��F5D��DhNtznZ������..D��'�V����_2f�Deb!)D�(��J	�+�x8�!�_DT-�4B�	�N	~��$�p�b�"M��L�B�I�p�b}s�B��~�|iJb"�l**C�I�awjq���*��Y	P�5=@C��)A}h���I6n��Q� HZ�|w�C��	>Q��Jմ_��U#'����C䉬<E��ڴ��)Z�8�t.�ľC�	w_蝪2(;`L��˱lӈ��B�I
���a��!�����וpC�ɘG2�)V���D�X�4kӁU��B�	��!bC/]�;����5�Ε :�B�	Nk̸�f�&x�N�U�X�f��B�I)Ɩ��EO<1%^<cP�#1�pB�	�f%��5g���AE�UZ�|B�I PG�e�m�f5�UjҨW�B��C�ɠ}������7���s+ϲf �C�I=<�X�fB�2iP��A��ALB�ɶw�BL�C>E_�Xu�Vp|ZB�ɣ#���)j�Z�:���gW>B�	X= Qa(�&����֩�=`��C�)� h�F�	B�����	ӠL3"O�Ub%ڦD^��[�ɛ�:�
$�'a�]r1�J
P\Pd	1s��3�Ҫl���O��!'�%հ<!�A�;c`��l �(�d�r�Jm�'s��1SK_�f剕[ 8�1��[�0�p-	2~{��C�^/���h���c��`o�	�������c��CC-�!]��ɡ1���GŘ�hG1�H���hT� �$���R�B���"ON+�fñ<>�!�͚`�����O���!�n�,8#g���I��ּAPf���Y�g�S��%@s�߂��͛pF4�O�ų���rnś� O�U�$q��7N�9R���>:��	3v�����P�,�ax���)2ܘ��'���F�:��ĬL(�hO�1��ʍ5 ��!Z�౟�!�N�ThHh��aD�z����U�������E�x!�J;A8�ǯ�mb0�Q�B=k2�@~�r��FR�g+���#�����7�� +�;anG�1��x���P�LS	�'�l̈���S8fH#㔦0�`-��']0���C���(��e��|�T�,lz������� C�<m��:`G˟90h)�W�:�Ol=��i�	:��hƪ�X)��KV�z������d��	�����e��~�axr�T7�����(��bb���hO�MU��;�hp!Y��n�(k�H��c�\Y���Y�}���^
�Px¯�Vrx ���z���j��?i��b����'���n�>�━X5$d�4��L�7���bqGAy�<iV�1{�z2��C�qKr�p~�$���=��'J&�Hb��s�6i�� @�\8z�9�w�!� I�N ��bڨ�D� F�b��ȓK��pJ��	�@?H���`���p���Q��ń�fm�����%wZj��v:����C#��Q2��*m>�<��q��#	�1�6A�a<@'�e�ȓ]�ޅ���N�r��D�0b��|�ȓ[�	�W���k2�1��ǭ�D��ȓ8�����>"�ܸ���]��Іȓ,�l�4���\����GJ�]�ȓIv����¹3l�1��˗?0��ȓz ��II�qZ��-Z��`���o�)Y��T��\�K���-�ń�]X����֩�Z5��1K���ȓ>��)C�ձ],�i�cΦ�@��q���Bo\�"Z���vg^8*��)�ȓ%��@�B�4|�aBP��;>Q�X�ȓ#~`��f��pA��yn6���]��L� ���$<���=���ȓ8:���mE&�,@&��uYx4��g:�3��ؗ7���_�sS�B�	���\��<D�>�ⵀзMԖ��D��$zj��ÌB�@��r�K=(0��2m�/�ybKY-������-JF��㯝��On!�� ��V�?Q�H\�RiD)07��&z�6<�A"D���w�T��R��#��i�Xݡ@@�OL����Ő:���N�"~:��M+��T��C��ew�0 Q����yRE>?�^u����cL<�`�R����T,�y`q(��˰<9�!TY6VI�"�� eR�b�/�Sx��J�o���r"�űa)�*b�\�jN�4���^B�	�Fi���1��3y����~}B�=J�;�|$���p�'KzZ��%�1��l�2��=xT�ȓ%���@_�1�$pc�������(��Uy��6e��D����@M��
�`HB獘�pN�m:E�/D��+�'ȹ@\�y�&�.Q~z`����<a'͘-�Pѹ!O��0<�7#^>[R��E�F�r��x0�Px��h`�M~?��3!�B	�hBD��4���e��fX!���HB-q� �:����%HB�R5D|�)&d\��0��O>h�[�i'XSTl�K[�m$~} �'*x\Pr��$;� �{�H�&YO�Dk�',,�	�)ސ@�>��O�>��F��6�v}b�$	U<~u��c D�8�I-4�6���!�.���RR ?}�où#VB1;�$�~�� �]ѲʏzB�P�2�ֲG�p���'�����H�Dy�­@�w�`��6mƧ?1Ѐ�t�W<�A��?1Ǧ����_̼,�gN�Q�'���fe�	\�q�H�04b�i� �E�R�~�j�YW"OvDk�e��\^�������'fD9Y5_�|�fΞ�qOQ>��/\�6¤�����Ppx�0Ƌ<D���Y5+�!� ��`�D�ӧ���yrf�"�C��X6b�돯�y�*��sY��!�iW\a68k�a�/�yb�_t[Б{�O_RwK\1+&��-%ȸ�p`�2XC$UJW��\j|4��=4��	g+G5=<��4I�kN8P�ȓC:d(��:5���c� 7�}��}~zԐ	Z�Y�"��T!�"'��P�ȓk�qj'�eC�=��
W�#�v���r�^�Ŏ��]�|�̍�y�<��ȓq� ���O+]_.y���E�6&��M[@tSG�ɵ'�4�(�'4	��P��P���	/T<%��^;d��]������O�@.�$Xg�V�&ć�(:N!�lK�UѦ�¥+�L�X���m��X�Y�f��-�������ȓ2ج��O�\���"n��:'����ti�@'&^F�K%�Z&WƔu�ȓ!T�1���^8Pk�b�>M��ȓ,{*9zTL��"ܬ9s�"O;MoB�ȓ~�@ة�F�|�%�TNحr��=�ȓAI�`ˠ.��n�|(�Β�.Y�ȓO�����>k�vh�OC
=�*,��,S�qy���UeЄ**Q��P��.l\���m�69�
� �%j�<�7B��,"��p��s�n�x��Z_�<ᅤܚz7 |�A���H]�<�W��2�̙3�k��^brt��g^�<ɗ
�qֹ�V��u�Ԥ�4&C^�<�#�:C%�0��N_;a�:���[�<��/]�8M�+�3!?�x�Č�S�<�+U2��	�Q ��4�SfMN�<9��W�hVT�"!$ظ`�)�Q`E�<	R�H�`Q"�1�o��)�j���F�<�`������֗^;�b�Jd�<ɢ���}��Ds�G6%+,��e��g�<�(	1^N�x�7��,9*��Mb�<�U��q�I��(�4*O��I \�<Y���?;9���1fQ���]�<�f��(D���Q�k'`��%g�]�<q�	�#k�p�IQ�*}u!NCF�<������,��OC q�V�0�j�C�<fnV4v��c,��n�t�"{�<��X�@M�E�&����1��%�{�<	b	S&f�(34�[�x�F�q�<q��V�l�"m�a��|����n�<��!M�%>x�׋��Y�H�p`L}�<��B(�V)k��P�O�F��7)H{�<Q�E?�0��`�.}�$T[���u�<A��	{�}��I��qBQـG~�<AU�фq�@Q�!L$f�X�eo�m�<Q"G;W��h3��v����$�j���z$o��z�~\�e�>ĭ���eK��eM�%�鸢
�?Y�D	�[�V8Pa�++��>-%>�0�c�"@��k��)!Z�с��E�;Te#Dʸ6�J���Z�x\���@/�N�K�ώ+C#�q���/@�q�<��:$"['A�*I��OZ�9:�曒1B��a�Q+k����#cn�-3�X�6���V`I��0|Z3H�v96��5��e ��+��15�V\i�C�^r�\Y�H:���'p��I�)s!��P����p��A�	s!�+���ɑ(5�� �E�ӌAQ��X�e��
�8Y��>���'��vm�*1��I�p]>5+�!	�Uޢ8����n�U�G�by� G���sD�_1���TVXKf'8z�ܓ�
�*/J��H%A�uybo�`��(�çb0H삥H��Fd�� @����}!.O�!ã@�jJ���O ���PY��N�ѤF&>)�Qٚ'Ēѳ��ĨLh`�R�"~��9��Z��ʋIy�Pj����x^�4��h� uڬ��,Oa����R�&q�f�ͮ$������KY�� �NRjW�	�E^X��}r�~eE�?i�@I�RB�a�n�QWF���Q���0������,f��q���b3��95�d�	9��%p��Sꌝ�Ac��g?�O( � щV�
��K�*�L��R��T��Oj��$�B�)]��$>���˧i]*��@m��\��&oKV����ƅ���2�(hӴ@iu�H>��8墵��g�A���??a1։X�$��J>E���Ǽ���St���3��s��� �y���EFX<�!�|��iՒ?�@��W��e1H�رl�Q[T)��,��}�d��h�ᓋbKj1�t��m�H<���m�� ����h3F�A�l�U>5h\w%J?p�f��*3\,h	7G&�)�O���"��O2t�`D� ��#|���(Y����.�s����2��8BI45K*�	�G�'��>�ɱf]�س$�J�L�*� ��h�bC��r'гw�(
� �0�"Q�(C�	{�\�I� ۭ�8��n��5C�C䉑D��=a'�OYGT@8�%�*bAxC�	7,�`�ʢ��+>ׂ`�ҡ#zC�IUL�kQ��]�r`�F��]��B�	�m.I��4hM>hs A���B��:-h�m3h��t��s���N��C䉬 &՛�	Y�D!�Bh�,)��C�	6��ͩ���U9�(�@��cĚC�I�d"�p+%E�:0������ٜx�jC䉐Z�}
� �(VDxx"e���w{ C�	*!�x)0E�!xz��Rlю6��B�	�O����Bn�.NbX��M;F�B�1�-Q��/48x[W�]>e�RB�ɑ2r 8�`�^�C;R�أ�A��tC�	�v����cҠ �ri2����e�FC䉜!���P��W�q���1��$�$C���vF�)9�$%Iʖ!0�B�ɷ4M@(@�>���NaI�B�	�X��g�^Aܭ13�K�g��B�ɢ`t���=}��d>q�B��]8�2�A�]�Iqf�5HB��!b<h壄�ʎ%�as��H��dC�I�߬k�/��	�Z��1��	��C�əIR���7k�i� �qN#$M�B�	1^tF䛓��R<��)�n�@�C�	�I-�}`aB׈O�`���ӌS�B�ɴn�p�4aA�ZfH����%��B䉾`E�}�fd�0	���f�W�apC��	R,��C,`9[�C��C��x�xf�7������#��B�	�Sp���)T)<�B7<D�B�	���h���e����I�o�B䉪h}@�A�&c0`��Ӏ�("�lB䉐~��ISc��K���O�>[W�C�I�S�64eI܂k�.�0�MH-�C�I�tw�0P�&�=|[2<�q��	��C�I�4p��
�k�� �,h0C/
"HC䉰(&�Q�E�/(O ���
5�C�u��P%��'i�4��a�*Q8�C��-Lp-b�6-� ���R�wEFB��?w`F��p��=���S�a��x�B�'Gh�%!� ��a�DD;LΤB�I�"�*�2�-{��9�Ӹ��B�I�h�V�:r�ٛ|T�#��C�	%nV��сL#��I2�eݱ-w�B�)� �E�g�)��3�X�+Ϙ*�"Oƈi�;�p���ښ2�ʬ��"O��[΅�
pR��Y6 �,���"O$՚��i^
�Qa�Y�{h���"O\B�S��TN� =�=�P"O
�s��� �D\0�J�Mx��0"O� ��+�$�By����uk�m�"O�-c��:o����hJ����"O�5Ce*�h`�A���Ma��L�"O�傐A��9W��9�MT0R�Z�"O��G��+�FMN�(�˦"OHA{B���zMꜣA��A�FPxa"OP�PcLڛ5�#:0����"O8�G�b3@�V��t��y�"O�t�d���x�J�x�""Of-Hg%N/�{�I�zإ �"O���T��= 7,�����e��]��"Ob٩dM:�VQrt+�:%����"O�ȱ��U�����
Z��U�g"OL��F[o⊴�#��(8c"O=q1o���V�(U)]V�p���"O
	Q�Ǌ
�\X��B�7��d+"O^$2�!���2�Zև
$g0,��"O\��!��B9Bh�D�΅l=j�5"O���B��#`��e� ˃�X
g"OByS��4,��"�.��ȁt"O`�c�_zm,�(SҺr�JQ:�"Ot��vI�W~de�2dO�*�ы�"O0
 d������"���gҴ$#�"Ot(�q��Yr�!�wkz�8az�"O��@��þ0�x���TP����R"O�s$�F�2~R��%ƈls�\A"Ov������`�Y� ZT�d"OH�)��؃<
��Á;?A����"O�`i񅃞c�f)z"�8 0Ѳ"O��"��	#��C��G	�z!"O�!Aˑ6�<Tp���2g�x0i�"O�!аF� b���U��u��x
P"O�I7�N�"[n��P�I����٤"O� �v
O�*_.�An�y,(0G"O����
���[�H�k4���"O �׋Ё"�V�S�e�:V��"OH�(���<gv9����E~�Q�"O��1B��$:_���T��֔Ɂ�"O��Jƪ154E�'�x�La�"O �Ia�֣d�X��t,��H2Tk�"O�l���G}��m���V/K@�Z�"O�x��D��u�Ë˄$=���7"O�Q��t�=2��I .$Hq�"O"1f�:}���C-p�2aG��y�l<3����(�I��1 p�B1�y���uJn� c�"E��T��!�y�/R��`�
͈::��o�yBH����$�D�K�6��\X��S�Py���y�@�X7i�+@��
`�G�<���$� 487�X�o�B�jtF�~�<�$C5FU�}Yg"�;F/؂���{�<GH�"2Ա�e���_�H���(n�<q�-�Y<4D�W�@m(���q�<aEEE���)�(дUP��	��Ro�<yঋ0��l��.ӧ�Bd��k�<�d��}n
�:���N�*pGf�h�<�R�G	k������:��!�oc�<!��{�.�H�nW�p�ȤP`��Z�<� �$(a��S
�@
�/�8O �"O�a�̕�%�����7�*e��"O��3b��X�����$W��X6"O�p2�FВ��E�#O�R�xx4"O�;֬�&}�>(�Ű|���1"OJa��Έ��d�q�����D�v"Oh��ZqFN�`Q�:S̉r"O�S!�5x���Ӷ�؆X;��83"On�{�'Z]�I�G�G�12Xɱ7"O\\�&�%!��q9s@��I0J9Yr"O���*��sJ�PeO4!I��v"OT���O�$n�z�s�ϧUK��"O<}hV��^l>i���[`��"O*5�`Z�>�(�	�	��~[(���"O�$���=4�^�!S�_5EY͡U"O�����O�+����h�}JƘ3�"O�T�$�]+[�k���*iC 1�"Oj`S���	qgz�c��հGAN��"OB��2ɘb�u��%9�Q��"OȽ �υ�w\�ٸ�
��@:I��"O�,��[�3ղ��P��
3n<��"O�\I#���n��`��;u"( "O��	�d�	X�=��ėO'j��7"O$��B?XuC�`yD�E��"O��k�"<i]�t�����,-��"O�����8c\�C��Μ���e"O���a,�= -0	A��.*��Kr"O�[bn��x���ĄAX̡�"O����>Q���8I�A�T�cq"OLC���Q�NтThҖL�`��A"O����OX���#1�Ȳ|�>uP"O.�jS�G\h,�A��,�`��f"OtP�Df�V��Pp
A8lW.,Re"OX�iPm�6�иz�ȏ h*��;�"O(VZ)Y��UH5�D�xL�`��o�<���y� �C�'I�~w�Pfe�l�<�1��*L_����ƒ�q�HݩiRs�<�ؖ.�B\AP � uXf���Ao�<��7Rv�{e6 ��-�Eb�<�"a8S��A�L`��@t(a�<�#A�C�2��(�r���DFZ�<Ts�����U�sC���7È[�<��!�c��)B�
Me
���V�<i��3��%*a�D��e�R�?)�C�	!�0����n�Y�G琐�C�ɿ)BN-����<9Jd� ��
T<�C�	���C��P$yBk�>��C�	v��	�D��J������C�	�nX0��E���f��#��/|n|C�I�%���C�?h�(��򅂝�8C䉇��E;��V�Z��0 ��@���C��q;��"3C4qwI9��J�Z�C�	�	��+bh(&�`�wިB��0;�\��#��p�L !�ʅ�Dd�B�I�H��X"$�:Yf��"�!#A�B䉇v��,�$� �e��4�3ǆ��]v	�u�#�ATN�~�j���Bp[ԇYG�s���?g����/��)�Q���.�@��TJǜL�t]�ȓ����Y2^B����N���ȓ �L8凹���:��:IL���c^����6������y�<�ȓm$2( s�_6�Z��Ro�r�*H��,\2�/I�M꼢�/�X��S�? m��Ɇ�e[�ҶJ�n���4"O�Ai։�"b�ʀ�t`�^mvq�"O���fhB�7>�ɶo�AY`P�"Ol�(�!��]�Q�.كY�D��@"OؑP�NT}Tά��<9��袵"O�Ic��G�&f��9QG-l�\�H�"Ol���ϊ~��� ��۷��!r�"O�z��I9_�4p�4ǖ$/<,T"O�=1�bA6�y�C��\�� 8�"O���sǟS��=yF
D�Z�=z�"O�tZc(J(?�yf�Ø� \b"O4(y�$�3!�}J�Q�p�I��"Or����2A	,�� ,ΰ`B]Ѵ"O4���Q�P��D�m��a��(D�4��$U�мR��	H���
 %D�4�@`2���"��2a:��!�%D�d��/>0@)���=��}��$-D����7�I�d�_�p�a�#+D����&H���8�6j-f���q�=D�$)���!R�P#E�
�,ԈwB:D�lӖ��'6o`pv��92j�R7�9D� �`k�Z�,j���sz%pF�=D��ʧ!�9�,���*R�j��亖,<D�d���   �