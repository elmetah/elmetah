MPQ    ŉ    h�  h                                                                                 	J=� 	���S&�r�?v����GY��>�u5Z�&n��J��R��	�/��f\�ل�k� ��[M7G�cshg���J����Wѕv�o���H�f��>��'�+��g*i;C�� ��Քr�G�>u'M�3�F�ŷ��9`u�r1�-%'j��(�� �N��t��	��8h��"d����� X� �婻������+	�Z�Q����'y�Bȭ�X|�TX��>^�@����b'7�i����ƃ��u�{��e��9@-�!�@�i�<(����eyÁ��l�墆v�02�;(a:��16�Į6�3�,��!�җL����Z��m^�P�`�b����{�Ms�kv����.�kb�գ�(�a���Y�2{�6�N��
��O9na0��:ƏN��q�c?� �-o�����ۜE�r��7B:q>^v�/%+/�C)�7{�j��'�b����Q%[b��9G�1�0-S��L&E������2��4�g��I��\�w��X�6�Gb:�D�~k����$[o�N�}���A��*�SᵵP���N�6�D��3����?�	�<+{H���,�/����l��D�p?z��!|�v��0���(4�}�dA�W���,�L��&�kղ���is+*��)��B�=�����A��H+��
�"![��(��`�j�9�_X��=�X�m�_�nU����UN�ͽ	so1�M�F���;H뭂X9�q�P��e
2�x>|t*'�?���h<�2��C/��� �j�Xo��t?7ڱ���F��=�jd�;���ڷ��@�-�*�i�GX4H���x�Z�1�D���}��=��)PB;L�3����ޙj�>�b�J�n�#�,�jB�n�q�R��[�w+�*F�<g|�k����Z�x[�}$��SrR�k����]:�T{~��+z�M9(N8$0�1���Jq:*i�ԫ���^��w#�`IM8_��ϟ1��ˀ�7o��YM����Uٻ�����JdC��
ӧ5"=�S����D��O b5���ke�)I���A�"c�S�6P�\�s�!����v��w�G�Y�R�>�h�3EW}�е�p-�z���y�"~��^_5��+���c7/�����}��U�tC�,�!Ys�"8�;�����̵�,x5�e)nO��m1!S��.�@$�/s�r�Zi��C�?���
6�Y^�	���k;�����g��<���Q�~�3��q�jh��~�-t�Ѩyo\#'�Ƚ	.���T���qte+���<�'� ���;�!�R�	���1y���u�M���넛�D��N����[����l��A�z�؞�,�^G[%��h*��B#%t����qHh�v_V=�����eW�_���e��H֕c���p��8�"MY�`��\J'!�\+����)\P��Ֆ�8\R{ځ��b'u�JmT�_�[L>��$"÷�o�$����/HU�5�ʾC!m!�.��ۍÞ��%1�s8=�4L����D�\iy�CǛza)n��**��tYLl��p���4)�����$�tq��7���<c�{Te�E��`Zw�K�_�E9X%c�
Z����Y��%���6{��Y1��Q!s偽F{�Bڒ1�"�χ+��&� i�f���E�x�!g�^d�^�y=�f���v2��)n6XY�C;�Ms��:Պ�
�̈5���S*{1u)ykQKX��IZ�ډƠ	�����]�_ l�A曉ԕ!�Pmw�?�ma�?���m��]�
�F�^��9�9�K �Á� ���UJ�+ԝ;	�9�ۓ#����~�QS�7}���{7"#0#3��m�I(@�t�u(����-���5�l@�&q\Ͱ���c M#��+��|l��,����i�ـ�k�U�e�����PnW��,�?�gį�MZ} ��A��M�=��1g�,˺��������[ÖO^��b]M�/p��lܸ�?f����o�n����̦�`=bT������/3ԙ�=�ɴ�^\5����$��%�4���?)�E�8J��g�}(JN��:�ө�5�o�HLl�D���@ʑ�뛉��S�s`E~�w�:���ik=r��W��	5�4%�/���"���d��u�����j�\���Up��sz̫G���� ����m��2�i�7qaH�҃��V��*��A7�U߸���yi�yfDp�M��@ we���#M;p��^#�B$�5~ɿ�-���K_�ރ���W��;H���r�c��{A�U�9�k�[���.�TT�f�&}���o�MXQ˭��p&`֖�OizC�,s<%g2�+%���V�L��#�T[�D#���п��ֿ�;w��ݡ��3\v��Jt�'����r�^�RG��)8	�$9�8ـ['Ǥ��E�N��kf�����/�3.KS��wŗ� 3Q{��1�!�K�(���7Y��h��W���/��e��C����ug�ϸ!��*�4�]��,|�]f��ֳOwkڿ��0�l�����o����m�tM���|���B�!�9���m��ɻ���=�r�����?$�W�P@��)��lLě��pך�^5�W���`O*��[ ���.эOܫ�j���0E+ƭX{�;TG��403�f�"�߈���Pd�k�J��'y��
��Ϛ�m����Dl�R�������v�fр'�z��~��3Teǵ��M@���}��0�g,"�Z�.1�y��q��^�WQ�f1�M"{N�Q�&��	�����!�;���;��4�d�� �����]�����YTR�����?=Gq[�E^�xXa�D˄�IAEs0s�Q؄�I�y5k*V^>_$��cӹ)�H�ǈ	�F�Ga�ȳ���p_�6_|�9�5K�זY*Y��f�c��33K�9kV����>��~#l�w��K:��)�!g~�C�����T��鱟�xW���9mH���^H�a<7�������zƀ�uAyP>��V�^��pC<�X�~8�:Q����#L�j��NV.��r��Q��M���ɡ�w��;/���6�;-� ���8�hm�������\�?���	��<��5��h�i*�}'�R���z����e�|پG��>�_��l��/�N6���O5���Q�-�|�������,�E,s7�Y2`_K)ಞ[������M������U���hʹAd4pӇ�W�Bީ6����qv�f�ZWCG�	�'�C5���sÔT�:�Z�@�{�<�`��R�7BY�p�?ƞ�'u>x��+%��-��@�$�<�۫��T��� �6�m��r�v��b2hn�a5D'�zv����0;�,+����9�)q@��A�mY�A��bJ���n�M�MIkQ���#��Rz~��pd���a��SY>�	{��N	T
�O�9iH;�).�	�(q�,���̀�^o߲�f�4E�`�G)L:,[�v��h%�fjC�@{1!����]_��8n�[>?9b��1N� S�Ȑ&��~�~S�[���{=g�Q'I�0���Q�Xk��G�)c��Ry~ͿV��-�N���eZ��R�SG%��8?�I_�ğk^3_�ߟ�	f��+�M����ʓV����~Z?5��!���b�D0�)�cm}`�T��'�mٚ��&"4$�-���+e<~��t��=����+b�cL1�2��.��c0��&*�4T_f�_�'��s�̌ڥ;I���0}U釩͸�o�a*��K�V?���2c�L>S�a�e�>x9Xt��R������J.��2���Aj4�j��ߩ75|o�\��X�>dZ����Z���-z��dQ�G�)��i�֓����G���k۸$=�.P=	�LT�T�A��3���'�Ie��g�Bu'�q�����2�éEԹ<�eɸFE���zc}���>r���]��-{�9j������(Iu�$�A���{cq"�\i�*�|��^�BN��IHe��깡��P�:�rj���ۓ�^�ݳ�	UԳ���J&�%5���Sݹ��,Ov�w� ]���'!k +I�"AU�5c�+j6����@!�J��Lqw�@�Y7��	R�hd�-W��ɵ\��-��T�W�h"9F\^z0��HG+��cr5�x�Q�x*a԰�}C�;!tYg��;���)���g1��'g/����OxI�1<$ĩ�@�l�/���w�d�񧞪��Z�6�$�ً���;��ᝁJ�����O:>���(����x�EB��Γ��0+ѣRvo�R�'JO	I��Q*������Ue�Ց�7��]҄�<U���-۵aW�}u�ൈ��F���󍟵��<��D3��G��|C3z1֒�'��G����#
�]v�tK(�L�(߱�'=�b���WD[����G樆8��d.�����s2SM�,3`��m\�M�ͩ�����5��hd�2��R������k�xt��=�z�tL������q��ыP������/��Q�� W�B.m��ۋ�����%���88��4\󊣩g΁w%yq �U>�n�e*s�YG߱��sw��F����"$y�Q�����տC� fEe�,
�6Z26ᖚ�E��c�=U�GR7��F�|.�!�{CM�YL�Q|$�s�_?F�` ��1��[��~d��.i��~�@�3x}��g�Y��=���xl�2|�n�sԣ�;��Ms�aA�%E������n:S�Sm1)|�)�ZK3e����$�	��i�2._��.A��\�PH8?3��AM��/��\�
�F������JWK;�z�^YQ��Q��tz+��	1�t�z#��I�Y�[�����2#(%7�#.>Kl���(\G�)uÜ��֎>�n��'̡At��+�>VP#�w�����w�V��� A$��W����r�0|B�7g�N�?��GWW���T�Ƅ�Vo �RQ�|�`M�����rg�-E������ɵ�cT�q�_�N��]�#Zp۩slf���ƹ��� �ӻ��~b�d���/�+i�����ρa\��f��}6ǺA�%�$ݝ��?�>����΂9/}�r���r���!�59
�HGZ�DMƲ�����[��#3s�NCS~��:���if�V�n����$�U4��ܰ�tg� ;���'uR�je˞�/[oU��?s�«�jS�f: �A\<�ۋ�,4i�hCa�����VK�I��A2�)�R�4�y�`�yD����wN�	նd�M6U�﹧�Bߧ�~���-;��K:�˃( ����?�6��2"�cXqnA�G�9k��[�zw.��;����E�bm�o^s+Q���Y`�&�O�Y��e%bx��`0saE�V�n��#��U[��A�[��к��1�;2�����37\��v�K�ᐢ��X~G�Ƀ)S�v��� 8�+'Qr��F��D�@��;.f����q���[�3�2���/��F2O�8�,n��/���һ����(՚�Mq���g�
ʈ��Me����(]�gI�]"Z�ѻ�w��i�|#{3�ֵZ���J�lJ�BmET���s|G����U��T����El㤣n�(!r\i���e?���I=�D`l��7��,�Ն�5*L�O�:�����:��ʃ������E��{Xv��T^�}��N"�����ZB�g9͎FoIJ5{ny��"��	�U���ɘ/D����:�K��[vp�a��'L�fz�%���MeB�(Yݻ���O�0r\,}����y���q*J;�2;fl��"Q����dJ��,ŉVm�!G�f"��0T��c]���6Rbp�ɟ�=¡�[��䓳���ߵ�zg��Ms���Q���I��kA(>�j���)�	������a�+��>��p:�_O͇��"5ש��d^* f���J��3&��k���x"�yz~���DK���)8:C!���C����G��dk���j-�Wc4(9�l��v�Hm��7�'���u���͏ΐ^>��'�ً��aCwbҥ]��5	y�	S�#���	B�ɓ�ø������>���$�w�h�/��j-�@���. ���s�smn�n��.�����ڏ�Q��{�q	��C�e�s}��a���v�H�E� �����ѹ�e�Z��S�6�����O�4r? �����|�W���z����EǮ\�T�,_��B�Y�n<�����{�ZE4Us�6h�3�d�ϼ�B�;�6�>���Pˠ`枡}�Z�Tn��'/(g߸����*�TN���5R3����(�`��b�7�h��+��ƹM�u�J��p�X��-,�2@��a<���lڠ���E���:��bv���2�a0����\�:�2�Kc,��#�����dg0����mTK��a�b��΁�Miąk,�ǣ^��3�u��5,Ń��Oa��Y��&{��rNU�
�9dO�ׄ�U��1Mqm���$xo�a��$E�2��:6:��v�%!��C�-:{lC�ݵ\|�X��쓪s[��9}l1�U`S���&�Q�<Sk�ú�;�gV�sI��a�m?rXFP�G�a��zHVt�Y���	�
N�������ZS�G赆�j�D]���(3Q���	�x{+�@d�(a��e�����^��f�?�!�Iy�݈w0��_��=}�E��_×����&=�ը�z�\�_+����_`à8u�i?�d5��~�'� �S�"@֞���}A�/9V_�
���������UU�$#��k�U�Iͳ�2o��¼���qV	�x-�'����e@k
x4�,t����J��Mȹ(H����!�j�g��j�7�fg�;���s��d�< �����AW�-뷥_��G?^��)�֮�W�P#-��8[���=)�P8*uL_��))���בX$�$[����oB `q�
Egp���`��<]�B�!攧���v}r�=`1r�p2��w]0TR{Յ&�)�1��(D��$��qh`q="�i���W�G^0Y�2IC�s�E�s���"�U���{��}�<�Nh�U����s�JJ�(~�@g:5XlS���g7���� X�K�ti�k۠pI�gAнc�#G6ƞ �!��c�,�lwiY>YR2�섅�h?Y�W�6��s�-�L�ϲ��"��C^�K�Ǧ+�S	c�!n���sn�`&CMj�!�_N�T;չcd���ͦ�"ve��O3�1W��$�f@�7/�4���}N_�X�����L16��Q��8u��;���8��H%��~��\Z�C�/�g#^ <��	���c	ў�o'^	d�	��}<��_ea��2#�H5`�?�;W��E�ې��Q=vu-�����Q]V�H� �rɿ��rB7����z��~�"vBG�����x�kt|!��'ty���="붵��W�v�qS��������뮞7MF �`�1\ ����3��b �g��dÖmR=���(%�S�����
�L4f���O��S��~s��/�N��(�8a�m���_0��v%g��83qZ4����d|���y���0;n+��*�@YBr'�&f����Ƒ��$����gƏcx�pe��e�lZ��ږ��1E/�Vc����� ���&wW�vi5{���YglEQ�R-s�]QF�R7{�1�� �=򧇜��i�l���xXS�g.�ŔX�=�ĉ��
<27n�n:X�Oh�;�s�0�����|p�<8wS�HC1D6)oj1Kd���ڿ��	�*��\&`_�K�Ajԋ�$P#��?T�u�����J|�
�kF���vd)��Kv���PB�ya���+J�d	)~��-#��Z�����P��-���7�D�Y��c�7(�.���u^j�����ɵ^��w
\�Pͦ�H���#����:T~�r�����Z��f��v���}��r'���8��^�W�����%�Cs� ��R��MO��ݧgPO��DB^�����u��L�P���]���p�Vel�T۵�ֹ
X?��dӖ�t�X��b�I����/�X�Y���;\+�hس*x���b%Ht=��V&?��j���Ν�}�t��ʕ�u�5��1HBh?D��#�w{��f���~�)F�~F�:3��iaϥ(g�ͥP�?�4|���"<�;��H�u��v�j ZA�J�cUf��s�i����-b� �����h�AFki�]a>UO�Ĩ�V<���4�A-�Y�n���2y���9���~�w�Y�Q6�M1Z�L�B��~��-��(K9Ƀc�*���1�1��ac,�AZ�9��y[g2.:uW�?=<ʷ�g�o�BQ���Y`�ւO߰­bx�%]�+ǻU!!V��:�#h��[�Խ�^�еF�̌@�;�Z�.dC�C�3b�@��]x��܌��IGK��)ne��8�ª'=�{pu���]�j��򥭾.����m>��·�3�	$�g��A�Ѥ�o�j�Jp+�M������M
��&w���dgs�\�,��'�*r��ڻ��6]��,����w!	4�76�N ȵ�2��%9a���m�S�����|�%���o��>���s�c$�r��y��[�?�|N��qX�_V�lB+�謶���85��ԭ��O�◢�Gi�"e��E�����J2�Ea'bXq|T���ê�������I�BB掁��J�&�y�	wI���lY�� Db���������^��\�N'�ܘzsz����e�t���j��� �0'�,�,i���syѐwq���E�f��;"��Q��ￅ!�b���q/��&�������.M�]�L�u�YRf`��Ld==��[~库��Q�zx	���˶s�TuQ��I}�k�Kb>�Ѐ���)���>�_���a����-p��_�>��o�(5�z�L�D*Ϣ�f��"�3'nk�`m�&��t���-CbK���)S�!]W<C��@�3ҊӤ�M$�Ů7W�g9������hHH�y7����o�p�:�+z��p>����T����C��_���ٸ0��d*6#���#z�D���Ő�H�~���Eٿ��wTk�/�/3H��1^A �Gd�@�m	��ۜ^���Jo��{������F@�c�}]�i���n��E��V�����4�w�h�Ǝ�҂�����=O뷅�w����|y����3N�K��Eb
��O�5_fe�/���4ĝ��/��S��$yUch���d������QZ�,�,�{oF��g�Z����`�'�,��s�����T�� �6���� ��˒W7��Ê��Կvu4�3�\�5˓�*-���@���<9pƫ'�y��03�,�ӣvr�v2��2�3Ua+���0a����ƙf�,!!��chb��}��+ݭmOܣ��b�Y��鴒M�Z�kc#����|�pL�ƃYla#�uY4wo{y	�N�A�
��m9_v���=�6q+p�I���aoU�͜�lE�$B��k :���v�8%�53C��#{����P�Z�S����[��`9�K1DLS��H&�e7��G�Ki��jg�I�����L�X!G�Q��o��>\��N+=��[��u%S����!�n�?{�U@3��%�j	\�+�S�c�9� �j��ǫ�Uo�?���!���Xw�0��|�?�}����
{�# W�}-&X �#��7D^+�$a��k��3���ĝ�_���e�{^�6���ג1���*��_��Mq���FÌ�$����*�U+�ͮ��oB���w�-�����G[��M�Fe۷�x/��t;eL�p��&o
������b�W�xjj��~�7�p�����ю�>dP���y���|�-�C�Z�Git<�y
���|�����գ��.xI=�)�P3kL����ʔ���ٰ��j��pM�ݙ�B���q��Ǩ�9�{P�<�h����Z�fI&�}IA��r��;�f�]�0�{��d�K�Y5(?��$A�_�,uAqX��i�l�2��^k���I>�砲E�b`6�p|h/Ԑ�?Q@9^���U����(�J�K�[��5��S�s���?v�߷ Sވ��˛k�N�I���AK��cm;t6���D�!�ƅ��G�w$�Ym����ؼhOW.���Y�-���C�"���^����e+~��c�J;ŮS�nҽ�fCoC�<!��]��H;����1Dʝ����חv�UO��N1r&�ğ��@�Դ/$t4�C�LZ��T��а�6���z��qs�;6;T��MU��Ԭ�L�L��^�!����U��D��	љREomQy'���	��G5;X�"5�e����-~�������r���z���k!���u�e���'���B�����m��:jb�M])��*zg1c�g�Gl�����|t�`�:Z�'��=���	e-W��S�,����bu����nci��*�M�3O`�
\[�XˍN]��ː����è�򖨞Rؖ��z:s{�{C���^�L�=�ȵ��5�f�hύ���/Y�J�fp{�S��m��ًyљ�OZ%PS8.Y�4�ԣ�M��<�y,w�X�nfbv*Q�9Y=%Y��x�e�0����$o>w�p/V�K&�V��e�_��Z��8���LE��c�����V�*R�r�����{�tY�W�Qr��sv{�F,�7�{-1���Ϙ���W�6i���6��x3�gi�^�/Ľ=ͣ��.�>2���nU��L�;���s3 ��[Ҩ�&��!�S[]�1_�2)��K邰���Z+J	}�t��:�_Q�A7�1@P�t=?�ѝ{~�6����
D9�Fℓ��)���K��ԭ�h���-�f)�+__	D��j��#d������xD�(���/V7S�Vt۠��R�(�Ѳ��u�W��̰Ï$v��C�w���!2���!#7�%�լV�mP�=�"��W�0����s��έcu����ܕW�Y]���̄��7 ��$��(�M���ة
g��ٺ������Y���'T2��2�]7p�#�l�.�p��%G󱁅��q�ও�b%N��{/D:h�nܩ�_\��؎���0�%��U��L?:�]�i�θ��}�#��bB��Z��5o��H=��D���2�i�"�(�zv�i�~���:��i\�������=�Z�p4�zZ�y�v���®uy��Ejj���eG�U�<ns�����r��}� �?��X���fi'+�a������vVwi%��A(4���d6��W=y��a�v�lM0w���'�M,��orBU'�~5�-1�0K�փ�j��(jN�,������c��A4�J9al�[B�.u5��7���
���o��Q���Q%`g��O|����%Xd���/��V�����#Ce[Lg۽���а���簠;�֛IW���3�{�8���A�רV�oo�G��)�Cμ��k8j��'x	���������}��`?*.�Ni��*x��33(�͡�<v���`���g�e$���
a��ވS����ɻ�g�Į@���kr����u�*��Ce]7k���+�w|P��h�i�a�P |� ����vm{sʀ���|����s��Ɋ�x��V��Z�ȶ�G�r�^���9�?5Z�����z�Hl��4臉��K�S5`�U�>KO;�,����=�q�����k���k�E��`Xl�FT��e�졷$�Pӻk����qJk�y�H�z��U����D�#&��������l�W�?'&�z.���ye8���6�Sl)���0��,3��_��y쇭q ߘ��n.f�T�"L�Q��:�%�"x���L����-�?�����x]�����X�R�{���=�b�[Ye�)jH�[��ƏZ�sa�\Q)M�I�Kik�v>Wp�4\r)��Ǚ
�w�a!R6�4��p�_��z�
t^5Ogק��*�Y�f�]@t�3ܧ�k��ͮIY�o�W܈�?Kk�)n$!���C�XFv0�%b6��� PgW٭�9�{�l��H#� 7SS��SiJk�ѯ�F�D �>�Kb��Аg�4C��O��+�贿!�#}bD�]Z��n�y�g�J;���ٺ��w���/C�?c񬤬&  ^��m�<���*�m1��hދ��g����S�A}�(i��Pc�������;��@ѯT��c����k�G��OF[9�����|�a���熩�E��O�J�z_\4H���#��������׼��#�U�IPh��.dE��Ӹ�l8��=u�V���r?Z(�$���'�P��.�o��X�TDz���H�,�J^�)���7S���ڧ��Q�u��ɓ7Z�����-b �@��<��3��E��ѭ聧�8�Q��vm��29�ia&������1���,��֨>C��ڳl��ڌmJ�bR�-b{5���M_#k����^&#�kk���g�i,a>7CY�x�{T:�Nˍi
Rj�9Z���:�:��qFH��Y����o�Xx�7E�6��X��:]q�v!��%�9C��{����돱�N���I��[N��9�J�1���S_��&1�1�r\c����g̩xI��cz�X��GN2��'�jw��g�G&�NFb��c�P�?S�-k���J�:�rİ�3���0� 	��j+r�@��]&��4����􇰗?f�e!���Ӆ0gc)�:}1���N�~s��8�(&s�=՞m���+�����s�.���%ڨ��o������j���h�̊x�%�n_w=�F��ĲZ�K���?���U�,Cͩ�o�~��2[����G�n�)��{�<Q�ev$�x*��t�d��+ �A���3�ۯB宒�bj���y�Q7F��]Eѩ�jd˽��T��Ϸ�>-KP��U��G��z�4�����F:٣�.��i^
=_��P.̟Lu��� ���ܑ�N��ڦ{���BFnq�BIG�c�j��>=<S��ׇ����j�E}	@5��Vr>�	�)?3]&-�{�}���9PH�(:[B$�儓�qs�di�20�/�^���q�I9�x����N��Ǌ����b!�{V�݄�eU�[Z�)�JP��v{m5�Sn ʋ�gD�HK N��*N�kQ�IRUA��9cHs�6<���߯�!������w��<Y��S�zL�h���Wi�l�-_�-��9�h�"j��^���#�+YOXc#���IĨ�iV���FXC�'F!�˔�h;��څ��8d���"�O���1�W��R�@��/_�>���U�:��V��5�6(
���W�L�;q���R�鰍���`g�=\F�y���]�G֏���#��&�єo� �'{s�	��Ü�j
3�N]�e���(���%ҵ���-��&��F���3cucXC��m��H��Q��65*ɵ5��(���-��z�?�xG�&o�TY��/�tr.����b$=X\"�A�WU*���@�� P��(5�I�c�$�M|g1`�_3\����H�K��TI�N�Ã���U�Rs5�����,��6 S���0L*5 Ȑ��p��!r���L/��G�!��n��m�*�TcÊ'�%��x8)af4m�)���C�ȆIy}�����n�:M*��Y8�F�ܪ�� `ߑ�E$���K6��	����(e��d�Zc����PE%&9cg������&m	�,Z4{t��Y�b�Q�jsQ�%Fg�m��1�2���8��0i���k�xJg��o��O�=Ȣ߉�2��np�vEQ;;�%/sn/N��ȍ����*�S��1z��)e��K��x5f���	x4��o�_��AR��ԁ��P�^�?�Bɝ�G{Ė� k
���F�&�lU���K�Э/�L������b+�4�	_x����#?Fm�
벆E�#��9�	7��S�Y��(����Z�u�e���q �V��X/h�=e͜���Ϸ�#rL�p%G�h� ���r(j�K�8�l��������
��Y���zWh3b����軄9 ����-��M�A^���`g��;G�.�%�Ԥ�������]��p��lwMV�+�@V/��wT�L#]�Ε�b�r���ӓ/���)�� Z\!q�i��kz�%~s&��</?����$Av�ӈ5}�˛=��ӕ{`5
��H8��D^�%��b��=l҉�MZ�߫~�0�:ik�iW�7޷��C��ua
4�+�Tޕ���6�~��u]�,��j��r����U\�Gs�ƫ3'�c�� ���M�Ë��%iB�ja4���z
V�(!b=A#���$.�e<,y�t-	��G<�w��Շ9�M'�<���NB�~5�L-�+�K�L��?����9�'�K�C�c�AOވ9��[�8.�+������s��o��=Q7�k�2�`B�ZOUg����h%S
��q ��3V�,��# �[�]V�,��Ы��BA�;cr�dj��3����������ڏ�*�G�� )�A��S8E��'����w|���E� dx��Y.�7��c7[�x�K3= ���|�7H�IrKEĞ�� �CbZ{V ��. �\*�ɶ~�g)�[+E� ��P���q�]�?��w׷(ʭ��T�������R��_m�����|X`�.�Hɥ �����5n�يr-	ϡ�7�?����<#�ٕ6�l8��b|.׆�5��έ�O��A�GI�Xb�;���F"f���dE�wXg$-To��� kȡ�z_��.����(��;Jޒy����E�φ_U��zDX���}�����s,o�R��']��z�$�5$�e�����U���J d!0�",�5x��cy�kq���ø�f�z"�@�Q�fZ�u�0��̇�����2���{�z���d\]�B=�+C_R����=3��[4X�d���]m���֨s��QD%IIs'�k��&>K�����J)����J42�a<r��ŉp˞�_ �ҽ�L�5;p�G�*E0�f\���<3�HckB��I�W�j?��O�K&Ul)���!S��Cqf?�=�� �1�{wW���9٘���hH�|w7�%L��Zf:��2���>����J#(B8�C(����$�&�9�#8e�ַ��:tT?o�2,����ٵm�w
��/�*�~6�'� 9$$�m?����أ�Ȟ����������C���k�@�}��`���S�Y*��Q~.�*��*���>�T�uƂ�8���X�O��pLk�*�N|oT��{v���E�!�E��_�"벊�$��������o{��CUDP�h�a�d����s8@���Щ"�)�1�֞R��Z�I����"'@��������T�$p���k�g������R�7�V��\5h�
fu*����	;!-�G�@�P�<�᫝+���Jf�"j�,�#v�@w2�xVa!�
����k����	,�>L�
��a�cmE^��Bb61r�{�M��k������mhf.KF����aY�8Y*��{/��N��
�]�9U$�וZN��Tqa�Nw���t��o��A��tE�h��.5:�v<��%���Cp��{j�݆Y��I�`�j[	�9�i�1:��S:PA&l`@��C����L�{g�\1I.�����~X��NG���Kǳe
g���d�Na��Q� +2�S3�*�W���5��!�3KK�K`�	R��+M������6�_���9��?!;�!K:�N�X0BafO�}̇�� �>�������&�L���D��uk+Q��0��)R�z��O����q�Wh���O�ΒgA�� w�_���:���>Z��#w��R���UUNͤruo�r���� ��[3��܃˸%�w6�e�hx%�St����
|�\���أۊ���͑�j�tˬ7����l���_dF��/������-��PiRG?��+���҅�u����ۤd?=���P)M/Lp�@�����z��W���9�S�NB�IqЎ'x���?��L�<�뷸����Ч"M}WeN�r�U��D8�]�I�{f)<�گ��V�(5=+$�����q�n7i�_���^�K2*�rI4Y��V+���i���!^t)�=#O�����U�Ӆ����J�͆�5�5���SI�6��F��^� ID7���k
�I3��AA7~c#˾6w8m�zj!��]�=w�c�Y������}h�1W�D6�Ȅ�-�w����"%�^�\}y+4�Wc^����TK�d���j�C~��!�1��Ǵ;fd�����_��cp�,qOd�1��fĕ�@k� /�R�yQQPڵ�
���F�6CFL�p�'��;�/�����������\��������������(W�4c3я҄o#Ш'6.�	���=���4�U�e2�+�#��Y���pX�����pǎ�!a��Wu�j͈��O�bmA�y"T�Qb�0!���]�h\�z���zG"wY������t�d��%�ߝ�5=�D|��<?W���������R�x���$��_�M�K`�&�\'�����I����^��-�R�Ձ�~y)�2��͹�f�L�L�k��������l/�D��_���~�m�X�/���z%8Y68$��4�О���]���y�f�����n�2X*��UY3���7�����ёe�$e͠&f���Pzeϻ�v�OZ!�`;E�i�cBI��3�F�`ݙh����{/\YY��Qh�s,�F��ݷ1φ��N3����i8�&�,E�x��g��4�e�X=����䥄2hk�n����u�;]�os�^�Ց������MTnS��1�ld)�X,K� 1p=*ڐi	s�o�m��_Ǌ	Am�����P�h�?�՝F4�Q�[��
��uF�*��m�]�K'g����e����^0+{*!	z%�`.#�n�Er�!������7�f��u��i(��3��u/�l��R9��V��;]�����X�m�#�|��O�c���-� �fP���F��?��#<T���ҹ�cWÉ*����A󄴈0 b�8�h6M ����gas�u��IƥOln�ݡ��:7�]Tʴp�#l��}��<"�[��w���'��	3�b[�̑��H/�����A�;*�\�zw�D�]Ǧ"%#�����?���ߎI��r}�T���]��.J5��	H3RD�����;s�X\d�A*���~��B:�iR{9h��p���<�4���/���z]���u�`��,GjQ����1U�/Ms[�|�n�Q� ��B����rS�i]m]a�rE�UtmV���(	AH��� A�y�a�7X�"KVw:��"k%M")�%�+B�&�~P#|-'��K�"�5��^���"�B���cD�AjPo9W��[�M�.���m�<�����doJJ!QR?��2!`�>O�r��3p�%N���̅lMH�VuF#���[�sE�ǗmЦ��̝�;.��r� 3�3��J�.���@{�%mG|$H)�_Ƽ�`g8 �J'�A��L+T����{j���M.�@���c��S�`3xO��8ꯨ2:����� !����ٿV�4��p�����ɱ;�g�]S�g�4
���Yv+�8�S�3]m45սw2?S�h.����F�Ӷ_6`{m�a��qX|��]�������~�L��c��r�ӽ��U]?봑���ٰ��l����=����5�#@��~O�֢#�s�Z��}��!���=�E2��Xb�/T�"��	H���ҙFhk��R�2�jJ��y�&�Z���A�y�5]$D���X��7�ǐɅM6'�pz�8H�PpFe.�������ɀ`�E�0,�����/�y"ֱq�&��"fX8"��?Q�F���h������5�����{����1��n]��j��MBRNa�5y=���[����1�K����(2sזXQ_�I�"�kq,�>�ë�jW)�Mk�O�^�nnaW���*Jp���_;R��@E5�F��]ҷ* '�f"*c6w�3�	�k}�������e!�>;K�ր)�^%!ΌCL���$��[�a�ӂ���fWO�9�<��b�Hٓ�7������a�t�<?��/�>J��ŕK�GCc����/.�!)ɴup�#�x�1��ɳ/����:Q�T�oٰpLwe2d/��$��9��B /|_�m�T�̦�#,��{�Y��]�n�.�Q^k}.�P��b@���C�B��E/�ѥq��R_�?��U��̼�O��+���E��|�=��V���:E3�"�@ݸ_1N�E\����r�J?>�F�@U�v�h�[�d����.�����ѩ�J�\����Z^ۻ��O'��/ߤ�i��T:�iС����6c��S���7	���L�%��u�����÷�D��-���@���<J?ϫX1�����bg�b�v�N2oKa�i�A�+�&3ܙ�C�,��9��Xi�P�y��53m@O���b�L��:�MU��k�T��JA�Y}a���Y�����atVY��R{
�'NA��
�q�9P�����v��8�q|�)�R>�O��og��m�UE̺N���:��lvWH�%\�CK��{X��!C��D�����[�d29�1�XS��&�c�������[gB/II�M�Y5�X�9GĂ>�憘`�����LN|��̴D�dSn�>��͊�0���f^�344f`D	��
+(L���[��?���B{�fHm?ܮP!6���03�k�}g����J�4z"��F&�"Ք����>z+�q���N�$1c��x�P��������hFC2�֊���!�_-��~O~�����AS���U�W��U��W͟�oS�z¨z����dWj˓�>�;We�]�x �tLó�5�w����.�e|���j;�o��7�O��'���yd��_�
�N�--�5��K?�Gz���l��%̅<�5�f�y�ߊ�=��sP$�L������Cl�D�.��r����kB|��q��U�����S���z]<I�ḍ����}�����|r�7�_Q]��{A�8�����J(0?p$RHo�][=q�rri|!�����^��ńxI/&n籗���牁��@�F&�E���ݺ��U�kM�ߎtJ�sۆ�A5HS$zӋS}�~Ι D���಴k�0IN��A���c�B�6��9�Ef!�����wU��Y�2��p�@h�$JW��s�c�u-pi�,"�^�y� �+��c����_���w�
C9eE!��{-;A�HP�9�n{b�򖗇��O*1�4�[�@F�/��ύ�WK4��ei���/6^����S�\;��&���{��ɬ����B���'�Sb�c��ݞ�Ͽqъo~��'�C	����5��K��e�{^�Oh����+�<æ˽�%��0`=��u��/��Y������46�l%�ɫ,��m���2�z8����G}����0{���Zth���K]����=�M��X�W$��]�p�/�}��K��ui뚏�M�.�`�9\l�Q˾�t�1ǒ�&�9�`�Y$HR��C��0���׬9+�L �d�F+��VW峍��j/j�A��Q��im�q�
�6� "N%��8��4#4�P%���z�ys44��n4nK�*"�wY.�V��o�����&ڙ$�'��G��/��'ۣeʙY�~Z�a��!�E��cϛn�����c;���3{�/�Y��aQ�L�s�:F�>b�=�1���ϩ����NiS˴��>#x�6�g�� ��=� ��?��2#U�n�7;��;8��s���,`��7䨝+S�[�1�x�)[�Kz������+�,	n����7)_���A��U�w`�P��>?@����@=����9�
uylF3���b:1[2�Kb�b�eo7�e��w(>+6@�	��y۞�#�%���홲�����﯑7�ţ��O%&(b��nGu��7�Sn�5w���f��c�͒���C�#�U��vp�^TT�N��u{��s�b*�w���^�Q�U�����W ��]M�	�r�/%� =�z�M�>���o!g�ɺ0���d~Υ�S�øxw�u�]��7p�Jl-ƥۡ�C�v�?��t���D�b������/U�W�$��VdH\�)�`���H%���ݢ(?K�����`�	�w}
S��i@��5@�H.�D	��c4��slމ�T櫕�*~2�Q:���iMs���������7V46�
0�'d����u����ϥj�4����UR�~s6�㫩���� ���d�-��ix>�a*gڃ0��V(�P-A�����e�y���vk��y�wu��ս�'M�Y�	B��~k�3-� �K��_�OJ���?��H���n�c�VIA���9Ҍ�[���.&6�����5�)�|oIQm����RQ`��rO˝����%I���'+���V(���`#ԕ�[����b�7СJ�����;�	�����] 3~��,�1��Zg�ȼ7���G7�)ڝ��b�8�Ŋ')�ȅ��c�|5�֐^�.�i��Y��.gE3��,��(;�-Lu������� w�9q�1D9�9�6��]ɬ�g�٥qo�O	��<�����+�]Ihոëw���#�/���(�ӑ�q��mL�����|��뤪��۪��_���
��Oq�rc�����?F����T��˖�l.y��`��^51y����OL�뢽V9ގQ[�1�������6�wE�i�X]�NT%[Ö�k��n���y���+�mduJ<y�� �"����a�P�DN���3�s�r��b'|�Hm;'�"z_P�k�He�rI�os�;jVG+0;i,D�����dy=-�q�.��y�?f�D
"�IQ�Fn�+���N���w�v|��V.������|]��T��weR	}�PA=)t�[�5�ڛ$���1�(?kas��lQz5�Ii>�kL��>�����)��IǪ+	��har���rp���_vC>��]�5�r�׸}*�=�f="�(J3m�k��p�t��``ܙ�XK�xY)�7!I��C'^~�+������Z�1�6W
�O9���+H��57*ԕ$�\4���k u��>2�6�@(����C��_� �ϸ�����
#��H���0��
9�4c�����٫��w��,/t��� ,�@� �f$�M�mu���ǔY�~��6�/|O��
$�/��K}��8��)��C��%��`�.� 0:�����z�
���^��@#OW�	��`�j|eG��1W^�7FEθ`�;,�_m_q� Vr�39��xh �%#����Uz�h�uXdVN^��!��
;������'��P�Z��;��4�'�}b�_����T����|3�ݫ/�L���!7d�͊�JU�@��u ٓ�Ȩ���-37e@�&�<���W��"幁�0����v7z2
>�a����Ϸ�� ���,�M�ϓ��������m;`�c�b��d�U��M��iks:2����ީ\ƺ��
�E]Fa���Y =L{�MN|2�
#�Q9KRk�KG_�k��q��Mm�Ҁ**oAQ���E�,�iq�:��vr��%�S�C&p*{�βݼL��?�$�Z��[��910btS�Sz&�ڙ�CZ���<��[g�!Idm����X�@SG�Z���f5[��xG(x?N�Q��G�T��oS�w�����+3�����3�<���	H�<+�S�OȤ�l�4�ʫ����W?�B�!9A��Dq+0����d�}����"s��-Q�i�K&���:��'9+�u��f� �0�0W.F���0�gm��(�Œ������_��-9�'�������kI���QU��͚|o��W�c:$���������n��`�eG*�x|zt�"��\����7����e�@���C�Xj�=j�j�7W� ��~V���d<�u���*�h?o-��F56GՉv�e��5����LF�A����=0�9P�BL&�����k�'�e���T�kg��B�qƆ�.;ǔ�֩��)<��7�h�,�F@��� }��y00ro9�z�i]��{��P^�!�(+a$��4��qĖi������^W]`>�I*��$��N���ܔ�T9���,n#�U�U�#��:FOJ���	�5KmS�f������^U ?*��;��k�E�Ii��A7(kc��I6�>Z�?�!�>����w�)Y����f�h�g�Wa%��/[-z���yd�"���^�~o:+�c�/9����Z�����C�3;!^+z�;vz�B��	�]�	����m�Oڃ�1ުIċT@!$�/�V��~�F����"P���)6yQ�f�Y�n";"���#�x�~ah�q�knK���d:��W�g�e�0���j<Hх�4o��X'��	�$ǜ3ˀ�T���ehcI�*�/��C���ƽfh��� x�=u4�i���|���#|чM��&X�S��(�z�g��	k7G�w���̷��+t�1a�n�~��5=)vx����Wf�m����J�Еnɳ�ft�՛;MM�(`�\����yU��L�#����0Ж�;�RD�	��)� ��gvm��L��(�!r;�!���N��ن4/�?�R����ܦm~}g�����;O6%n�y89�4~�x��%Wy�!v�w�nR�
*�RY)1y��)�Q���Aop$[`S�܎��7sm��eŗ�,<Z�ʙ�<@�E�P�c�k��G���i^|=��{�#OY�C�Q^�s�2F��>��1Ŏ��[�C��in!k�"X�x�&gU|�ś��=�_�ߚ�2�^ n�]�T;�as���lM����SG��1ˤ6)֗EKU>r����qh	i�[�#�[_=�A��~��Z'Pj�	?{r*�|m�v���R
0$�FN�b���6'[K�g�� ���ﶼ��+�u�	���V/�#��a���o�W�W�75J�e7?�X�{�� 0(=='���ueN��t����≲��&A�K�`96##�7�AO��Y@���n��LzᜌM��y9�Ra�Ι���Jm�ȱ�Wy��I���$T:���Y :��ޅMV�����gփ����?�E[Óo����]��2p��cl����\i��C�m��ݨ2��\b��푄��/����Z'�q�;\�����j����%O��؅??�쩒U���$�D}�ɛ�as�F�5�I�H)��Dov��M���@����p4�~m��::\eiH��� =�t���R4����g՟bmg�O��u���=��j��џ�U͢�s�����4,D ���^Rm���i�/a�{����Vc&��Aܰ�5
V���Qy#� z����<w���X.�MS"��a�BA��~��s-��K\ڭ��������T޳c��A��49M�[�w�.av��e��"g��+�o���Q�Y��y�M`�%�O���i�g%D��ǂ�)�	=VCe�ug#���[8 �����М�S��;�{�ce�3L3Y_LgS��d�N��X���G��)��^���8�{'d����w�d�1�q�LƁ.������	c�3���n��(~ĤZfKv:���4��(��-�tU��-'�ɧ�g:v�,�Aj(>��3��ɸR]�}3ճ��w���s��Y�<v`�l���pPm�1؀�w�|i��_�0�����t��Ʋ>���r��#���?��I�m���v�l�\?��"�7�I5��
��!�O���x�wީd���̫׻��q��EhJKXX��T�δ�Q�3�#=2�<;���N���(4J�`�y����[Ϸ<�kOD�u�R������݆�C��'n��z<��h�e$��Jr?�?h�h�0��F,���K�yX��q��TVf�)�"���Q�fb��8�	�������!+�1���+�;�5�C]����<��R���k�o=�dF[Ť���k��%X��1��dsM��Q�mI�y�k'b>�����Ҥ)�/$��3c��a�V� ��p\@�_�TR�v�&5�3�I%*vt�fX&	,�3H��k����[$����6KW:�)�0G!ĥgC
�2Slґ���w����W� 9*��X�H�!}7?\���[W���}0�	>M�8��6�ݛC��Q���	���+?P#i-='�l���7���o�7��<$٦֐wW5//���椘�� ʾՠ�mgW�¢~�٦���6J��S���e���}d�����j����)�{�ћ��ύ$ƵP�������bO�(I����{X5|�p���Z�r��Ei�ֽ6��_ȭT��o��N������ ' �`?U$�h��d���Ӥ�I��F��{��8�� Z�^3��9�'Q"���s�05fT0��W�5�A��ޕ�b�7�d�����[ڹu�.ړ���˺�-���@{��< k�Μ��=⏁��ƣ��vY��2�P-an����ӷ������9,�zM������V�2�m6�6�c�bg䣞p�MK+�kN@^���`���WW0,� D�a�o	Y��q{�=#N��_
��V9Fצ��&�?q�,��˳�l$o|��ͣP�E¾#��B:I��v�P�%k�Cw�{ΰ��Wv��:JA쵴a[:T}9��1��S�/&�����t����]�{g�44Iw4�Op�Xh��G:S6�f�V��ә�3�N��v�0���S�zb�(�+�&�p�9�3|e2��	�-[+ޑ:���a�˓��4�y�?R�K!TlD����0�~ ~&}����v���  �$'�&�.�Պ��~0�+���u�O���U\��� �����y�� ���8%���_�"��ش�0�Ɍ7�F|,���U&sL͕1o	5����&�Z���I��(�qe� x��t�������.�
�H�VӮ~"jq�n�eL&7��y�t����d�?X��YWϣ�'-����AKrG0_5� N��P5w�2�B��)�U7�=���P��L����q�k�B)g�:���F�Ն�bB���q�2�6w�Oa��7<? ��CK�����P��}�[^_��r*[鮕�]_m{�좳��:�B(&�$+ړӔq�� ir�v�yJ�^�����I% T�g�a�	7ց���KĐ��Dg���#2U�����JJ<�b��#�5��>S�s���H��� :Ϳ����k=��I��DA��c��6(���KZ�!���N�3wˍ�Y����fZ�ha��WUK���8-u�Լ;"V`�^7���]�+�Ʒc��ŵ���U��-�=C�"�!1$��;�.\��ʤ��p��=0O��m1�[���g@��[/K���JEmAHP����w�6�������}�;]�"���yƃ�̸�)�O�����I¬B���k�j�ٶрwo4��'g;	���� ��I��ek��%�js�ҡ���@���h�۲0.��.u�b|���݄s���T&Ѣ�zɡ���u�?znEb���G3(�@�x�<t^�?�I�/�N�=ľ���W��Ī�1�e�K���w/��XM�u�`�;/\"��4'��g���@������r�R��'���
:2��"ӓ�7�LSY���z�\��ؤ��Cz/ j<����ڻlm�?����v�2%	��8��4����ꄁ4�yi/d�R�cn�۱*Xp�Y$�W�H�ѯ�B�\$$ָȠ��֏r֚�]Pe�����ZOS�W�mE�c�!w�䵕�1�Y�^��3{`7�Y	� Q�	us���FSc�^�1�B-�_F_��k�i��I���Qxz�zg� ��6��=�����`�2��/nܾ1��;�sZ���b��X��^�FS��1��;)Qg�K0��!�/�aS	dȋ�~��_��A��/�mu�PEF�?�s��_�V��l�5
���Fi�z�X�<K�ƭ�����/�-+��B	��%��#��S��C����������7���s�E�%(���Vu ܶ�̏���DU�	�͈R��;O*#^����G��TL��^C�ZO�Xu�-"���pi�����ÈIW�LA��?J�%�` �o�mIM� ſ�Rgr�������������n����V]%�p�>l��������p���Ӹj了ʱb,E��/��J�Ɍ8�\S������W�t%��ӈ?Oݒ8\�?]�} ��y�Ӂ 5v�zH$\�D���م�슉��"�K��~���:�A@iC�-J�g�/\����4�R���
���J��'u�,D�vCj�R����hUH�fs����84��4 ���`{����i�@�a ���_xV�eY�<}A�	ߐCΗQ�y>�l�Uֈ�7�w�6���Mg�6��B��~�x;-���K7������/��H���m�cu,A�f9ȗ�[�<�.��C�>͵�}T���mo{�dQ�~���`���OAT#��%?�B���~�V^��Y#��[sv˽��З̮��;O!����x*�34%��Լ���N��6X1G���)z��ī8��'��q�,�r#矌=E���.#��O����~3)���	Z�#�o���`1�d�숍�/ y�ޯ�=���ɢ2[g�2K����g�a���F�f ]>Җծs�wC��ʙF��<;����G�(	m�񧀷*{|Ĥ��F���c���z$��׈r�󚡎o�?�6�(2�w�l$`P�·S�r��5g�d��j/Ou��3:��u�'	������i�EK�XS��T�a�����>����d���Jr�y�c^k��r�~��@�DDZ���Ő�苎���>�Z'�t(z����e��-�%�m�zZ��0��,�Ɨ��uys;�q���/ �f	/�"S3'Q~����!ѧķ/�\�l瀘���f����]��\��,lR�Ǝ���=u[[��S�P���V�� !ls��Q��iI_��k-�>7���;�])����`��r�a�a�����p7�>_�����5�*��n4�*1�'fsT��3#�k.�͵ہ�V[��O��KW)�I�!?�C���m���,8�y��VwW���9E���zHj��7z�,�Z)LR��M$��4>h���6����]COX�V�۸�,��ֵ#$�UB`��&�{��m���%�١9Mwv~/�{�i��o �6e�m�A����4��ڬ#;e����QS�@7Gyh}�D��������=M"ٖ�����[���ٟ�&;�����Ol\G��'|[����(�N�EЄ�1*Y_#��v���i�ܝnqa��J���|U���h�	AdaY�_�j��E�[4˝h9�>�;Z/P���^�'�������K|[T���2��S��el��R/7T��H���v&u�̓~����{-i��@v|�<[.��$�X�-�D(��q�v���2@�za���R!8�W�v���,�9��ia��s�ͮqm1��ԗb"`g���JMƁ�k)f����*�KRޚ��탻J�a�M�Y`�{��N��
Yl�9A ��p���q��lc������o���>/XE�p��4 :��v�k%~��CܝN{	�\��l�5����	[��(9:&�1&GQS���&X�C�y��}O��6�gsg}I����=�XCGuk ����Q�¿.��EN���=���vS�r��@�!��w��37��� G	>�e+�d�����������'�wA�?ʏ!o��:�.0���;�S}8JT����E��߅B&�d����YY�+=�썜Q��!��sJ��}�;���]���M��;���[���x_>l�M&�K�i���t!���h�U��͐�od���8�.x2�Նf�$�ce}#8x�t]A<��u����a������*G���j+�`�q7O2�X���0�d2�������4-R}@�<��G�TT����k�(���+���)ې��=f�P�FL���,��]�p���ĳ!�Ԇ?!<BMl�q����S�
���:<�qh��m��X�!}��~���r國��\�]���{��ƌMW�x(!h$c�_��a>q�>�i�wV�T!�^�TX�ZI M��4�Ď��J~e��j��~݋��U��L��eJ��܆�]k5u&�S��ʋY�O�� 5�e��k� �I�˴A-��c�j6cŗ�攇!�:_��7�w��Y���mh<M6W���4[-p�/5"�^R��e��+���cJ�0�P���P�vԈ7GCj1!L
u��;����?����^s���hOP��1-Mā��@��/�����+|<<�v�5�2��6�v��\U���~;����YW۰tK�'�{��� ����L$�'榽���{RUo�M�'"Y�	!)�)V,z>��[e��G�@t��u�\���\��ۍ`���suj�f�����Bg�e�4ѽ�R���o��Tu�z	C����G����c��5��t�~*�$}q߉*�=_'յ�l�W��������d𲳐���K*M�I�`Ԃ�\} ��q����|�����
��Rz.���I�����O��R��L�����_���c�(�э� </{�9�ȾK����mt"���eñ	C%��8i�44����}/�O٨y�\��-�Cn�S�*��.Y�������ǴE�w�u$Q1
��~G��Y��:1e���kZ
���r��E��c�T�D���sT�=���{kUY$z�QTVs�ΒF���t�1��Ϻ���*�i�-P��*xUqgˤR���0=�}��P�2T�"n�?t�G�;��s�[K��y0���9�S�y1]�)�VK�s\f���TH	_�7��T�_�I&A�+i��cP ��?��ϝ�&U�V4���8
��(F�1;��j��p�K�ŭ6����ed��G�+gA�	�(L�e#�e��1��(��
C P.7��2���(�2�-u��j���F�2���Z���m���#����w`c�Ox��_�*Zd��Hy�Ӽ����m��&2蹾�W/#����Z桄��� �1"�TtMM���źUug͸��aۥ��jX�;�J�I�-�&�]�p�p���l>���[��ǁU�c@ӓL����b�	o�zK5/ffh�Ќ�ɧ�\�0Jذd�ǒY%�!�Ϋ�?\�P��@�Z�7}{6����Ӽ;:5_�HJ<D%�����7��\���N��&چ~�'7:pGi>>a����?����4x���cП�������u갲�y�j=���vUÕs��8�Z��j�] �9��I�^z`i�q�a�b��CV��y!��A
���&��4yY�@p�-����w&�AՎq�M�'�J�B���~��-��K.z� J���5���8�
Oc0�A�X�9C�[d!�.�V���TN����:�Fo6!YQ����ot�`�%�O|�٭�z�%:(��8�g9K8Vy�8k�8#e��[���3NfВ�	�;
]��x�@�3J�u`Tf�����]GhN)+��w&p8�l'�2ԅ�9��mʥ������I�.>����U@����3dl�����Bw��V����������깯�c�ɝoFg���F���\�����7�?3�]�F�թ{w��>�T9��ŵ2q[�"CS"�m�/����|�����u�,��j���|bZ� �{r4>ꡉ?Wj���
���l��M��׭x}5:���ӷO]�+������w5��n��bkE�kQXN�ST6���į�Y	2�2���? َ�JX�y}bW�]��-p���!�D�^���YW�#�'3���9kt'$~{z�K�����e Ћ��)@'�0�u,U���ny��q�ԓ

�fDT�"���Qy�<����.���̂��Ӈ�2*�k2�]��z��OR:�����=��<[{[������J-���|!s�YQ�=�I�P�k�<>r����)}��ǻl	�]qa���f�pLH_'�6��g�5�B��?*�APf��O"�(3�L�kiFV�P���Q��ܪ3K�|)��!�>�C�������Y���
�B��W;9`��N�LHE/�7� G���M�����x��c>����R�A0CO�r��F�I۴�;#�R�]Zf���k��e����;�ٜ��w��/�� p���y ���K��mF<��]���z�gܣ���I%��z�=�}�����̌ D����ٱ[eё+K�I*�+�H��P���6Ohϑ鱄B|�#h���c���E�k�,�_~�[�1�]��%�����2��UKQ�h���dg��po�穉Z�xW*�yOJZ�a��ܣ�'��ߐ���f��T&Y�����˅ �ȕ�b 7uc���GƑ^:u�9k�Y\�0\-��@qWe<�h�D�ىs<���$V�sa�vϘ�2�՟a�������Ǚ#$8,~��`?�<��hl!m,S�td-b�������MA�k�f�6�v���M��O�vq%a�K]Y�!A{v��N-��
��	9</�\����?q��h��Y����o����-	E�Bi�zE:��Hv��_%��?C���{D�ݍ)��0d��k�[���9U�z1��S���&���x�x�B��g.��I����E+X��G����R�\L�/�����x�N�1���LrYqSZ�ֵ^�,�͘�ғ�3��Ҡm	�\+�WX� S8�=�9黦Y��)?ȽW!�"ɴ�|�0�6	v}��@��~�����4&��Հ&�4��+xB��7=Ǡ태A��<��V���:��A��v�9�n�`�	\_��fj�{�f�q�-Q�����C�U\�!͋��o��9��I�ƭP�}��V����eP�x\�t� �� ����<� �����"$j����[By7h9+����Kn�d�@��vy����-���7�~G�iӚ��ֆ�( �����c=�\P��L7����x���0����c�zҩB�D�q��(?������8s<5�B��l���I�_�}����r�����(]�,{�dM�T4�8(�$��œIN\q�oih��/l^'�1+@I�*���3�-��В���ݥJ�&)U���K,�J��z���5���S��'�?�_���� 0s��L��k��1I��A���cjbs6�����B!�腿��wA��Y*3��\��h�W���� �-k��ϊ�f"̇^m���:W+{B�c��
����K�����C%`�!g+�v�;� 0<��)���m����aOQ�1/;���s@���/��㍀2�7܃��y���o6�Re�״�n�;�����@�o�.��!�Zm�Z��?�'������;r\�v��o�Q'ݳ�	<۳��KU��Ve9�Z�
{� �y��/[i���y�h�<)u�)���3�)�� ��؅ɗ���J����Sz�`ĩ�}5G��n��_��P�tTU!��"C�ċ�=������Ww�R�I	��U����k��놀�M=`��\�F�˪*���+�����å���EA�R�l��8����ט쌹m+�L��Ȳʷ����Kv��z/ւ7�����ڐm�$��vn?��g%? �81-4�uʣ<0��j�My_�D��Sn�*��1Y�H��x㯂򌑒�$���m&�����E�e�Q^=4�Z�Ľ���mE�c��ߛZ��g�fON,4{־�Y?E Q�FCss�%F�c� 81�
�H�t	�i��~��d0x04gi��l5�=�<T߫}U2<�n�';�<�s�*�՘0&�L���Sxn1�~)Gf�K����@Mڗv�	ZR`�4I�_nɷA��*�c
TP�y�?,�@�M���vs�"�[
a�F����N����KN���э���PU���+"׭	g�Ǡy#ae'�l�(���Y[�"7pʵ1��;S�(�ݗZ�xu6W���8�U�40f�~?����#ԒX���J�L��p�ԐO��V��N�p����J�Q���y����W�Vz�S�u�A��R �ݤ%M'�bŵ7�g(���(e��N��1�$��a��][��p�>gl�7Fۍ3��P±��F�nN��0%�bbu��/��X30�y(�2��so���N����@��c�{��~-��I�)��mQivސ�#�f=\�$G�Ѣ���Y���}atlf�&��;]���{��R��k�*G�<�g���@e�fp��K�ox允��(��a�
-���8"p,Ś����	���S4>��50��O/RZn߱
C��z��Z=NR�E_�!�^5�g.�s�����1�:�,� �Ĉt�lw�7ZmgCDl�}��|Zu�y~�A�s<_O�tX�hjZw	�(�c�����/��AC}�������f����Q�(W0F�S�7��Y&�B����$(�ݕ���Y�FĠ Em���,���Ķ�6F�)(&�M�������T�O�c"N��<��]��5H�����v0P��G�O�h�B�|����3ԣ�ܕD��34~��1p�i�n! �`jPC��j	_��O���N�"nz�HM.��63�D�|!�(ȼ�@*N{����o����8��ݪ�6�}��AH�9g~䐧tJ1|f������'�˅㔬�]z�➨�@��狵�?"=W�GP�r�(˲ME]%{"�<b/��o.���7��l��{�Zp�O��������DB�e���7ƌ�<������n��-�_ �#*D�Q����[���<���5����~� VC�8�	8b��s���t6�j�0���9�M�5�i�i�ހu���-�̤pm�%=w/�����şq/{&����DC���q��'RU�3�R��2 X���T�����g��b�� ���R֓��kdvG����)�|R�/ɽ�&Lo�V�0��sy<��:�߬�!�Qg��>���-�Z�g}�yC���_sK�|��X��S�[�T:.��lC�a]��/�7�w`��-5P�S��_ػ�Q��&UdM�o-5�?n��;`�/ۅ}9��E/QD֍�	��#��-��#�я�2/P����TO������o��d��?�k�d-\5�6�	�\-��Y*�d�ۊl�Ԣ��]��H���Y�n�_����nVFϥu�x�s&�-���2u���V/мw�nA��Sr5�
��!�ȝyIi9
����@z5,�EC#�:�a�ov�ȃ�^���.ZY�Ź��"}�}?8���kZS��g�ufͯ�o��R�E#�"����4�b��=��|3[F��oRf�t����mhF �J�IG
h�|��!@p6����G��@N�7>seIR?���!�v&�k#p�$W�M�TQ7����ɦ�0%�_ѭ�\#�4!��!@u}
4�������>�#C0��U\-�B:�!W��`]�kTf������]��q���Y�׆��XD/���n���8��;0�r.^�Y,��܉E<)!�h��d�tq�r����/�T�	vAvU�	>ܓ�Fl<�3l���O���k������z[�7�>؏e#��P�
�os3����9�(����GM�݄�����e��֦$H����.�(��*�&����S�ţ��$e�r�*�(R79j]6ƅ�?�dg��Z\�#(W��p��G��N�L"G�mN�+?5	�D����DO��<Y�P�7YpLL����=~�R����Ɨ� ����^��n�&�jj���2��3���+*�Ch�q.׍gr �����M���2xUX�E`�8ω����'�l "�(%e�0�e4�}��Zwk�;E7�������˟p�����y��(�EEZ�n���?lу�e���AE��ZJ��W��1�מ8=N��<�B���S2 Y���F�9�%�Hc��o��5��\ƁOSf/�F��[\̧\ʴ�/���| ���?��h[l�	�T�[%a.����cl��75��v�w|h��6�{��AY�K�ª� }5��L�����f�?�ߏj���'F���f��s���ș=�?�رn�I=a۫�����霗���H�b��1���e?���vNu���{��sh.�2o�u�:���5���* v�P[T�h�;*J�FТ.�q�_��҉H�gKԯ���H[�{������-�bH4����=*N���5���k>b�Bo/�Rn�`!w,�#��ٞ*v���>pN<l���Y@���q
��awQ��|��X�N?���Q�ld�Z���(q)��'C(�o|�ީ0L?Ȣ�Q�rZ�-�#E���O��+#�,G���Ep ������}08Zf�ك��+�ð �6}���Qo	S'�%C���V�*ڜ47{^�6H�?�q����|�emHW'wNn�㣔��Ld]�m�fh?���D�����xо[����9�nL�/l�Z~��p �G��)P�A�U{q7^���h�j����%$�59�����w���׏c� ����h���u�xW�kE�V�Q�bͬ�)b� d[%�G��'kf���Z�Z�;�H��^u�Ĕ��S�l�ҧ;��(�6�Z���?��l���gtǴ�'���t���s������=8��m��GB��2��6�YOf�F�V�%�����Zo)ξ�p
�ƃ�=SX�����[��\�KOq<d�'� �@/?+�h��	-�'[��G��[8���	l	o�5rv�v���h#Lz��-��`Y�~��)�gDg5uH{���Z^9��]����5�,�'�Bo�(�s��Kw�=Y�T���h�a���/�,�^o�Բ�Iӽ��u�&ka�a�Ҷ����\��#&J���Wg�V�~�_�{D�X�b�w���$��Ü��lp�T�`��_���d�r���X�^��9x3��a��l�b������N��e|'fI9?��~)���H�����ֈ���iX��Rض2[��]7 2C��X*�H��϶We�$Qo!�%.��� ��E��/�;��\zU][��� �l�O�^/	����o	HK�Bz͔���ˌ�!+/1��O}Y�,�����̀���pXd��E�b�3ԁ&�y�S{f
�E��.�%w��6d���>�sd6��Xש{��|�[ .�OW6�9@T�3_B���8J)ݮ�{�� �S�)�����U6�y��v��o��cuD5H�y>#8�H��G7qUY����.'���&�e/QH�Y��cGȣ��,C8�1}�<�I\]i��/���4w�`��&A�O��	�B,���<�_���JλVg��ȖL|���bv	2nN^�,ۃD�Ze���K����ޖ ��{6�a�����Ѓܑ�Zu�,Lh��5������+�u���/�^�Y@c����{���oJ�ZE+��6'F�k���6��;������I�J�����׸\�����M�^����S��}�ݗ��칐(��q0p�2!�c�`�	Ix�76����\��g �_J��q�J7���C����OKU�L�8��#�㦭�߈:/'yXH��5��Kh�����Ȍ\
��%���f���X��}�d��w�I����;�X.�%�p���������V��cZa������`��w�'�6c�ۄ�r�-2!�������,Q�ʐ� ��M7���}�x��|^�nT_}���f��BM+ٴl�S`ƫ�X*·�ΧǴ���f�F�K�v�x�m������/��a
=۳oUn8i`1�#����f�^��?��ji�H�R�h8�QU��%��;��A�Rv�V_��^��og�m8�$}NۘIAu,�_���-�t-���Q%g� �l�rS��������A�7o&�^t�\���p-Y�֯����`/�K�A*8�u��ђ*�h�Y�ӑ�z�������)l���Ŏ(��=�N��A�|�gym�̼,8���_)6�](�j?Mu!%�zv�8�v�Mc)��n��P����j�Ƣ�C�6��P�U+�v���IW��f3��<1������3��԰��!'�|`q=���MjЩ���Z��n�eMu�}6Z��%=�M�L�{a�^��3����$X�6�Ӊ���H�#gFw��N��1������ֱ"��?��E�]a"V�o�"�|����"����n��f�˹��]�)"��^/[}.'��7H�\�1.��k�O�8��gwB��8D�x�e'�[7-	<׋��-6�ѤqFe|��jD^?j�)���³��� n�57��z�eK.V
��ܸb3GJ��Si�,���&M��U�45��0����ܣ�'�'�3�Lp���=�Q�ˮ�ņ��B�1��ۘ���=V�T�R-c}3�%2�T��U4�b�Q�f��Og �YR�ع��U�d]1^p1������������m_h�}s:0���y#ҫ:us.�5Y(Q��+>�m����`g��y*�ɾ|��KpkU�߭xS�dT����V�h��?C7�!`-H��JSUy��3��GYdT�-��n���`+�Ʌ�n��Fh'Q�E��0��* �-�����0��B�r���*��\���s�N���4>k��z��5PVLp�t�MYQWИ�Q�p�I�oc�}H�"�
��'��N�n<SϬ��_��&_m���?k2�I��-@�WBNnhBSy�z��㞟U8��Di�i��û�=m@�WEv~�LÕ!���6dx�*b���Z���1	"�4 &��^Z�g�5;fT�o3����"D�~���R4�!q�)|�oF��o�@�t���x� �_CI.x�
��<|4�!ǰq�m�Nš�g��7E��I�j��<�?����#��$��|�{�@��S��|�Ǌ0�߹�46�#�s��M�u@2�4�N��KC>Y�0���U��©�C!H�7��I	k[�:��9��$���^�Θ�b��ΗX�	����Q՜ݗE;�gn��9�K�r����v�)Hw�h�4p�[�Lr�y��['���oKv��U��>%��M"ޱ���s���N8����`ӌT=>�W#�nP�xo:^��K�9!$�Y����Cݫz��e3e|=v��IF�y�:��*�*����[	���
��re���*�7�[16M��?/\���>��J�EW����7ʣY��L��<m�E�?�wwD'�^�k���C52�O���7L�V_�_�B޹[�[p1��5�@���e^�A�͜�j�
0�Y��z���=h�JYh���9�T�� +MN�mO �:�Ux��E��]�����# ��%����~j��,0Z��;L������������q����z�(�3�Z�%��Al���,����7��ᑮ�5E���H-����8D��P�B��L���YT��F;�%
���$o���gA�H�fS����r�[��\��V!���� ��?�!�h�	2a�[��t�-���xl��5�}�v`��h��퍘���Y+��Ѹң�/25������W�$�ˤ�&�F�C'M��Ms�sn�"xO=^8?�e$�a�m��8��u}��4rV�����,�)�(��vu�$�����G/.[��V�:��Ü��(#v)��[[D �"��َC�I��qf��M:�H	���(�Զm����B�з����5cb���=*u��ή��%�b�91o֕n
%gw��!���g*�ώ�E a<SOK� +�w�b�Jd�w�dB|�X��u�8�{�Qq�~���Yf)��������,����?πBQ���ݨx#��S��G+�� ,��$�l`������RD��8:�
��+F�gT�}��<O�&rc�F�.�8Wx}]A�$���)H�ޒ�k�s}9"E����E)�])�~)�ߔ�`Ϧ��(����)���"CCB���1�*pߡ����'�1YJ�p�ib��̅z��G찫k��~�~_�]�?5F�\��M'�e<��d��+%�
�����X�t�uF �W+,�OX�w���(�&A+� �6'N�T4٤W�um�$��Wˠf�X�=�k2R����
U����mgmBtt2�Y�?U�,>c�8G$)ȱV��A_��o��3���T�αus�G�	�Lg������إ��!�>(�o8Tx�q����i��#r*���N��2!��f2x��ڤBr���΅��H�Ct��������h�!��'��
/�1�;�t��M`NT��S���-��U�-�o��K���$��b�mC��կ�A��j���r���B��yp0��b���λnt\ذ��ݯ���>�]t�p&s@��M��	�J���V�a��INR�@-d��
wȷ߉�'��?[�	�ګ-cb��d����K���#�(��G#�dpǗ���oc���"k����t��|=c�~, Xp՜����s�K�a����b����}�=���8��$�|�[9!��>��*�//�� �ȝ�{J+�$պ`E\r��4��1�i���vy�Β�G��$W���>䷶s�z�P�B~��o�P�h�צ6G%zÉ�B(Z��kŚ����~�?�c-���5ĺ�M��>/�y�s�ˤjKPA��ʚ��i�g �>�k�4I���	j��	���26���U�ڈj2�w�M�v����� -V2撕��L@D��,����<�xF���҄�~�Fxr�U7Y�,��nW�1C��s�K�)�GI�Y�������+�f�j�3���4n��M��j�"@s�Q@&\J��=�3o��Ϭ��"msD��V=�	N�K@��e�������18ࠚy�{�����Ҝr<ߒ��TS$�+�h��)���GNH��=Kƕ���$��������:9Z}`x���1�{�L�������cV��e=�~N%�3��Ÿ� ��������q�@���4��X�N1�3^C `����Y?�}� I� ���i μ���|���=u��Ѷ�D�CRmͻ�:�ՙ��-Fw�hhu���:w�G��Fi��O�?��Y�!��gPKs�ۢ�A't\�5�}I�OJ�T�F��?����)/5L��7�\�m���w[��%1��,�V�)枋n������z=�Q(2X�f���l����M$��l��E�<�����<��U)�P����7Q�ո���5X*բ��@u��jP��K@��b�L��kݯQ
Q��(��l�8�e9j������|>��t�D�2Բ�m��C����	�_:HX.���XRpd�T�i�p�VY�5�4tl���b��;40ְ/c'U��y�Xk��Hl�iH��O�0�̩OW2Yx|�U�ok���� ��d�|�ӤE]t��\�xq��d��
T#�i;b(���
�@)mEp�=
|3�Yɛ�Ȋ`��F��3ԩ7����3�9�/�,"8MJ���9�$T�3q4}s�(�X�y#N���,,Z�Ѵ�'����h���VI犊|� S9>#\��:�J&l��*��gYP�{��k�	_�8n��	J�#fa�������Xi)�%�|��Z�٭� ��*|��x����r]L��q��:�`�����r���}�~F��Q�Se��:Fo�	gPL�n#�(������ȇ���ZF��8�i%a���"�VA�s��9��&l��Wq��r�{O�m�a6���_a3fS�B�5;���<>�M��-��"� V�`|��H;�6�;}ʦ�'wx�{�MLS�s���V�ҙH���mͶ��ֶI9f��ZO������ j�@y��Ƿ��&��p���z�HґQ�n�IS���PЖS7y�Ϙ���7AK0߀;Ʉ�r� E��*\N��>��6 m�ޜV���K���۬sX�ᛵv��!��ۤ�TV2$;�`h�'�����«lQ��
�~�(VdA�v4���,}m֕�� Y����)�/B���./
>;G���6}8sBBK7�OGvN_��W��*���
F2\o
���������d�D�32W��\������9�51����Z�dR-�	�4��>�)Ճ�ݾ9BiT�1�'v�?����y-wٲ;e����pW���k��`��nY�ߢ��u�����]��.�f�R_B&�����=�Jm���	���r��WS��X�������֛�����s%@`I�r��ײ٦�i6H# ���?�5�#�������"Y.P�Qo�O�/Z%8.�� q&�/^Py�=�wL&E���̻�v���L��kD��7�espr�ta&�@Ѳ�8N3sW{qO�!�!4�sхa���Žc��ܯ�M��R��c��?M��2R/��q�oM�T�ѻ�RMC$��	�fE8�g'w�=�>5��,T�?�60�6����4_�+U(��'L��,Ԉ�y�����]�3��|�4������t�p�{��w��̥lڊF���3IuRD��������X���s����+��n���Tr��P��"�`�(�-	_����m������O�߬�zo��'�B�/{#s}��Dz
^ч�EÆ�С������BH	��S��T$���yS������\��Uh�
���� ;��i�P�*
�+�ha�A��.Á8������fW�?i�Qb��;�/�`��C���D�[���R����y�_' R�P@��,�C�9�o�Y��gZT�4��^��P.� u��+�ŀqA�m�+Qۋ��M�3��y�������j�)I�xK˲�ӫ7L�%�)�[�L���%��}��/f���$I,�{��a�ǆo���hPȫ�S/�$@�u'^c�� �Ѧ���dS�b�"\�����t"�^#�C�IOp6���j�H���6Y��^0�=��(�U���H��;gr����݇�;Jߓ}�.�?�8��R���J�vWT�VED+_+�i�y�����w��F$�/�����l]t����_��'d�L�K�kb"9%�D����l�d�VW��O�#��Ҭb'��9� ~v���e�I���[����Zի�y�c�a�DP	 	��A�3���De�!�$^'e�]9�.��� �xE��z�hH��)�z�[���7o���N�K��)#ǜ��H�Hz:9�ߌ�����M+|v�<����	�t�M��c2KX,S'����b)��n֚yL�f7QtE�Lt.ԏ��\���$��!�sQ�����{�$R|��.�J�Cp@7_�����"[)j��{�� �Щ͖���9bU��0T{�\Q���3b>uyߒ����TjU��Թ�'�J&~E/~B�&��dvG�C;���i�~T<�
}]��&/�N)4D�K�&���\/K	0A���w<����p����K�h5>�����|D	Ǎ�N����p?�Z���xf��w���X�{C�N����Il�^��Is�h�9�5�k���S�إ��ҽ��K��5q��^ᡣ�J>A+%^q��Ȃ^3ԏ�� �BK����n�pRJa�˯��C\�����EԤK*3ŢР�\未;��Y׷(��(qݜ2n�M�M�+Ia�6
���}���Z�_W�q\���C �0�nu�K�I[L�����#�����o�/t5�X5
��­>K;�?Ч�3��<v\��%>��f�X��&}���nxI����2U�e�%1��X�G��E �v�~���/��)��w�Bd�Կ�cӎ�{�h-�ۂ���	�;Q��q�*���5�8.�el!�	VG��=�}u�uf`��OC��a$��Q���8*[�˳�m�T�OfLlK�)�xy�y�����a��D���86i�Y�0��U��8>�g��z�����cR�袱�u0e�h����R�|I_�;?^��g����dH�N�,z���%��t��Kz�g�:�l���r����:A��as.�t�s~Nz�D�壬H�[g4/���A�+��5�o4��v,�s�kM���q�����֮��^�(tG��ے�neH�4pMm$��,k�X��6ZG,(���M>$|�v��tc6n���κ���ǰF��/���c='P�F��+�V�����23� �)���GLi�`L��}5�!�M`~Rd����j6f��pX�b�^n]MB��6�a������`��T�W{N���D��>���)6;5��9,H��yg��!�;�71��:������v�_����w]�?��NF�i�;����"��b�[�0�!�ƟI]��"�c�/H�.��,7u������#�O�����c��YD��fe��B7Z��<��X��<��'2�IM�7��DK�����&��P����)�غx��VW�%�=�b�ź�����&��5"��Ra���Q�}$�r������`��p�|�=3���h]�3���M���v���Z�j`u�!B�R��U3ǜ�Ƭ���� �Oۖ�����6 �r�Rj?Ƿ���d
�^�����Z�͐
/���;�:�����I0���y��:���"��Q{��>AB_�^��^?g��3y�BҾ��K]z8�l��SAGTN312��u���c7�r:`�^I�ES��+�����&"=da;W-��n��`վ�'Ց�s��QX�\��Û7.-D#���V��(�����-����U���m�o�k����z�5�6���*AtY�����t��9I���xjh���� �O���n���Ϲ3��"F&����� 2�b����X�$t|n�o6S������[���M�1��iM�u��Q@������Y�_���*փ���Y�ٗZ�!Y��3�"�/y3�1�Zgֈg��if��oIv	�Y�@"�����k4E3��Qp�|Ǡ���)o�`wt��[�X� �,�I��Y
'�|!{�!T<v4��h��ԑ�7R)I����}�,dM��o#�=$k����肻c��9��~0����;�#+-����u�h�4�R1�C�1>�Vt0��*UpPw�ք'!���"kh�~��}�q�� �%u��@�XX���|"��ϛ����;D���l6�Iן��ܝ��)��h�o&���r�$�H��hi�vռ�U�+�>p��Z���?���3�;QtMt���ߛ%K�$
OW�}���T]��&�.�=�n��,�	3�r�H�S��K��*�C�̷/�Ɔ���5@���r�Κװ�'�S#~y=�}���%�p�ċAo`�PșF���Z�w��'�q$�F^p�=@F�&�4��!��4�"��uuk�U��5ڪs.G�t߉m&�<J�6�87�W���_�G!2[Fs�8=�������7��Q�Mf�%�}�}���0Ê�O�q)IڒCB���M� .�5L�6��'5�{^�jjY?��L�'�P2�4��tU&S'
/g,RmEy�=����V�]p�4/�J���Ə����e��I���<*4Fm��q
�R-ۗ�_�ug�J+ss��Р�K������6t>��W����`��]-G���jt�+�������<͜��.z�3�ُ�+B�r#q񽵮��z�ɒ�� ���l�V��{cB�S��Q!�T�q�󒂏�,�U����� ��h���� 9sSi� �*�p�����A}j.������W�i�ߛ�.;�$ܺ^��Cq%D|0l������72'~5�P~(�*�1C�T���E��*�T�>�a<^g%sPlIu��d�y�Af~�iq���&��1�R�f�
�����r���x�yժ*�Jɭ��-[E
F,y�%������_�.�TIj_��!�хj��"���թQb����Ru�#^E�Y�Ӣ��dtu^��Dn"����v��/^a�PC��Xp�A<��T:�5[Y�{ƫ�l�0Ld��-��SnR�_vƹ�J���݅i�J������x}�c���Yh.J���W�4VC�*_��^��G�Uw���$]i��gi�l��A�묁_v��dEM3�Mc�iz<9���,�l�c�=����ݙ����'�y9���~�D��	�G�t���$�'ҫ�f�!c��� ]:����u����Te�K�$\���.|�� ��E�2q�&�]c��z s[���V�˲7=����'���Z�dH��
zx�ߊk1�B%+�?;�zey��q������v��v�X*���*8b��EԬ	-yJ��f�K`E��.L������_���V�_s���zN{���|/|.8K)AK@�s_�L���)h��{��C Y_���pH��_�U��.��������� �|y�����R^�Uğ�R�'��i&|X/<�����3�S~�Gӥ}������-<�;]��/���4��Z�d�Z��	���ʑ;�<�$v�n3Φ]��;u������W	��eN)�ۮYZ�n��6s���6*�ˌ�{A�&��������>O�\{?�^Zh|�5P#4��a.�����P���p>�����f���JW.�+#V����c��"ΏȤX�@㗍�#�J�J=����\]���nӌ��g�Š�����4�(X�闃�(�ʀq�Pp2�����UId�6�
�58��e�_Udqfݶk��C>z��l�>K@��L,/��΋2�b|J��/� Xsa
���^K��g�%�_�;!\?�%�Gufc�&X�&}��bk:I&���*W��c��%�<{��7��Y�tO��Nd��K��Z$��Ē��cQ�F� �-�t��{���O"Q;v2��ٸy�����;��4�Y�{}�3lf����MI������=N*Y�����.�ҖfB�K�M�x7&������Z a���ZK�8���u�ݗ��ѹ���P
������tR�ֱ�#n����	��AnRA�._ǂ�^�5g����of���Ly�,8��ˣ�OtX�I��g�'�lEwX�N�-��$TAFܮ���t*w|��[[�!�2Ι�b/�i�A���@g��u����������%B�����������-�(���9�,�"���xmb�X,����6ش�(���M Һe����_�!'c4���?+��������-���!�P>�{�!�#�TዔM2�3fP
�g�*�EM��m��m!�S�`|�r�C�j�}H�!���`	�n�[�M��Y6e��e�z��Һ�{�;�������1�o4u6y9G��&Hb��g��yɵ1�Uw�m~�!�5՝󰔾;E]��:p&����� "�Z��ـ!�D�'��g(]w�`"f#t/���.�[73�L�|[��,B�O���ҤN���D笑e���7��<"���~���+���hҵ��D�n鴜X֭Y2��c��6������V�%���b��]�Ŵ��e�I�<n��Ӓ����[a��c������ip�B�=I�$���3��ǂ#��������(-L韦GRؠ3�oń�}� +�� T���I���\ +uR��[��#�d��P;�ެ֛�͎s柁\सI��(�30�`y���:@�ܬ`j�Qy�>��gM��,m�g�o�y���GHK�w.�j?sS�R�T��p���s�M��7V^�`XO%G��S@���M<��d�d_M�-��nOmZ`V�Ӆ%�=�1��Q֛���<�55�-S��J��@��
��ܱ�I�����>5�-&�kM�}6�5�S�[F�n	Y�l���� ��$�:��;�������6�;��n��Ϸ�����&&*����-[2��6��R伢wn�S�o݀j�Q� (��oR�iK�E��1@5M����Woo���3���UFU�n�Z�V��| K"O6�]���v�Z��g�kf߆Co�����"�X���ӓ4u�����|J̝��]o�QFt5��?p� �L�I��
�6x|_��!R+���l��7PgMIp�%�|3�jɃ��r#�S�$�(��&�Ż�u����[Y�0��ѿf�#ӵ٨:�u��4��q���>$H�0��OUn�@�!�t͊2-Rkf0��L���� �C��#ܓ�؆�X־������ܜHM3;���DIB�Γ�]9�GU)�P�h�Cı��"rw��ޡ�f�v��]Uh��>�yҟX*����><q�y�^��K�Ɍ�>�'`#�y]P���o�����9�s��D_n٤2�VfM��pe��F��+�����:��*���������&O�e��*jk�7��6ش?v��D������W����NΣ$L�m`�>?�L?Dr:!���NfZdV}��0L�k��P�ޤ���������L^�^q|���0cj|$?�D����=����U@/�bq��r V������%�-x�[�E2�NṤ�<� ^ �I%w�s��?���ZI��;WY��W�9�T�q�BTp�������(#-�Z�H5�Ϲ�l#t�2m����l)� |w�8]_��*8OT��qB�ﵴ%W�Yߘ�F&ۛ%U�5�o��Ɓ W���.S�<��X�$[���\\��v�,�_�M<L'�CZ*�]X��/}�~4&]U�H(���"	��8���]<Ȑ@��KΊr�J�(�ۜ�0�4	i��N�\Aے3ZT{�Q�Y�z���{�!z��|��+������C���hkUp54)A� $ܽz�6����m�c/3Ղm�AჁ�J;ص+�<y��D̂@2M�������c�q��J������\A�S��G�m��RǗ�	ݜ��v�{u(_��qK
2P\�o�
Ig$V6�����q���{_��q����_C"b��z'K$��L������W��H."*/V<�XW�A�$��K��Љ���C\y�5%�.�f�g�X�׍}{.A�F$-I��G����W�%��'�:��,�؟��2���uD��>J���v�Bc���x�-!� �_�icm�Q@��o�ٜL=�=��W�k�E�=y�}WuEf�F�Ǳs�a���Y�!�[*�ML��+��6�9f&��K��<xA���8��>}1a��i�>8�8�d{f��A
��x��I����8�7�NR��� �{R��w^W���nR��;_�.t^}�ogdA��7kj���3�,����Gt<���ugy Cl�l��2(���*A*�@U�Ytk��)�?����6�}�/l6Ayf/����m����=�MK��	,r�F
��xyw��|�(�BB�=���0�mFY�,zV8��K6<(K(ܦ�Md�H�I�*���3�c����z��/w��E#Ƒ���P��l�V)�sL�1�3�9�K�0��qN�H�_;D!�͑`�XA�'�Bj�\��t���Q<n���M$��6�%���?ϩ^���6�1{p�/��횃��΄�I�6]�ĽHFk<gu�?�]�
1��n�Qw��RՁYu�"^�]�H8���I����� �9"s�:�=��(�U�(�][�8"ʒN/j�.4?7�������O1O}��[���Dˬ�e��7�|<�y���д�@���(2��Dm���X֑�6�2-}�����:� ��]V9�NZb"�멅/�ɗ(� g�7i@����_[ �����'�SpcT�=-?�:����$qF������� ���T���*LP�6���<���Ҕ�d�3��܎���L���{���8�!yw�`;ʩ���j�S��HG�g��n�`�M�K�6����������i{�m��������6��6 �B*��H�7�gX鐠��1��Tqo��U�D<۔E��]3衞�K��2����z"vD��������G�K\H]�\"�Uc/�1�.�;�7�m�CY1����OTp�9�3�ߜD_�e���7��:<騌�l���cN[A����D�W�黪�֔(���鞇(��]�7�V]��'rb��,�z��,-v��Ig�Z�H�u+�B���X㙹�V�_\pƜ�=�[��]�{�X��T���p�$z���fזR�G3L�M���+�gR����Ӗ�P��� �|<RO���<9�d/���AV����͕�h���(���^�04y���:�u����4Q���>�A�S��ۺg�y�� ���*K��A�q��S��GT��L����x��W7���`��N]�S'~������d澆-��4n�\�`}f��,�1�*Q��㺂�4��=�-il��V0�+O�	��Q��઺:Y2��u̔��k�]d]6�5�^�B�l�W�Y�n,�t0�B,	��7ϸD��/Ԧ�L ���n��l�>��1jE&q���2��仏�Y�i��n��S�~��{�gʄȖ=�iRM���n9@Ӣ_�#��jԕ��7�H�=�|h&���Z��,�CE6"�����VZ�Z,�gn3f�o����"�"�힇]�t4j�����|,�ҝ�|6o��1t��Z��{ %iI �`
�4�|�I6!Y�����`�Kֹ
�7׾FI�J�È���ۚ��#�w�$��I��v����u�^����0�n��@S#���E�u��4GR�h��>kK�0�/Uu���{��!Z����T�k�L���a�6���j�@�*��׿��X�今a�c�8ڜ�q�;	|K�k#����D���C�)��hE�d�-}�r�d���mBvz��U/Z�>UƲ����� ����Y��2S[/�2���f�>Q+�#|�7P\h�oLH��x�9�ו�+D|�&��� h��eN����%_��\o�ASS*�჉��u�,3
ӭ�Xe�"�*���72�6�F3?Ir�����gW>/`e=,�k�)L�7mgR6?n,D9A����U��:}˻���ZLEK����ދU�mۢ�`o�X�jr:�^�����j��]�+���4n�D=`��B`���.�f2} }�����6�i8x��=E��hSWͣ�  ��%~�U������mZ�N�;މ~;<{��1۟i���n���(�f�ZH�Q�V��l��w>��:&��sJj�߬�m��PT�8ֲ́�3ZB���L��Y��Ff0%��ܥ�o@��g���ZS��_a[�!Y\#���Lg�>I �:7?�c�hT�	�o�[^��,(N�$T�l �y5iw�vr�<h�f �*��תY=���#H�~��5lP����P@.�l�Ő8go�cŇ'��x��Xs�����=�u���6jlaT׿�F�0�U����RĢ��JX�����:\4v�	�ט�_��	.m�X�n�2:�6�n2@�)�Nv{�U[���i���|�Л@Mq����G�H��౗�H���1R�T �	���Fbmb�����O*Ǿ ��@����b��o(�
n���we]d��f�*�0�׷@<%��2�N��>���t�w��	|��2�ǷS'�@QCP'�����{)�`[��ț9�";C?a��Q��=��P�#>���h�+�d�,�X|޾�2Ý����DVY8S�Rٜ�+Q@�y��}��<�2pD�LF���8���]ӸWʚ�)Z*��R@sS������ׯi3�t�f�`%'��A3�?ܓ����CU���8#i9��sE~��P?1���pwX��42z�%��Pёc��~1�/]�Z�F����t���~t����}�Y
�?�qX͔�ÀFr��+�vRX�tgw0�ˠz�A�=���j�H&��a���mY��iJ������BO2$����+�]������m��2��(?��>��XG��G���M�U�5_����N��	�Tmum�G̈́Ly{�����7�!nҨ�}�Tʖf��1�r�1�59ڮ)��B��!�'1fDxN�,��r1a����p�ܽ����N`��|���ztb*��5�t�g9���^M�[�b���ޘ���8��-<����8�6f�bQS�C`Ձ���ꠧi��I_���nI0Ңb1t��`W�t�i�xz�g���A����忴o����@h�ȉ�ɹJ�[��S�a<�N$>=-�Z�ߋwZ7�B�/�[L8�=�c4�d��)S��N(��LG5k_p�"*X�c�� �4��-/RtJ�=�8�~>��p'/�qP��$a��1ʴ�C�0S�=_0�J�����LB��P���|a�/�Zܚ�~{\��$'��E�2��
�^Ci�_u�3��X�S�Yb�$�$k��ȶE��b�)~��:�����Wu76Y}��N�B����=�	���Q~,s�c�5����_i�ؐ�Hy��h�vS�PSH0ܢΥ9"e�P�؆v�dU/j`(���[2�I�q�㥬<�jD/�w->�vB��e ?=28\�A@%D�n��>w�V�0�
�Vy�X��Wbјss�WYvD%$0֌���1Հ���+� ��{*G��uY]Z^�"+ۊ(����3�5}4�I,���˟a������W@x�b �3؃e��[�t��Dk���N��@V�e!��ҩ�I1J����М{!G?j�SҮL���������\�h�YP�c����_�u�#K����
\�������9��Zx�%���^eF�G�>�I�����eOm�Nw=A�CIq����.`{�J���ԛ�PH���ZN�k�3�8�`R}����ϢLI�Y雩@ �9�?:"��V�uTQ���ز��h9�M�^:c �0�v5*�AByu��:��eG��F��O���k�g���g�E����S�\��}�O7=T�wܡ/�1����)����&\?Z&.���I���Hg��&� )��<n�4��)�9z�,����϶փ���[����~�����[6��x�N�ZU{�L���	�t(E1F5����a��j��K�h��4���ӝ<��~��'ܷ�=78�P'j
�<�Z��|m���uĄz��' ��P�Ns�f��X�D�W<a"�k�����։�c ���ۜk*tlZV�����'0D��O0�"xu�V�:k���sۆ�Mp(|kN�EB���x�d�}�
�%�i����\D���,�E)?�
U�R�5��e�6���fIҬ��7JD�����E�,*2Mc�捤$��.q��ɰ�x�2�O�t�U,%5;��6���6�����0W�#)@���p>������~J?���c�@���`���k�1@����{�Y��Ӄ�$�)X��Y%i�[��Q���[�������>yr�Dg�ʫ�:`KQJ���r,��r~_jH���+�ʯ:��ԟ�)`LR�+���zi$������"$��נـ�Y6a���"o�Ӕl�|9|&�"I�K����"OLB�a���޽43���[v\;h�<�����Ә�U ��UиH4�韄�;��-���׍�y�L�_�P'V��H��}m�A,��z9qE�ӯ��*��ci�3�簼�3'���3�pL2��N�k���'�xS���I��lԵ�ٛ�)WA�b����B�=�j�ِ��##���֟�moVwӷ�Jɔ
�1�f��&����&�����V�(;��h�${���U��D�Q9���Ҁ(�����ʴT��}&�}�ا6�	7�B�B��/����
���z�V}��VB$�(O�Nx��W�ܾ�JѢ
�q(o�/mֻvd��b���W�P�\��w�K��Q71k���\�dKj�	���wN���񚾲S��&�1�{2v�Mz�2���^F�a�����.�ƣ	!�ЙhI�9P��}L����)'��Mi�][��-�_�-&k����=B��R��	��r
�S;����G��>��|Ķ,�ɿ�v�@���r��V�K>#�".Q#����8�[�4,ݿ�)��f�k�w�Pc?o�R-Z�����f	q?�.^���=tX&�=�e2�/�:�%�k=d��P�}s��t�b�&"1
j�H8&%WT�?�L!M,�s
-��[+��6�Y�u8MamĎmvZ�8�ԥKd��qG���M��kd�M�hk�����Q2�'�����UZڥ�?d���G$����S4XݙUA��'��,-�~y.^#�c�+z¸��4���33 �
�̥ɕڎ9u�Myz%�FȻ��,[nR-���ax�P����aTs:�ؠ�����m���O�����[�	`�l2-�.F�-Ӂ�&_��ߠ���3���zU5�j�)Bh6#���ݯz����<`���=�VB�����_�T݃���Ӣ��wӽ��J���Дc���1� ��i��*�찜a �A�i2.��E��s�$��W���i��/���;����y}�C�RLDW��X/��zwj2�'��P9)��E�kC���͞�=�>TV)�\z�^�"]P'�,u����<�AA������Q������9��8�骱�b.�x�Wk�L��2���I[�]��7%��n�>l�	\�I�>��Ltр	Ԓ}�]I�;�l㯖]wruv77^�L��n9��_�x]��[�"6�5ff�͉;^�:�C+��p�v��C)���w[Y��ҫN�X0'�e�h���ښ�_���`�ƕ�ݠ��JF�������V�5�T3J���WM~:V^ _d�����Hi�wM�$X���¾ElV�Ӎ�S_���d �뱈-�(C9�N~���Pl���@#�.}Q�t���K�'��59��~O�� Ԋb��:e���O#߫K��Z��r` �D�����+��m�eS�$������.׬S ־�E�������>ٝz;'/[�k�QTղ�;x�D�E�B1v��Hq�jz�<��%0�=[�+U��5������J��̦�ܞ�X�NZ��Mzb`��g׃ye!�fpt�E��E.��֏Og��Z�2�0�sJm����S{q�|
�.s���q@��Y_h�
���0)�X{�� 4�����o�U�P�	�X�U��	���eydD��.�U��9U����#�'��p&���/�⥰�j���Gn�����`�W��<��]M/?4�~9��x/��`�	�����<�4w�%V�!���uv�2T�g7�	���N�h��i��ZaI㱨K��ɖ{�
�ǌ�"���d��wX���!h�V5����WT	��
��S�D!�����x���J��Q+�������7S������[�C������J��ӯ&�I\XoH��.̤D.(ŻS6�MB,����/(���q���2GG)�F�}I�*6C�Nt��M�_��qؗ��7�C�V�
9K��0LI�	N��LlyEm/My�X.�+��K�Kt>�� jv��\��%�O�f���X���}2LQ���@I�ղe/i��x�%���1j����?������<���2����OW�čg�c�-�t	B-ؔ����)��VQvd���Ǜٳ���O^�m�" ��B�}�q�f��K��i���y>���3�*t�m�4�����f}��K-�Ax2%C���ça�����O�8��fҿ�x���̃w�@Zp�s��R'i��wb��ע��)����R��_�B�^4gog�s2�JP�����E�,3)���#t�U�dig0l *���1�&\�AA�LL�t�L��F��?o�����E/Q�A����h�`��w�������`�<�}����GJ��	(m� ���'��F��dm��,���A63�(�=\MQܺ��,^�5�\]�c�ey�ԖѺv��ǩ�\�HkϜܢP��\���/��HTm3����"�`qdϙ���!ƿ`\.�>�j�	��ܿ%�{�nGN_M��6@�r�)�˩uFh�-ri{G�]��{��wU�J! 6��/>U H]#�glc��4��1�:���h�@a�؆O�Y6�]�'S��}��b�����h"
.M���h�`W�_�K]r��"�[/A��.�N7��WI��g�FOh��͈y��v D�{e�L�7�]�<�l։ 3j�wg&�|��oDD�Z��-��(����o��:�q���h7V0���~b�2��@���@�͞w8��n�+��Xf�V@��kqe������p�ܜ=����qCH���&h2
���{�#���z�KR��3` ���Ê{P,�H�|��#��/½ e~R�|v�Pv>d�f������Nͩ�,���뤓�T�c��0H!y�:���TQ�&�>z8(�gn�g*�Zy�پ��KV�:ʅ=SzbT� ���x��H��7�D`�b��S���(�ڥ��d�K�-��n�~X`˓�@���|Q�⑺_��О8-��w�Ln����%�4!��$�]��;A�a�(�Ik�'��B�5��|�3H�GY7� 9��W3����c��Ȣ��;"ޅ>n"'��Rh����[&�ѳ���2�;0�#��}��nN^S��eO6�{v�*Fifh߻L��@���+Vn��ﮕ�c�\��Ź�,��Z&p	�WI�"��,�Hȕ���Z@��g�Tf��Mo������"*��q*�4��j�*S4|�ޔ��9o�t�_�z� 9II��@
 �h|��!mBZm�h�tX��M�v7�PIk�����W%t�.� #=�$�,�aMۻ�V=��P��C�0�����S1#NF��mhu&6<4[�8���(>]M0��$U�q���!!n�ЊmӾk���G� �J���jU�>�x�S�bX�������]S�C9�;6�����|��؏F���).�hY����2r���A@{����v|UC�[>�@���<��������4��+�`���H�zq>���#���P�+/o`~���p�9��Ƌ����F�ݑC�3�
e��1�0y�_�ʽU2*i�����������>�e��*ŭ<7ƌ�6��?�^�����0�WRL�����pL���m{��?��DMݍ�Q���+{_϶�$�Lٓ��l��潁K���l}���^�?��_�j�*:�U��x������%�]���z` �������x���EmE|�^�7�� ��b%����2�0��Y�Z���;��[�R� ����#t�xn�F�(�&�Z�}��j��l��R�H��3Շɝ��q�����j�8��l?<B߉̴�<�Y�5�F��%0d�p�oT{܁�\��nY{S����s6�[)+�\7�B<����E ;��?��h�� 	�j'[�<@�@8@��fl405�~v�� hn�c�>n��k\�YQ��·�3���5 ��	�G�����Nh��L����'��^Գ� s�k�^*=�r��J�ta��٠Zw����	+X۶�^����5��N��v[l�׬T��`a�.����a�:�U��4&�=�v��[��������/!�q�ó�'H/�t�K�\9�213�h��Н��Z)sb{��'��*[0�%<�Q�b��no�2n�^kw�Z��
a*�o��뼕<���Fl��]����w��|�Y�[�U;^�Q�K��#w�?�)3Ta� R���޶��?u�wQ6O����#���|(�+L^�,����R�wñ9b�E�oj3�8�ƴٰ V+�A���k}���<���ج[F���8=�9]�wh�.�=)n�f�n�s#4�/�����C�;�$/���`9���~���S�'�.*�CiD�����MNJ����ͩ1?��p��Q�4(fz��3�xБw��~��]۪tF�,৭�{�����m�x�
�N��Jw���hFR�+���XswD��dA� �����\[�:����m��},+�L3����:2�\`�$��������m��82�9N?;��>	S�Gl�$�ׄ���_,яP����T�9�u�!GaƆL��W���K�!�B�(ۢT^�)�+ Y�,?�I������VE�!1gwfX�\���rEh1�.�4���Ϯ)���b���$�ߎz;��I�����ǀ���MFNv�,�r������-PO5��_��J*�b噂Ct3��КӘ˧���]��MT�0�:�b�N�tDti����+�����U���*%��a�V��@|���?��J�Ǽ�k�aP;N�˼-(�i"%wn�щV�6�*Y	[���Q�c��=d�����b~C(qyGIip���>+�c
��H�
��&t^&_=h~R�ep�CA�,bDka�I�H>S�Dd�=�c[^?�zQ�"U��o�dp[���/-Ӌ�._�{p�$�mgE�]d99��Xi�F7����)�m�d$=5&��9�ٜR�v~��s��N��뤩6m���o�pB������q���~�~cӖ6���ϯs_8�$ty�Uq�
��Pg���vܶ<����K�d���q�x�j�����[2�����@hIjX�nw��vVKX`�7 S�;2��ߗU�Dd�>�R���ꟺ���!���P�,R--lMY
�8v��T��1雅k?��4]�N�G�lEY���+o琪��#3Ko4�MX�3w�˳�4��7��N@��vå3l����3���cD�T���N�e@��Ge5�=�=1�1^-��_��{5H��������xa���d��*�h�ٮ�������^�	G�K���q���&2��ԛ9@{�x�������r���ۈ1�][�lS�ec�!Nh*�W��f�Br�����C�4����N�B3��`��o��cK6I��=#6 �������{Mu�Ӷْ>�)e<�ag�:�y��D��\��U;�u+�:��G�9FBKO3���M��t�g�cc	��g�\�TC}�D�O�P�T����aK��n-)�h����\�R�B
���xW�i��v�0�)L�n�>��?jz�(���1���j��Ĥ|ȳc�璮9+�E�o����b��UNs`�Rݝ��<�@�%�5�="� $0�|�j66�K�Y������#��7�z���I�D�O8��Wj�O{�n��|��W�=����Wq���Ǽ�"�	��@H�0ˑwR7���:� i�VV�O�5@R�x�Z������"Fc����ZkWd�l'L�.Hz���0�/�O}Sxbx����k0��@N��<"|x��E�ݪ��x���
�*
��Eia�u��-���C�E�7�
���?����Cƽ��l����x7W��IQ�<Q�,��M����$z�*q�B�Ξ�ߞ���כ,GB�Z���x���N��F?�0w0�f�j>I���̭;J�;'Ӑ��ԍ���as�k�<�����}��	_�(�,�Q��X�@[%�x�� h.�X���P������Eer��ї��:��TW���S;Xr�X��~�d�����%�:N{��k�L�Q�N��g���<v�촍���<��ŘX'a-��"�� �Y�H9�9W&ґ}��X�vOY�Ya�@Ŧ+�e3����p�;:�[<d���Yӥ�t �T����H!���,��;�3�M2��a��L��9^HHV�YH�H�ms��<�y9>�$�@���7��A���f������ؖ�HpWS�`��x:�ԯ�S�~�6���5�3���A1�H�������&u0��j�3��=m۱:V�g���Q�Av�~����1�u9v�S�����V�o;&�dhI��j����1Q��w��)�(|�|�\Y۴aY�}ӫ�%�۰�^w�Ϛ[B&��TT�
$O�8}�NdBq�O��|N�W�����
,��o�$3�]��؏dva�%c�W�>D\�yĩ����,�1�� /�d8��	H����Cթ"��v��R1W�v@���z�q5N�	�a�T��e�v��F_����ө����V����:]�=S:�0�X &��3���=���E	�p\rw��SH^��k�����·�ⶹx��+��@��}rg`d�X���;�#&�E�%�����s�F�3f�S�Pp�R���yZK����0q̧y^��t=蒃&+̇r8W�ܽi�r֙k*˚��js�ƀt���&�Fwu�8�JCW�u"�PG!ڭ9s7���(D�ţ���M�ގ�-ŀ%\���=ZIhq����:��x�oM�G�֙p��I�-�'���dh%���?q˳��_��2�4E�QU��'�N�,���y����p��������4�0�����7�p�����N�Z���Fg��pPR�G��?e3�j���$�sG ���O��+��቞�	ۈeh`�sm-���:������,F���&�<�z���78�Bne�#p��V�z0�����ʆr�������WB.�����T��m�:s��� ��Jxn���h�0m��9T �AQi@�O*0�L�N&	A%M&.)������N�W�}i7��'o�;yz���WC�!D$�Z�Š�ۇ���'&��P&���
�CJ��ȕ�G��;Tc�C	X�^��P�u�.��+)BA#���w�)jut&N��Qﲷ;�v�(���xqF������_4����[����n@%7�V�4�V���+I�j���=�-�ϒ� �6���4�����uC X^�N2�{���0A��_�H�"ç~�b�)���j^	Z�C8�wp�%=���W�݅#Yw���{�[0���������I��jT�a긳@Y�-�yJE`v�T=�%��/`���J5y�W:�2V�a_����Ԅ��JwZ3�$�K�::lC�W��GT_�d�1�����)�9�q����l�q�> �[.��A�Ƹ�!'��a9R>�~�e#�?V������ILƼ� �Xe��6��j� �9���t?��>eq=I$�����.$: ��E*mĲ�8'�z�.[�`����ߧ˿1����U���H>�z a��2≌�N�+� ��";�C���G'���ӷ�Ҋ&Э�/�|����'�G'��kPߓP2?<���]HSx/m3�4�l�8������	�0��S<<�G��3�z:m�:^���K�� ">	Y�-N}��ۂ��ZD ��
/�Im���{��������`��ω>�� �ۭGh[�55$������j����c�]O����]�@�s��J+W�+w���u?s�0�ӏ�����a�5wa�Jsկ�Rn\1����OO�]n�������|�Y�k�[(O6Lqo&�2@Q֤_��IWYB6��S��>��I�_���q��(��*;C�f����K��L��;�����;݀/FUXG$3�
�K����y�]��\i�.%���f�p%X���}k3��6ǃIz�r������T�%�b��*���C��Ȕ��"T�e5~�.Yp�s�f��c����*-΂�OSNQ?�_��ٌ�C�
�wN��[z��-�j}GF>fr5�ǡ@����?r�1��,*�:���R�&��f�oK�Xcx������.T2a�6��.�W8NAk51�1�͍��Z�9�����Y�'��R��^��q�B���g�����$R�,�_��^mm�gTA{����ZX����,����0�t,vC����gi#9l��U�"�����A�nEBKt��О�/�q�uY�m�\/
��Aiq�������m�	��w@+=�����<�6g��ht����(���-Gr ����m6��,j����6�6,q�(�lMT$�9�p�P���c�-<��U�oh��cƁ	M��_�P��X����稠�!��3�4��;����7���U�O\
!�`�u�VXj�uk�����f�n�c�M�(6�T��L��N`��&�@{`�����sd��J�6M����H6�ge���M�j1��уA�8u�F�qh�KJ]��i�����{�l���"c�-���˟���]Ke�"�k�/Z	�.	N7P�Э�� ߸O!����6��o�D��	ehD7���<v:����~�0w�����	Q�D]��r�ց��"�x���j�*<��8V)�^��b������8~��p�'��s��O����������I�pS�M=���*N]��9�aό��2R�␊�hs��\VR�!�3��X�Ɗt֔�a����%���� ?;R|�η	ӛd�Z���ݬ��c���U���(��O�0$yb��:�sD�4]�Q�`�>Ӡ���� ��g�Fdyi���D$Ko�rʾ�HS��2T �DQ����G!�7�n�`,j��SS�ءVۥ8Qd�L-[	ln���`*=Ӆy?3�UaQ*���5��H@-��t�H�؂��^��z$i����g��be��8�k�_
�5/�/"$ŠYЍ�A��ʠ��}�|�=��ꦔY��`�n��N�*�%�&~6t��,�2۔\�|Vż��xn�X�S��7�>T��t�x�C�di��	���r@`�����̫�Q�`�d�U�	�)mf�eo,Z���Ц"#��j���l�Z9b�g��Of3��o�H��+��"�]>�*s4���#�l|٘؝��ox��t����	k ��AIm$X
�e|3e2!�hwƣ*������4i7�.�IDzɎ��>@ۚg�#�ϲ$=��}�X�l����Y�0˵~��]#��B��דu���4����d�>x\�0�bBU���h�/!璗�`k�3k� "��CÙ�R��wi׬��X*�{���%�b�ϜO�;)� p*�1��o�)�aho���w�r����Z9��RvgqU��
>�=��K�Y8>�����M�wd���ٌ�>~`<#I��Pɜ�oY
*��{A9�Py���-'��*3��lKe�0��
�}�x�]���*�!��m.��Y"c�z��e��*�7ߩ&6,�q?�%��@l���W����x�vL��#m�¥?[��D�����7�Т	�8d-�H�L��V�>~'�xlݽ�� ����%��C^�X��̗j�e6�F��f
�q����ϸ6�v�sb� *�áLG���Ux;VEDv5����� �o%�3K���w�c�Zl�;�L��+Y��ۏ�wQ�P.����(wO�Zu�ӿ#�Bl�aK_���n����0��7q�����}+i8�o�E�hB�/�����Y3>`F�*.%�^i	Zko�ށ�p��g�S��Ҭg�[��\�P��=�y�� ��?�Fhh�	�q[K�����Ql��5�$�v�h�#�w���F�Y����P�A�KZ|5�3�ӎ�Y/�e��Hs�Ž��'���Ԍ�#s��w��==�U��9��aa��g�A��ת�qv ���'�����,�v��R�eǸ�9+�.z�:�|�[B�Ķ�v���[�*D�a�������H�!qE�c��H���N%��D����a��жn����bn/��]�*�7j\����ub͑�o��n� �wRD!��+R*Ï��<�n��?�v���)�_ww�|iך�����Q�i����X��)lHhM|7�Uڜ�OK?.�Q����#�󇢵E�+�"[,-�������jK���oc��8 ����FH+>�|�`}8��<�B����F��8V��] ��ʇ�x)�����sܗ��
(��!�\��]�p�S�Z`�8�����|���CbcO����Y�`w���m1���pD����z��F�D����~O-]TMFħfxO�T�i��㡋*��
�a��^����F�Ư+���XL�w=ͽ�'�MA�\	��s`�Lg�����nm�Y�v�+�eU��_x2iJ��_��y����m�x�2���?T�>B�KG�/��P�l���(_��5�v���(�T�m6uR�G�d�LY͙+�>�z�!��m�!Y2Tw���d��_���S:�V�Z��!
S fQ#��aKr~q-��Ǳ�i��9��Ϡ��؀߇��A!���Q����9�M߁/���K�o�$x�0�-����
"B��7�b~VYC-����_H�̺L��:���fg��_*0_�~b^T��-=�tB	��H��ݎ���sŴ�@l@59���~J�W���wa�lNi�-�_�zyw'��/s��#6�[� sڊMc!��d0��Vʨ�r�(���GB/ p�=�wS�cr9B��ā�Z��t�=AL�~K1gp��x�ei�t��aZ��0f���4=�`�Wי��[�m�����\�ʩo9/��_�%{i�X$�BE;%��C<c�i"K&�Ճe��$�fy$V�����2�����~O�߯�X����6f�MÈe�B��*r�f~Y-c��Ȑt���l���=/5y�s��cf}P��"F�:�o�����]���3�=��;�jM���`�/2���>��	jQ�$w�k�v����S� �'�2e�:��D=j�K��v֭W��fu��9��Ō���Y�\e1V�m�o1"^Z�Hl��5k��G���Yʏ2��|+��ߪ�O3�Y4�+�����l�e�a��6@%����A3�D��n:�����D8W�|dN�Px@�en�bҖ�1ל��]#{�y��.�һf�ߑd��3˥��W5h*�蚐n*���p��xJK�i�����3�����9��xf;�p�X�k�z����������e�?N�aů�y�?��;�U����P����"T�#��N�l&3�_�`�}>
��|r�I�R��t� md��l��p��u�n�ң�B�?͚�*:PD��r<���c�u<�:��G�rhFH��O��V���0,�og�4Z��f�`�\���}�ɨO	}�T6{��\�V��)n����\��{���6�I�z���߄�))%Rxn��z�֓�z��l��f0��h�}pwȌ�+�LD����~ؕ��ۭrU���Y��v�w5Nt�)57gS�yt���j� �K�w�ݡ�>����P6L���H���987�tj7�0�'g=|}r���4�1���L�W��}�\P(	P��H��~���(R0�L�S3i���V{{5��`�)M1���z�~��MOc&.��X�Zk�؉l�K��6��l�0�(�Ov�x{����k�Hy𹶚�S��|1$E��|��xhb�Cǧ
�fi�l��b.{��W�E��?
�u0XO:n\T�x#���J:��x��zaT��V�'���aP�w�D��_����᫇' �Q�i��.*8�۲�ARk�.�� "O���Y6W`�	i��r���;D��3��C��ED��
��h��4�[,�'��P��\����C���ZΕ��_T��VTY^�;�P�2?u������A{�&��׋�������t��?8��U�\��x���Ɗ��@���zV[ڪ�a,�%d��9��C�I��n��z񣒷}*ë��&�S�W̉u�+9^��4�($��Y ��������"��G�/�#^��C���p� �}D��j�vY��^�H�^0a-������̅�TB�NQ��@�j�Z��J������2��V��N�7J"J WǴ�V"\_^���T��L�wB�$R�V����l�ͬ���N_��VdZ�-�����9�R$��
�l��kz7�(��ݮ� �ţ�'ay�9��~�{墊\u�����ɔ�����W)� �z���)���m�/2!e~�$�B7���.�� P7�EW~���o�x7�z�L�[G@��K�<��&Ϳ�&8��Ҳ��X�H��Vz-<\��܌7!&+�`ԯ�9���|�D0A���_VxXW���mb<���ݯy��fj�E.�5�	��TB���s�M���o{XA|D�t.�7�Q@��"_���)�~)=]{��* nM}͉!�)'U�2C��ϡX��8e�w�y�>��8Uç�U�v��l'&.�&Q�C/�ג��*����G(w��S���9<��D]�]�/�@4׬J�nf���	����&{�<W��C�������=��#��!�q	z1�N��Z��xZ��㫫�
~Ӗ��n{��=��|��\�E�0;ّ1��|;Th�52�G���O��坈����f���`��4U�J"�+x����F��qv���jv������8AJT#����)\Rm-��P���D�uGߗG��=�a�LA^(P?�q�O�2��L���I���6=|fJث���_�]�q��� )GCso��A2�K��RLA������W?(/��X��K����Kn�h�:x��o>\jB�%�f�пXg�}짊��˥I;ղߨN��!,%����k)N�D}��I�~��i4�&�ɲ[5	�ć��c憈�o-�$i��-�I�Q𑆐`��٭Vy�K���)i������#%}r?fS�Ǣ`�����t�rh�*.K׳.ז��zf���K���x,M�!�]����aj`����8��{L{��2����z��h娜`R!X:��0�#m7�hn-���R�c�_�H^�x�g��c脸�;@���F,-_��8�t�f���Qg
��lZ�� &���[A;����Gt_�nQ�?�<��6�T�N8�/��A����E��&U���o�@�.g�څx�7�����{�+�b(��ɮ��c��4�m��,kK��R6m�(-B�M�䆺ڥ)�5Ԃ�1   N   Ĵ���	��Z��wI�+ʜ�cd�<��k٥���qe�H�4͔6Z"<ɑ�i�6�3{�\2V��<d���fJ>@,o�$�M3P�i����d��f���{�9ݖ<Z"��5�����@�MC7����O�5��4_@�,F�@�x�cB�c���'��l�������.O8kq��8 �"/O�!�k޿q��	QǊ o"��>�P�޴4.��O,�Ӧb���u%MHy�A�{<:1aO�)1[�A�΀�H��(]��'�n�	B+�C�'K���=�XUs���X%�h u�c��'���ቨr_�'|P
�g�=-T�8�F�.��Dڝ'�!Dx�_�'k<|ku�ʣ,6��À��+;��@a�5f(�"<���>�1���"�D g.m� i�d�i��Ѡ�O�8�{2`S�`z
��1EDx��9�M��0�2^|"<�G&��\ᔰU䄎׸-�iγ
m�I�>a�L=�2�`�F;� ����*}�H��ӭ-XU�'U�]Dx2�JA�`��9�e�QJg�%�=�.!�?<"<��O���`��3+�����_�* �)��@�O �L<Y1N��=LdY����`�e�ÉMd?�%+=�B���<�1��UVU���'HD�8#��ʟt�O������*1�n�q���y��5jb�
ED^'�U
D*��d?h@$,Pi����$��xr�x�ݠp_�Xh 6'V�h˃�&����$���u� ��G"�E�P�-�W����u厭-��P��̜��y� @� d  �                                                                                                                                                                                                                                                                                                                                                                                                                                                                      �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   
    �     �(  g1  �7  �=  CD  �J  �P  	W  _]  �c  �i  (p  lv  �|  ��   `� u�	����Zv)C�'ll\�0�Ez+�'N�Dl�^T�9O��Q�'��(�bE�f��
լ�( h�n��%�~�#�)�t�6��7�5b�ͱ�~�e�E��?i�Ǉ�?�K����D�Ιx5 Zce� ۲l�.q���`֨S����� .:��թ���uB� ��t�'�:�+U��ڰЩ�̀��հ�.ءD�0�Ă�O��v��$|�#�ѦX�D�<��ܟ���ӟ�J$��E����Ɵ6bx�4��՟��I�M�1��0����O�柆�d�OX1af+�;�,�+!*�06N�O�Ġ<y��?���|���'@�͙p�rP�U��*l�lJ��ԋAE!�_55"��f J�82�	��oε^��	�<I>��'+��^a�$�Id����DC�	=B�14B1�?Q��?���?A���?i���'I�,��"�|���v-��;����[(��ep��=oړ�M���K!��"vӰoZ�M��B�YHE��X`Iy�	ε2��!q�II>��V�ǜ ��˕�~��g$��j~)b �XVؠ�[ܦŋڴH���O{�)م#�҉(�!V�<��i3V�)�V�A$��kL	cUV4�b��q�84K2�T,<�8V���)`7�Ħ-Rݴ\�Du��<F��8❢B�>j!B7if8ċ��ގ_&��B~�*�l����zo�9��+��P3:���
2ĝ�~<4ys�����-#˞)qg)���yb4`u�rnژ�M��i͇&�5:��_�|7Hy�'�;�@}��k[�!
(�A�hG�a/�!0�i\PC3��1L*Ѐ�����'��O8��C��C5��Q���]���I�A�O������(d���M�Ο�HJѡd�
��O�^Кy�4�'�I��D����p���$u�ĸ���Q&�+�1�jU�UE�.z,%S`�V�3f��	=��Ƞ`�#�P5�2�B����%"��.��ZH���	��O,O|q��'����8G�T�O�� :#

/3J�����OL���O�㟢|�'|>������'5���D�Q�����T)jL���H�"�q	�&~�j���h��eV�)G�D3�nM�Vo(hᐅ���/��8�f"O��0KP�Z�B]0��3L]JP�@"O~��e�O*� IR��/T�y�w"O
9s�Z�8����r�Дb9�""OHa([z٢%�T�;��2@"O4��ǁ\�C�X	�\�k�'����`:�S�O����O�3�����y[T�1	�!�גNhXBSF+�ř"�
 p�!�d��H�	Dޞ��L�Rh�p�!��Q�l�P�R��-I�z(���J�b�!�$��j�P���.V?J5�򀅆�!�	y�L a�!A�65���1$��I8{���D6W�<���Gv�~X�D� �!�dF�J}P�A`��"E����@M9�!��=YQ��	2���?)ڱ`w�Մ�!�$*�Vt��F*F�~���郇�!�D�'X�J��'J��r�(��}l�y҃�u�7�1?�Ǆ�ߞ0�� i>I�`m�ϟ�'2�'_b���86I��
x�$ܚ#�O� ��+�Xk�5�p�qlv4�b�'1�}���J�T4ڰ��D-��)�\��e��oJpzgN�	�0<��j�ԟZڴX��'V�-#E��C�D�p�
?^�&@XP�P��s�S�O8|1��U�9���PQBܭh(
���}��D\�N��-{%I�q�195/��?�H>�5O��:��|Γ�y�,ǋH�@��]��AD���y���Q�Ӌ\~�0���.�yBΛ9L�ڥ��kͿuJ8ȉ��-�y��������Ǐo����D�3�yB@[/�%�,�`:Eaԩ���yB� %2A���H�^d�y���u)�f�'�B�'�<� �O��3�'�b�'���##��� �>H�>��NU�/��[q�?���#���#���h!]>���i��'�~���/�L� ����Y�r���k�.܆��'-ޥ��Ejg���m��)������h�L�󮏲8e<�P�$�6�`�:��?s�6�ey2�ՙ�?�����?	�#�%h�XZ� �c�h�,�sϓ8^�O$�#]�6 y�L�T&hy��]�${�4f�V�|�O���Q��
�D�i<������}?.9��Q�O[��]�`��ˉt>���,	2���h�#�1=��C�	)�����ܸR�����L����#����n}P�sg�@�}Y�Իr����z����e��U����P?)
�b6D�L�`�! �LH83�����};Ѐ/�DNĦy'�̉������O�h�ߞ-���k7�N�sZ�]5��O��ā�
s��d�O��
��H�3�¹c~�cv��M� �L�R�ˎ����F�50��+��'��!�H�\�0��U�5T6�)f ��@����xy!F�aaxr� ��?A���dЛV�I�AD� a*���qb�s��'?"�'���!�ٕ�pЊ���<9��EK���8�l���ӆp��1�Co��?A)OFl�B
N��Q�IҟԗO2�-��'| <���<aHe-�j[j!�F�'��۞m��h�Wc�M0ʄpwW̦�'��i�&D�Pa��BB�fe��:儍&8�I1���v�G���ǯ���H��l�#(	7` ��gkx0�����ra��O���/ڧ�?9��@�|"��b�
�� �+�y�%U&r�xk�i�76�A`p� ���O6�E�Tj��`� (x��9Jl\�a@N�����'���3�����	��x�'�<%(TI�:R`��E�0j���Z��@F��:<��d��L#�p����Ds��� 3ցY:H
 �fy ���l����s�'M��I��!��Ϙ'�|�:G ��0_��a��M�d�r$R����������'�ў�����~^���f</#�q��AM�<��\8Oͤ�@g�uId�i��My��?��|:����D�zijؙ+4�T�%���V��Ĉ�ƦM�Iӟ���Ny����?|��ٹ�I�$HoL�@��C�ę������� 	4B����ڝ1�6@����w(4�J)Lx�*㏎�j���G;(�n��dN�j��)[w��gH�AR�b���,0��'E��^�'ћV�M>Q�,�2�b^�P�|�"Ox8B6O��`�)R�̃-�DT1��|�CsӶ���<I��Ø��O���ӍU'#�@��蝗a�l�������O����O�4���!g�Ҝ{6aT�ki���FJ��m�=]�4�efK�x�L��d�>R0Q��fզ:�@���O�L��B%��Pn1;�&�c�'.9 ���?��OT�,Ш�U"�P.I���ԓ|��'����	���� G�C��1�	�e����5��0�jS"	�N0X��6�?!(O0��qG�On��&ʧ�?��[�:*�P1�T|�>h�@���?��3��(��&l���!W�	]��)؃T�<[4�"Cd��3"F���ər~TtK�ɕ@�r�C�I�Ok�A(����v$z�L��Lp��O��H��'����<�7Ddת�'��� �P(#��b�<ᧉ��.l��(ʀJ�Pի�C�S�'9D�}�7��/>f��:1��9��b��M���?I�f&`�Iao��?���?����y�:���˳.��n��](`�G�r��V'�@7�٧2j�@r��D�1V����)?�(�0 ��|���+w��u�uo�10e�pr��9�3�	�^�ꀸDcXm�X�Q�ev��$"?�f�Zڟ��	؟x�?��/��s����c�'����r/�2�y�N�xw$�E���FU�1�V���j�����'e�ɺH��y8w	��G��`�!�1
q)���M���?1����8��K���T��J�M���zSIU�6@��Q�G�2��`J�)��sϓx ���b��P�e3w'=Y��LB5䚄mK� #b�-�M�T�'ؒ�	��^�J�ԓS(ȢC�@� �!� �?��i^O��O��� ֍;�����K38*,Q�W�<�g�v3�賆Aٓ{vđ:&l@R�	,�M+���'[p���O7$ t��[=L����PͲ	�'�T���3h�� �c��zM���'*���7�X����a����'�T	���hD P��䋸G���	�'�`�+ �"s��MI�[�o�$(��'���Ț���H�Nõj�\#��dǾC^Q?sg��>⒔za��=+t�:�m8D�p@�̟d�d�7��Wl�3ä D��h���F�J)���Y�,t��n3D�H����;���w.��N�2� 2D��[Ԇ���a�ǥ@�!j����
;D�����;N�G$�*p�����O��F�)�'��a��쐆`\䚧Nj�=[�n2D���@>�ma�L^>�(P2��.D��@�]�A�@%�c\�����,D��#wh��Q�^h�B�1T/T�� �>D�$�mR�p�����&WJa�o!D��*���-<�|�w'�o��<m� B8�X�+�!CbQ��@-b��Z�d:D�� �����P�����_�+�<!rp"O�D��?�n`�'N.W��K�"O<}·�ܫ{I�- �%�:j�thf"OĔRc�E!ĴXd��>�|�S%�'S�]��'���!`�](<��JՠJ�X�
�'s4�6��9�t,b�5D��$	�'�IYv!	o��C4 9�,�y�'o~5:��G|��!�d��-��`�'J�jAӗE�����G�2z����'v&�ң/Z>6�H"[5&������dM"6@Q?�bi� 8�k�̶/_\�X�0D�$�OڝW���vF�':�41��!D�4��!�P�ݡץj��1�f>D��` ˘�� AA#�,<��C<D�`٥�ՙ<��)������xh�"8D�t�ү�F<f<�` ����'��O�D�3�)�BYiQTJ��k���$0��Y�'��l�U�>��ђ�m\-q�Y`�'�������]͖���͘V��D��'���@�ȧk=b���I�H�L ��'�� �WEX7�
��F�;Of|�	�'#�e�w�XL��e�$��q)O���'�'�vj�-�)D`qs6�Ƣ0~ؐ��'��l��GT�j�n���*ߠ{l�\b�'�,��smV�ekFB
��s��P
�'IhGoG�h�����,�>`ntc�'�6p�v�\(|��NWT���(�&��QԂ|Ӈ/ �^IT��DȄ�"f�مȓ��5x�˛0ޮ��0͞1VF����{� `�	�YzA��F�*2����t�*��ܱ|G�t�vm�PO�!��#y��ǧ��:� ��O�$�"��ȓI�6���F�jVn�9PԘO;P�G{�����!x1H�,�x�P���3`,�,��"O\�qw)��}[��C�╊`"O�)��[��#�(B�^��`�"O�:�@eX�i"�EF0�0D�"O�����r�����6G_j9�"Of�#"��2�A���iW�D���'�̵Ҍ����h�%S�H��Pۢ�[?�0���Բ6a׷6���e�����ȓfΒq"1��q̉�%
�SN����IzR!svN� +k���B�8�L��0;   �U.I� [1Wz�ȓ-�$p hX)��(+C�(JO�`�'Z�����ɋ%���04;�+�W�M��$GxU
�խ,WfHI���(.%�ȓ�(ԩ#	D�C2<epC�K����_֔�k0KV*V:�$�5����ȓp�P�bY�n�p��g�ɕj�����	*�	Ss�(�!��W&ށ���t_�C�I�E�̭�f� ���X#��D�ZC�*8�D[a��Ki�hУY
�4C�	�
����D��×K>B䉐y�b�0

�@Un|���#2^C�I�G�Jy�FW
0A�����O��D�=�Z,�~�#��[�j�;��`JPڤ�S]�<���&�zXPo�Pa�3P�Y�<qS�ɣ&���R&G�<6$���jV�<�f��l�V�3��M:\^�Q���\O�<a���H��1HE����6��N�<a����!xW	�2���Z�j\ǟ$���"�S�O6h�!lN��d�,Ϸ{�6��E"O5J2�H n�b��*�y(\�"O� X�[7��(D�cjЀ.a�}��"Ot���e���x ���.JU
٠"Of�$&�^���"�ǖ)_>v�؇"OP�h�~��i�[8�̓qW��#��+�Ov�22��+�V0k���14�u�"O���Ƃ
mF�`@�,���q"O�X�1EF�M�qc�%�m)	�e"O"<���R���:���}7�Q �"OB��E��5q�nP�HU("P t�'�ܭ��'�!����b��Z�Hc��6D�(�m�?8�`��%O>!o��Abg9D��aOH-�c�@��$��4D����D�%���H�͍7?���AӠ>D��Q�4���"+0�\��>D����Ϙ�-y��� ��Ytq��!ړ{N D����ig���7�T��|�!F�.�y���+��P�T�����D3�ym��5.4�2��&��G�U��y2ID�H(c3*N��G���y��6,r�ؐ���Hޠ����7�y�$V�.�;7�BFԨ���H��?���A����X� $h�Yȍ��A��	�Bi�&�3D�h�6#6.,��Jk�\���3D��z`(!% �B���:o� 8QN7D��`R�Tq܎$h4�Q�*���.:D�K�BȤEd҅bb�ɮW�*�(.�!��[3uѕ��)�V�#*Թ@S創TX����S0u�μ��M�	�&Q����"@!��IB�98PLR�M�r��d�"BC!�$͸p�s@�S6ԞpB��u%!�$�'��<�"�R1T�̅�q
�'/!�D�A����EڝcԦy�GcSc"�}�����~�ޮ]��I�H��dRQ��7�y2���=0��Q�r��4����y"i��'��T�à��X�4�q��y�Ή/w����O��L��eA�n�<�y".�n쐨K�׎L}℩�d��yB$XNȒ�Z�I�I+�Ւ�j��hO8����SLi�v���a.u��k�T��C�I
&*|�7���f���#4�LC�Ip~���7Fү�$���[�KDC�	�	�ڌ㰏	*]�mA+��#K�C��5~> �F�E�  ׄ�2!9$B�I�*�ec��Ǜ[Z�r���a!�����y�"~R�I �V0��P���8��ԃ0l�(�y�CCN���#�Ї1�u�w����y"S�z��`3��.-%���w@E9�y��Q(X� ��d��|�q���y�e�y���%'8�"�؆�ڛ�y��\`�$(����2�N���%��dU�qk�|����_�
�Q�JR7tNa�e`���y�bZ�&z���11�LQB	:�y"��Nk��y&�Ex����˵�y���"���!�kݔ�#��N��yb^�)gFh�qgޭg�h� &Q���>y�ɎM?�&gʅ'��!�Fϫ�������d�<A���8�H�k��\�(a}3b��]�<1G��)�<X;�g�p�m�WRV�<�R�/ؖɀC�#tY$C�FS�<�mɏu��E�aN��2�\)(C��s�<�r���W�$����r8�T1Dj�s�'1V�ی�)P�{k��>��Г�e� ���'�~Mh���o�����C׶8J�!�'�4tQ��ud�9���J2�h�*��� X��fo<Q�`�AE-�@�*�"O��K��8>��	+lPk6TӒ"O��v���A6�E���5`a"����'�������SŨ6���Q�s�T�����"k����P�k�р4`/,���Z���B	ۧQt����E�z�<t��F��1����EPl�3�?@+|H���dy��
��Zq\��c�B:b$X�ȓ�����خ{l���I��tb0�'DL��j�&y����fLk��-3�Ņ�H�V�0"�T�l�HcPIP4=Nr!�ȓ��aA.���x���(n�D�ȓ ޲g��'X�<�z"儤,�lP�����fE	<-�tH@u�8S9����ɇ,�r��+N���Kr�ģZi���cZ'Z^4C��+|BD ��I�G�6�h� �'f�B�ɚB�@)��g�EC�S�A�S�B�ɤf�A[��ߞ0�!�I	>�B�I�E�����90��(I�J�)g*:B�	�z ⳅX]�j�I��F?p��=�7E�Ots��^{|�D�@�{7�X��'�����&����]�rE��'�2���1[0ε!6�ڏ�>��	�'�=�dLN7V  A���!�����'2����vD�F�F�g���'�<b�B��q�dQu)��_�����)֚�Ex���8A�Bݺy41�P�4#�dB��7\V�H"�Ċ�
e-@tLT/K�BB�I�Cc�-+�L\�W8C�̒�W% C�Izt :��Q�B\py"�O�o��B�I8#���a��0:�(�`f�_(LC㉔:�TbaGH�H@�r�K�K~0D�ɡ��$ץ��$֠ n�?	J�ׅ9���Ʃ��rn��b�Pgy2�'��'��]`懃:dLJ�*��/�~�4�8����>G<����q~x�A�	3h �\��j��b��\1��V���2�l����Y0��bRC���O�<Pf�'B�]�k�b\Á�2vO�n�c���J��dk�
O���{�D�#)��]
!�Ov��'8��:A�^�>Y%�ā�Y?\�J/O�����Od�$�<�+�D��O��{���Uh�@F#:؈��	�OlABM�m ���)�f��)�,��� $$�5���0ĄY�*l�j-*D!`��pl�E��O-�蟌 jfH:e�,�T^�g�Z��c2O˄��?������4��Dz&�� 0*b�B6!�Ny�tL"D��:��>k��T�%@Ι"m2Q�p� �}E�?ݩ�Ǜm��Ⱥ�@��*���O��ܕ'ςH���vӬ���O��Ļ<�'/��Q��Lӏ`ڐR%��
I�H�A�Ծ�?�3��2c���?U������6(���&�+�����JY `��Od1!���J�v@!��?#<����1ޘ�����d�BT�I[~R�ѣ�?A��?���5��$C� ]�9i�KG�"�4�"Oh�iq꛸Jʖ�� @˶ra��  �'X@"=ͧ�?�*O"� ���O1�$�tn��'�p��H���09c�OZ�D�O��BѺ���?��O�P��b^��0U��F>b1��.�T�K�W�}�����'ؒ2 �ZJ�r���i��&� �I�h��(N�r�/C	8����'/H�z�!�F4���MZ[�=JuDS	K*1��?���S(��i�B�/��p����>����ȓJj�L��N�	{�(R��; Dx	�'��7m�Or˓�E�������O��?I˦9��'[6���9dk�4W�T�dN-y���O��D׫~�4h���/ �jaX����S�:&�W �h���\�H��t�IR`����4,�T�M�p�tLA�IK�8��i�kf��#E+�O�%�1�'��Y�l��%$̑ �d|[�J�2��IP�����ǒ��9� %�Z�P�c5�O�l�'SR��g��t�����H��.O��*ZЦA��🄗Ou��@�'��	�6m��y�慴 tdK�
݃b.��-��
Q�K�P��1S��O�F̧ � kAc�f�f�{�)�(#ۀl͓>[oҡt��;q+E��h��A)p����-D�[�3OȐ�'�Ҕ�����S�? t4�R����xg˕F�.�0�"O�U$i���%�֖~/���	!�ȟ&Z�h)��Q2�m�N����O�˓R�V�
��?Y���?�-O��_�e��J�eB�y��cS��)0�8���O�X8�iC+&
FB1�?#<A�FB����dQ�Dwd�v��d����t"��2�AB�\����O���A�
sP �$� �ԙ�� �O���5ړ�y� 	R
�s"���l0`�O��Pyb�#���Y!퟈L�V�z"��۟�i��4���D�<I�NG]N�J�d�(?X�u�.ɪ��P4sQ~e�I֟�����$�	�|*cJ�>�	C ʼ ofl�EÅ'I�Z�bt���$0X3@K��<��4Jp�S�W�<o� �b�M�0�����&O���0��)��<р��ӟa��Z�ξ4���	�|t �a��ԟ D{��U�I��� ?��Ek���!�zB��!si��@4%�8�iwB�"X=��CÛ��'"�ɛMKX����$l>=@�'M�*+�����!��$
�
�O���B�O���OP|9� T�f�t�	�9!���i>�8�`Φv�؀���!4�H��i&�1H�h�7�� C_��*G�ˁ��i\�V����ӎ�>�Nlr�e�X2����j�O��D5��A� ۶�@�O�3v�=F
��0?���L/{�41���Ξ=O¨a�sx�T�/O��+�IS=H�h��BFv�����O
�$�Ov�?�'1
�CD�R�|,��D	����1Ó�hO2%bV�6L!:`Ν�t��B�$n�.O� ����+�:��4�϶:WR5���V���DJ?���v�T>�ɹd)�Y)g�S�5�)��� Qaf�t~�	 }���!���ħ/�bI˶� H*�!���	!�4��B�)}L���F��'ݚ�y&L߹Knq#�� �DM�S���	���	0~���'�X�9�aA'��G�0!� �!Xd�	�w��'D��2��	�2,D�P���2S���@B���t�����5B�-�=�N��Oz$nZ@��$@��;@l��#f�NӺ�%8���O�`G�D��^F!����"0P� ��_�)�I�S�pӧ�9O��@A���Hb�̫FHh�n�=�Pi%���"δ�'M���OR���	� a��E�M�%N�8T�[&e��J�^?A��Da~ʟ�D4L��$F*��	�#�)%�8Cf��(@���I[؟$��.\QP<��/��C��C�.=D��J��@(p̩��	X$#���h{�b��.�$�v��O������*V!;�
11*�wn1�F��>�O>y��T? ��P6G}�ȁP���Rp0��v�4D�����)_i65�O�v}"��T�/D�:H_�zG M�s�C;���Fm.D��(���a=��I�`��r�7D���O�m�T<s@,Ҏ2������5D��z�;@�+��QQ}|!��b2D���d,�%	S%TG0�p�.D���㟛5����2B��)<�IĦ1D������/j�A)�D�:,J��e�"D���5��B����C��8Q���?D�@X��ET����"y����H<D��IFl��#S��@'n�2l��ꆠ$T����̜(>��A��/-�����$x>|�"�F�1v�་� 
 H��� �B-\t�L���3?,<D�<3�i� �C��dl��B�4N����>��$*���)%W��B��"���@��N�,��̒T�[0&� ����įw�@�Pc�,_y�U�Ҍ�t�f����*;�c��(����艵B՘]!�'�f�����J�I<<Px�	�C�*�4���?A3������1K�,oi�i�G��~�bC�'�ʥ{�眪=�,��'��J�@ћ5Ҥ\"&�*=B)F���[�Qք�UJR���%�ē?����	���F���i�y1e���&`I����?q�6�Z�a=$�X(�lX�&��h+�E���C�8OdiDybe1V��!P�!\
*b蜚4`���M��Oz��ā� �x��h��.DV�Ѷhρz�!�ď�hEh���J�[&�šC�T�!���,�����5��i��NX�w!�d4i�䲱*R�Ε���udĄ�}�<���_2&��DjSV�U�8��L��Ec�(Uƪ剐�sH�����d�+�lQP
X��r���S�? 
Yb�
�����M	�k�"X;P"O��F�TP�����υ �Biy"O��S��6 �0K�kПo�9�t"O��C�J7Ux��a@+�+8��"O�] �	Y�IQ�m�%e�UW$ɓ"O����"P�i,x ��Ë(bـ��"O�t�%�h�TX3�g�$^���"O 5p�k��d�l�2�K�t\�0�"O�x��V*K�D��ӯ8C�iC�"O��I5k��&,�<%
��>8��"Od�ʁ�1��A�_�6�P#�"O�JD���K\�����$K6��"O��t��f�(|2׃F;q�&p��"OI��'��:�C�:��!"Op�R��S�E[,�+��� �E�$"O�����`�<��v��	7"O��PY�����Џρ ~�iS"O&)p�
�[tt� ��ZG���g"ODkQ�A#\!bC�J*����4"O�J��C+(��!&`�h�"OF�#%�*��(� ԀW>��f"O6�kP�C�%�5`��wAX}�"O�0C��S�t��� z%Ȼ�"O�p��ƞ;f���2�A�M��2'"O~ {3�Ƶ#LT�0lAy+p� "O"�!�D�2�Tz�銃l�-�d"O����MJ�%�^h��Y:6����"O6q��� �|�4I��QP"O~	�3N��&����^u�Y�"O�y(sƀ=P<�7�A�Ǡ (�"O����%���Q���&ǎ��"Orp�4@7��BWZ�Z5xB"Oڈ�QA�5&Ĉ@w��aiU"O(�4�Q�3�D��,�6E��qhC"Ol��&e��.����G�Ÿ@lru#�"Od�QF���{�Cb(�KAЄCE"O��2�D24�p0>B�A �"O��s��N�w�%�F�B,B'���"O"�����L�a�`�R#���"Ontڒ-©h��p )%����6"OР��Z?J�����	�!I���"O����N������	&&B��0�"O|�Ǧ,?$�A�a��[��Ӕ"O����j�
�,�;�+��lM`�"O4����]e*�(�Lݮr-`t� "O��� 
�x%Ҕ�+�tIK�"O�m�D��"U���h4�;�J���"O<p�$E�D��  "iL5~��(�"O`��Q+; �\�ϟD,�K�"O`q�ca(m>��g�6� 2�"Ovp�+B$+�4P���Ԛ�LP�U"Ox�����M�Z��EG�r���F"O�HC�K�P���*� oub<��"O"��-��	D�4Q2I.y��a�U"OD��V	ղ{�.�� �!ZD�x1"O��(��тlHj �E8@�雳"O�R��*\*$I	!�̅DZ\�9D"O�thu͐)���A����p�\�'"O��I����(�¤sd���H���"O"�H�L[0>��4�	.}����u"O4L:[�����܄Z�j�s�"Or8���j���I�.@��(Ht"O�<Rmڽ+��D��6'c4p��"O��ۦ݉W�}�ԧ0]xM�"O� ܊`nʽ8� ����Xp"O�� Kӊ�@eJ���.w�T�A"O%�����$�c!��&�͐a"O2)ik�$��ԳB�g�*��"O��R��56 t�k�aЬg��\�"O���'�4�d��p΁)m6m��"O�iG���i�m���	s�"O��j��Ŗ��}a�Έ�#U<�q""O�l�A��H�D{�+�\D�Йf"O쁰a���qӾ`H�*ܹ`?j��"O��i�E�)x.�b��1s(����"O��C؂q�I��J�2H�E�"O����fԩ7���z!/޶Z<��"O��`DT.º�;w��dcp���"O���$�K�!~T	Ū��zL8�3�"O��Q�l\9A}�-[ChR'U՚Y[�"Of9��e��U�J��Bb�ad�Ih�"O��cO�� r�9
CgZ�z�>�B""On��$�B�	Ͼ�i��4[�����"O.��	�(Oq>�cD�פ<�B���"Or��a�E���!I2�ʥ�l��"O�1��*^�a����D����F"OdM@���'z�fPz�-e����"O��K�䋙�hm���Q%/����s"O��@4iC'�����Í����"OR�hR�-�^���?|N Y14"O���4F��0&Z!i� HF�t"O�q�v���rJ��q���-�QX�"OZ *�I��麁+q@\�\���V"O:d颅þH] 8C��d��h"O�}��7P�Y���6$�:�"OP@zgE�sfT<CVj��r�"O@�	�"XL(�M�E�]�n.i�"O"�Q��L�Z@*���4�a��"Ol��ˀ'F�u벇Tf�j���"O�����-%ax���cJ�ryB��"O�Es���3�N���@�,:
�a�"O���/ߤ�d���M�.a�
`��'"���T	A	����s|E��'u���M�U��֮ƙYXJ���'Ү�r��oR�P�uB͖��K�'�@���E�I��e��$��'b(���-�ɳ�Z�/�A��'�qp	�3Y����v�!����'���Ʌ�M��� �&����
�'kTI ���`���A�>t�tTI�'8V��Gi^���٘ե�5m:��'uZHXSF�	"M��f�Ҏ_?�h��'㎨;�
�$<�AJ���_�d4!�'?1���'���:%J�9Q�ȁ	�'�BT�h��nnX�Y�Mm���')ji�0jsܝ�+:H5ځ �'�֝�D�y����ȥv�4��'�UK���l��Q	�X8rB��
�'zT�"�O`B���i�.n5X%�
�'�ڽ�QK�8��B� U=`1�)�'���p�Ûx�4P��a�$TA��'��P7��]�Ƶِ*
+[�P��
���&�і��@�+�.�`�9D�`��T�2������T[�"Ms�%D��' �@�H2��<*�1sD�0D���E � 7��C��ް��t"D���Bɨ"9�aI�(�$R|�#�O D���욽$�24�DMZ���?D�� x �M��<'Ba�TA�;(��B"O�p�+�$� ��*��Q�"O�z�'WQ;~���R�l��ؕ"O��
`�@	���a��ұG��y��"Oj�XC � m�Z)��E�D�1�2"O [�A8B�r@DcS"i��%S"O�1ffF	Hr��E��H��XG"O��ס,(�8���+�ܝc"O�;C�G�:�y�Ɨ:0A�]��"Oh	�O�+h��,�ue]2/H�*B"OL���"Q.s$�Q#�#E f+L�"O�b��i���p��Y/4`a "ORQ�_�$�
�'�!+��@�`"O�}8��B�_2�%�g��[���3�"O@cv�-|�x�`/�ZaT��C"O܄������RI�ŀ�aX��J�"O�=��F�"7Y��`7oC;es����"O�m� ���(<Tx $�g(�k�"O��W�C�T�D�M��F-�4C�"Ov���!`m��B��%
��U�"O�7�,A�v�q4����"On�����6Cryנ�O�x1�3"O�e{��/M�t�i'��`i����"O(�z5�5��3�ϛ�t>��w"OZ�pܘ8�ԀW�f_�d�"O$��Y.�ph�S�~�̰�"O�d;�J�-+��I1EiKX��$�U"O�PґȂ�,Ҕ%�զ�5F|�#B"O�.4�8��!� b�D����!���'_��*��m���y�o�3w!�dȝ҄����a�f�7� v�!�d� �L�KS�(v��TY!��!�$^?7���D =/�����:'!򄗉5[A	9+�dI�nW_ !�]!��e�'J�e��-:eAG!�Dt|�QpoS�)� ��-D�O-!��%�q3e!��W��]�Q�L�!��8v�pX �ԓ~6��2�ʼR�!��F�X�ꌴ>z�I��b���!�$Nxe�10�g��f\��PAm3C�ɆyC����<��sF��
w��B�P����TMݰ��0���]	��B�I7%��`�f]:��H�X�1�pB�	��"l����Q���2kl:B�-<�j�)�KIp_�%p����#�>B�$
!��$�c�18�iX/�:B�	���[��۵f ԙp� �&HB䉮��'g�;f�n�X���'l	�C�I-z���ql<C�lxy�	�7��B�ɞPT`�!��8�n�` �j�C䉨=��G)-=�B��U"I�\�TB�ɓ+�B0�-��:�ق�lH�i B�I�Y��T���%s�Dy�13�C�ə^��`s��ݦ(��� cQ�L��C�I�K���s��:n����
�rdnB��9ft�xP��]4D���R=�6B�I9q��[�c��I� ̙��Pg^B�#����)R�Wԑ��<�B�	�R2jŕ�?���v��c��C�ɛ:���U��;[�|�Ӳ�r��C�	�ozZ0�HI�'P0:�dɎ;�C�V.�0�ˑ
~�m�GImt�C�I�7�e�-B�����#����y�ER&o��J"����牂K�J �3c .�PePTm�6 R�C�)� 0��kɒhW��I��ȒP�j�"Olm��H�q�rR(Ѳ2G Ȳ"O���j����ؔ�>A��K�<Y�C�E�.h��MY#_ˬ��h�^�<�a�#�l���i�	i,�q�Y�<�`"�z6ݠ�lQ�%'���&d�Q�<`$��z! ��'Eyvy"!HE�<�]����;x	�]Ҡ�ߎ!4B0�ȓ+tpx�@�� g���lJ�.��0�ȓ �8�C� ���j!��)X�W9ā�ȓ!0<J��L l�V�.Y����k#D�p�!%��@�ВcnN\��[fh"D�*7N*lH�dk��=9�	.D�DRvi�PCh�!�f�i����!�*D��{�O�^�"M˷L�H��<��*D���/�q�J��b��p�(D�@3��RX���� fD;��qb�(+D�8�FT%-�L�i#��!����aL)D��C�߹[tj�a�#\3X����'�*D�(�Mۓ�֬����++��[�,&D��Q�U�(������hI��!D��RHJ�T�yĢ[����%D����A�	K�A�7. �a��]p��6D������r��e�7�֝T D�L 4�D@���@�i�����m8D���拎H��d�rnG) H��)0�&D����eR �U( 4C����+$D�D�%�>'�|�� �[�8U;�g,D�0��L 1[��;@�m"R����&D��!U���m*.h[S��X�<��$D����_��\�[p&��� �."D�!:?(}k5�=E�v�
�:D��;�/:%,�pF���a�-9D�$1��H�^sFD�w�OX��"a;D�#g�B�M�=�P-Օt^l�	d�3D��Θ��2|ya�d��U�>D���Pb�>� ���U3��m���7D�0�3'؁v+����*�W�J�
�+D��ۢƃ8KB\���^	_R����!(D��fl�]�2��%Ȱ<E�U�"�:D����/����%"�$����&D����i˕5�Hy�%��e�@ٳ�o$D���VmC��ɨ�A��%�(�F$D��9��7vw ��a+/*/�e�/6D��`F�S�颂�݌f����U�2D�,J�S�O��(;��,C���S�+D�\+�X�&D�ik��ѱ��5`p%D� �d͕)ZL�[2н��"D��"�l�.��Y��*qԠ��u-"D�H�6��>�P��,mxA"D����I4\ڂx��Q�V���!D�X2��W�A�X�k )�jt(AA�!T������¨���Z�;,���"O")�b��hj9▪D�=T"O <�Qp���I���`���AQ"O��J�l!.����0��]�~1��"O��I6�G(߮�Ҵ�՚w��1)u"O�0K�M�!e�nLQ"h�,KP�"OK�6:�"11���p�r���!�yBM��oYZ�K��(d<@�"� �y"!�����c㙹a���J�G"�y��ёNF ��ҦL�t;���1�y	��'���hë30�0A�LO��yR�Q2��b�/�5z���Ŝ�y
� ���q퐑W:6���&��ܠ0&"Od�0�.ɚ�(y�c#$ֲ횠"Ot�: ^VN���i��;�"O����J
�2��)�ʌ�g�~a`�"OQ
C�DBdTx'�آJ�$y�Q"O"L0�+�)O\[�*��"�B��"O�%�T�ΙE�n�rv/^(%<09��"OD9{ �֩C�"Ȓe"���"O�x�`C�g~��)�VB���"O�8�ƙ;c<�
D���E��Uq"OF�� ��x@���W�H�J�"OX�h�J7PTn�ҧ��	[�8�%"O�,���ק%�
 �1 �Xs7"O��C�A�%y;�8벇�1e��d�0"O��7E�6�h5hζm�
Q�"O%���̞[<��D D�$9��BY4�ɂj@.O���8D��l��D�A�䏣 Z�@Y6*O6pH4�R/$���Xw��O�\jd"O~�
C�0G洠��e�)Qx�c�"O$�S����$5�A���@��� "O�[f�kx��D"�@쨋0"O��[�LƩ$�:D�Q��|t (0"O�m�%�F	�*�P4�1Yڭiq"O�
WjX�T�jq��Ȥi��:�"O����G� q�˦(��Iy�� �"Oj��s�ţ|�x��v˿g�9� "O�E�A�K ee�xh�AH���5"OBQ�P�H	A�����+�N�PT"O:m�F�Ͷqob��v	�ou>P��"O�HH2��6�N		'i�l�T��"O^��%HGʙ(v�к_Z�!�"O0-�C�E#ihః.]e�� Xq"OL�YÏ�\z�,a�FR�?=T�b"O��pG�е��[c/$mn�f"O�TC7`°[84�^	
:K�"O~�83�1Ʋ�2��Ӵ�L��"O�+6'�9��Sď�>wL����"O�����M�^�B��W; d�z�"O������ r�Z���#'�D` "O�]{cb�g�v1K�#�	YmD�Pp"O��i��UO�5J�`�b<4�i!"O�|�1���bI��d��\*~irp"O(��G�Z4���������"O�`x�O�=�
x�'K�s�i+q"O>��LWXTc���K
��d"O�z'�O�j�~�9��Ѹ4}�1C"O�uy2��X�V�����"����"O�k���r�81s(�+Rj�A	�"O���Cͅw�4�h�ET�fh��"O�i!�@A1J� � PxH��"O~� ���`|��H��4=D�,zD"O���BNڮq�e�1�1:[�sB"O���DL�{�:�ѵ��- %�1q"O��B�J��%��H�N�v�ֵ�E"OΔC�d��\����E���T)�"O(�:ԥF�D��5KوeO^�� "O��{R�׋.����G�T��Q�S"O����ݼ)/��戤U�Du`"O��Y��Q(Z�h%y�Eȩ$d)�	�'G�5b�(M�I"�գ�8�'K�t�1���eb�	��퉧���
�'Y�8`c#��w#.رW�\��P9a
�'d�<���i��)0�/�3TVq���� zD�7��R� ���U�4��p�B"O8X��nXI��L�#j�!<�B'"O�j�I�H&.ȋ�땣Y�U "O�	v���$z��S`X�re�\z�"O$�KW�Z�#�N���L'(Y�<��"O�!�G�D�h�x<9��c�.8�"O$�`��?}�d҅�.K��T*�"O@��Ee�P@��	kX�l���"OT���	48rH��#��W�F��"O\��@ŗ�z��#�A��"��5��"O��`� �>�FR�)�/T�"O�YC�iP8$ R��4F:8x�"On@X ǆ5jK��;�薆+D|�*�"O�u��&J(7��Y��M�CZ��"O��"SMH0k��(r�(FR� �w"O6H�!C�K��c�.�3rWd,��"O���Pa�,e�F��o/��L`�"O�xkA�p��p��/дC�6��"O���fU�8nH�)aL���D��"OX�v� ��ڄ8� ��M�j��#"O�Ec'I�35��*C�A ���3�"Ox���A��/t�Ay��VV�:Ȫ"O�IK�Nc��я	��|H�"Op�c����N �]AEA�m>�5�s"O
��q�ā$�|���A�/;�P"O�q��P�z"�uڔ`;4D���"O�1�Z�>��ѐ��$n$���"O��؄�Q�8}���vbP�9�|��"O��kW\q,�{U!D��9�"O�q�Ċ�!:���Ta�_�v<�Q"O���#�T�crZ�u�h�k0"Oȑ��C)}5�P2f�����غ�"On���gͮ9��$)�C'#��b�"OR%
QM�;u�d;�b�)����4"O��[ N�;4^!f�+��X�"O���^
n%�t���� m|���"O�i��#�?Q�0)��^�'Z�tˤ"O�$j�o���l�0W�ر"O@فI���A��ur ]�a"O\{��D�W�P���X!CyV�"O�U��Ί[���(�1K����"O`E� F��^~� C���Q�"O��@�'.��crl��,q:�"O�y3G	��hr.���i#����r"Of�z�AG�&���N���h��"Orc�F?fв��Δ!�f�a�"O� �7!X�?d � ��:��p"OR�a��� `-rg�]�C��U��"O^�+�eݠL�fh�ե��=Z���"O�@0嘐&���ڤ%�<NEV%�"Or�{P�<^�A*U�C�'P��"O4ܡ�h�����P֤D�Q�ȉ�"O�L���ݢ`�<�ūٍ���[t"O�e����~�����꛵�F�۷"Oz]1��޲[
�� "ɍ�~(��"O���h��]R�*�HG�-�ؙ�"O8y��-��fGf�v�_�n�q@"O���Ǉ5}^���]kZx��"O��Vb�=k��#�'���yg"O�#���(�"y�f�V3i�ܨ	&"O\���O+1k~��7IX�@�ĥy"O�P�5bC�G�4�P���q�&�B"O�|�I� ��4� M͒g�h�"O|T�p�Yc謨Ӥ��y/��"O� �}��O�)~x��dN .~�	%"O�)���U�6.�YbQǨa(���A"O,����_-;P�hro�l�x�k$�Z�:�~ճ!���A�t�/<OTxzf �6��A	��S������"O����LH.
xc��ʒ����d"O��y%��^�f%c4H�I�Xy�"O*$r��K+TTq��dN\4�a"O�y�̰g��,)��C"6��"O| �
�>i�tucS�h��`"O��qw�ۼ<��TXT-1a���1"O±	���_Aĩ������D"O*q��!�R�S�e�4U�2�i$"ODTw�J({h�h��
�9�����"O�Iw	O�yl�ը�
��E Z�V"O��1�L�
����&Dr���"ON�x�(�=[ǄQj̝�6wn�A"O�)��^�k_@ ��*Ӕ%g��"Or�)N;�N<��K(HZ]��"O���ǉ�r��	 ��wq�%�"O�eK"��,-�jgK��3�8�"O�d R�=`�<��U�^ . �4�',~UXVbB1{+��t�O�n>)��'��bfFH
M���C3v¦Y��'�"I)�0�ȼ9c�H)[�z���'^�p!��)z�P�3h��RQB�'��4s�*��kk&y�bң}q:��'�d��U��"~�i���@9u� ��'4�p)�䉣	*�	p���qu�YR�'!�0J�雵Y����d��d��x�'����oBR�0�A7gZ7J����'��1
EN��n�����>�<ĳ�'�� a�ƒ>q~*=h�%#RZ���'�D��U�Vj&�@� �J�K�'�p}ɰ G�(∑� �M7����
�'�b�`�^�q�^u�U��WP�)�'���%�e���"��S�����'�阒.*Yc�����w�����'-P}��ǙD&l(�B*�6FRRT��'�=8���&�#A)F�/�`@�'��A;��͗'1�T��]6-��,��'vB�z���UNPA�G�-H�ժ�'��5Ə
ls�(JpG�5I HS�'T0HW#ڼ�����Y>�Ę8�'��h��M�hpL� �n�"�'.n�q��gtA���4	dd���'�(� �l�.%yl˕�כ����'I pS0�]�>k��
�^�Pܺ�K�'/�BC��1}t�Cc�]�6�xk�'ì���,��w��Q҂�1lj3�'@)��1r�|���˄4]�F���'� �A�nF�V��;R慺[�zI@�'C��kQ�ϳ���I��#�'��BP��8kT)Bt-̻p����'
��9W��/
XM���n�̴��'����2lR3^B�`ƃԟ9�ɱ�',����eP�8�pucN�1��
�'b (A֮!m����əR��{
�'DNI����ڠ;�gO�����'J�02�BlJ�QAI��v��'�\�
fKL�3ŒDq�N4af4��'�ԉZ�-��(�`ѡ�P��&ѐ�'n�!�f�gO^d�A
Q �,E�	�'@){e)Ow�"������(t��'^�P��ϨY2��L�vzp���� �Q#&��bS0�R��[�Ԕ٥"O`��͔>�� �#L�����"O�M[Ď0N�n����@��qh�"O.����B�_j�#NK5_���u"OLjD��8G�:=a�MԈtN��t"O����s,��e�ÔnV�I��"O�qKR�	8Wu<*#�Z~����5"Ovx)
�y�@��4i�+]��<�"Oĕ��!h%���[W� `�"O���V�4�ԇp��"S"OR%#N�1i�	zjrA[�"Ob �u��#k����H�>f.\�E"O�e�#�f�R�!fǝ�	G���c"Oh1���hy>���y����"O�AS2���rG4��dL�y,Q��"O��;7H�m�^���@.g��`�"O���B���Y��5i#1�fMSD"O^�(3�W�&,��+��̫?�|hcC"O\ءU�4^�\ HRI�D]3"O��J�*}Hd]��G�8XD"O�M�F�H<*������1���`�"Ox��NՈB�����8Ү1r"OA���
�,C�ɱkZx`�S"O����g��S#�#�ڌ�"O�����+W¦Б�ݸ'�<�h�"O�y�D�1�$QrAd���e"Ol�bV(�Q�\��!��U(�"O@�I'�6PBa��ŲQ�i�f"O��kU�Q�C(4,�#@�?Q
�"O�d�5�[�:
4�FŢ!7ȝ��"OtC�o_u���х�W)^#ĕ�"O� ��#L'.���Y��p�
��"Ov��' �;���iw��<�,�r�"O�ЂdN��Cغ ��m���	�"O0�Ҫ��vHa��Gֈ=}�ّ�"Ofdȥ�P�dV����g�1:Sz4�"O|��`�\l���G.Oh%Ѧ"OrL�w ܳqL̍�3��.j�,��"O�t��)\��0�I�Zڨ��%"O����8�P���źS���"B"OD8�B�	]���d�O�H���"OL�{�Nk��)��IJ�|hBQ[7"O��vc����%'�(Y��"O~1���*OC��Vd�}r��)q"OVq�5�΁l�P�a⡄�S&dK�"O�b$��x3	�����#URh�e"O�R��9l6���+W�2F4]Zd"Oj�p�mɛC���BEZ��%����y�$p5 [�JR�ċզ�$�yrC�v�l��0��@�`m�W���y2L]��mPD畋6�H!�6�y�nG�N�����Ð1�0H��,��yR�N�9%X���"y�a���\5�yr�T,�>}��/$�R�%'�yB�ú���A��	f�:թʛ�y�eճT�Ay�B���b�D��y��Q�[E�D1��
y���d����yR^�҅��5���*�εy��M���]X��h�@�9>��Ú�m�(C�I Y���&��"C]8h�gg")xC�	/}"�N\:R@��W�RպB��;���q��b��"���e��B�IƦY�d�� 	�4����C-.�ݡ�)%D�xP�+z �8�@�l.�PWE D�� �d�ѠA3yG��qǮ�3\��Y�"O�܉�'Lݜ@��Q�>=<��t"O�j��(N<��Q`��=#�mA�"Od�)��@0�>Đf��v�c"O*�!6�]�Z��[ŭ�<t2�Sc"OX4��/hrv�"猟> ~��#"OZ�A�fO]!$���-C���p"Op�a�bOv1"��X���X��J��ym�1&M��Z���<]=@�o��y��8v;� [u�PY��iԭY9�y��1�8U���ڝC���3J��y��%$x� ���_n�0��KK�y"��~X\U��AUx�t�����y  k�j��P��wy�����	#�y�
��4�@A�߯9[�0` ��y2L�_ѐ��"$��b#\��$&Ԩ�y
�F�.���eA#���e��y�n2zX)��)^*�����y��\�XϮ	pU�ӄ�ih��S#�yb@�.G<)�`I)!�$�4���y�G��a1�aP�@�F�����h��y�e�/ADoʄ>� �C`�Č�yB�R�1W��R)�3�8�Ѥb��yR�-c�d�2�(�����.�y��Q�L��Q1�@�0L^�S����yr"X/x�L��IJT�I�#d/�yB�T��$(�oܾEK:�S⎒�y����n/;�X��&���y� Շ0:4	M�h^�Z��� �y�l��)�$��TB�ZK.L�@�:�y2B��z��$�	;T.�`{wKȱ�ykG�Bϲ)c�MЈ�&c	�y�b��d��I��3m�X�Z�"V�y��&���3�5j$�93�̈��y���[�J�c��]� C:}4����'H����D�0�%;�Q�pk�$��'�j��$AΔ )��@,[cQ���'�|��`�v�M����׬q�	�'�HD:��	4D�V:�D��%
�'?���PΛB�ᚖ��8i�<�	�'�*���@&?���a�FI�Br��'ɢi#���:T�%ٲ�D�Bv8�x�'���⣩��F����`�51l�ʓR�PѺQiK&Ld� 1���?���ȓU��2t	�EB �li(�����܀3撁3.���H	}~U��/��ؔ�O���`�˗H����ȓYbJD�1%>q=����K�=���)d2$�#`�*fd`q��G�
��P�ȓp޹�t�ײ>��LHAiJ&�I�ȓDMbpX�gV*i�� b��Ʌ�R�Z���6;�N���.�kX
X�ȓGR,���)��D��I��9��I��f�E�gcֈL�Z���`^�|�N�ȓ{��В���W���W�͆v�H���~�|yI�.V,�Z8`�LLj)4X��'����3�K<�s����-�@�ȓT5��s�![0��܋����(���ȓ0���s���)2`*��v��܆�H���C53�:�v&Џ\��4�ȓ9v��{��H'q��sJϷ]Y���ȓn���Q%�
�v6, ����ո��ȓR/��B��X����(������5Z85�V���z��������4Qx-��S�? �D��F\�a��Q(r��t.n��"O �'Z2���(��P ]=����"O�3�DW�j���kɞ�*OB#�"OdH��tEzI2	ʖ_0$9P"O���,W��e3�M�uMx$��FN�<�7h�W��h7�� 
7�J�<�	��~�$Q����&J�ð��G�<�v�Y�O�<���i�O����P.Iy�<���]+L@�EA6�L"�v\{S&�o�<�aNQ>+�h����e�b$��Yg�<�� �B]��ZQ)�,�^�*���f�<���G�%�q�O��īFk�K�<�J3M�����*Q�p�� �F�<��O�{::!��FR%#5�0W��g�<��Jٸf���d�[$h{hxU��e�<1�o��Q��{�g��i�䁋�@�F�<A���deȅ!fZGp�CÅ
�<��E��@���j� ��u��|:��{�<!B�վJS��Zr��1;�\�`�f_�<���D	;F���*<<�<`P��r�<A��WcX��:Ӎ�#!3� H�n�<��M+FV���o�!?w���ᅝt�<��K�,;&m1�K��	ː� �(�G�<)'D��R��	$�A
`����Gm�<Ѡ�[� �{��ʍ4�^�:q���<�тʡ^D�UCA���5=&�Ҕj��<���X,�8�R=1���x��Vt�<A�G�o��(���K��<����T�<R�T1}�Lu��;Y�(�+GEQ�<���J%6k:��EG8&02��P�<�&��8�^�����.0|2<���L�<�fi'J�%(4�--u�4�S	�K�<�ҧMb�l�cCl|���	%��q�<Q$'�������o0
���d^k�<�UbڜI�F�Њ��	��ȃ��1D�����"8��Q��F�1���.D�,����*qh$����>V4��6�+D�@ a��~��IQej��.����s�)D�P+0B�Út!4�)���uE)D��9@d��kW��j5ˤ����%D�dr4GF�0�b���E��a�b#D�lSucZ�/x����k�A\����%D��B���B��$��f��Uf��+%D�*c%�.o�NpP���V�fa�C�$D���FmSn~}P���6{�h����"D�ܫS��:%�X���R�9Q�q�%-D�L5��
����
j��e��f+D��yGܴ4v'�*pC�ѲaE)D�,U��
s6F��j�=Oa�y�g9D�L�&e�+8Da ����JI� `�8D�H:�JF��C`��fD&�y��:D�������<�U) f�:DYB�(8D����� V��K��ТX �8;�7D��G��	u�ʹ#��L��`�c�8D���b�S?v���AJ�hа�1I7D�\ZA��%�f����p���+�?D�l��'�Y�8����& ��h�w#D��r��}��0zwG�:�x�n#D��8JW��q���3�R��"D���+�o��P��.}b���,D�� �
&(gXt��/
(��%�ve(D��2��re�x�Ώ5bK���>�yB��1?��y�7.V/BE��B���!�y��1Y������D?eRtyओ��y
� ����E$+����4D���"O��b�G:�|y�	W'G@�D:P"O
a�t�XXDB��ŽVxl��"O���+�? ��#ꊡgM����"OB�����_�����ȈL/��H"Of���
k�:phǇ6-����"Of�i�Ȋ�R�������O�D*�"O�\I���1!0��B�)����$"O���n^�#��I2i۬�{"O*݃WFO9>�����k�6i_�l��"OPdP���FY0lT�X�v�.ّ7"OB%�b��cT�(�d�Ƹ��"O2�@�EP��7�}��`�E"O�4ITo�q�^�j�Y�a�����"OFAn��}����@_=zX�x�"O��r��)KiD��$o\���\�"O�B�/_=2D�JB�_, A!A"OhUQ�*P�$apY����u- �"O^MB�&D�c+�)��)h��0"ONU�pfަT8~��f����Lj�"O�5Jl�
B�H*��N@N�QW"O�l��ח�Μk�Hў���"O*i� �85g��g�ڳ>%�"O�I3�
]
���2k�p|,�"O8��E�[4K�D0��L�{����"O��X�g��Ptsfi�$k�<m��"Ob8�@kP���Je�]"X��i�"OVĻ�T�B�����:!��"OPA�zz�p��1.d-�"O��p�KI�=$�Ƌ���K�"O>m�%ΐ�S^��aɮ
(Ļ�"O6|�7O�g�&u1�S"�i(�"O1ۆĄ,l�����++���"O��b/� c�5����+2�N�Q2"OL]���>���x�J��?x���"Oh�q �=8�+�'��,q�ٱ1"O��
S(�)�L��F�����[E"ONM��l�(�^Y��&�vZ�#e"OV��NP=�*hXa� \�"O���smV��v��fț�1�"Ol�+<��y{�J]j�D��"OU(7�f�)��ѹ�DpV"O�Ma�-˄N\��fB;0�� �d"O�x�&��,��9�g
�����"O>@Y���N��Aֆ�2�≛d"O���A��0�y��G��>a�"O �R��[�/�h<�M��m	P�{4"O�9��_�9�L�A�	�q|i�"Ol	�Ql���<H���U`�Y�"OD��Յ�.�n�Sbf��e�ذ�"Ov�k b���l�c�ܓu�le��"O�)�P�� ����c�A��my�"O:܉0�� ��HC�J�#bʬ�2"O��Y�C3"�dP������i�"OP\s�P�&���(1!ݞK�P��"O�C4C�V��(�r��+�bls�*Od9!U+M�+o�i�E�:?�S�'�d�yD�X'Omz���j�5ŸP� "O� �C����&�!@
���Ջ�"O4}�uA�P;BD8㨍""�h��`"O  C�_�x;(�c���y,�)3B"Ob�RsE��Jl]KI]�j"v�"O�AJg��=O���p	Y��5"O �l�C�b�D�@"Re<1p"O� ���H
3p�a���D�-al}�"O�m��	�JX|IU,Z�M/�$�1"O�L�k��Lq2=+��Ww+�i�"O�m����>}Z��W���>�xy�"O����\-d+d�A��$�p#�"OZ���
ۇ�8�#�Y/��z�"O�H7I��q��E�^�x��"Od�j`��7������.|%��"O�T �N�B���"�I�=����"O~�q���߲E���nF�[�"ON(��*@�&��]�F,Ƃo\,a�"Oح��� W�İR�E�BU8�C�"O�0s���SnJ|�I�M��})D"O4�G&��o�I9�H�'L���b"O�<I�]�P�@�ف���pY*@"O\<�b�06�
�
��A�r�Q�"Op$j ��5s�u���m�1��"Ov���#�(>1�islY%!����2"O* ��V�/��)�Tj�'j���)�"O(UQ����l��@�G�C�(�b]!�"O>�#R�ޘ5�u��E�V{�k�"O�ժ��w�l��B�5g^us"O��@w�ċ4¢��@��'yq`i:�"O����Y-f��R�˜�WW�5
�"O����囓0�z幱��c��)c"O�5�B�p)�d&`�~�jE��k!�d�!��-��k7ܐ�"�I�!��ȁ}��cv"-�����'3�!�D�-�!"Ǐ[##�ޠr�GV�'Y!��ąx���$�ʼ&��\�r&�#2!��z�\U:��"^ވ�)�"
u!�$˞b5E��+>*b�he�8>!�_*j*��Z�l�(��Qt!��u�R�J�L�5&���+�;D+!��Y� a�e����<&0�kӈ2�!���Ak��":�V%��!��?t<�4�	.�.Ȩp	�-!���WWzA�"�ې:U�d	$��i1!��_�Ku�i��(D�8�n��O!�$B�i�I:�,o;��Wo�G!�Kh�j���p3b�I��+!򤛩|0��$,�-j�tt9�P�
!��[<	���b�%��|b��E�۬	�!�Y�0��:s��g`�yۇ�g6!��Z�>��M�#�J6M����T�)+H!�D�2<�	+J�&��Z���&?!�> �n�����*��14�Q�!L!��4���!A#�ZHy2҅u!�D��qOH41fU��8��%��|!�D���v���n͐$��`ǉ�Y%!�D�� �6Q ���>�W�"8!�
�%�f(�H�m� �(dh�)(�!�C�A�L�H��ᖩ��N�!�D�?g��� P8z��1�7n��^�!�ę�Y$�����&��ܓ�џz!�$�? 5jX9�������Ӕ�>5�!�d^5U(>T	��I4��d��<!�$WA-�p����Z���8C!��ƑlP�R��J$n���p�S-!�!��6��0�� �iW�����#G!�d�(a��="�j!L1��{"�O�!�^�eb|�� �ְ'l��!��To!��4F�> c�푃"�����V��!�d7;��x[3烿$�>����\��!�� ���ZJ�\��RNX�HG !��"O�hKbN�w�LD���AGB�)`"O�t�`薡c&�����D�)H�"Ot)1��L�.�d���h�;�����*O�� GE�;n�xz�[�P��!	�'��|xW�Y8o� ��ڥMM���'�Q�c˜��F�C�<EX@��'����v)�:r�9�+�@eP	�'d�my�o~�ĉ��;��IY�'UV��T��9h����3��5@	X�'/R���Ǜ�5C0lЂ	w��D���'{<T:Ձ���5է���E�is�1Ira
h`�`���h�X��!
�l�U��JI�a��
;^q����w�!�!��OO0$�!mT������4eZF )���UvK҆����k7%`�F�a�E7�\c�P� �ޮN�����)j��ڴ��!�I��M3 �i��s��(�A���a#T��W/�;���4�O���%�O�eɴ����f/�bGTt�P�O"�O��lڭ��O�2�̧a�֜:��{n����7DpY�(��E�M��9F�m2���d4J�Jg
�lڱ! >It6�xu��dUxd+��P9G�ԁ�U�';|������"�K�m&����C�2;K�@	�������"�����I��e�&Iį���V0Dt� D�
f
�d��j�-~��!�\���OړOP�D�O��A�"i��&W1s,����G�d��I�4F�Obf��<x�*Q��ʶF�����CP�M�����|�����$�-�3�g��`y�'�պ_RUE�%~�����OrVB>-L�0"�J(��je���:xK����5�fd(!.V:f�KCU�'��a�7.
BN�&�fU�éU�a�8ⅭG7%I<�i���ZZuA��l����=��F�@l�����A��o�R�!�Вs�K��xr�')�T>-�R,�95�! C�ŹK�QХ�ޢ��xbiG$)^.A����F��������~�pӜ�lKyr��	m7m�O��į~j�`	'k�6y��ĝ}8��@�&0��v�'q��' �p�^ R����D��I6�kR���|�BC��?���T�g?D m�v�'�f�b�ʗ>�B�w���@�E�v������d=�8z�+Ɂ� 5ZAe�r:��QU�Ā91b�'c��6��+qfꔐg��f֊�z� ����IM���h��׮#�ْ�L��h�b�v���p>qB�i��6�w��x�'M�5�n�9P�G�_˚��~bA��e6��O��S��x�ϝV�\ݹ���3�4�q��=Sk� L؆{�����G"1`d:�!��OU���1pأa�IN:���JqH!n�Af� "�C�&ڌ���E+~O�`���σ�F�Q��~�1 /��jA�4�Y�1���E*�QoZ�U-����O~ԕ����i�*��d`�����Ò��4��J�O��8���<y�}�
ǣrִ���M�u�~��	��(O��lПd�I�M������P�k�NE�t �Sx��@�n�
��'֤s"n�<-8�'1r�'��J��
Ta�|�u�E�Ro(���"@��]���K�d_���c�*���4���$X�l<�T�1��=Yb��+.SUP�����U��d�8B�2u;�S?��ٴk&�
�-�<у����3wJŅ�g2X)�'l��S��?���x��'�X�L��AF���<-��4
+�	R���'-�̰�!�Y -���0J�+5�����/s�l$oZB�i>���L�I�ɺ�j   �   ]   Ĵ���	��Z�t�ʔ*ʜ�cd�<��k٥���qe�H�4͔6Z <���i4�6�<�TԇK��,���I�q,�m"�M��i�F��D�J���PEK�=������0��1Ï���M�A�d�2�O̨ٴ4e`U�5��nzneP'�R(f9�'���1�.���q-O��qo��k�<(Oh�:���*soұ �dV�O�r�2)��P��-O��I�b�[%�?�ɤ3eR`�W�MW�|t(fNM/��`��e��'��u)����4~ �KW?2A�1P�@8RJ/u�u;k�E?�eeD�P�?}"J��l�~	�M~��
S�qĢ�x�-[��n1����<�@�5�sv"<9c�Xb\uA��B%N־t��J�~�T�%ቕ*C�I�lS��Hi~�Cd�!K���'-: Gxr��xܓ~��IՄ�4�!����FG�\o8V�h��� �Q"q�Z�	H���$�,\�28ya$7�	����a���1���;P�:0���H�Œt�<�H5�����zqO�l!�,�v��)���[�"Ԑ�x�	4/�����y5	+�PB�K�Ϙ'hP�Ex�
�u��%}y�9����	�pH  �?�*�I�5��hE�xb`��l[7(2[��Q󴅈�^p@�(�OP4�-O|�雡4�1��q� m��~�MK�j�*���wv*8 %g�@y�2\>�� 4}�i��|��J<�
/�����Դ4�2���"�0TH@"��s�	 7T�"-�^���/y��DM�]_�����b��B��1kp��  �OV��?1��?���ܠ�JaJ_�*����u�P{� (����?�(O��np��IƟ������a t[�HS���X�����$�g}��'0R�|ʟ��2d+[�p���)>ԑ�U-({A��3$� 
I�i>��7�'"�D$��X�#ف:E�T	T#�^�9���Wşt��؟t�	��b>�'7-�4�($� !��"�p���V?��E�!��O&�������?��^���I�O*��K��LD ��*E'���	��@����e�'�R�q�#�Qܧ
NDR7�Z�D� �s�g����$�O�$�O����O��D�|
!$Q�!p�)���U#2L��hS�n��������'������'7=歷��F��k5�墎�\��͉�e�O��1��ɏ \մ7�}�@)C���X�s���    �    L  �  �  "&  t'   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒�"O2�*�Tn�)PgOT3Z?`�%"O$�27���]�h�QB�E�V p+�"O�h��N�i^��B�K�]�Ā�"O�����Q�z�Hd�ACx�U��"O��#w����P����>`w8�u"O +6���~���"-?���c�"O��e��)Y������FH1�"O8�L�<4�*���Ɍ�M%z�!�"O�I)�n�~�P�"\�'��j�"O�� rU+xX��⌚N	8!��"O���a�Ґl�<t�VkOp��2�"O&E�b���D�4�*�d�`�D"Oڸ+eŇc��D#��.�2�J"O��I��r(�y�3fN��Cw"O� �����O�əf�0Mn��"O��S�	�g���
��/8��5�"OT=q^\�i�EϮV���W"OH�h�Ã�x��Ӑ�ʉl���"O�0{Ei$R�zp��)!����"O�z���5�,E\����r�"Owq�s��BU�-pRaCd`�ȓOIP3�&�XA2H�+*V�ȓ�N�8v��i'��c��������8�lQB�ʇ�^i2�鏻e�4�ȓ<�D��t�æ`:T,�Wg��^��ȓ){�1w�9��K�O�NrZ���ª�A3A�+��(��O%D�"��ȓ�u�C��k�L�C�P�0��	�ȓr��e�q"z��`H!) |�ȓ_Qh$�f�_�>-pi�9G�4\�ȓ�������6���vA��_��P���
�(�7Q�J��3b���X(��/�Ċ�o^�m���S���E��m�ȓ#�
)�e KT��B`-�~H���y4�!(�Գu�B��D˔-2 ��ȓk�-Z7�N�@���9��.[l��w�:,Q��Ĉ��uy�N�-m>l-��~�F�j��"`v��C�T,.��ȓ-�Zq�S怇�V$P"�ut`B�AZ4�x��2C^DMx��ӚI�>C䉪V&ɫ4惤 ���SOT�Ls:C�I�UU�EA��Hp�蘣I�&��'&���`�%�,�xc��%~v<a��'� ��D��6��)��"thT|��'��0bOS�[��|���m_h�k	�'Y� gc0�\Ӈa��p,��'5�Ј4$�5*��������C�'�T��׋ͺ{\��8� C�i�TQ�'� d������č��̂�'6&��Q*1���"I�:P�
�'hZ��%mМ&�0�s�g>5S�I�	�'�&�C�ƒO���01�_>-��(	�'�J���̈Z0��5���
	�'.��v%N(.V�*v�����#D�y#�.{Э3�͏YG�e ��"D����%����2. �x�(���+D��*Ί5n���aq"N�H$"�bG�4D� ��kôa'���s�G�"����5�1D�|�ϵO��M)��u͆�9u'>D�h�D�V�U���d�8q�z-�S�8D����Ǘ���	97F�p��:R'D��*C��2b�8�3��Of�p��!D�L��N��A�^Q��b_�/Ԝ8j�O$D�������YkB! �g�+Xx�M�� (D��a����(:Y��-�t�Z�Q�!�$[~S"�0Dj�v͎`���U:9!򄇪D����o�� ���"���dn!��Pc��� �t���;�iO�0I!�R;$x,4��n�5�H���!�߫ ��Q���r�A�.�~�!�D�8s�jdi��J F�;$��6�!�5<��X0b�-Zo@P 4�29;!���Cx Y�D�3R3 �Ru"�gJ!��� �&i�#� &���E)x�!��C�Dك �i<�i��f��'���#���%��e��/l�<�P��8b
��Gk�'�*xS�#3T�(�%eߙ�^%�$L�A��Y�c@1D�� -zVD<7|�C5U&Y`��"O�	�!/^|�T8���=Z*}��"O�P�E`��3���2m�j�hp�&"OLź0.֚U��X:R�[2/��XQ"O�A�i޼`D@2 �|el((�"O��sRŎ���H�'�9���	�"O(U� � 0r|xS��Za�$"O�6��#`n
!���-w�p��Q"Oڕ
�ʐ�E0�d����9�HR �U� �i[gEfX�X��/�e����2G�(%:�{�I;D��%�;?TPvHS�co���3D�4{C ��"B�����ΖxX�0�j0D��eM��{⍨� ���.�(��,D���S�݂)��c�P*Z��W�)D�����L�1���kBc�i�0�P��;D���tM3T%XEK�K��D�Yq�d?D��A�T�h@�*4ӱ4@Fx�7=D�@ɶ���&`�C5�Q�L'� ���>D�����%#���0T�O#n���z`>D��yuϓ0���CҮ��Ȼ��;D� ���%CqԼATm�` �`�5D�dQL��c�Aˡo\��4�c
2D��"���l������F�F1t�4D�4Z�;|HJ�Q' !_&P�/0D��uN�x,���VG�� �`3D���l$ &�)�ǮO[��y�*3D�|��b�)"��"��8YUk=D�BE���� aI�*�t��L:D�ˆ^&N��
��J-/�`�Ӗ�7D�|2b� VȖ$�0�<�tM6D��A%U,12s�[�8p@Q :D�|�Β|笐ӂ�׮H(��`-D�\NV�P8��%ԗ>�&�Ib� D��BC��z,b<�g��,IC�!�&#4D����_�bG�DaT��
Fpt0��1D�8R$	�E����苦7hLk�-D� QT댻Q�R�B�
\�PJTPR�/D��a7��|Kt��E��.RUn�"��,D�D�U&͉cX�-Y�Gݓ�:�
��&D�<��/W�0��'
���8��G/D�0k�L�� ��#�bWy�ժ:D�	2ǖ�\Y���O&O�)�F�>D�p��cöy�]۰��15;p��g=D�;Ѝ��:Wq�ׄ۸=/"8ca�:D�`�"�$jV�z0�ˬO�Ę( �7D��ۥ��?L:�;�����L(D�x;����m�>�J�^$YE�|8�'D�̚��&Bֈ�S�[..}h8��N'D��!M(Z�^�֪�7lp�Y��%D���5&(#�����L�&�V5��#D��"��r�Z��@HI-&Mja��?D��ؒo	4��B���. 6F�ǩ>D��S0�� ��1�$B�y>i[4 >D��c���$ ^e����QI�ᑑ�0D�h�@:[yжJ��R�灏 �!򤌤d��|jV��6]�	���[dr!�DљD,���A�N��^�8�db!��G�'it1{ �*W~�:d�Q!��D�R��69i�:�nS�U;!�$J-Bҡ0�� &hTĘeF�Z�!�01q���R�s��5!�$YNM{w-Ǥ0I�Õ�ϐ3�!�D1~w��F�;k�T��K!���p d�#$	L�MQ^��j�|!�� ��{��L H�`�@�[s�i��"O�I�.W�x�yӢY�DWde�@"Oڍ���[�$�+���+ZK�i��"O @s���)9�^��׀�8N7x�"OVx���޸w�)p�ڂB%2MH�"O0h�
_���ŃMp�<��"O�e��M�Ɇ�JV��8L1 �"OTE�B���P�f��c�2dE�5{�"O�5Iũ�Z��cÀ�>J�D%"O� JW-��4����b�S�3�)�"O.���$sf����)�h�`P�P"O�IK������T/Z՚��p"OP�ҳ��K�� U�N5q"�ZD"O�e���M4u�\�2��'WB�c"O��s�h���,��L�1�"O��+�%�@�vj�B+�.�
q"O�9���d=6�#��V5�rI:'"O.0�c�Z��4<��o]4
�@X��"O��v	���8���Q��$+F"O��-`a5"���vU��ț#i!��m�l�S��dzܔ����m!�D�v�̤1DM�H��]b�͢}�!��Њq-`�7��"|��d�b�!��F�?H`՘��sN��b�	q8!򄞲V����&���AO,>~!��[9��m��aY>Z�@�C�.�Y !��ӤW��t��$ЪQ�����ѿV�!���y��`��΋�Q��x0����U�!�dM=Wʂ�S �/�,$9�k�$l!�ƫB���DM�.�v�)4�ɦM�!�$�S1l���T�+I�Z����!�C��f욂�ާ'=`�9��}!��2yq���� �x+��1��P�I0!�dɷ^h�q��&����K�~�!�D�*���2d��5�B% d�!�D*&>��kC9w����O�!�d�X��0��bJ�yKV�0k�!��F�$Y��� ��K��,	0Df�!�d	y�ڐs��̩)8�IIq�_'�!��H���`��8����Aq�!�䓄u���Y�h��AZp-z�HL��!��&�A+���RF�M�6.�N�!�d�D���F�y(l�R�Z�!�DY+�U�z�H �'�!�_�Z1b ����&L`�Q�TF�06�!�dP�Q�n�Ae��RQ�f�?�!���t
dH��τb>��3�d��!�dV�e>��Q��CFdZ��C�!�K�Ws.����9	���nܡS�!�$V�OА�hT�	b��xJg��tr!�d��j��$Av�����ɱI�!�׬J-`@r�B�Z"�-8�L�L�!��Hpp����R��[e'+�!��TP1���6IvЁE��.1�!�^[V���v�� aBt�P�V�_C!�	-� �ŋ
 9峧�ÔV7!��LHl��LC1 XΈJ.�'
!��ߋ��� D��QQN�b��&\!�D�d� (�7�?HZ��
�[!�		2'jH�`�Bt/��WC�9T!�dֲ^�0
c�ڠa ���$��7�!�P' Q�l���x��ܪe�P
�!�� V%�� �nA,�L��'�!�$�6���B��=�d[���K�!�� ��ɶ�8&���"�M�$�)�"O4Y��dڬr]Q���!*/%P�"O��Bn����7&O�DT��"O ���#-������\
��S�"O��Ñ)c�X2W`�&pP����"OZ��ee_�8�ı"�5PA�ME"O� ���ق\e>t"#�+~@�@"OP��C�+hN}��Ӓ,�x�"O�m����4��,W�|҇"Ob�s���6��Q�0�� AlLL�"O�0�Gߖ���JU�8wh�Y[u"O0�y�e%_��S���!=��z�"O��£I�3"m�a����̊+�"O�d�tiE�2x&�b�H���)AE"OtiQ��?z��ѐ3e��0�Lz"O���V쏯1Rb<�D��C����"O`��IGKT�icb׍f�ԛ�"Ob=R���� ��'ґl!���"O�a#�KN��:��XM�"O�������!��(���`"O�K�m"m����oU�2�P��B�<�V�Ϛ�Ɛ6J�S�mB�/	B�<��C�TK�IJ�c_�i��3V��~�<9�䄩Y�e� �ʾy�|M�S��x�<��i�?�Ѐ���Z��QP�DZJ�<)R��6'$�ܻ�MK�M��Q�D�<���Ј)N�X��ݣ�"�Y5�@�<!��9w`�`�h�+����T�<� ��.�]���Z(}��@�7��M�<Aţ/&��p'��*���2�F�<�b΀�|T�qB�_��|r���D�<! CY+[�N�*�+~�P�#-�|�<�$���U����խa�)��Iq�<��.ƫK|�{v��>���bFw�<���+�&��p���%d��tOk�<�M�'�p�b6A��Qh��P��o�<��F�
)H%��[�K��؇D�D�<��ł(c�x�/�x��T0D�GC�<����TI;�
�+!,�k!]|�<��F:z�=!i֥9J�=��%	z�<��o�ACL��N��h��q,�]�<�ֳt1��[aߤ��Ç�XY�B�	�ʈ��7�X��rȈ�O�h�HB䉶�Ps�N(�8(p"�1,rC�	�#��H�ѢͷXr�B�b�Q(�B�I$h�8��@��1	�O�S
�B�1E��ƫt}�]J���
BhC�	��q���ڰ�)��'TH+�C�	<j��%f�>��AԆǚshC�8=���� -\�Cm:}bҢ�l=TC䉵�~���/Q� v>98��	�zC����%��#�g�
�A$�	�C�I�q�X`#�Y)o��|!�ǿu|�C�I����Al��a�;&�C�I���������m�#��8�C�	�j �*c I�K~P	�К5Q6B�	�P�tQ1�!~Z��@�N[zB�I=�H��!�\�"!X!�6�	�	�B�I$8�����=�܄s�I��pB�-0�����N�DE�Tx�!I.T��C�I-B���&��Z��熛�S�C�I0RE# .Ũ}mX\����-9[�C�&(r�A�7Ğ�^
�E��/H�4C��7#���Qԭ��c��g$��	[�B�)� �Bр�Ur.�*� �\���f"OLəgCZ/h�&�� �B�(i��"O�P r�L4fb�"�Y��:t��"OL(д$�2X�BR�,i� IF"O�|��bϬmO�2�G�s��p��"O>���Z46�J�ȶP�a��"O���r-��F��߳EJ����"O�� ��@$x`���e-<��"O~\���?b�D9�,��)���"O�����љC��y�r@��U(��S"Op�����N�����[�M�"O�y�AC8X����hJ�����"O�ز�&���,���E ��"O�Q��  �P   

  �  t      ](  �0  7  _=  �C  �I  <P  �V  �\  #c  ei  �o  �u  -|  �   `� u�	����Zv)C�'ll\�0"Ez+⟈m�R~��8˔�DBA��a��/60yfN�%w��U��&��*ADu�mJ�+Vi6�;n�$QA��<�Dћ��n�r�rgȓ��V�J�����l t�T�-�O
+~u�7�S=3�̬�#��L�s����<�D�{G�4ӧ�4��r�BL5i*��DÚT�z �	��:�dIM�0�R�Kݴ�|L����?��?���T��?�~!��ˑG�Z���?�ȭE<��\�X�I�+F� �O��D��$��A{��
2�� *!��ln��d�h�����Oh��B/[' �	׾MD���?zhȞ|lE�Ƶ��5�QjP+�!�7ns�JvB̔T���C�x��I�<H>��'YREq��Q�d䏰�Tu8R��w���qAP6�?9���?���?���?�����v�KhR�kC$��m֯.�^%2�� ��v�h��!oZ��MK���&NnӮo��M��W�����Q��`)#�1�L��#�	^>u����\Oh݉Ƅ_�j)�a��>~M ��(LV�����m@ܴ{��O���������X��\M����5,���� ��n�1�90L�!?�S��LYr�̛)%���۴o�$f��t�_�e�t�#d&F9h���r��R�<(�7�¶Zg��o!�M�Աif���E�3.P���Δ$Ё��oȿj� i`�%�@��
Q��3��٫FM�� ��k��,n���Mc�E�����F반Q�+S5*��q�ë�EM������(�ؔ0P�i� �%�!GL4����P���';�O޹�`�Q Rn���tŃ�x�N���-�O���	۟����M͟Dѫ�
D0.����̰v}rQ�6�'��������������R�@20�Tl�p�*��������|9Hd��蒥)�����5W�hX�B�N�W���)BAXܟ|CS
�)Y>�A6�øt��l��2O�@�B�'2���#�h~d8���9#�1�?����?����)��.���'$�*g� �s �<Z�R��O����gט(����'@1]|��'�'N�OX͸f��Լ��LW� �yQkě$n\ɓ(�V�<��FQ�f��\��(�o���e�[x�<iA.�5?5@��Q�s����a��O�<�&�(��B�@�'؈`�KPS�<�� �$4�R���7�>��'*�X�<��e�TԈR�J��`�F�Vҟ���b7�S�O�R(X�&�[����GJ)T���"O�4��I�>
���f� p��x"e"OR�����Q��@3���	R&"OD �gď)`��у%��P����u"O��S��&6B�CTTM�P`"OL���-�=l�t�r�̸1=�(T��(��4�O��zqj�$A�q�����e"�"O����j�$= L�9n2Ջ�"OZ��P�Z�h*�1���7?V\�(�"OĸjP��7����� e+Nh�<y6����,C�o�r1�T)�"�Jx�[2����M��O��D� �^��� %NJ�u�f�2S�'%���|�Iɟ�x�nZ�N�[s�ft{���O�a�`��Z�Jt;7G8�cA�''�m+�0 ��\y�hR5�BH��08` !  ^�j��w�ӿ�0<��؟H	�4Q���'d�̱Q�A>lZ����DN23.�P����Y�S�Op�\s�`4i�
U�Փ�YC���2���Q��Z��X��:���6�?AI>����6�T��|Γ�yfN�Fh����(I����4T��y�H\�}�*5���߹=z5jǊN��yB�6P�,�*���4�p�9vɄ��y��B��x�@�ԅ8��hUҕ�yb�.	��G�Uy"dhJsn��y��xc�HS�pbd0��I^5.ٛ�|2%��m[���'��'B�	
�P����M��)&g���)��͎ xX��44,��cg�����f����XR�	d"С���
G7J���O��5OZ��5��� �HdWŖ
���wA����Pk�6)��ٓ���|��6nM�!S.O>�hV�'G1���'d�	@2{�,�x��o�ذ�А<��	�ly�O*�k6{�@��E�߁/p@
�Q��ٴ}��ƒ|�O�DQ��P@���W.�x��@?2m�1
�e�;j�0�IU�L�F�
[C�Ҥ����k�,� �C�ɟl/e�T���$
�.��`��8�s(8�x�TAQ�vT-�E�%^b�q�0L�}��$�r����`�:k�t��b��O�� @�&D�d ��"T �h�3ǆ:w@�!A�#�$YŦ�'�����2��h��s�H�
�� �S��Q�H(�I}y��'���'�z��a"45� �r��?(Cn�n:� �E��j��T��4��EM) ź�D�'`�l;"��
%�����P7-���4\��j��H��0� �]axҁ�?�?������Z���9�ɛ!�`$��FϚK�'���'hR� ��%*�ʹ�FA�5CA���
��V�b�촣��h+��� �ͼ�?�+O$L
"e��$?E�O)���=��,��#ԥU��4�G!�=6�2�')��˶JA(i{�\+&4��n:§'��Y(�$˘��"������'P��K��փ!Cf�:��\�?l"}�0i�.X#�5*t
į9B�x�s.K}~"��?����h���䗽a�=�F��8$!0��]�C�	�v�]�3j�;C�n1�g%^)A�V�?Q���.i:0p�6��x�JY�&��lǟ��'	
q�6�O��'��Q�p �OI�@ڌ�cCD�Jaj�F3��y���&=���O�xb@p���y��i]U�M�`Xą��;��|acm�A��ߴ(�P�ATH�g�n&l��6��%r�l�bb��`>h��D~�����?A���hOBL�$�S2F�+���cF���)D�@���]�����Ӝ�`]�Pͦ<���i>y��y�a�+
Ӗ����ƦB�`Œ$���u��=h My�^�D�O���<�|BL�]q����^���T�KRҹ��!M�y>t�2��9D/���ĉ�z�Ɒ��G���D�	u_|���ϓ;����c���N�T���I� vh�᧤ϔ]ƌ��$K<J���g��O���*ړ�O(7��1��P#���,E�L� D"O&��F������L�|�VX�I����u�6�'��I�B��K~Js��2M&����L�2ND���R�h�'r�'��LYJ���wf��7��d�������7
Y
?�ŻuB��W5�T�=O�Y��S���=�bnļj�$n�Z�rͱ������	T4���N%Z��'N�	�t�^���ƛ"D�]��3��O��эs���q� &�X��t�� t}�"��O�܉�C�'k�P�2Eg�;SH ����' 剟Y�%�	C�S]���'8 q
�ۇP3z�� gP��A �'A2��5���O�'�����٦#|��(4��Cޛq���Y��n~��!�����Ϣl^�`�)ҧ��p"�ȗ- $,L�P�ѣ}
B��'GNX����?)��)v��㡌�O�R�(@��l&��È8D��r֩� ��W�ٺ@��%�gh7�%W�>��G�ޭ,�f�� %FQ�g��ۦ��������)h(��1������Iߟ��I�c'�ϜU�Nhz��*,��M3a��9E�lXP��	=�?AP���$�
$�|�<�F<r �@����a��#��9]pT*Ć���?���ϫ	L\!�|�<q�._�����J�h��:�h�ڟ8�'�!����?����ǘP~��CN�V����	P�1�B�'%��p@�oL�����3��A�'�T#=ͧ�?�)O���ъ��!�`sv��
(sL�iR�ݶ+���cP��OJ��O�������O���"�D#��!d��w�daT#�>J���R�i�1)�A��w�	�%K�;tӌ���@L��p�aA�n�r4o�) a{�훠S,=���ȸgإ�E�͆ �q���?ُ��?v/r��cK٥|JR�Ir�Ė:��͆�p�i%R�+葒�!E�&�li�4�?����^���4a΍4���VO3��H����yB��]��ъ�F��2�N��مȓn�d��V���hh�h6�*K��х�3}�̣$/1R�(d  "��Fa�ȓL�J���@ug.m�� n�Ʌ�PC�u#�ƞ)cQN`{�E��[�9D{�����r���)�ĴC�\�g.�u1�"O���h� �RIc��Q�B����d"O�����ſw3ޱY�B������'�Vmے�կ~~B����s���1�'�B���&YXR��!ޗ��
�'���
�%��ah�.C;}��9��_��Ex������LS&�ֹE��dc���.�RC�m�I�� �Z��HЁ[�0C�ɛa&v�Pw�ćC,Ҭ��k��k��B��[�0�)#���j5�Ј=n�B�I�m29��AAb���C�uI�B�I���d.ŋ&�*��n_�C���k�d���	�$j~�^b;�����C�bB�)� FlZ���):�Qjg��2�2�"O> A�V�8��6fC��h���"O��$��:z �%B�$��q;w"O��C ��5
�x�E�$`������'b;�'?�)�Q�5v^�q���GOnͫ�'�@9�S���X �ݹ�e����-��'a�2R-"!m}� !^8t����
�'�\�[ā_-?�P냷�VAC�'5�\��
۳1�Z����&Pr�'㰐����qK�0���d�SQ?��qT�/�v}b�A�J�JԢ��&D�̉ѣ�Y�����k36U*��+0D���E�?.����.G�����-D�����%[d4��닆o����-D��@S��TFh	� ��6����'a0D���b,A	N�>��֪�i�Mp%l�O�i3�)�;�Qd"ќW� +�L�#�����'0z	��T-p��=µk�:!�n](�'��R�ډrl��8� W �	�'V4E:ȋV�D��Ч-�Z���'A�\�2ß͜�ae�W�x�65��'<����JI?N0��qb��w�р.O� :��'E�Hڃ��4A�j�����in L��'Q(t{��1bz��#�ΣX���'�1f���)I�vV'R���	�'��a� �$�9�Ḿ6^L��'{�HA�n��Bi�W��6j|9��I�����\(⁼{PuC��ڔ"�vԆȓ&��0K⨀�^ٜ�	f�C�o��T��jbN�Bc�(D.8�  ڊ`��مȓ8�Tq��.-Y>�
v���	t ��ȓ>�*����Rj��:�I�)bH�ȓ�QXe%�S��8j�DNv%&�G{2 _����@(H�AϯR��kS�@,nM���@"O��"֠ފv���aU��rCr���"O�x;AL>lD�h۲�X+�
�"O ��HR)YSh�DFS�,��qB"O�`c6�؅D�p���+[Jƍz"O��(�
P+K��("� 	d,p��'S�HI����;|��J�e��S�%�(2�ȓ-���q(�<Qe��[i�1@8t�ȓF/�` O��R���ǍX�7�Q�ȓ8�~080lڿİu:RfG�f����u�[0l�2^��ae.�G3D��:k���T�	<�  �#Ʉ^o|��'٢�5G���0�F+i�$�4��)8�N�ȓT����bA�;ak�-�$�=����3J��m���������11`��ȓ/���0%�$L�x* �H5`p��ȓjȘ����Z9~ $�a�X<?�΄����@0��Fw��Ǿu�~𚳡��|B��h�TT�``�'C{!.�z�� D�PY�
��D���[[�(U�#D�HkC��.W������6O�:�w�4D�s��S5���5�K9	cd��0D�\�!��1Ͱtcvʎ@�i��� �|蚵F�Dm�~fX�dǗW�@pȓN[/�y�B- f<���gV�@涀Ȓ@���y�BY!G�>A�%Q)M���3Q���y�'��;s41c��.��\B`��y�Ȉ�|���o]�s����T�yb�G�0w�9�-��]hU�G�P#�?�hEL����¸9�E�#d��LK�AV�{����6D��2��6���j4m��$4D�� ���� %�����+6j40	�"O��J��X+��,�0��gh�IS�"O�I��F�Y�F����Mt�-�D"Ov	f���вG'�Qn�Ш�[�(q�$!�O�����0� ���B�wz��P"O�!���ґo���'P7
~J�0"O�!#�,��`6D%*l�"Ď��u"OT���o��AԱ@SD�w����"OZi���?�*8Z�a�t,��v�'��<Z�'؞t"�v�Аe@�5q����'3p��T�Y������.�LM��'fJ5k�m�V*�]�s�p��EK�'�*��Fe�F��l8F���r��$ �' ��z�Q�X�ce�ޫAkĈ(�'S���M׬lR�-�8w,����d+JzQ?�X�
�>)�ݡ�F�>�U0�� D�@s7@��l��ʇ�(}o���* D�l)��=q�`#ՎU� AxAE�+D�Hb6'NH[�m1��؍j�����*D��k��G)v�@i�#�(��P�t�(D��zw� ET��!��VZX�tQҬ�O���)�'
�@���|X8%�!.�8���''`lA��"1��w"��6|�x��'���!	�՚,��+���p�'9�pbbj.�®1(�h��'� )�Q���R���J�Q�'�������<P �a���W��0!*O��Cp�'n\%̆='��h�@�8�p���'��!�
A6y��� �Ց.�l ��'1(:Ŀ��S,@�p�Y"H��y�㏓���M�&4as6&­�yRǆ�}�� �� Δ`@wg�%��>���Z?q3 �����H7V|�iæ�c�<A�N&!J���^�*��T��Ny�<��H ��83����g�a�U�x�<��`���\��"P;a{d��u�<��g�4���ݴC�J��f�r�<ٳW�f�Aӡ��Zy����kC�'��:����
=2V�2���V`�e)݋\!�D�k�N4`
]쥹pn�4[�!�䕤d&(���-(_p���G���!�$��1C����/��T^<1�A�K!��[d�� e��!s�58Ո]�-�!�,�EP��JlH�Q �0vk���O?Y�f%���CAHXom+M�`�<"V��B��M ���`�<�u��Tw����^q��u��N�V�<�dȃ�y�l���,T��X,�u��H�<AP��,�t�����=�H�b�F�<���;��FC�hu4�ACCy��ǲ�p>���Zd��!���4�s'�e�<cQvo��q!c��f[��@�,_�<��Ԉj~��P�b�="l�����AE�<ai��@�T�hR�ĶT���2�HW�<��')P<Q .�6-�F���o�kx�x0�����5Ő�*�5�OW��}b D�L�b	���
!�S7W�vi�`?D��*f��_:nt(r�V;d9�G�>D����@�w�ų��40�~e�C�7D��A4�J�?O؁���U�=�8 ��5D�����($��eSV��!g�l:!
4ړ/�^�G�4ƀ�,OA�N�D(yH�8�yb
[�	0G-yR��8'���yb�I�[�`��I�5xl��6��y
� ¨��*%���®�X|~�{"O�HU�YB�<l"Í�lx�j#"Omy�D4:F<F�T�f��J��'�������SY#���]%6v�X��1k��%��o�$a�q�;�f`Q��Z/G*I��_5t��H�<.�<��*�*=�� ���A���"/�B����(zm��ȓv|�5ѧ�68�qeF 4^�-��sD���5FF��(�6@���0�'K�Ly
ap�ӎ{�}�L����.X8�3���b\4�b�Ύ�|���N�p%R��ʃE�R@�螬7<�܆ȓ]�sg$W
/��m(�l�%Rd2���
<x���1M*� ��cZ$0�!����O�b���8`��H*x'����JR6�
C�ɔB���#+�=S�)P�E�"B䉧V\�xaP&�f���B�n	�<�B�I,w�©I� ��@��;�a��rF�B䉴m*��s@ţgz���F�.C䉆'Ex��dD�Iv)�s>\��=�S�n�O=��Ȳ
L?��V�
�3���c�'��{C�Ǌ>�Νk�W�/ںܓ�'n^��A�	&�q���K!)а�	�'�� Ц�^�m�r��hESp����'Q��*�=������M���'��Py���<#���p�ŕYd6l��h�5Dx���	_t\Ȃ�G@��<)բԟ^Y\B��[Gr�C��R?s�,-�/ߵw!�B�I�D�(�%צU%ș0�)
�;o�B䉴E�P��� .,��9%L�\BC�	�giN�!g��%�YX�l��^�C㉋i�B�ʁ��Ir�q��oL� �ĝ�I+����#	���&K��I�B��4�@P80Ț�B-�c�ɟ����O���O��!�"'4�g&�O����i>q�2,Y����Q�Nz�8af�)�&>���ƍ���H���Z���)�?Xn�bcbXB:��yd@�%�����O(�!���bx�glC1�43�	�$b��0?��BD�&u&l�u�j�0��FNEx�`0)O��� 91��T[�n�א%��Q�`+�l���X��Ay�Z>���� IS`��,�ĭ��*-kT)A��0�n��y��U�2��+v��,r�S�O�2"Ìҳ&�0�8�AD�WQ�x�'���"��tP㗛 ��?�p�K�'3 Լ���g~:xQ%k�`*B�O:��5?%?y�'�r�b&9�(��@�S|8�a�'2FDЀ�6u(.�a� �R�b���dXs�O�q�5Ma���+J*Wjʈ
��'���4N�)ڴ�?Q��?(O�IS�p�l�!�Ҕ]r�t�r`�L�U���O��H��G�>h�ax��Oq��=1�G�x�����LD���A�O�Vɱ��0^<��b�.�j���O�Y�P�˭:{X�{���Z̨�@ᔟ����O��$�On���'!����'H\�0�F��T��y��Q���ʷj��]�e�"!P�X����	�HO�i�O�
6(��UΛ�[�BA�(�1"-���
ɠ䛦�'B�'�)擇+��A$K�\8DigH1hh	�A��E���
Fꦉ(�.�8��u�Ζm�����ټZ�P�r
�>H�@�8�d��9�Hu�ϓK�@��	�=ƀP�`M	TJ��b� �;O��������?���I\� ��s�=|����2_�C�I�:���BV@��aXY���o���'��I?Mb%p��D%R�C㒌�����t���o��!�I���I�\fd�"��.�m�tܣ��|��'Q�G���7(�[� mp�h�J�'!*���ܖk�Fźq�^�:��?Pi"ڑ�F���%NV�%#�">�7*M�h�IW�'u@|ꡩ��L✽�&GϨtY��'�a~��4C�Ȍ2`���0# 9j�� ��>�Q��0��?,� 1S�Gެ\�ި�&��<!�̌�y����'P�I`���'Q����c�����8���15�[�A��B�(�"+Bw6�8�'�O?�i �M&)�b]����x�n�3
a�$�q��T���H
���4D�4同>,���b�Ri��
�Ʉ�y�B)�?�������$��� �{���I��KňZDb�iP"O������,�rQj�g��g,hy[�퉸�ȟp݊��ΡD����hK���� �Ov�C��X����?���?�,O���8S`p:�B��C4�3"�H�wA����O��'�N$3=B$x#�?#<� O��/�h���䙌)k��aq`ؘ>� ���7 vm�Q��%'��O�u��\�g���h|0�V��,����OJ��:ړ�y�D2G�Z���+B�q'v�"���yb̟�S��Eˑ��lm�=
O��?���i>��	pyFO�"��mC�O�" �j�kӷ>^���'�2�'�bQ�b>�CM��]��EB N��%�pP��%p��Ag�7´R�炜��<��OF� ���ñ��=��hE�!A�\d�G/��H�����<)T�G͟��pJ H��j��n� �'&ZßE{b��7:��d�¨�8>1<���I�
B�	�Y��!i+<�����`���"S��'x�>[x���f�$c>�+�śj;�%8uJ�'&�:��OPФ��Ot�d�O��R�/�z@�9�nK���4�,8"%@B�#�-BE)�#K�F�q��p���t�	�U���qO|�S&�4?v^� ��,�
Ѓ�h�'t�D���?ъ�T[�JIzI�5�ʙ�7�µ��$9�O�u`r)�!�t����O}R�a �'���`G���
7Wa��A�K�",$0�'�R�'�R��8?	ǌŖ\D��ۥhN�Ux�r�C�~��F{�*��!�T�Q� NYE˓�6��'|�v�x��ģs�T%'"@k�z#=T� �'פ�I�T�lӧ�9O��W%�(���d�6a��6;3��lR�{Q
�O��'>U�r�_-\�ƨ!Q�\�,q�%\�*��:G��=��<�w�A<�t� V��8fײ h4�P�b8�O��O�ۥ�>��[?5�F�5Qz$qA��H��C�O|�Y�>��
J�O:��RF��=8"@(�@�ղB��%���'c��{L��#M��H�=}��h�4����	M�~\)��P�V�v��t]��aE#})%�'��*2HL3B!Z�<�H"��Q�S��[�
.�S��'��,P�Otq��m�,�t9� ܾ)�!���${�2�q�X��'�|�D����:����tE�$oY�a�K��?�C���`�L3?��y2�נ�~��]2vR�`���_�/G\ԋ�����?I�.�O��`�K�\Y��gG8=UjE�"O�]3��Z(8�0��� ��6iXL�v�i*��|r�~�'~�s�"��A�&@��"o��
d����V��$�,F{���QR"j+w�4��R�S�aOly��"O��1A @�A-2�#v��;�ܠ�"O>�zC�����B79g!�"O����>0ߊ���d��iG��"O�Q���}`�=:��	+:�Q�"O8i�!"ζv�U��
�i	��Q�"O �a�䵩w��)�P5�"B���yB$G�`򕇘5W~���1�D%�yb@�P�� ��
�QGҀؒj�y2g	,Ӿ��g=_�VHJ�!��y"�����S�I�(KF��6G]��yr�Uh��4DD�+�&�f��y�fS�|�ڱK�"��#0��i�����'L�]s���Z��G��+WVD�;���0I�� 
E.Ⱥl丩���3@��Q�A[-$��k�%B�M��N�O}le�A,ìX�h	�a��)|�l�Z�FT3�
�*�)�_���2ƍ��ܐ��؆H�Q������bF�
\�HE'\�4�9��MT.5W� [K>amU-,`���C+9(��KB�<Q�\�/�(<��H�2.��1OI|�<ɵ23D<�"��R/6}Bt	�E�^�<����$�r�@1��6+��b��\�<1���1iHmX��[�D��T�YR�<i����.�2w�+V�h����s�<����8'�>̂.�#y����ao�<���޵c�Qe��M�l*� VS�<A���.�ƬI��0X=��qE�X�<�t��Z�X	e�N�?�`���XU�<��LIq� �JÄ��mq�/�T��L��8�Eʋ�SNzQ��a�9/Z8a�ȓ0�6Q�Mܤ6�D��+2Q�=��S�? ��	� �񉄧�-[�ya�"O|�2���"��]S�6/[��q"O ��Vg]+<y�tRq
:���"O�����;	�r!�R).�6	�"O֌���W�Od��)�3ژ4�T"OZ������@C�%
�'�@X�v"O"��r	�$;�nX�N�%�����"OXԥhD�&��$�H(��"O�5 ���T�rC�+��d1�"O��
���("�a���b�P�0"O� �5Ƌ>m{>麂���,�"O��	s�\~Z���Ň�+; F��"OB!Ja��
up� 2�J�Xm4H��"O�`�dN�,P�En%XkZ�"OB�;G��e6��9.[%qw�iX�"O���t�6X�����-ݸX���@"O�<x�Q-���0J��W�r�Q"O���#I��S�� ��Ì��\+Q"O�)�m�/h����({ߨ���"OLh���|7JP�`� ��"O�賔m��GQ�� �K.�,�6"O���ѠM&pa\���*Q��:�P�"O��E���E��D�7�[��T��"O؉H )�+��Z��[�4�
yy�"O��� KG�48�����c�>���"Ozt/ץ �P ���;4����"O�P2�G�W�&��/WX��-�"O \cEHJ����6��x���aW"O�D��*�	3.ā/��"O<rtl��\��!g��Tˮ\�"OT����|2�%؃���ZA*""O�!B�������B���� H�"O"���J�rf8� da��M�\U��"O����$��
FG'~�Y�g"O(IբO���R�_C���"O���cLB`El��T䇀	Uj�`3"O�5c�5����֘h���s"O~A�� �#���.ʛ]O�tS"Ozl����sҠ��f�(FN8T"O�ܨ�# �+�*��KF�45<�g"O����c��bdt�ȧO-�%�"O����R5���+%�A���My�"O&$��/��XQ������&"OA���ړ@���� g��!�q"O�ԛ���9��#hֿz�����"OJ`�D1VB��BgΌYЪ��"Oh\�6&�:�$SV�@7n�D{w"O|�I�'lU~���.`�4#"O\LRaEX�["9��Ć&U_��b"O�HW�s2�;t#%r*`��"O����֞;�6�@4�P�0e��!�"O�CP�ɀDK�(xd�ӉB���K#"O0����>3,l<��IĥJf���"OF0�&�ʝS�2uP�)T<�`�7"O��z6#�=��a��f <��UR�"Oؘ
���?rФ pgF��d��"O�}낉EU1��1UH'��H¥"Oڑb��B�d���-I�nqɵ"Oh-ё�Y��9��J2� �"O�,X�k�A��x ���t��Y�"O��7(��W��-Q!�J�9�:A�"O�aߧGK:���u�b�p�"Ot=`�Ǒ'Q�P<�!hM*�Թ�"O�@0WbLN|�R�銺DzVh1"O� �+��*+HT�s(O�o�D|"On|@�ņ	�Vh�&

�F9"O�4�3Ɵ�v��D��.��3��[$"O`�rAd�*�z��I�	o�x{�"O,�Yf.-�f�2��-g:�Xf"O�����ҡ|`�Rc'���p0"O
d��C6(��G �B�q"O�`I�(�3^+ā`��X5u�ꘓ�"O��Q�)��=
�n�H��C"O>d�C$Qٚ  R��+B`]�r"O����9~���]#J:��`�"O������43Z���"\3hh�"O�y���M=i%�	:d�ө:V��r"ON�8�DM2T���U���,�"O��0@J��b9ubdQ��#6"OP�y2b�bZ���A!�*Jjј�"Ov��T�h��t�M�U)$���jĖ�yB�� f����(9c!��H�h ��y�-�?����hV2Z��3��:�yb.��IaQ0/��"&t�qꅘ�yb�R;���I�L�/쵐��Ӷ�yr'�>\)D��5mI�f�hA��3�yҠ��`!�
�яul DT��y��S�a�~� W�6X:�TnC�y��L�E��90�L�s
��s�6�yb�@3h���!�&���ȕk�5�yR�#b��	��~�X�um�*�yD]���22��A�䜩D�P��yR�-O�v%Z���	*l�j�o��y�I �+�q�M� Xݜ�1�d��y��<Cx�\ؔˍ)8�N���C�y��<in��Ú2#����+�yb���vB���'*Q&3F@�5	��y��
	hy��/Z�:B��%��6�y�	�2��RC�=*��3���y��O��eH�)g	��.I926x����|c���	�Bϛ�ɇ�pH8�gi��RO����]�b'�`��\}���]$e8��&�5M����ȓ,�z!�Fa�4'�@T�J�XEz0�ȓL�r�ۖ�W��`,c"�^���ȓ]I�2��
&qG�Ia�R ԅ�'90m�"�L�t���N"���ȓe��X��͖4^Ǿ�U��*C�t��6!N$Y�NG�=q05�`��H��܇���q{�Ƙ:;�$�å�4�^���.~�x���RL�(�.���9D�0Xa	IIw�y��L�`1C�$D�,5 ��ED��!�S,h�4���"D�be)nd�|X�R&<\��?D�X #o��;��X�`ݖ	����o"D���"�R�e�X4�'#�aǸ��ӆ!D� �eþT�b�%����#�3D�HA)?mQV ��E7���B�2D��zƥ1��Hk*C30��l�P�+D�����
'P�������(N?�P!�*D��"Ԃ�H^:�#!���֨���:D��Ð$<�r8т"�"�X���D=D�H��
���pr`�P�5�|� �l<D�lȒ��%o �}�E�Z����:�7D�p��L�>9������}t�Q �'4D�ȻP�G^ak`?���ӥ-D���v-C�\ɖ��Q�#lp�SV�8D��j��7�x�kL�G�$D�� �z��O�"TQ1ۇK̄Y+�"O�1� �tG���1��*��1ر"O�]3S �y�`���x���"Oa��$�:9�T�,Y�X@"O�U*����J����唉]��"O�y�����i�D]�B���ʂ"Op�:���:W\3�Dֶ�bhq"O�l.`.\�)O�!��p�D"ODE� I
�+-l� HʐfH+5"O�AasGA.e��z���4�x�"O����iֻn\$���Č�=�c"O�|��P�����.ʊ1���"O�a�&j��8Y|� 5V�~��@"O(���VT\� ��)Rm8@"OB��R�Y�w>آ��K<r"�0q"OLQ�����
�[DF�s|��sb"O<q
�k��H�� �ΚSi�4a�"O��цhӵg��=z�+σ)i��j"OF�X0��8��@l� AQ�؉g"O.MᷥU4���!e�FF��	�"O��YT��_�vH��
@cx��"O\�w��	f��5"D�)��"OHк��p�F���ȏcM�!��"OJ�1$`=LefKS����9�r"O���oK�z8��	^; ��"O�p��h�5rN����H�R"O�����	����C��T�~\��"O^�3�I0K�̥#���u��$C�"O��č_ɔ�B��ٰ/��1��"O�H��#�L�X�ɾ@�0��"O����G�%���C�uʠ�9$"O���TSZ�	
�832"ORT���'IV~��c�)N��D"O��x��P���̀�d�����"O:ݫǎ�'9S:�'J�.7�NA�"O���� ���
Y-M�X�+W"O4�7��s�R�Y�(c�)c"O$����+yE�;W��	�Li�"O�	�0�)`��#'��9�tի"O�E�� ͯD�Ys`�������&"OJh`@�"'��訧���6���"OvPP$d���`���`?+���"O �a�+{&TȒ������"OT���Ɩ"q}3���Y	�(��"OXź%� ���s�N;Vd� "O��� �<GP)kE�PPըiy"OB��⛜tcxm���0g��JR"O��`r鉗/��ՋZ�J`�� "O���c�?n9�zp\l����"O�hB7g�6&��{'�ճ �
�W"O����舃`(��@H� $�NՃ�"O���6�X:�,d�$��'��I�C"O���2�H���)��+2ݔ)�"O0p����`���b�Hu�B"O���%C�p�������n�4i	�"O���Zk����`(>?J`z�"O���Ӊ��u���U��%.�H�h����@d�4�B��nԔd�q��"��'�v�jŁ�>RT�����@X*�H�'�b�I�/RJ�r�ʄ�ހ
t��'�"�����/��
d�Q,z:^	8�'�pB�O�$[�ŀWBT�q���'�"P�!�����[�?��	h�'�Z�QD��6A��!�Qbذ<0�'q��ࢫX�#T�b!��K&�	��� �5I���.i�l�%���"��V"O���2�ɋ4qZp	d�χ|dj���"OV�����8;�2&�5~>����"OM��J�H��
/..^�a"O�A��F�Ik���@ߺU(x3"OQh"'Q
*����G��	�朊�"O$Y�LS$*G�4�G�G�\�,��"O\1���$4��ڲ	�G)F9h"O�T�%��6?RJŪ��>ZT�U"O�|ӑ��387�C���B���$"On@V�P�1�,��MQ��(�FJ�<��X����f�M<�2K�)I�<9b�&~ǔTk�C@0`�>�ȅ��}�<��]�v~�9I���1D���D�<I���<��u��O�i6�����_J�<ѵ�N1����L�J�ș��Hr�<��E�c=�����v��hЧ��O�<YS뎘oAZm
��ECfA�d�@I�<!tg^;m��m��Z$db�FO�<M�;���IH�Xp��FJ�<Q3+�7F.��C�U�������@�<���ވ:`����W��F�<CL�\n�0��q�
P��\�<	�b�'|h�H����>͒1!f]O�<A����x�d�o"P|��
I�<��_�9;�D���zL2�� ��G�<a��еBe�������)#R�@�<!�FώB�@D"R��4/�Z��U�<�7B#b�=IRϔ.u/D�&#^T�<��%F�D*��E����	��H�<�'�@�|0ITf7Ji�U�;T�T;�GA]�
��e�No�����5D��be�D5�N`����"n#�x�3D�����'�x4�P�t�B�A�2D�(�����8���U�����c�<\j!�d� �\�EŎ΁�d��D[!�d
𲁋���/�L�T�dV!�D�&|i�f�Ox�H�Ԉ�!�d�d�r2@#w�LHB�#!��<&��a�*�9H���
�B$�!�$��7(�H%Ƅ� ��}�'d���!��%gJ���G����d�$x5!�d� ���G�
�lz�P�a�"O��@ߘx᠐%
W�Z���q"OF�1R�
	(d���IA[��-#�"O.���F��ACǯ�S\<-"O:1�-	
!'*DQE�S��)2�"Of0�2�S�}�h�*q�D"&�$��"O\ K�f�z��q�!e�nA��"O$�  �B
���X�LΤ�+�"O�uYv�� T.�`�.�&WP��"O���B()D�]�3ۈ)�䊲�!��,����2�L���1�V�w3!�Ğ�A"L�yb�Z:}��z
�/!�dZ-9������c�z=��c�"OZ)�7-No�XE9�o��+����"O��)��Y����`'I>�����"Ob����>e�h��U(x6�
�"Oh��BR�eӎ�0��W�x��.�!��� �2����f]�l� ��P�!�Q�|�Hբ�jíY*Ua Sw�!��`ĸ��u��@k��#�C6�!��]�L�:T*AU�Kg�&�L��!�D=� Ȳf(P2[�d���%N!�� ,���-H�����ZcW<Ͳ�"O
<#p��&y�:1 �+:�a�"O,����4?�x���ڥ9DĈ0�"O$"2P�4�40�UG3r�X�cG"O\��t̉�k�ʜr��ѴN���k�"O�tQ$�O���y��ѣR^���"O�A�7%�!�I��L�1x��V"Ob�b�n�t0�%�޾g�r��"OR�{҅���S��C>蠁�"O�V�d�"y�	ʺi	�(;�J�<���Y������7(t� u�HP�<�$Ɂ�G�^�aO1o$��0ABo�<)$G�*TJ��ߊi �0��Vd�<�#��@`�=��Ц�(�MMZ�<�4(ׯF�J�S�ˉ$���r�g��<i5�[�_�����ʤ���<��ٜ����<x��cQ�~�<Y�ڢvt��S��[��ċ��C�<ٶ$�?-� x��K �>4НS��GC�<��ޅ���a��:��aK���u�<)ѪE�(E����6&1����^s�<9�M�{D�ш��~T8�E�U�<rÈ:x`�9�ǞWu��c�%]X�<�o�8�<�Y��-6�0��m�<��C�$
��ivK����� (T���2恧~MbAFM��bu���*D�����(aT�Y���J�\����,D����O�-4����e�+���y�f�r�E��ʣ;�L�CA#�yb 2/����Sd6��R- ��yRą*�$q�ƯZ/9:u��@��yrCE�&��x0�kY�4,X��p���y��*V�TCJ�`���@FZ��y���aG
��1'�.6`������y��b4iW-C�8?���UF�y��8RJ�a"�fz�@�mR��yB�V�,G�xW�#lu��$���y�K�$@�i�P)I	ke0;į_��y.΁ �0L�&!Sn3�`I7��y�кD�^�����=.�ǬS(�y� �:�|�$��#쉡F*�y"ǁ7X)l�3��	�!C|�"FON��yRWI��\bQ�/]h�3,N��y��H�s���@��M�b� ����yB���nm20���R��|�q�m��y��Ύ(0�E/E
wZ��J��<�y�E��Iؐm)����p���x���	�y�C�
+�bmC� �pt�ȣB��y� Μ.X"�۴��g~�8B�ʒ�y"K��\I�2�A�4�>M�%���y�.�%6�pT3F��'�V%P�C�y���v�"�ҰK���5yA���y"��7~��H�$��	���F��yR�[�6b86��t��0YP��.�y"�;B�L<ӄ���䦉��J��y�c���Ba3��S��@x�3���y�ǁ�U �ؚ@���@iyb� #�y"� U$���!�.Ҵ���_��yB$F+
�q �"9ԅYBJ���y2�
4]^R�  #�l��cBeN��y�&W��� I�v� ���M�y����bԘ�ʚi��,h��Ϡ�y��.,PM1SW��b2�S��y����!H�t����+�֝�����y
� ��ñ�S03M�5c��Ʈ�@T9�"O�0@#�+A*]A�M�#�t��"OH�/ .P�Ѓ�@���ڢ"O���E�M�c��q�4���#�"O0DbWj� /�Ra�"�����W"ODX�ֆU�A� ѩ��+5�8Q"O�-�o�5.�S�*�?�L�s�"O�bg��^��B�(B�xT�v"OP#lȁ-�Vm���Ʊp;��S"O>���;h�����%1۲�z�"O�ܳt�\�'Z��3���(�r�%"O��I�BW�v��� �՚V�\D�"O��0ӈO��r�r�DA'�C"O�ih��ݨ#l���f�#&�q"O���F�F2�rZ�D�x>���"Ot��s�ǣI���FD߽ Lҥ"Obt�䢗�?Ҏ��ej�z|d�A"OR2Oړ k�["	�xJ�8"O8� S�Ɓ<�:�n�#��)D"OF��c��JL�'� �!b�w"O&az���z&m[���*R��С"Ot�Q-��m������e&&8�V"O�y*Abǂr�xH� F�u%�8�"O8�d㝧���(�S�\�"�c�"O`v��d�D�U��t�|��"Oi��	�~0D�R`	��p��"O����a���U�Ո���H!�D/o�2��AIZ�!	��+��p1!�D@"_H��d���<�e�+� g!�D����%�"���lġ#l!�D%R_����A��g#��*���m5!�D��$�X�*g��Y-"8R%��.'�!��8`Nx�!�� x��2L4K�!�䉺c��h3Q�6+��Y�rmK�&�!��ن&!Z����U	A�L�����'=!�L&hP|[��àQ�ఁ`��z0!�d�G���Q�NC�nU�pb׫k!�$�<�x��蛃�@}(fh��.!�$��C�*��MH(4��3���	|!�[�T������D�a�����M�??_!�4ܴ](�K�4]���[�#��;[!�$�>
z	{�X2.�dY��on!�dPo�ʃ*�̾Y��-�jk!��Nwb�i��L	 5�`S/�f!�^�2��pR�L�_/�<9 	;O�!�ā6 Wؕ[�kZF|�O��!��ە�.��V�/9�\�(b�@�!�A#!�>�:`G�A�"�8��Ō3�!��
}����n΂O&���Bǟn!��D�G4l-���C e�iѳK�@}!�d�kT]�]
A�Z��0`��w�!�$����k���i�dqł(D�!��Px̱r����9��	�!��-7�`��e�2�J�3����!�X6ɨ�?m�i� B-2�!��φ%H�����5����� Q�!��Qn��-JԢ�S���g'P1p�!�$�qJ͠p��]���	�e
!�!���(���b#L :�*4���%}!�S��ճCl�V�C���G�!�V@��a!F !����dW#�qOH�p����q�� �
!20�`b�|2c�v��P,�8FIPC؉�y�n�'![�$�DC
"��8�-��y�-@+aV�3elI/"���0�y
� n��*�/H��mc�%P6Q�� �b"O~�iF�׻`'����T�>|L첶"O�`I���.>| ��!���\�Nq�"O��h1��D���A�JO�h���"O,$Ȳ����W�)8X��D"O^5Q���J�AMܫg�)
�"O4���'H�4 "�Ī3�z<I�"O�A���C� 50�hp�6X��"O�D�w���V�T`�
�l#�Ѓ�"OPػVJ�?b��c����R�"O49�#a͝>y*�z�	��3�ܙHG"OP|"4씦~a�ֈ� @"O20d�րl���(�a��A����"O�M�'�	=ͤ��e̝Yy��b"O���Df�[�,YQuN���Dq�"O^,Q��E��Z���&Z���"O@����y
��`�"OTP�ƣ�#���$�B�r�����"O�%c���rT^�*"�H�0R��t"O�D�7*���لCCI-t�"O�����(Jb��@$|�4��"O��ӡ^���#կ	\w�e[�"O��7Х/m�9�w�ӊ1���8�"O!��@Yv�^XjG�A�D�bH�"O��k��.qe�Q���:ua���`"O��1�R�ap�Ñ!B�.J63�"O�lj�H:N��x�FF7��@P�"O�:���U��	�A�O�(�>T��"O�'�Bf�5)�oܧ2w�IA"O~y#1%��r���� O�(@]��W"O��J���)�����NI(I�S"O�XS��=��p��7F��"OjY0�
���� Kwkb�д+7"O��	C��@����dL�5_<�9Q"O�8cB C�x�6U�J�q:�G"O�´EH*����i�	�^��"O$u(��=�x ��= _:u��"O����B�;���j> 8�"O 9j Gч{��<$h$FMa�e"O���C�a�N� ��L*se����"ON�����;ah�!��H�^be��"O�����bC��ʀ�-���7"O���ʱ_�䁛�B����4"O����%1�����A$c%�g"O��AgB_W�fQ�V�z���a�"O�i��
T��b�eݍ.8�9"O����	��R�CW	m,�"OD9k#��+�BIS2b@�x�
�"O��8��"-�9B3 G�3�ƹ*�"O<Z��S�>,��O��<�tx�"O�tS����`J���&o�`�"O0��e+=�t �m��!�x���"OI��*���q�F�%����"O°)W��A{|���D��\�7"OUS@��9Xw���ΑV�~�Y�"O�=�P�����MJ��Z�xQ""O�HʅC�8�jR쓼t��p""O�k�Av��XANNEȮ��"O",�'*N5ev<��,���\�G"O:y����:��U�G��i���1�"O,�P��Z�p��ݫ�#��2��Q"O�1!�f��_	��EI�:a�<(�"O�q�D^�C�����Е"O����Ɵ6}1H�#%�ܯsA���"O� 2�3��	�V���M."xq�"OB8f*OX�����>��A"OZ]S&&� wb]0gς6:�e�"O�hs��@�h}Zd/ǌ$����"Ohi;G*H!k�>�'�8R"��3�"O��)RH�1��Ȅ �9�0��"OT\��-)I:��ӧh�;��Q�%"O8�v�	pe�Cr�R�S�j�B"OΤ�P�کg@�cԥϥI����"OҠQoQ���h��6��̚�"O.]Aqf	I*���QAȐN�:d+�"OH��J8w�b��Ə]�L)�"O
������x�'nQ��X�%"O�4Rt��J�� �@F[��#�"O�� c��HC����ٰ��"O��b ƵX^\�Ja�<)���"O�)�b��2�m1B����G"O���B�L=^�R�Q��S���m�"O�u;���~�8lÃ��8��yBd"O�4I���1�n8����kNve��"O����%مa!܄�K�
6L̛�"OƤ��HŎG�B �R7�Q[s*O�jS��5�2s�@����A�'�cc�߭>pF��A�[�z����'��{1�ūrb���5��oA�x�'&�*5#��$����d����'��I	U�	�$`b5�O#I��) �'�.mk�"l�fQ����:B��3
�'���K��E b#���s,Y�4p�XK	�''�Zt(h�@y�+�!u�[�'��=��(�SJ�S�S�g�4h��'e|�Ct�/n��)�� \�Q��'��$�w$  >t����n�Ѹ�'!� 
_�G�B��2V6}�'g =QEdY	6
x8�e\�.4H
�'.�	{���=�@-x�H�%v,�K	�'6�L���7:��Paf杖u��'�������l�j��a�xͪ�'���$&����\�AF�-bqb�'�.8q@��.Lg���M�7&�F4��'��J5 ���{!�"�$�A�'�8Y#ǝu��$kR�8�,Z
�'h�Eٷ`�}s�M
e�0Ӷ��	�'�\Y��/T�B ʡ��vF(���'�Z��%��֭ ���n�� �'RX�22�ԉTh}	1k�`j��'����Z�>�4K��	^5z�b�'Vz����!Ax���ǯ\�^�z*�'5<����J�c���a	Mdwzȓ�'O�5ۅ��/g���"��\3�'��x�ӭ��Dx"E�1n���'�$8�1�	?�F�1��5��'�T������3�)1!�<��'^��;E�P4Q�=c��0x�X��'kظ(�ZW`ʜքE�+�tp�O¢=E�T+$b�L�rD�ӐdM�H�g�T��yR[��� ��Rk���u�ȓpڙ����t{���-�9MxA�ȓw�fPi���7>�j����ӵX"z���+S<0��U�Y�*xҲf��,��5`V�I�A��yF8����ܭOwpȅȓ.~�C��/%�Ԙֆ1z�����wb}�hڨw����+Z��ȓ*����`��@�i`�Q�$SL��S�? X�B%�(-��4A2#��P�"O6�٦.�+�d����Q��Q"O�	�dlZ����Oz*���"O��x4�P'A�2������P@"O^(��FSM�t��2��h��lS�"O뇃 .V����͉E��t�"O�P��j"6�>]qEL��}�"��V"O\ixc���^���
H�2D"O�X03B��بƮrjJ���"O�5Z���� �.�sEh0+�p
�"O^Db#�EM�.��"�гi&H@3�"O�EuB�=b���r&�K"X|��"O�R�^�I�}qQ�	V�l��"O�e8W��'!��U8����""Oz��U���:f$9i"��V���
"OJ�i���,�č��͖)��i��"Oh�`��' �@	av�Y�*l��A�"O.QY@��L��s�+A:���"OdP`�X��l�1�c±#(���"O�90��.gP����7O��0"O�1�H�0�Q�t��>�" �"O
��q��)T8�����+3��'"O>�%[�&���V�H��E8�"O���cș5�R�H4g�r�dx��"O�l���h��u3�FRzp�"O�� �B�M+�A�ReߏHY:X�"O�%:��͕f\b���dx� ��"O�52�J;x9�3!��-jX$"O>�KH_�`:�ա2�D�b< d5"O�}h�+�yd��*���,YȰq�"O� �ٕY[,���֔aM�\��"Otp��l�j�����G(����'D�TH��ؙw��9
��]�p��9��)D��H�υl�����o� �I�'D��{E��::��D�n��9����� D�����u���!g�V|���rd?D��)wmG!�tC%��n��pH�c?D��`f ��s{�؉�D9A�g�;D���WJ�H�<�uE�.m�(xPF/D�<�TC�gB�0�#�"W��R7� D��7�B�(����kI�%^�C�
2D�0��Ϛ�r
P��ň� �S�1D�j��՟ul�U��-΢<� ��G�#D���UG�>��z���}���q�f D� ��-I��%"P�5C9��Z�=D����E% hc�)��S�Z���&D�T �D�i�ZՀ��W[��IKA'%D�����Ua08���R�*��<�Qn.D��xË�;o���C@x��j+D��"�*�u�J<�1o�s C+D� 1�m�T��It��$��l9��6D��j%��8�@�؈E�lip"3D���" �@=�"��@���2D�[�J�-̮)�qh�!j)��*2�/D�T��ܲ���߁e%2��&�-D��;�ø* r��qk^|��*D���fc��B~N��&O޽ ��H7#&D�4�ԂA��f^�I��$�r D���udP(�'	��X��t���<D�8�dՔ4��1(���4C��C J9D��1��9@�P�ӰaX�Z�:76D�𓰈��#�b�*h�"MхN4D� ��,?<��� u�aR1>D�ԁp/Q��
��a�>$q�C�)� �*5��i<����Y#2Y*=J�"Oz�1���6�|y����3QVZic�"O�}�O�+Q��p4�RHs��"O�$	T�Y�阄��'�,Th4�"OxQ'��/tNt�򧖐S�nTɁ"O8��F$"qo���fF<L{��D"O�)uN�a*�;C��<wpv�0�"O��ҧ�={o�e+d�>R�^];�"O�G�SW~t�RF��Kрɡq"O8 �$�N3�)����F�)3"O~��Z�O���11d��Q�F���"O�`�@Dʙ�
��#N�v� "O���,�^iQ�lվif&�"O*ݛu�J46���r��-M��)�"OJ)p�t�MY�S��x�����y�E̎d��+ .όB�d�*נ�yoB�,a�q�$O+�(�ZW&�y�̊DG�	G��~�*ٓ�e�>�y��O :X�@��@�|�H���yr��&��z�'\�&7��S��F:�yr`�x�h5� ̐O�@�3�_2�ybO�F��M�c�	���F��y"��I+�USa� tL8a�lJ �yҎ��EL����Ѫf�@�tMC �yR���>p1p�ބ\���g�5�yR��U��H��%��^D���1�Z�y"�D�=�=��"�&+� <c�N�0�y��}�F)�(ΓX.b����yRo�1��82d-X$���q/��y��[�!��8���$�W��~�C��8Y��, �]*�3��v�C�I�cw���VgD="��'����C�I�T �5��@�&vu�7
��!�dB�	~ٞ@;�a�.�JI8���5	`B�I8�z���ђ1�F9°��(B�I2Zw 0Y���-L�1��*7B�	$tAk�6������j��C䉜���paL�'h�q�-E� ��C�	�#.����j� 6ŝ�f�nB䉭8lp���]�t!V)�'�i`FB䉔�`�"�±h@>	���;R��C�	]~��JDώ�/�6��`��S~�C䉾�tU3��mx"%�N�F��C䉧c	�� �H-b���#�Cͫ(I�C�	>U����F�����lʻ~��C�I�s�HJqA�w�ܼ!r�\-�8B�I�dO�)Pfӎ39�C�l�5#�B��0=%�Щ2ᔲ�D����	�"O ��8B���*��[�R����"O���f�t�ʽ�$΀;>�(�u"ORYhq�����2�
��"��X��"O��h%n_�V�,�◯�0u�^�h�"O*	[���	����&O�	Z\)�"O��ےkI4l��x3�Mʄ&ٲ��2"O�}#r��W�𘁡
��E�8耳"O���V�H�K�<�X�3�Rp"O���B�#"����F-�t�iE"O�0S��*5�
H� �Ӷ	oh@ѡ"O&]�mC�I���k��߰tO؜��"O��9�L�I��m`Q��&?���"O���f! 4+�f�H��ڸ���ó"O.�A"�T.�m�Ffr�l�+Q"Ov���.+08��D�#I��С"O�92nH��I 6���M���1"O� lD9�n-Rc*�3z|�D"O��9��>&~��)I�[Nt�B"ODd�e�W�f]D�����3OX�I�"O�@T� {�Y��k2_*J��'"O��au��b��� ��l�r�"O�]����'����K�6��x��"OJuP��1r�b��Cb!g>���"OzP�Ư� }3(:6k�u6Qh`"O����Ke����Ծ6l��"O�Xc1�ɟv��h�G�7���'"O8p�A*�`�x�'K�7�6y(R"O�U���$R�~���ɑpt�#�"O	�GE�~nPp�Ҩ]e����"O}���[��6�(wh�8cxdk�"OhA�գ9NUf!�#�V���|��"O<��C7l%3�'�|�0)�G"Ox���Dޥ5/�s�)��X��"Ot`SE+�Eg���i,?��zP"O��3��/f
|R�AE�|�t5Sg"O�| a�ΑJ�p`���"�(�14"OB�K�Oݳ7.ؓC��Z�B�)�"O4�C0(h�N(���#f�D��`"O�l(�"��6pi���oʈ���"O2���K	\��4�A�F)@�^ ��"O&�Q�C�8c0�T�0���jt"O���6$(�|���2fIv\+7"O|���ѹ+jԔYp���$~�p�"O�]i�"��g�m�f�&*l��"O`��SE@D�{V&��o&iX&"Ol�G�P��8\��&�0��K�b$D��K��Y%��ӳ�WJ/JJe D����GM�q��0⥄��GQx��K?D��ڕEE�'�8ҕ�(�t�)6A=D�`y�GQ \�Hʀi���X�Q�g8D��8�Ȳ�|�홌~�&����5D��I���&>a�e!6��h$�?D���aI'.hx�s��$�*���!D�D���ސGG�Up���2���A��3D� ��L��[�6iWG�:^�r��?D��1�GF�O��i�g$�oĪT��#D���M��tf�m,�8�D�>D�4a��K�3��`;�ٶ�J����;D�����4<���r-��@�"K��9D�P`�/S:Pu�uC�AōP�
F�$D�paH�&�ft9a問D��Ѫ��#D���c�&P�Xڒ�ԜI�6�@/D����/+fM�58�%S�MJ��cO(D�4�A��b��Ѐ���S&)D�� ��1QyHhda�1Q�����&D�T����W��ǯŧ+���W$D��p��P�u~H�z�!����(APj<D�t1��^Y|h\iץPQ ����o8D��`�_�yĉ�aiۍP���%�1D�� -�~C��;�'�7� ��*D�(�g+�*���A����J�*D��e��.< �$��q/� ��&D�"�NF�/�LXc�j�=+�f0B��(D�l����\�8���� (�YO'D����y�5K��>%��(
�j7D�P3���ZF��hB�
J�(P�	6D�PA�*]3q��dH�^L�ೳ�4D��;���"�P)0�?H�D��8D�lpT��/!ī�ׅJ����6D�4	T��
��U@�&�:=�n`��l5D�� �` b�KF�=�f���x�U��"O��3�	���4�C��	b�BU
t"O�x�"7e�tN�o�B0"O��#���d".j�����f"OJ�3���7<Wf��oR��t"OV�j��)x@`X��A���L@�"O���OɌERF����D6Hْ1�4"O�|��Bٴvl�����/�pq�W"O��h�&�5g�zx�n�;*��M�Q"O�A�̑�|ZBip�l�>���V"O* �b̯3�vq�T��,Q��S"O6�����6+<�� R��l=pDۂ"O�e
��<�~����O�H.4��"O�42(H<,.�k��#Ct��#"Odr��[U��	U��N^��B�"O�ɣ���K��\B-�&�b���"O�)�&$��}��i �&Z%p����A"Op`S�!^�Q���Eh��� D8�"O��K��G�$LC�&ה}����w"O�QCɟ)�$�[eZ�~��P�"O\1xI�<� �j��B�vp"$"O��a�-���L��%M;|�C@"Ol���#�?�`R%N�E��Թ�"OH�їoQ�k_�)P�%�a���{B"ODY�u�E�
�&�*�΂:,ई��*OH�r0����|)�&ٹx��K.D� X3 ؐF�iK j�7Wۮ��a�'D��P5)ש
��Y���Y�q4$8�'D��tꛋt�̉��؝340���/D�h�aF�3D��00���N�<��D,D��0�F�Q������`�*e8��>D�̹�{�T�i3�۽>��(�Wk8D�`�`É�W�KV_�v����)D�T��iZ�L��Ȱ���� #G%D��� �	E��r�WS��'@#D��93`?r8*�;��T')Q�0�?D�(Y�O�4|'v,��됴-j����)8D���cچ&�ؑi$�Й@�~���i9D�xbJP� 8CV��	J��$	7D�ȃ�E�<��0K�
) a5D�j�a�N�x"0�̠B��(D�r�
�#�~�h�+�-cc��K� D�p�ٸe
B�[%`.|�`���+ D���@�P�
2RQ��j�i�(t"qJ(D�\:PjT.=�֡��eH����#D�(�Dą���!�t��):`/D�d�1ƒ=��T2�����(�ק,D�Tj��O�& �*C����X�(D��3j�&�Ɯa7h99�f%D� 0�e� s�&�Q+R�?~�AB1�#D�����U�2��QF�,I�tXɀ�6D�xr�I/ �rd��!¿"���E?D���	\�k����3N��R#��t�;D�����:V�6��g��	~�c6D������{��AҢ�
;%�����'D��9�B�63[h���N�@���5K#D���V�ȃ �>L�GDM?��YY¢?D�l!wjʮ"��l�n
�f0��b=D�X�%nO.�@� ��{C&\��!&D�����]�*d.�Se��4%+@��1D�,!QA�V�����3��)D�@{����
z!���N"	86<D���P�=Q8I(����6�°��h8D�\Q1�����2"LΝ	2�9D�� �,�$�2%� Z�ԒS��h�q"O��a+!2�fDI����'"O>�92��9n[>u Pa�0��|e"O�E�"ŗw�E��S�B��P�"O��B(��`��܈�#}�"�ʗ���p��sɛ�'J�_?���e�"CŚ��@���`��7�+[Tv)R���?�w�<$+F��*r�ڹ��
bo*@3\���l\$%�N59aΥ\&D���Q��HOֵ�e(q�|�S�V4:r������|� N��QBB(��at��ǗN�'�pT ���?9@��D�i� �
���!��}��.*Cm[���O��"~j�4c��p��a���t[A�����ˉ�d.��O��6m���oZ0j���3Ѡ��\f@����A�H֞���S��X��iQ��']B�O��`y��'�·i�H9$�̢U!� �5! ���x+ѫ�u��[G�XA�h��,"ɺ�H�O@�S�?Ѯ17�
��$˵����td^�ﶈl1p�؈�@'+�f�k"�+nr�s����ޙ���Q dTFr�D�4�1��iy�8����?I�i��s�$e��I�/5����Ũ��pȻd�ON��,�Of��rY�.H(Px�I�)Hҍ���O6�O��lZ��H���]���x�0�Vp�$8�'
@#L5���?A$,^�_��p@���?���?������hӄ�I��S�6�n�E�/D����F�3_��r̚�nԜP'��_���4��@�)�/y�q cAU����`�ĝ`�8yD�:x��C_-��'"�����ޅs�2h��ސQi��9��C�\��II�\��Of�&���	Ο��'�<�R*Y==���'\�uے�؍�$=�'&�.��A�{�Ɉ��8<�
�b�qӠXo�r�	g�X��+���O�0��5jH�$����3nb�H&$	ß��	���	`�� �I��$����Q���E�#�ݺ�e�iF��K�ˠu��U
�rX:�uB�&#���	�k4a�2]�A�\������Av�U����-f�d̹�o=��yPg]�(˰#�}�oʲ�?��4J�(P�@�V{�\c��ȪI�$���O���*�d7��R8N��]zcaIf�~�aǙ*�qO�tK�)�IYŪ �6I��,� ���y�]����M����?���M0D��i���'��;�4��� (O�̥:a�2A�X�n[�'p%@(�fD�v' f�q�B��8D�̧%ޠ��4O/��(�4É���Dz�K
?���4H�	H��S��֎5���Ӹ&Y��ھ_�8�3,V?J�#=Abl\ܟl�I��M�����T~1��@��a��ǟ9#�6�)Vj�O�"~�	��̢CnQ�>�(W�W2$8`�'�7�\���lڊDt�(��L�[Qn�rdE�*B�����jZ�ʒjW���	r��K�]�R�'�Fń5�U�ө�I D`��Tn�X@�iz�R5Kʑ4y�)Cė���|��'�5֧�J��5a"FS�G�n���h-�M�Co9*����א)��u8�B5��>�X�cm@)Ë�k��i��-�&uF�7-�� >��'����"|n0��%`Pl�Yl�	[�Iق��P��jX�D��*�>8o���*R/��Ps�:ʓNT�V�'r�x7��[;�$���C�D[�D���љ>�J=$���퉟t�jp   �   \   Ĵ���	��Z[vI
)ʜ�cd�<��i*<ac�ʄ��i�)m�@x�a�P�mڙX"��xP�MPy�p$eb����4\ ���b��p��IhPY㒩D[���1�N��z\���SV��+<�ɋS���{��i��,1Q�\�n���۰�Թ�0��O���A����M�]��P�#6B��A\�0q���%y1��̅g̐��]Jʰ�P�T��;��|9�B"ΓN:I�A��؉ɀ�Y`����nM"v���O�@��f"z��'j�Ea�DN��~BF�:��\S$�5���#�΄ �~�"ș�y����Q�<�Bf�,|F��P!$�<�L�BPD��<9`6�&r#<���N8b!Yf��oP�AbJP=5 ���W቗>
�	.� �1!	�6�x٢�� �'�nEx2GR�=� :���Z�prHͬMj�oڿA������I�5 ��P��`�x9��KrCr��0K:�	�\D�l�e���Kצ�>jslY� 	�?(��bl�<Ib)<�FI��) HΟzEV�y��*;��L@6*Ԯ�x٥�	/Db�d eh6��#TJ�A�	�Ř'�Fxr�V�ɲ~6M)L�r��r3勺o�
��`m����x�M��\y��R�=�-� N�y%�����O*Q�ṟ��pN�$}�b>JTe�'e�0�`]��*|h\��@�P8g�4`{��Iq		��wEp�S8�:m
�зϑ�4�n�������s5#ݏq��'�04%�݉��'�H9�6�����'ڼ)���S?�!�dދ	 �  ���"O���t)!I<(	�@P�N�N�Xa"OH1B�ks�r���-$THpH��"O�X("͇�%��$�Ɓ]tބ� "O���$B�D��O#�>���"O�B�O�;���9ǌ�<]�Lk�"O�<(Ѩ��\Sl��6�L�7y���`"ONH!E�]����Y�끹���!"O���M�
-��
Y�md����"Ocf	%X$�ʦJ�6l<P��"Or�;%�ݔR�y��n�	�`"O�GEC�.��V(H4SV$<I�"Oԍ��(��ialT
QS�q�t"O�5`C��0�< k̙P���C"O|QX����z|����O��9w"O�Ԣp�L�G���KƤ!K�4�"OZM �'�{1`��6#�l�j"O�m)DO�к ɍ�dc�Q:c"O�YҒ�E$kl�2�#hP@p�&"O�)���Nؖԁ7�_:@�]� "O$Xz�
�]�.�c�OU&;P(�"c"O/<H4͂��->@X�@�K��!�D�pP<ű@���	(�aq���!��Q�j�����>=8�8�/�(SS!�䙜5��۶��Y�Ƞ\�Y�!���%�[�,�,�9����B|�'9�� �L����Żlݰ�'8��KҬE���%ϏV� �
�'��$��C�N69*w@Ҡ!4"7"O U�2�Gp�BIPu�5/6�� "O�|;wmF�>T^���*D6'+8� "OPis	�.!���$'
IC�Q&"O6y��Gΐn\�����F�T%��y"O�p�aHM!h��ǣY�7�9�E"O-y0	�+��Iql�p�s"O0��c��s�~%�eN̈{+zMzt"OD`�u���j�����{�6"OQ��)|� 8dB]}�]k�"Ozr���8��
�JD�p_�M�a"O�\�CN(W����ٌqX<��"O��֍٫{#���C�	|(��W"Od��`�\(<�e��	�z��q"O�u!�h'����ED�$
�R&"Ot�X�!L �hXAc9 �|� "O� ��4)U2Wp��b �S�,E���$"O|�6c�'lN:�� �  *�,��"O�|I�e�-�T\u"V#��`G"O@m�U)�lR,��f�n�M[�"O��z�τ&�1�)>^4 H""OB���Jvd�����'_fӇ"O6���K��e+j@�9u?
�at"Ođ�U΂X�~��E�U0>q�6"O:��G��8W:�{��B6���"O������B��d��7F��Kc"O�ի�fȀ)�d+�$V]�� v"O�*�*��B��j�	�_��mH$"O�p��.N /�.I`'�.q�){w"O�$��ЩX�nͩ4��39�ֹ b"O(rԯP�dte�T���D�j�"O��ʲ�R�[b ����&�J��W"O�M6_^�
2#S�|�n�jS"O�
d׎uv^Lc�Dĝ.�0�B�"O���#k���f` �K2����@"O6�05hF;'R����#8��uC"O���eFG�Em�9��R/.�Д�$"O��*햨+��:F+�:X��c"O��C�b�;�Z9j�����,�T"OJ����-nЀU0�A�WItyb"O&tĆ0z�������f"O`�BV*�3�f��G�*tF�*�"O��; �.;��#�FƼVQ���"OAIA5Ba��Rǚ#$>>Ez�"O�m0�C?Zt@�O�]�h�*"O�)Gg-f^J��s,�!\@��"O������
�RԒ�)Z-e�$�!"O�a`�)�(�������(k�5K�"O�5P��~�y�7���|��e�b"O�Tcb���"Z���隍n�t�R�"O�����E>^v�(��E#,��,��"O�u�6�ҏenqX�$;J���{�"O�	����s!v�KP�3�(=�"O�X�4�ع nҹ��/vu�I�s"O���
Zg2a�1!�DD��"O���Db�Fel�{��06}�g"OH�bē��\B���$�&iB"O�D#�)+`-�!�=;�x�b"O8��E-ܐ�4<�� ��V����"O�����){��m��n� xa�9�C"Ov]i��;{�uZ�h��1j�"O�ɀC(!c6��#N�%U�.�z�"O�0r�M�)>FBH+T�N�a�$\y�"ODD�S�NSP�L�I�e�l�Y��x"�i��b?ik�V�`�$Z�!HN�.G!�$ѣEq�S"����Nl5�Oj��$B�i�t��1�M8�2�[��%?!�$	xj&��@�(-��-��+4!���2��Pa ��y�qSO��r!!�DBzwz�۾�:�y��!���W�HRU�N܎xۇMS��!��	���s��f�
�I�D64�!��;A���p�"[>n�3'����Wx�P�B���X�
����¶d>�O��m�ƅ�Յ��$��D��x9����G��h�i�'*�n��#�O�&6(��Lږi`gO�(ex��;@څn$BՆ�=rҙ��jX/d��b��q����ȓ�\1��2M�
�	�E��M�*=�ȓW�V Abfٵ9%�U��`��;-��S�? tHE�P�YJx�R@i��O(V�w"O��+![�-�:}9s至CB�(�"O�	3����"��8�X�V��Y�T"O�@Tj��"��-��^4L=�mk�"O������2�Zh)��̀x3Hl@�"O� p��8WMdDmտu���G"OdY9'�|H8�k	� ��a"O&5�҃�������q� ��E"O2��s.�
Θ��`�P�7�B\�IJ�Q��'6�X�dB�.�@�ċȄd8<�ȓo?數�C�lnle�e��VX.$�ȓo�Cw���"��Q��>T5��&O^�	�=�N��Ꞑ|��9�ȓ3i�����>#b@��g�]��%���B≬q#P٘����~xi�&wbC�ɶزe�uHװv�PA��,2���0 5�����@�=YU��g�T��a�'h���l��h����T����x9�'����7��h��RW%~���T\���'�>E��'xʠ��K@1����F�X�^���'J�~��yB���$���݄q��ls'�.�HO��S�� sqd�-��$s��xqȜ�r��B��*l@U�v`O<,hQ�'��2(g���	1��'Q�?��BK:.�X  ��=tq�+LO��h� �(Q�TZ�bU�$��s�C)�d{Ӳ#<Y�y�J��,�j��c�-��$� .�yB%B�8��L�F�R��w��
�y�	� ��j1)u�����0<9����Gq�e� �?U�hԳ���
S'!��ܐ9�\ñ�F�!��#�BL	!��jG�ɠ�� 
�|���8�!�[�RZ�	 ��2\M���ׁt�d�L	D�'��Ց��B�dJ���7�̋���<��'#1��@��d�n���+e+��@`�"O�p�0��D�^���IɲuV�����in�I�<IٴHO�?7�G�a���4�J3&����p#�L!�D��cW���D��Pّ�b׹y�Q�����<;��m��!O�Fpr5#��B�	1x���``$�=+:��6dߢa����2�S�O��0�σ|����Fa�<ݎ��6"O:�k�G�r�����ʌ�40n��Q"O��v�T�cL��D�u�|����O��	R�$3�L<ͧV,�5#�59M:��$!�&���	Y?�T��(8+���cE^7cl�}!*O�$�<�hOq��D�7�F�=�T��6��i|����'^�~�$}��J�
d�P	�%B�MbY�<�
ߓx�ԭ#��n��@��.�Lm�D}��S�y�"4;(� A�:(:4�H�,4�B�	�a 0��W�v'J��F�"�xB��;T_*��@�=]����� ҂C�IY�i�u$\<7��R�!�RvC�I���Il�>�qR�d��_:�B�	,d�@`SQ2"q���C�_�{�b�LE{��tI�k\x g�B*�pt:'"֟�y�L�<B8Ę�GC(��$�&'���'�A��	�4{�;3�
fOn�h�i%)��,�S�O��&�P��d"�/ʁ��0r��ĺ�yB�D�HG�I@�JD�Q�����~"�=�Od#=���F�2PB�@� ~��YG�U8���I�8��'j�X�Y�N߉;!���2g(�D6�S�y�81@-�-ct:D����0*��yFy��j>��!خ-����/��C�Za!�#<D�|����,����g���%�pQ	#�8D����Y��:��f-T'�$�d9D�� T)��̒kL�`�	?<�L`4"O�JCa�=' ���e�S!H��X�"O��Q��� f�p�T�
�It��x�'�`��NK�T�Y�)Մ�A���?a�'��y�����*N��P(���	�'��){�VNتa �ϩ;�.5���d&��?%nڮ"���a7�T1*i"��p���U��B�/c,Z�Hr�
�$�X�b����"?�Ӫ/ڧ#> Җ�Z�}V��3 ��/"�Єȓ%M�U�p���(&���D�s��<	��퓋}��i���G�O����
T8B�	�f��D�BC��$B���F ��O��C�d�\i�F��$y��Mr�S������"?��O>�q�� z-ԅ�#��w��ĉ%"O2�;�KG�������V��}3��h�H�>�I>YE��oHp#s-��>�~�(��V8��Dz� L"FW�0��F��T�x��J0�y��'p� 0��X�P�K���O�=�O�� ����,8(eِAԴA�'��d����a&ԚŤ��2�}��'�����͔�y��ec`��� u��'�R�ib/C�|�����}'�=���.O~�X�9C�D�AP�-[�H�"OXH��/	q��b�,G�{��ʤ�i��$�"�X�dgN=S����ʟ�5.!�$�1V�]�&R7x?�EѧFԊ!�3���8��C�r8��ʶ��8�!��2R6���*�L!j���cU<�!�ȥotz�!��;	�T�68!�
��}�U� ��� 	sB�-+-!�+#ZD�II�g.�p@��v{B�ɕ]4"�� +�"K��T
D�[�����9}BE:
k�pc�݋���!gT�<�!�$�1:�ʢ.N�@4��P��gɡ�dٟ<��q'���]J=R"���y$��b��H�E�m��$��5�y]y>��
g�XL�fș�D�:�y".Ȇc#� �W�Tv.�u�#�yb#�*s�)Ѡ�NG�`r�	ƃ�yBǃ(k�9S`�ěB��h�g��y�@,D�!Γ
7A��ZD� �ybd�(!���!eO�~o\�B�f� �y������k���.~)�؋�.Ł�yBD"x Fa�1�M>�HU0cL��ybmSbA��hSl9����ǒ�y2���J`DU6/��"(��yR��#v���./����1#��y��	?��9vAޣ;Qx����	�y�"��������-,a���y�\�-�j���MU�*�4xw#�<�y2hT�CD
܃�MYX��+����ye͕Nz���Æ�|bl���E�y�I�N�l9��	�j�����y�1 ����A'[$�Y©���y�훈Ҭ��c�<�|5���-�y�kP�ʨ�ؔF�(eYа&I���y2�lQj��aHҗavl�Q�MM��y��W4&x�лGF�9Hn%�$Dɇ�y҇��مA:&�8,��e�XvA��'oJ�$�49��׫ )���K�'�V�9u��;?ˌ�@��Q�8��x�'�Xc�ʺJDa�����xJ�'��E9W� 9����٠OgZ�(�'��XۅJP$pl1�G�$H�@��� �ӦΗ�A��c��-{�r�"O��GY�7 �D�F@ɣ$"O�a92eد;�<��j��8(z��"O�a�3�C X�:���
-��Qrs�'�D�y��@E�6�A�Z\d�{��zA��O�3r��(�'��X�6@4s���أ�ռ!�pH8�'d�8�� �<)���%�1����'&,t1�[�I@HÔ�Ŭo$L��'�ƵB1�R�i-��sG�\�,1
�'�����ΨP�0E�B��+Pݐ�j�'K�H�d�8���{��P��hb
�'�x���RT ȑ�,KC���	�'v����G"d~��:�qK�&L��'&��� # ��p3@�^1]�6�z�'�b����%��}w@�bv��
�'�����[�d�h��3_��e�	�'�&�� �	�/,���siX�S��
�'�2�"P�J�M�i;3̀$�n�8
�'�&Ԙv�E,.+�L��`X�I
�'��I�$$�6f"�C�D��:�	�	�'T���#���M!Q#F0@���	�'I�m�u�ٯ)�I� ��+:�r)9	�',����U�>H��B`��;`)�'�����X�zR�Mq!ǀ;$�ف�'�$D	��Vyil� 2nT���'��p��H�N��AZSh	2;�vآ�'3��e	�LY��zS��jځ��'T�d؁@ң? |=Q�V�y��Xz�'�&%1$#�C�P�����qƱ(
�'����3_upt����F	n%F(��'���X"�D�:j���#)C�ȹ�'JVT�L�X�Vd(�`�)��\��'�j��$@>+D�98U���F���'��Ɂ�8^�x�*7�z!ΐ+�'��	P1(��\�#�	� �de�'����#c��~, �g�6��t��'f�}�tJE=b��B�3��9�'����'�Z���c!D �._�D�'uLH�V�f�\t8 e�.$�P�@�'�nH;W@	1�X�c3�F����p�'�R5+��V�'�H��q�ǆz�lb
�'��;�� ,n4�C����y��@�
�'Y��8���(���)�J˼|�y�
�'Ɏɚ�M�b��Y�g*��E"
�',��HA�mKr�*W�4|-�pY
�'V����_7�䉰�l��kV� H�'��@I�F�e�KFA�k�̤��'�$a�5.Tmv��e��/bA~���'?��íؒw:q��R4"4�h
�'z�D�')h��GP��!*�'	D�y�k�*qC�+�/WzސK�'	�a���˒� ��p�.m`�I�'M�8�H�q:F�{W�Ҥe�܁�'�TȠ�*R^0��ݗe���[�'В8s%"�7������?x��Z�'7r�j,\(�R����Ă2(t�'�6P�� �z�l�`��ŀ 4� �'��PסU�����EI	���c�'�<���Y�g,j`�@$�Jp u�'�[0�b�0	�MS�Fk����'����t���/�l�����A+�0A�'"��QgG����xԀAo�	�'�8� ���g�ܹc����6$ܻ�'�$`# .ɕZ��#!�JRr��
��� �����VT�a{��ؒ �ʤ@0U�T����cJa{b+ĳ[�>�� ��lPY���͊�p>IE��6(���̖.�	y����k�b9X��GM�`B䉂EU	�)��Z�V�#��<�B�\��B���"�ӌ#���zg����O50��'䖌s*P� �\��Y0	�'_��*bC�z��`��q[�3��	+p%<P����wY� 1�E�� [����G0﮽+�D�EU.��#j]�e�0D�"Od��ꌔ'�8Ab�	��!~��n�K��LA�MӥE��2��+L��.R�1V�tGxRB��7�Jxy�AL�F��xV'��p=s��>.���7�U�8�k�H!K�4���-�Tm��@бe�@9��A��(��䕺i��xb
�#Lb(#C	�ArqO���ԉC!=��eK�'P]I��L�:��O:0�N�R�ք�wk�"�'t*,"M�?^^�G�=Z�$G v��ԻE%�Y|��Å  �D~$82��t����y�)W�3rv�v�Q;W��,i5����y���\c�JL HB� �0�� 2��6��<���4�a�#�x3Q�M#NI�$�O��R6ON~�0�hg�K\�I�G�'�f��CQ�+�>����} ����S@ʁ�sN!�nYu��.I8h�d�<�L�Qn��0<ٴ��d�5XebD�1��m�L�1��y��L܎K���
��XV#J(#3��N������N�#>ic��a�f��Ђ�=I��Y�QB���?�E�z4`Ѓ�J4f��3�],z�ǀB;��d[�a�?;%�q�e�y	 H�
J5��B^Ƽ�+��z�d���΅66���t��B�<��Ë�6��p*�}Y֝�RI�X8�H;���f���/K9uR �0K�heT}���U��{U�и�̗*�V��(�GƼ9�D�>LO� kd-� e҈pz�χ?`��%2�-�.�6�;��V�f��3��R߰�I�6���Fh^�$�џ�h��> g��H�Jȯ95&u��!#�I�.�PAű@j�)i��ǫT@�S'�b�gM�\�~��	@BX�D�ܧHq�8��'���ë�D�d�s�O
+o��j'
�9��P���?q���Ҧ�)�u�B��>���UO�)B���� �pZ� w��#�yItg_<� dҝ�d@�]"w�B�ɖ��)T�H����d�׼i��QI5�T���D� s�L��V.�*��d lt���dXI[f���*#+nџԩ&N�b*(y�U�Ϊg���I�� 6^x�2H�"u��<����.y��PCWy⤆�0b��92�'b&����n~�[��]�43�3(O�=�.P4su���l��K#�ݓ��ڀ��1�J�Rɇ�"��t2�O�,B�`���6*�~B��
s�Crf]3";�ӓ��U�ֵ'�Ѱ&b�Cr�2=��@9Ջ=�i�>���BR�ڄL��`&"��M�bq�����@	F��u��o�̋qM��¢�ٖ+�[~4�fJ@�ў���K�h�x���	H��,q��c�n�����8�"�?I��D� J�A���٨\h촲��ө#���;u�H�E��z6$V&!�t�z1�ν�x�g�8����
An��[�E���$>+p�����WV̡w�D(on�ѳ�0��3?j:�y���'h]N��#Gu�B�	�6ކ�p�E�B�py3�^�S<�
#�وD�R�t� �7W�I�Q%3�i�5U��b.-8��� M�pQI�k#2����`&9�@��+6|�Y��큨9t�*���"c��n��B���`�j��$*o��d�G��,�����_�"�x�-�1y���#FSx�F�p�	���� 4z
�Q/�D�1(�C�I�!�%��ዺc�m5nպ%��b��K�ɽ-�f�P7 ˄,�c?�kB�%~�4E�P�N�y}D�B�F+D�@3ի�k�@�f��풝��Tu+ÏAm��i4��1�~2�K�ʃ�|��a�ᘍ*�(D���f
S�)������7N��r�A�O4��2�(4�A�(�-�<r�քp�UHb�Y- jxÌO���Q`F�3�<�p��C�z�ôč�l6l�YP�E\2H��OJ��&*�'"JX@rSƉ�=����I0?�b#հJL�������*��4aw�I�"�l�;����y�-��F�ZrR�+G+�r/��R�޿jӢ��<E���X��0	�	�	�>����=
/r0�ȓ�^�(���-	;ą8��&|MJI�'r�#!�W>M��y����%9"�{�'C/~�&` �5�p?	e�R�vt��+TGȴ,L4��6"ܪ5�>���-D� 
�b2"�`����Gy��+D���� "���LŨXƬ J�)D�\W%^
� Yh�B��0/'D�4�5.�q��9S�Ɣ�ij2Pa� .D�0�'땼;�4C�'����=Ҋ(D�� ��i䋐1f�<��*QMD�9�"O���U�ͧO�T���(�zB䰡�"O80�S ��~;P)���OU9�(� "OT��Ƭ�I�\+%��#P���"Oڵ�����-�fA�'���$�P�$��xpm�Óo�HU���	��L�&��'{����m�@�+U4DP�X�dP�>l7���|����'Sp������A�e[�0qNpi��dǫIn�eR4����'EҲ�H��. 	J�x�H\ݬ��ȓ0
]8���.7QV��ƕ 7Dj�'��\#]S��OQ>-��O�RAlT��#rJ�QPL-D������8\h����%����Te�9��II !{��m�3�/m�`�z�Iٻ���J����d��n�x�y�.�]���aa"|®ك��Q����$��B,)��S��B	J)2D��5��  ��Qj����0�!(1֭�RB�BV�B�	�!h�}�e Q����JW5h��8Hy��+B*^Y�ҧ(�,�R%�z7r� H0Aǒ�@P"O���6n ��W)�`�`����~��Ҕ3�D�8�/%��䈤�Te�1E�=RN8r��&0�!�����]x���0���� ��!����W���E8�����hX\��[2x�d��!N�%��xbM�o���<yF�Z� x�P��[�u�:P{�jPt�<13Ğ�5�&��1��]c�D�p�<�#L�&66����ɡ��@v��m�<釯׫}V��T'^�U�������m�}���xC�6O�Q �z���咍O��a�O�qSA���ussc�?�)�D�9T�^eʀ?�O"$q���]�hI��g^r���I2+x5�U�:�O7�]Z�O�3����a藲Q�dY�'��H`2 b�0a蘿Ue���,O����f�Z��O��|AhA�;b<��	�O�<��@\�<-�^l�lD���1�c��@�z`���>�3NG0����J~�=yG.�R�j���靝7��-��M���P7n�"��<�g-��x{����a�1V�8�Xr��}�ab�S�(ݢ�[y޴a�&�Х��O\���i{�m�N|꧆�B����`ƺ_�r9gk�N�<�����\2��I��\JyRI���2� ��X����5�މ�T��FL�9wb��p"OZ�2��0���'J�t��C�Z�d�'�8�#'2��D��L�vU����a��ۗ�7A�!�d�N��C�Ζ�i�V�;P��0�Q=�n���8�x��V�϶kL$��P�G�e=�xN�	?٪5�<�O�!8��aB4������b�<1�A��9�����όDL��@���_�<Y�V�R�ƈ��]	8�� ���[�<�aM��h�+��Af@ (f!NH�<����"��]�b�Q��8�AF�<��*����貂G��0����|�<YaLT\��D�d��O
v�#/�r�<�e���L�!і{����b�XK�<�2'ԁO�.�!tJS�@���F��H�<!%��$w���Pp*��[��Lْ�DR�<yd��Q*p��c\�s���J�<)��5!�]!c��P�1���J�<i6�4y^8�bE^�
/�}h%��D�<irA˼�;gJ@��I���B�<���֛�1���g�
��q�<Q��$�PAJ�L�:��e]r�<�d��;z �S�AݙlHQRja�<i4�݂_�����@��s���C�]�<��k�(h#<����ÈpM��ehWT�<��ƐF��]'�J�!��ɠE�^[�<!�f
ވlbtƓ��U��
�R�<� ڝ�&/�r��J�EJ?&}10"O@�^-ٴݘ c�u�~ap"On�T��
yvdM�p�0�l�Q"O��x¨D�?.��S�Ȉ"? d*�"O�<�$�SS.:�k�`�/S,6���"O���u�D�Xe�2�\�B����"O^ej6���`9r)�Q������i�"O�e�ł�^~`��P��`yj0"O- ��<xSX�oH�j�UAI7D��ɳ�S�z�^,�Q�_�e�^�`��!D��[alI�MRt��g	l�vi��=D��91K�?m㪈�5ņ�if^��`�?D���#��=��\$%�,�p�c?D�HH�]9 Z√�![�o�x�Jq6D� �_�e���u+�"�`�Hf�:D� �D�N� ff4Z0��>e��(׆;D��ct�=%Y2E��1f�%D�X��	��(��yb�j�v�6+S�6D�t�'�&*h�(BN�bV�� RE4D��!�`X�`؈F�--h����?D��:#�ũО��qC�+�0�H2F8T�<+�@��:��BX�}QP�I�"O�X'�	;Ah���6��/�|���"O(X�4�آ>R`����&_�ܒ�"OSZMߞ5��Q�0�N�в"OR���"g��3�*��
��	��"O���@Y���Q(��.����U"OY�u��X�AYUf��]���"O�����(�T���R&C��A�"O �E�6$��@&c].O��j"OZp@ [�3�0��0�˽&l�:'"O����D�b)f�h���)5H�c4"O����F�,��+��#"�af"O���3,]~��Ǐ�6-ɒ"Oy5I.(��C0F�W뾹��"O��d��`I�1�vb���T"O
�2M�<{�v ���AQԍ�e"O�k*�*P��X"����#g,�q"O�z�c^�������#A�Q%"O�|�GW.n�f(�&�M�P�My""OB�{�E=
��
Q���"[�	s�"On�!�L7(,��A�s�iY�"OD�pQ���+=�qȰ��X��"O�I2.�>+�<��膴'.�pp�"O��
���tr�t
6�ۗ2��Zb"O� �J�8�>�b�!��p*�"O��i�AD&9uV�!��T���)�"O\8J��+�xxX%BI��ĭ�r"OZ)�T�; 0�@	h&�:�"OH��j�0}���W�k.��b�"O�H���́�;�O�s�"O���ֶLL��;���#ft�Q"O�W_�j��E����!�L�u�<����3���0��,�l��5-�l�<!4 Q�_�f�B��.Y�h$b��Hn�<Y����y2@S�/Ҡ���oIq�<	f,���}"�KJ��9�$�y��O��D���v�XqC��C�y2)�l�Љ9&�20�fā���y�Dԗ$IF��'��.��4��y���-/���I
�R�te�2L��y��*�t3�X�Y?��0����y��D���qJD@\�]�J٫%R(�y2���v����`+K�:ݸ�A%@��y
� 8<�sO� gֱS��=N���"O�ey���;��t+�
�j��e�"O�a#��Y�+�H���fV+Cc�x�"O؈bE�;���iR�A�)�h�`"OV�V��$w��X$�3G�lݹ�"O&��Uo�<�`���ƽ �F]P"O�us�mG�5&ؑ�F�W�h�jpH�"OZ@2���6��aDCQ�"�0�'E�@t�H'��		�P�˥盿>�\ 3 �Z�j��B�Ɂg�z��b	�;,��lث#�rb��̘*!�xhF�Ӥ;����`�m�D-�[\B�I�v&�����Z�ڸ�0�L�{�48Q��9Ol�˓2��	��L����\�h�M��抍4��P�?4�����:&��U@��`\L��`�5{�^�3ª�pV���	`�)�$K�Q�v��4܎b����dR�n���]a����z��Ǎ	S��)r��9����'�>Q���*=~�4��g+'�t�N>����)!�H��C���T�˵�k�L���*OB��"OƉ(��]V�0�så,\����ꝋt���H%+C9�4T��E�-
���&:��%JtV���J�7!���I�8ͬlh�OZqC@A�"��&XlH�)K$O̲.F�9��
�	K����3F��<�r�'C�XS��8�Q�Ac�h�S�}�D�9(Ǟ�g0O��&%�rM����~ �pIa�,�0��u��:nd����iӖcɆ��;;�Xa� [�G4��qq	V�BF������hdcX�j!zPd�::�@!0@ڃC2���'@L�]�{���0���sC�-)d)� WwPB�ɝ`2t���5n̄j�P�Gl�	F�8*(p�1cM*A� �k���a6x�����6jȔB��Pxy��
r�ꬡbO��,��DY�̺�p=���K;9]N��N
�-��;��� -0\H�!I
eTB��b�=q=H�L\ ��ߚ����6_pe�A�6fŀ�)���'�h܋T��D���� k
�D4���-jfM�2 :�5�#�ihd���
S���s������U��FpC��>Ϧ=Rga߫�F��ጄ5�v�#�lZ#t�ם�U�fKa��Y�F4��OkB�u�m����'�"�j6&�pv!�$w�B�)�kG$9R���YQ
��d���P�y)��#T����(IT�	!��RE�.�剰��X��J�<&��@�	�0e���?A��(������SŞ�났��Bh�ayՃ�~>V��V�"%�"�X�����
J���r$(O�Phc� � er2����J�R�0����  [BRX���� )K�a��$6�b�&|�d���B�"DAK13�H A�7��q��^6I��I��.P�&��A�F����}��
�9j�@YBeړ�R� 9?��F@Ag�Ҷ���C�`���u��PðA�:P�m��I�VɕI�,h�a� a�"Pp�Q%lɎlɤlv���ŝ��隕-Η=���
sI4�vOr$g��4;U�`�ˌ�R�>P��6,b4�[f�@d�6A�q�(XW�u�
�'�����6P�%� Gf\8@,OpPI���`��Ш��$9�Dlc>I��@Gen��qf�V�{08��1D�Dq�Yq*�e�T�)�,!$)���)�"Q!Z!FŘ�) �A�\��Hݰ�	 ?9#� 0i9�BիqZ���C<1��!:��1�ln�Ќ���S�D�(�SK�2,����L	z�4�h�� OԱ�t)��mH��)�Q)�tˑ�'o�)iW�H.G�X\m��v�6I*�*4��a �H�=�~@q��ĭc�!�\.FZ��FR ,\�-��E\0&��O�}9g�H�w�091��K���n$�����V� F�ԃb2R-�"O��;A�-y��u�5�Y�!���Ύ�v����l]$Xt����h���S	�Qw+��@h�i2�ܣc�!��-�44�Ǉ�w_�l���+���zv<� 7ϕ.�t�剾>�� �,�&c�fpkCX	����D�7d7��!*��8��h����.Cl���DŲ7�Z(q��7ːx2(����)���z(�|�!��<�O���w��;&;89�3L[M�KTY�4xes�cF�1{T���U��sC%��0��(�Q�	-�4	QE��86Q>T0��ͳ��)�矘�c�ܖnԴ�
e�C�T�j}y�+8D��3����)�txrp��#&D�a�"?��`ƦTBD�
ϓd��tZsj
4O�f�����	*���	����K�	�<�D;R&雃g�;�!�Ē	��Å�@�dJ�98����	?!�� >�)�숪z��$��KJ�(6"O(�[QH�4EecQ�)f�� Q"O\̃f��&ʹXg�,C��h�"Or���ㄿKf��3�G�sB>��&"O���$O/�Q�AcV6i5t�ѧ"O�)j1�ѨQ%!Z#!�IL�)Y�"O� �&�w*��!f܏z,f�: "O�T�Qޡ{@��Q&תI�� �#"O�M��lޓ!�DX��T
C,$���� hy	�S�X�U �&O�ր�Uo�u괉���S�P�²a�< �-�0���Cj0�beEF�.~�����3�#�:�*dXԫG�K[�GR��_�؛�!o�S�q�4`0M�*��)�G!��J�fC�I�l��} Ԁ�����c��%Ѻ�~n4�gϏ��`ҧ(���q�`V�:�`HГ.ǸRɑ4"O:h+`G�c#(�&��!㞼�v��@���&��РH=БѳN�b��i���8)D�b��M1�Ġ�'��l�,,�$I_���
V#I_~�Ї�	32��=IEj՛I��d�#T.%Ot�?1�ĕ�Sc>�z�$�I�4X�J�yr�R(d1�uxCL;!�H�����#%\p���E�F�Rn�� a�Z�/�S�O
��c֮��`��"J�'4��'��2t��OD���'D2�v9�.}r��g��"���{2�$
���rs�ƫ��� gY0�x"��L��B��}b�����Ýh��`[����+�������&��"�Z����X��p<����Ct�b�'mW�R�2��dJ��s��TZ�!>D��b�M!.O 5XEļ5�xpؠK?D�4{$��>�l�AA��7MU2|p��<D�p	aτ)Į���-��&e8�[��;�	�3�%���'�x��aآ�<�[wO0I�H� �'�h�1��WI"PX B�(_=>�ɡFM9A��`��'c8�z0�٦~���P�l�-,�x����A e��9��3��'w|��򤖺N����Vj��m����eNx5���u����e�&Ֆ'��QP��Ǯ^Q�u�OQ>E�R)O�Rۮ�b��E��h�f�1D���ԡP'8�0���@�=+8�7@+��	�yB@h�/A_�3�ɏ7\P�2��1'�6=���?���đ4VH��B^m$B͓%�R�w��K�w'���	���!�"GQ�����BaDb'��O�u���\�S�*���RjM2cV��dGL
�B�I����d��1n���H	&��ʓH>ʘ)��� N �ҧ(����e���s7�чM�$*�8�"O�H�B�Q9)%��*���)�{���d��%1T�)��'���U�7��F`�1L��lx&�*!��՞2vABaj߯U��S���QJ�Z�W%����$�Ͷ�s�F�7�8�h����1��xb�8�hx�<y��P.)=ʭ�ŉ��6kxy�Q!�p�<�(S�3�hu��,߸U�� Lr�<y'��/N0 K�A��.��aaw�<G+_+|�(�Ae��7CR�5��[�<��*/{X�U�G�?������P�<)g�`���������ܛ��x�<�Q��B�=����B��a�<�jJ��y�Ӥс\��=�ΜG�<�VkA��V�P��֡ ��ĂB�<�#mïƱ��c$�c�$	W�<�Ggαk{�����(r���H	h�<)&㉘/� `�IJ%�lA҂Ze�<�t"��vv���G��,B��@h�<���7N�8!���U�PD�k�<�D��ZB���(�Bb�����]z�<ɆGT<U�\�06)�>���W [p�<���F*|�!ag$�0)R5��x�<� ��B��Z؀ѫ�S� ��"O�R�Η?;*���G	�xg�AB"O�KG�F�'�4R���g6~v"O$�Sr�>K�ܘ��	��!s ɂ"O*Ls��;;��%�ǡ��;Qa� "O���@"��d;JAaРV�-e�y�r"O��b��<i� I��5+�H�<9rJ��ˀ1�+Y�T��Z�/JA�<IV,��.+�ZG�M8P �G�B}�<a���:���0��
�e�GM�q�<q��;0L��:��	�c��Z�+^d�<��. �izB&ޥiS&-Y� [Z�� Y�7.��+p��s�n��(�-���i"'�3S�D*)D�X{�*Z/"h%c�N��˰�mY�<�aξM]��	Ţ�J��I�w�*D�KC&�T]�	G�<��Q3'K(D��i���3�*]q��I�v���&D�pH4ˊ!a�l��/�?�8�pB!D����W�&t@L���]���7�>T�P��:�ZaSƋV4`�lB��I�HO��Ivx�G�_4cZ�hc�ȸ9��ɽz����J�3G��S�'���O��Q���D!�6h��^�0�	\�YL�I�@y��	�1v��DJ��7"ql���ƭJd�k�$D(�t�'�(��ᓶz^�}�!ٍ{�t2P�O�!��l��E��1��BH	�e�3�	V70u�q�f�i���G�@<bq�O��@����<���	ç������ͥ��Ѭ���F��'n,�����f���$�>%>�.~���.B@,2� �����v
�@�Q�S�O ���*�*�䪚����p��O���P�'��좐&� �0�+�M.EsP�8
�'Q�tqAA�6�b\o9E��x�%"O����M�,���"C>0�HxE"O�1�cPj�a�A��0ި��"O���4�Vwδɔ��Ŵ�u"O��K& ��� ���ۗ7��C"O0L"bx�z��R�(MjD��"O�!�df�.����ǜ#1�[�"O�x�)	�"pUZ2)N$\�2���"O�����Ox�UJ'h����"O�D3&D��(�A�C/9�0#�"Op ��KL�����O�*#���j!"O"����ό<�r���NҢ0��ٳ"O�}��)�+��+ .ߦ-�t�"O�\q&ݨ�2�a���p��˶"O怘������k܊D��@"OX�����wڬ�� ]��R&"O�P 2�^y�pq�*�?+t���A"O�YѶi5_�>$�뇕o����"OEr�o<��Znb ���"Oz���ѹ&܁R����:htIKT"OtŨi��,�Ƅ�d�G&h��"O���+݀`e�p���3y��"OX���-SCJ@��e٬1��4��"O����퐷J�z�b��<y��5��"Oz@Q gݝX�ej��K$iD^Dh�"Oj$X4n��o4�2���?H2D	ar"O��G�Q�1�"mɏs0(��"OT}���O�]�4Y$�ؑ`;(���"O<`q
A�%@����.!(�"O&��g�^�sR���&.Ѽ#�"O4�aS��"tò�j«^j�A�S"OZH
%+L�%z`5@�ꈉ�͸"OD���<z�(�	�##�:=��"O�=��I� G�~��v�˛�.���"O@A�a�� :�(!2F�R��7"O� ����*R,+�4h:���27�TE2�"O��)�*�_�Ɓ˰EʬH^r�`�'"��ӦP�#��X"�",�d[�'�֭�v�Z`�����\$!�-*�'�h�dc�4@�P :)����*
�'�>T����A>�X�ЬW,���H�'6���g����!BŌ�Z�!�'&޸S����yJ]�.�~��pA�'D��"Mɲl�\1
��Ջ!�Hq�'�N|� �06���䍸O A(	�'���BC�G�1���(�b�HN ���'�����^�������;"���'��,jW�\�N���).k�i��'�Rt�P�V��r��u�F�#����'n�4�pD@�D�H�U��6H�|��'v�Y�Ү��?��h��L�t�z�'f�Qt�E�*ŀ�W&�	)�'qRH���2\؈��+ #R�*�{�'��Y��I /u���s��K0!�'L��*Ձ�P��vk�F�`	�':�m��K1 a��b1O�/:ƼI(	�'���ZC�&P�H�U�θ=�\9��'������pL�Ӿ���'�Ĕ��Ƭ|�r����u�t@�'����8��!�p	6u�8��'Fv��nלz.j�����q�'��P)���+\�֐����H�	��'J�%�`�2% �=��Z/B�X�q�'!�Q d��FERdTȲGW$��'	�hP�b��-�&��S&�G��q�'*�d�4N��1�đ���2g�v���'q:����B�y�D��QGڂ�%K
�'�tZCE�t���Ɇ��))��C
�'�T�*���>r���ǘ5"hpi�	�'���CͲ)�Hh-��/�jqS	�'}��Z֪S**�<ӡ.�#:B��'��j��M�N@d ��o�'`}`k�'&&�`5��F�зïTGL�
�'�^���Լ&�l�ׄ�Q���
�'K(��fR%^�
�FD+z��A	�'�*�86�H4I�je"&F��b� ���'e.�(�fݐr�Ր.�,UD$ ��'[>P4+ϓJo�]a˘=Q�y��'���9����JFhӡ.,H4���'e�Q�c�����b�_�;n���'�+A �ِ-���5�m�'Œ�AP+��
]a�� ���'�<�2�f2M�*��G�E6ABZ
�'d��c$�8W��E�M�33���	�'6�����1:�R@�3�Y|�����'���; #x�^��BJ�@\�,2
�'�<���C�x�"�R�	ǁ?�ب	�'8�p�!h˒s�x9�� \�A(	�'�.b��'mr��WJA�o.�ٲ�'	L��gmX(bՋ6 ��T���'�@ �!��L�,����2E��1��'/B@���p��h+���@���'�DA�W-H�:����z�  X�'7�hqE�FJ�ȕ��$zf�i��']J���d�:cg:a�]��j4B��y2D�4d�d��Ү՜|d���y�L�9p�jw��x0�Ӄ�N��yR�C�V�A�e-V%���c�H�yr�2b�={Q搃#�H���y
� �q��))z5>#�X Y���V"O�%h�BF0k	ڥ(��!��-c�"O-�d ��B�{�b@^d1��"Of� �o�`�I%��*=Qz=�3"O�}B5�L0?jt���;@;̄�""O�1p� �l��W����U��"O�m�"��.Y�j��� �(�$�"O���p,B�~�%�V���dV���'��t��T:��y�#�S�vK��P�'�$�b0�W�*LKS�вqH���
�'IJ�"��h��xE��h��P�'::ɱĪ*��D�I�S��;�'j~�#j�jG�]�7`�R�B-��'����U�ɟ��(�;�n�a��r�<Y � 4����i�9gO�����j�<QR�ĵz��P��ѮS�həF%�]�<aVo��&��x��M�#��ɗI]Q�<���̽)�	3�`B`|��-EF�<�`fʦ{�,�w`�x�N��K�<�E�Ӄ|� �d��'蜣�b1D����eU(���b� y�=D�x BL�O�Tlb�(6ڢ,z��;D��[#�
]�`����>/�H���M;D�t��a���5�Qb��Kl
( �;D��" G��n�b4�ȃ�u�Ľ��$D�ĩSD�3K�\\أ傉;�Z@�k#D��"`ü{�����.�)[�N)5D�xjs���9���R��J�nOv� 0�&D�������K���:�cGa���8D��Y�D�
�� h$�� 
)��5D�L�Q$W>vS<����Z�2����Dm)D�hr�EњPJIiF�I9ΐi&�&D��
�W���e����9�p��$?D��T�M5�v�bB�oSH<D�ܱ��OK�h9�Q"����Q�U�:D���
�f�z@����`��PH`�*D��3��M}��="��E+;�޴�1m=D�$�t��,@�
z��c�,���6D��CqJX�3~�e�Í�"2A)�K:D�8�צ�w}Te �П)]Ν;ԁ7D��A��D��(�GS�H����g4D�� �L�,O*^1$E t�0�2�M(D��Q���A̬���ٶ7��!�$(D���`�\-i�9`�%z@(C�%D�p��A�lz0���fPjb7D�4i�(�?_0��&Q�,�Pm!D�X��C�n.�*��9�	���=D��A�G�J�����	�Y���JF�6D��Z�ώ�u#��t-�	+�+��.D��+����[����LƓP�b+-D��9qO�XAH	���8�p�8�K+D��z�E1u?��$�)�,X(�G<D�術ʶ$�ܑ�v�]�*H٪�?D�`�7��0ut�:��Z�w���9D��X��"�D컐�D9$��+"�,D�H�dC�U�uH���,�!�#6D�P��c��������1yw:�C�$4D�ЀeT,
�R\���U2`CR8�E�3D���`�,[���U��yxÕ�,D�X�6EJ�x����BN�S��aS7�0D���!�Rs"�P Ά31�=�TK#D�`WFO�{80{i�e��9��.D�\q�@�7�B��gJ���, �i(D�( � ^EgL�AR �1�|��!D�� �-�Ȅ6/�^���H�~.@�"OP�+U˞;y�l��1ᘈ�~���"O�M��&���!�&K�R�D�s"OZ�w��Rd:%! , �Z8�"OҌ�G�R�y��@�aal�-H"OVȠd
ȴn �|K�ɮs��M�6"O2d VC](Os���I�!��Q�V"O�Œ'��v��DHR1SzΌ��"O����?JHa�fݚ2]ht!�"O8�Y��(�2]�Ě�EGF s"O8u� �tabxZ7��9�@"O��C��5�! Ū�)����W"O�2�lR�8���"�̪��R"O.��B.��F6���s���ڥ"O����OB�V�j�KE�J�~d( "O���w�͜w���a�W�<�jQ"O(���-KE�P�ǉD�t�L��"O�L3�.�$���JǸ_l93"O~����B���ЀIO�4nc"O���H��7��m���m3��A"OHh�ª����XRf��X
���"O�s0��"}l$P1G%�
l�0*�"O�<�A�_��5��H4av
p@�"O�2�9 ����e:9p0re"O �����V��j4��>BA�$`"OΈr�+F";@���c,)G��"O�4KW�[�_��z&#�
�v�r`"O�q����v�<���hҡ���B"O�ht�+���jL-
��\c�"O:�:1�[�W�p9#�E@�����"O�@��)�LH	u%M�J�2�"O���Anji�����$�Y�����y2�';�&�y����`I
7��y�M�;t�(�5��m#��O��y��%T
�j3'���J2���yR�P^t�6��	F	���
�yr���J�H��AN����
Q���y2��8X�6A����~�V��SbE��y�ʅ�.��$"I&'�a�&� �y�!3>d�	r�[&le�4à�D&�y�j5_9���G�gǔ����� �y����. `  �    �  �  �    _!  �'  �(   Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�H�!xn���G*W�(:h�.|&�t�BfE�C�V����5��8b��M�5P>D���@$K���x���1Hm�� ֡mD8�3�̕�Il2�"�JMz�8-�t99��'d5���!"ӫylhQsϒ�UT��VJ7Q&��&݅tΨA#�7z]Ҝ˴�USX�\8��!s��L�;u^"�z��9D�D�ҡ��[�z�{U���Й���*D�|!�*eZ�h7��K򺭁�*D�H�� z�.�ك/%��qu�:D���߅Mu� zBb�,5�f����5D��ڵ���?�i�d�R?R~�覬8D���RF�  hyI&h��D����&8D�P�gmܩS�d��wቀ`v!0w&8D�ܐu�lR���W+6�p��Sj2D������~(I���;�`5�#1D�h�ŇOB�t����Q�y>!05f=D��+!b;��)��p�X�(6�;D�8kC�|���^�gHP��6�<D��ʳn��v�Ȕ�-�IP=� <D��
�����P$�9v��!���y�B�9�~���,�zi�I �nފ�y����w^iZ�n[w 9f@H��y��Z3;+$L�RmT�7���h� 8�y¨�IFܳ��V8��&�ɹ�y"d�>xRLɋ�ˑ�Wj�ƌ���yi�$�����N��\�b������yr$�twj��0*e��Ā*	�'lp����=A��������=����'[ZԒ����􅛱��&;h��'-�@��Ш�D��)F�H9����'�@}���0c8L�F�
�A���	�'u��@K:ɀ��AF K�x��'by �,S��>$q�FX:�&x+�'�:�"��Rx�S��R.,�~���'�l��e�S�=���+��ܒ�'~v��锆P`�+��[ze��'K�Tj`o*G�^CQ'�7D�*��	�'�ڔjӬ�`Y���ň}J`!
�'����u"�Gw8�.� ���J(�y��kO
U�e�F�Sٞ5�%��yB��"�Ze06��2K"��Xd�
��y��CgI��J�2�u��oϪ�y�D�0~=���X�"��[����y�R+�DE��%�����1�!�ĕ�B���)	�<%�҅�7S`!��ǣVz,aR�6�Q�U�G�P.!򄇬��l�aeR� ��R�N�8{!�>7�F%�a��D�8�3�.�"<�!�d�68�uV C :��3ޝ2�!�d۾Tޠ�
��´h����F�L�!�+u��tB�!�H��	��%U�5�!�ď�<��E�B��\�d�4
�;p�!��?1��sP��/asR�����#n�!�DY&���!#�9oZ�8E&��z�!�DV�%ozx�ǒ�{�~1*pD�.�!�U�]H p�j^�u�,����.`!򄋣h��P+��*7�:� ��<R!�^�����j��+�$���!�ܪlk�u��$L��Q�ʺA�!�d�	pN���P�ndQ��J��!�Dߥ|���zeQ"y� ci��Zy!��W�V�ڝ1��R�Kwp!;t��1U�!�$�-t�"\z�-]cn��A�HLu!�$��x8���A�]	a�ٲo�
!�� �]#׍�*y���eY�Dt2H��"O�����%bD$�G"�����"O�9"��U����e�+��pв"Ov��)�+;��q@��# ��q"Ony�F��5��u0 �&z���"OXe����5�Rp�t�ɕf��T"OޘбIT�_[��
uL��LyBb"O�@S��޷
TxZr#V��HI;�"O pж�ݶ����QiC�G�B��C"Oz��kd`���
/*B���"O�H�jڡK!��ڕh��|�'"O��-��W
�-�үh
�y"O���2����(�9q}�]If"O��� �S��X4�߼ks�)Ap"O������0��9X��ͩfE8�# "O���L��ʱ	w��?PT�J"O����H��c�z����$.CP�h�"O���Q%L\`���䚁B�^|�C"O� �*ԁUآ�RPd��v��&"O��#��@i��uz1$Ɨ{G���F"OҸ�q�5X�%��Rv�����"O�\o��"JM�u犝.	Z""O�t���Іa/��K��nu^�q"Oh�S���&���A␡T�̈��"O�-��+ީDB`QqW�*��g"O������|M�m���P6�Y"O<�nԾТYB���d%�j�"O�i
���xpT��(M�jMa5"O�Ӥ#S��j₻o~���"O�}�G���]�ya�#Nئ�)�"O�I�@�5t���pPo=�Yp�"O��9�Γ^�&p)�ș -~a "OZ9�v�_�0��c"m�����u"O��[�F+sL��0L�k�N��e"O&�xP%ߧ)�@y
uD�|h!�"O,��	̳^F��@��4Ұ��"O�@@�i�B�f�bu�"O�<S�GW����s�.m�`[�"O�\�Vo�!T74� �
CYz9�"O2��ëE�*�H��
�:t���%"Oz�k:]~�j���% �@y�"O�%�p+

f����g#}��B'"O��{�jʦz7b���b̷#h��Ic"O��i�-�6�2Tڤč:K`���T"O�x�%#ºP���+Wj~�$Rp"O�e �h �]>��+��wq���"O�8�r*۾tr2 g	\`hQYs"O8��5H�{�up1��rY�(�"O�B�i-�8p
űBܲ���"O���;^X�91�K�^ʹ̒��'��h�]���G��1y"Y;��=m����"D���)մn�%����;H���o#�	#&���ٔ�G�OaЭ�G��?7t-���Y����'D�8K�-
�8�n��K�E@�����Y����FPy2`����I�w���Q,3dq�� 2)̀jΈB�	�R	DP�`%�'a�E�plȠ%n(�(�HL��\rID����S$U$�r|�Pb�,=�<A�F1,O�����Զ�x�������2�BE�¼A���Y�7�l����b�<A��~�4)��k�O�D��~��v����$��9<��!�'�F�O8h�H4�F�?�2�r&ʘj�P�'?D���ȶ�^��S�O�x�^���KD�o��mId�՞|��E����
���K�ҡ��	0 r�|�5����i�}Y�)\(���!���26LP FƷu>@���*,[2�9�$k3LO�As��iluC���!a�\����']�Ma7��$W��BD�U���� 69xVkÇjl�DB3�\W݆��"`#4�h3�#	]`h)q��wr~���1���7�~����S��Q���q�' sV�a�/�!gyr8a�Aw�^���4�lR�k�3j�j$��x�6A7	�e8��4�Ə���s����-*�h�k�B�44:�ԑa94�� �
o����LLC��
Or�����^�>Y#�����<Y�P(xf ��OF:y@`�u��E��q4Ѝ<����
Ӎ�.��P �M�.�aGv-������`���Ɠ6�I��a�+J�����±x�Z%�O>���I�#qh�H2Ȗ)u:-{��i�{���
0�t���c�+!�؊4����d�;Z8�1�f�֜"��Jwb�;~�V���K�.6h�k%��|Bm��]���`1�Ksڄ��/ΐx�l�$o�~h"��#V��|�0���l�M��B!�=`1܇N��z2�!�cCD��W���靣�<�Î�.e/*`�cI�K�a�%AV��X�JE���� O/!��/J�<�+d� ?~��u�
�1O~��q�3JEn��3�'mO&A�Պ_0'@p�a���vy�ȓ`o�Y��!K3+&�:��[�r�<�����52/O�6m(�g~�b˗��5�WI�I�$��*��y���/?L݀�͕�@�<H@ĢA$�M��헉[P����x2j�!rHW2t�����:)(&���I�/X�H�'m�h��ܑ;���c(W�9:�'x�Lq�o�4ow��Ue+����'!.�8WΟ��<8��V�4�>IA�'��0�Wm��a@��Y�(�
ni��'�r��DLǒ#d�H�F�7��'���ӡK�R�b�*��+)֌��'wLD�g�\1'��#`ŭ*(��'66�f�	2ʱ�h�?MDIy�'� ���ݤ���PAGτab�'->X�FH��p\j���)U+ul�	�'~��+���\�tq��K�6l0J	�'F^M�2-��=�&ę���fp9	�'&�z��z�@���z|��'���[�M���D3cĜ�>��Yh�'���g'�%p(�T�A�>Sp�	�'[�y�5 ��:?�T�%!�>�v��'��5� �#�D�85nN<�9��'n��zB�wxE��I�Bl��"ODU4�/:�9H���+R���"O�r���r��d ,Q�ب�"O����.ف
�v@���N-)�yz�"O�h{�Nՠbǖ%�!�Kq��"O8|P�,�&@_�U� ��"�иB�"O��q�d���Lpz*�){���g"O�0����@�Q#�!�H8��"O��C��+E2Tbc��S���!�"O�����O�f�l��*��@Pa�$"O@d@�c�2HZ��҂C�A�f"OB��E�@�F�+�.چ&`�5�"O�d�P�NKȀhE��OFz�"OZM�a�
?d4�b!E��;cj��e"O��p�O׍Hn]2be�$nV�Ȣ"O<�K�@V'*�&%���I�aH}��"O�`@ M�d�Y��ɛ,4�Fl�"Ol��L�(T݈ԛ�Ԇa���"O�0bR� ?' Epg�V��썓�"O�0�Df��qEjB����DԊ�('"O �:bN$�H��BRҖ�a@"Oĩ�D��Z$��
��i3�2"O@�c�B�(���8vϔ2N�Q�E"O�( &�T�o�Tc���K�9J�"O�c狎+�X$3T�b�΄0�"Ox���cS�p���%�X�fx"�"O� *d�'��0oj��W$D=e�t���"O�r劝�1���Y���LƐ�@"Ox8�Q �kv2��'&�.b�b�R�"O<�CֿHN��EܕZ�>��u"O�i��	���(4�Ɂ\B�"O��Ai�1�^LI��Z�yZ��0"O�
��?f���i�7%Th�S"O^h�E�?��cqoر]��R"OV3e��-v����fj��U�Qf� s��cU�BoX�`�m${G�,������=��B+D����8C��4������t���(D�d���/ l�&��b&D�D�F�/Kx-����6�p\�p!0D��J�(J��HA��H��9/D��33D��)���$@���B�5{���0D�,xP�x�DY�զ�/���y%�-D�,��oU�^�bEqr�)94�ٱ�,D��SGK�Z���!a�O� Q��i+D�t	���/��$�c���,\� �)+D�����T/Ԡ�6bW8%_�q)*D�\q�牤+�ĉ��Y3S���q`'D�D�G'�0e��.�Jv��� �#D��(���)tDɠ�"j��1�N D�t��G��^�$ ������?D�<�ALW�}*Q;,�>c�E��"?D�� �i�&�6QZ%�Af���d�=D�P��m� Q`C���+D�(8R�g;D����8x�̜ґ�L4/���S`�5D�T�H s�,�q�H��'�N� wN9D��R�͂L�����K�j�� �`8D��k��3R����P�^�'��D`�m7D��O��Vm�
d;0���6D��c!��[� !p��)� P��1D�(�@��=:�DX���F�횁S��/D�@hČ�9n�A3�G�?9=�1Q��-D�d�M&>�RLR���2�b�`�>D��XF��f���z��!��9�L<D�4�e��/ژ�ɃǶ�,\�f�?D��	��[�2ج({k@�Mح�ץ<D�LQCN�!�X��1k]�WcjyF�?D�4�իQ�`�����Y�`6f�qh>D��!R+J�8�iGk�*�81�%K;D���d M�ZXy�jW�*�ň8D�X���J�0��)T'��!8D��!�����؈�0��3]ޜ���5D����R�N�(�D�Q���%J3D�TK0� 'h��(�M�&u�x �@E7D�����)fH��j$ޘE74���o3D�p�&���_��X��ڞ^m0�P4�3D�@bp��?�X��G�Y"Ѻ����2D���amʣ̚�
'g�#M�IV�2D�x�iٖzE&q��Wk<v�1!�.D��)�-��p|��t��b�M�&j7D���.)�(T�r,��s)D��bF�?&M~�����iS��:2�'D� �f@K�
Q���3톃RZT<aC�%D��3�/�.�ȔXK��:��!�&D��Y[y�8���(p#@=1��F��yb��kFMi��N������y��j6�,��H�&��������yn�,jz�2'N�4w �$b��yR��O����iWuh��ՋD�y*�!L�~	K��8U0$4[�����y��M����#'� F���s���y
� �,0f PI>vd���>� �"�"O�<�B��}~l2��^) D!"O�� ��{��r�\�#���"O���3$�
M'LTT*E�U�-[�"O�$�@��.���s��3���['"O�#��I<ے`��lĭQ�"O�$!H�p@�)ѠK�=�Zᚡ"OL�;`�>NVX���
�3�"OB���#$�1�f �`y�3�"OP �0�#Y h��`��!3`nQ�B"O��Oǯ}�h�r����^2,�c�"O(u��h����"��Rp}Z�"O><�)r�p��Z$���À"O~�x�-
	l��xa6d:mРc�"O ˂Û?Fp9�q�
*�����"O6���F]A���*�OQ�4_�y�"O�]�� �9.Ș���
�|\��4"O:�&��8^�)��QN�^��u"O6������n�m
���/7&�"O�,��EHҁ��/�N�k�"Oȝ��E�yXj� �j�	l��X�r"O�`��h� �4�#�&F{� Rt"O��â��ZӨݲ���
S���3"O24)�,��fLjP: ���Tʠ�@w"OjtCsI�kp�IU�T2s�|�7"Ob=�MߟQ���{r��2R�� su"O2DA�2e�dP!�
�S��9�a"O2؂�F�Z����b�T �~,�`"O<)��K�1�`jc� ( �Z8�"O*�CE����:���͂�v"O���SC�+C����J5F���b"O
�Q��7������!X��k�"O,X�S��?���1�jA�%��"O��8%HM
7"UzT�O=-�i"�"OJq���ѓ,�JZM��iD/װ�!�I0vL�� �N.��a�K5*]!�ʹk�nh���R-r\h�k۷3�!�d�z��(Q��vU�*��=�!��/Ws�=Q�A���P �]cW!��ʞ,��?g�NM�5�U'@<!���ⵒ�n� {�@&�`�v"O�A��ҕ0FrĀ�	�PV�"O��+D*7B5�i���oc����'D��s���?q(�c�G�A��y��(D�\b��9{\��$G9 0����'%D�pk���8��틵�[�و�#D��a�@��	�T�Qs ��Iq��B�.<D����ܦ{}�TCr��ELА�ǥ4D��+�S�4����ĕ�Tu�(h��1D�4��_�VXp�ⱭΆj��h��);D�t�Q�Z!V�2�r�KpD�8	�:D��+d��!n'��SG�F�#�8D��B�!V1���G(D�1>.���"D�x���VE���3��G�ZM¤���?D� (tn �7���c���&O��P���;D��;@�J!�>��e� ��BR�;D�l� a�j+&@�Ţ&[�h|"�<D� a�!]�[��	o��Y�4�Ӆ	:D��Xs�C�M�@MSD�2<��ҡ8D�l�D@�-���Ƣ��D�@C3�5D��x�f����`���M�g��l(2N3D�d���P(xd"��H��4m;D�Y5 �%����bo��F7v�T.D�ӡ�@�V��c!�&����*D�� 1#����p�F�C�T�J��%��"Oj��d!��Z���2�e��]�8x��"Ol��d�\�,�ƽp���xF.�$"O�(�n��j�@�p��L��!sq"O z 朅=���0-�d,�d�"O�m��j,��cv�ёq�QK�'R<�2�1Q@0vk�8^�U�
�'.��c*��M�hW���p"O�t��͜>l)��5xo��R"O|�"�S��p���(Q"̛ "O��*6.�
*�����ZQClA)S"O�a�Ł]'f���#̧�ڄ��"O~�gɗ���P�B@�z�>���"O��҇59T5p���4@ �&"O|�̅�'}ؠ�C �t��r�"O����C:B�(X���J�Xelq"O��jԇM�ɦ�]-|A\DC"O��k�n	G���T�>�p�$"O�	���|�X�S����i+
��"OX��S��1�$q����Ė)�"O��X�MD��a�#�|Z8�h&"O.���i��}��8���@ވ��"O̴�~I��L۝2\�MX�BJ�<�Ā��7����
�N�į�{�<1WgBUq�@F�f� R }��	��<c��̥a�޵�dJ�6K����ȓ%�vⶄ�A�½rM��(�n���S����w�A�kJH�ր�,�>�ȓ}��P	R�s���f�lА��ȓS0��#h�h�p��$�BR��}��J�� 9WmE�"= �������,\��"O� 1wF( ���1�hD�M��ͅ�hT��,M���釿*�����AL8Гhˣ"2de� �7�P�ȓG㚔����|���G�[�
�����`�T�\�<t� A�_�|݆�~����$N�6�B�2�阭E�b�ȓ	�	 '��L��CR�L�s}N��������2���)�?
Ը�ȓ_�8�v��P."���B��6��T�4�[�
/,`���.X*s˰�������a�js�m\�4}��J���d"�J�qq�,�cDi�ȓN
�xb�),i`��lÊI�|��ȓ ����5̘9	�]�䧎�-�P��CP�-I�fK��̑�Я��u��k&�E����??���Y�ゝ+:��ȓ]������2m̕��m�}[�1�ȓ7�2�P4�Ȋxf���+�4�i��n9����W�`��aG�)�6��ȓUyM��>U&�� ��HMnx��>}:����G#XZ>��j�	vن�)aT`��K֒鮙S6%v�$@�ȓ=U0��a�D��<�cQ�	�F�ȓ��A�Q��P����k�8���^�R��CR�%K�lM�(�N�ȓ�
\��_cZ��B�읳.�d��v��d�sn��W��LC����t��:�$9j��f�-S��496�Ʉ�o� ��k_.H��ڃ�ծF:��ȓlF�m��P�,����C�X1��\�ȓd<����vê���#�<X$!��G�e�1AXe����+��U�捆�=j1���'*X1��C��&�Ry��S�? t�th�ii8��g���j��!"O�mpS%R�B52в!���)���˃"O$�rժ6�ʡ[�-͓A6�z7"O6H�D��E���I;8 ��'&V��#hڌ>�dK�b
�e
�1�'@�	��S�-��P �W�	��q
�'����
X?rAf)���� i���'e�!h�O�7h��۶d�&	�8 {�'��1��!H�kT�����FP��'���Ȳ $�±�cbP������'z����@�����Sy��'��e�QN�!��IR��}�*hB
�'�j�0I��S%�#W��l��ȡ�'��9@ ��P   $
    �  )  �'  �0  �6  '=  |C  �I  �P  �W  ^  \d  �j  �p  &w  g}  ��   `� u�	����Zv)C�'ll\�0"Ez+�'N�Dl��T�1;OV��g�'D<y�g�4gfD� .��ږ}����'?���2�O�Ey���l܄@��"4C}ݑ�+��?e�'�W�?��F�8?�X����k�&����	uV���%�}a
U�l��KV ��u!?��4�'�*��&I:M꺍1���"OZ��C)B?|��pL�O�4��]�Fk�	8�ΦuᔣRT�I����ş��N"o�@��`j�~��2�џ �	��M�3�ƞ���O �{�����O���L�;^DR�$�@�H{��[���O�$�<���?��#G�4�'���)����D�ř#�Xݻ6�_*%&!��h>\�xw�!��q��������<�M>��'*����^T�d��m� �
� �T�r�QaB>�?���?����?a����6�I;G���P���^l�}
�@�N*�d�����ش���z���� ��i��4N��� |�\��G��I���2<��a��՟
Ez���O�Ou��"C�F;�X��f��H�*j�XD Ԭ˅��|�ӿi7���a�S�?��S г�VQ�F��0�d��%��D��1CN��M�6��,dǈ�`J�?zO�ɐ��A����5)�=���iӔ�oڵ�
�A2.�WQ�	��D1i{xi�4� x���0d���Mk1�i�27�N�U���<��(��/=El`W���5�*;��ē�f��e�^?�	Yb��C\<ɢ�i%�6���8%��3��Z�jO�j��苣HȺc����#�-���3B^�F�4 �4`�T���ޠH-d��ߑ8�D8���'�v�Xgk��11.�z�i��'�
��'6�O����O�MP���ݦ��I؟���D�R�J�p+
�2�2-��d���$�	�\A��������'sƪq�6#J7 �2��'BS�
��a7n[+=o6,)s�*C�ĜA����p�f	�j�>Ā��^L:�k�*J�  6����Ż�C��]ʰ�w��HO���V�'�R���a�i��[)~ ��I�)5*��Њ�Or��O��"}:�J�Aq�}�%'��{��y�'�O���ɟGw
m��J�f �����9A ��6��;@p#|��wE���i3I-��1��9xd�S�'����g�
�IБ�*3�T���'��H�G�BNP��i �9a|@�']f�2p��	!��܎,UV���'�Ą"T��$7x������� �'T�CM�p�����ے	��	��k/��Fx��	E/k|�ٚd,�p��{dOM�	#�B�	�lL.�b�s�H�*A���B��u�q��W�
�a�V�F�fC䉄K�*8�f�ky���4&Ƴ1+�B��;%	J�I%6m� � A�.|6C䉩<�6%��aC9P_L�H�F�&5��r����	f�,��MF�35a���Z�}�B�əl\HS)Ż 7�ܹ�c؉�B�	:	��i���S�\�a�TP��C䉸���
�w*P�"B��zC�Iz�����/H�h�8�"p��d�-�d�l�Y~BD���GK]:B�{�J�7�?�(Ol���O ��@�P�E���1�r�����ȟ����J9�bq`C�6��Zs�?O ���	�hڽ�ea��#���$ڊaR�HZ���!]�HZ'$ժ:�ax�f��?!�iP7M�O�(��ʦo�8���Y��N�<y����(�Ա�0KF�|��]BgO�jon�:1�',*�$����B���u������|�X�i�+���'��.�N+D
ÆH�)�8�����Qe!�[7u��q��j��C�́dMA:KM!�K�7B��r������c$ �	.!�dב!Ɛ�GI�1s&�ش-SB!��$�@��wKɗ�H�Qn.w!�_pf��`mL�Ey����M%Pb6��O��d�O�!r��/|�����O2���O��.N���MIA� � ��9�����5F��;R!RtRs%��Y�$�� 3��O6O��b2/K8@��`�Ӊ5�A��  ��V�K����?u��P �\�f(1��	QPFQm}r���|(����`^oɆe�eÕL&�V-�<Q,Ο��|�I͟\����<9Da�&��\�`)\�"�ji�ȓp��@ �\�M��sB���H�U�'��"=�'�?�/O��a�O.Z2���ǔ:U�ʉ��Ok��!�Ot|9�!�#O��a���%�X���-��s`!��8y�l<���T ��y�"ʓ>�6ȃ4Ob,��U�E5�|3�C�/�摺vN<6�@.�OH����0:H��;�� ���c"O��z2I�6I;�q��L<_��,#�|2�n�^�O��S�Fܦ������
b���5�ƌ� d
��ߟ �I� Un��I�|̧CvH#s�!� �)S�|���� ��c U9@�桩"oC Mqv�;�e�'���fIC�O~�h2�K�3:�(�s���<8�b�Ƌs�"́��ݬFi�/�*zd��	����'�.��m����B�cA�:�jx��?������(���b7ͨc�L���/`�T��'�V��߉T6"Шa�^�L$fJbP�(X%��1�Mc���?�+��d2�l�OL4�s���sJJt���חr�"��O����@q�KGբ̐�I7�����E�W�͟n��GoФi6H�.��0��D�!kлd��5�ƍwS�l�Ҋ�4�̙�N|J�d̆6|8��P�J3)�T�g��b~���?�����O��e�k����Bθ	h��K>���0=	F��M�Ve#�5t���`�'�ʢ}�'R�
`
�sBKX�������с�M#��?Y��'��
e�P$�?���?����y�����������H�z�	��7�h����X
�o����QrP>yϧ��9h��C���d�N�3dw��t����d��1yݴA�*գ�����O՛i�t}lҊL�������)q�\|�s�X2�?Y�OԵ�F�'>��'�O2qJ6��q��\+yZ� I��%D����׌ b8I ��#��}�e��<��i>��	ly�hZ�z�4�q�]�c�̲u�X��u$!7���'U"�'���'8R3�^�戉j搨��N�s�����3�F���ȅ�D;.�ҡ ��?���+ 2d�#G��CTz�����E�Pݢ� �=R�2���;��9�4i8�"=��&��	f4mkB+T�{K60�uA�##�p��I���D{2�	���ub4c��xI�)Jd�U4C��Ԝ��.�'FŚp��*��
D6�Od�n���?�B�nҤ�5xW����\+$���*�SX�<V��H��$�fa�$kT��r��BV�<ц�ïA�썁�ǝ1�N�b�`j�<A$ 9��A��i�4nʥ��d�d�<aƢ��*�<Q��+��U���"��H]�<�@.��6O�L	�:,�Lx�CGX�'��m���ID8C��B�OM�C���o�OI!�$J�t:�F�Է�P �$eA�cE!�d�U+���u)@`˼��a���k9!��$�B���J+=MH� EO�w$!��;^�t����.]�d�B�<!�$+#qd�qe�D"-�=���⨉��O?����ً<r��`u��o��`8q�i�<�P�U2�qa�k�A��y���L[�<�)L#a�h����I�5B��A�<�3�j�A�7�]�&B4"�/}�<i"�A�i���W&t8�¥�|�<Y0��=f�k���=#yb�-�uy�C���p>���֡��P���ôP��a�dK�Z�<���X��Dݚ`Z�!��P�Q#�S�<D�Z7��h"A]� (�*�*FT�<I��!}xe ���9ju�S��K�<ɑ	��B`�HsgҬ�ڔ��Ex�h�Pk��l ��@�s�03�O�@]~AC�%D�X)!@�^�.IC��}��fi"D�,�@��$a�X%�u���~��$��d?D��Z���#AX�r���M\��)2D��V�I5c��4Xeǘh"����-D����L���I�E,�,/|���"�I�H	>�~r!�U��N�q����P���ˆR�<�� R�G�x	6L�{�*a���IR�<(�,��Yؐ+Һ4�PLA�/�T�<��h
� ��Q����{̥��
e�<aEε���-��G��]IӃ�d�<A�A�._q
��r,��Eu�ɕ�A�	�H?�S�O�Z�3�A�.Y���r�BՌu1@��b"Od�[a/��M��0��`��m}���C"O�����.0d� �0/(}�Xc"Or�j��-3���:����\�&�t"O�����J�r�o�=�hu�""Oh�A��K�i��g��qAgU���P�=�O�H2#�`�["�B�Z�l��v"O� ��A!�|K�P'��j�z�B"O$`�6�F� (����JR���"O�H����3R���s��@`X"OQ92���]c@l� 1.��a�'��}i�'ش\��n_
���
��f$�A	�'��p���ֹt�qc�ЍX���0�'v���nK�w�>L��%ٔIf�Z
�'�^I�惖�>��(�暖FD�`(�'�\p`�˧i�p][b�B*HN�š	�'t�Jd]�9�ND��a7k�蓈���"|Q?���WGn�����d�Z��c*D���V퀴p�4C�	��(a��1�(D�|Kf��l9~!��O v�2@&D��j�($u��՘�ψ�^�@��4�(D�	!�O�;�>p�íŤd�(ږ�&D���%n���ѻ�`��m�<��l�O����)�]KFH��g�hE� ���CQ%�8h�'��̈�nґQ�:�D];BֈE�	�'�`��/�^(��l��<Z��k	�' *i��bO%v�DXZ�GU0��U��'������Y�=�fS�%��K  Z�'\x0��
5B�C���J���-O*�Z0�'���b�+{R� @d*ǔD~�Z�'��0N�'Z��'�/Xp�=��' ��Ȳ!P�Do��XP`Z�a\,��'˲����8~&���CG%]R��'^���͒�u&5�pnZ�%.��Z��h�I@~��
,Y��00�
�����9]�ɩ��*;(�H��LI�9���ȓ����I�4SSG�*`��ȓ�ٲ&#ՏI��s�%
	vR��ȓ,�֙���I��r�z�̩��y�`w ]-5*��Lž�G{R�A:������2Hˎ/��as�+��y��!"O�� ��Q~hD��&�[w��`u"O^]��&ކZ����dH<_ �"O2	�B��>��Pi�
L©;"O�Ui`Q�08`25o�"t�n��"OFu�'+
*%����(�M�FI`v�'M\]����,_U�����+L@f��6��Q��@�ȓƅ�'��Sw�
�IB&h��q�<�'����A�43������i�<!��K2lD��WC�1#��]�SeVO�<�\ڨ���� "�Z�����E!!�V}V9�����6���ۓl@< ���9E9$����/gT,��.X�H�jR'j˂]�!��ԣAUԙ�Sꘁ ���h׈ȷO�!�D�B�����K@����܃Kn!�$��S��q�b�+8����|��	�'9@��0-��g�ФX��S=0^(�	�O����t�#@T�@ 8�A�G��m�ȓlH��%��vz�t��ɎN������8�0��>9�=gj�p~����p+��sn�5z���ÇO�$��[�^���^z��ܳVbS��	��T�&Ѐd�1rԱ����]��F{������B��h�B����m�V^=	�"OV�8��L�{��C�J�?�b�YF*OX�C��h�z�$�#�X��'(P�z�l��|0z�xU�4l���S�'~�S�&]�j�L�� vI}�'�8���}\��;�'Gz����LU0\Gx���.sV��b]8��K���,q9�C�ɿ�N�����G�z���l�+���� ����MR�i�(�faTO'��r"O��V���o��� �����U"Od�����t�&�_��yD"OlD����}D���CdvxфR��"p <�OF�!�	j����U�4<T���"OЙ�M��n]r9B��/3@�R"O��&���n�b+��J���1"O:xxL
wȽ����;J=��3�"Op�Jl�;a�}�a�ZC��� ��'y&9��'�f,B��<.��7k�<!2�R�"O�-5F>�
�Ã�\.�ZyY�"O��{��D�X.�YS,�����"O49�S��9Y�N=9�`ߋ6��i�D"O��֡˚;td���  5R�6�Q"O� "U	ǥ{�H��v��r�P,��� Uw��~��AW��Hw��P ���5�Tp�<2 �TW��(��g ��J�K�j�<�"�(4*X���nL�� L���e�<�7M�"T^� v�W!3&` ����a�<ٴ��w �hF�3$�@��C�<��D�KJe��m70;> �ЃZ����FK+�S�O*�y����met��],��"O@�2�����⤜<N�V���"OT�[�J��a0�}�VJ�5z>9""O��i�?��3gÞ�8y1�"O�����^�趧W�qe>��v"OJ
�	�$.1i��8d��\PZ�D�3K.�O�xH���,&�J�A��o���%"O y:�D�2�B}��C1�¹B"O:L�陌|�
h���|\�"O�@YE�U�z�b��@-� fI��"&"O��wh f|	���7"=�8���'�j�8�'&��ĥY��YS˖��
�'FEt���z��!"�������'z"��F� ^C��Ϗ )Y�z
�'l���� !^���`��(�J��	�'g޼�N �$�Y�"-S�q(	�'g���p&^{���0�Cܲx� (S����TQ?�7Ə'u,I�KD������$D��1aH��d���¡;�P��5&>D�䪧FBSs� E��tR�f�;D�4�g�̊)+u��A5�`;�=D�0/��Ow.5��Hݨ'�褰a�9D��*"�G� h��R	"�r�S�K�O��p��)��\i�D[2��M��@�Q�����'y�٘0�Z�#�,bU,D,�1�'Tp���C?=�=y���8T����'�ޥ�G�\80 ��@��/�x)�'-�}����	d�Y��)VEڡq�'���#B�O�O�~����9�̽�+O����'�|�F�_�T.��A'�*W�pY�'ݬ�r�.=ơ���#�LC�'�`s�EY~�����Ġ��'(̰Ad��\�DqV����X�'�x�SD�,.�v!,�L��;�y�:��0Q��"]\X>����T]tf���Z�ň]X8(�(�h�`(� ��m�<9�H؎G����[�g�̵X�Og�<��jD��.Њ�Ƅ;>f�H2C�e�<�i�N��q�1�9 h\2�_�<�6%�>G�9�@h���d����^�'�N����	����]���`!cG�!��:䁻��Hp�|�`��[X�!��0�:M2dGW��ؘ*f_!�� ��`�灝H֘�y�JRU"O8���%o�1��&݊ �
-H�"O�1s,�Jr2͈���0-�XEz��'8\�[����1(����OƘ�j� \XQ\��UI6��B�LL�Y2@l
��ЇȓM�)������H����	(���"$5��I�(6c�T�'ۈ�|͆ȓ`��AI��Z�rbЍ��Na(X=����Y��@��D;L��dμE�.��'����k>d�Vk��LnY	ci�;.=�܆�چ}�Qh�8X�4��o_�C��ȓp��)�ɜ�k�lyfMG[����l}H�bҡÃ ��P� DJ�̈́0��6��0a7,��/�R� ��J�LC�����03� �I�6&@yPb�CM�b��P	D�o�bB�I�0Ƕ��$�E!e%XL+��N~>B�	�(��=`��2% r���H��#�B�ɗ��4�3��i���v�	9@�@B�I5D|�c�[�lk�Y���}^C�	�s�I��H�8�g��]4�=�wc�O㶸����+PwL��3��,T�|��/fb1*  ��`y�CL*B$��ȓg&P����
>M�
��� �$b����J� $	�5M6��i�J�+b�� �YZuH�=�r��o�$k��0�ȓTՔ����B,~�6��Q
rp&��	��#<E����}I�Tg��BLa��R �!�5	���Cn�&P�qV;h�!���W�С���E�F �!xVcJ�6�!��;X\��KԏZ�����еQ�!�ğ�&М���#�y(a�?@����D��=���N�X���8i�s2.��O�����|�����������x�aA��8 ��P��?)Ô��?���?9��!v_��)G��>�l�Q��Pcb���@�h�t��/�,�(�g�֎׈O^���K�^2��Ӧ	�1�b�z�lr�ђ�噩&8�ɠ�Ci#����a,o<��d����O���&�ӐD���b�ˍ�������2G.˓�0?� �M(�����ƎN��AP�Kcx���dZ).�%�,A6�[�%�mm�I�bn���֟h�	_�T�UKR�'N:9��{iyQk��ia�Y��L��?��HR#����u`�'�ܽ����=,���t�'@⁓��ӂT�]��lZ� �q�ԉ��"�
�e���s
�^wn���~-@�^l/Q�Եo�X���r��'��������ӂV`��RC��&ᾼ3K s�<�A�E�c�*�p���i60��6HW�'��#b����bQ@2�쎽P��Ƥ���?���?�V�8�y����?1���?�ƶ���;|�Q�-R:��0�'@�Ş4��'�Ʀ�3ra�4���Yv���?��'��'
`�x���Xj��a��#wx�*��K� ����&�`1p�ød �SΦ↖x�+��r0�]�D���41R����d�=#B�'�r�D}>������P$I���!%l��Պ/D��
"��S�H�0(ʁn�l5B�@�O2�Ez�O%bP�@��ԹI�]sbm���
h�c� u��2ش�?���?�,O1��
�[��pa�5��%O���D��� (a'�M������Bx�`Q" [z�&%a��T!���`[13�jh$�fP��@�Sx�p$��O�-�֪ټHJ�R�k��q�\�e�O�=����&
n��3�E�!i��5:��X�P!��^_$P�� �'~zU�ڇ��I<�M����G�Z���~�MO�
�8�2��8�B�ꐯK�����O����O2-�Ѝ6y��d��/=`�&x�i>�[��+�#��
hޠ`0�=�]�<	fE܈L��q+�A���)�	=�<aA ��-�B��g�7�x)���O���3�S.o9��c���:���D�7L<��0?��	�I��,��׸�x��u�Dx�4+*O>p�'�&/�iRw�
d�fI2�]��xr(�����ey�R>����ȑ��ʏ3;��"��/T�8 �ȟ��A�����As�)J&��8��S�OF�$�$�=#l�ms#O	l\˛'r$z1 վpW�`s�ʵ!�?ճ��"3�.k� %w�!���a�4*#�Od�D<?%?Y秀 ^����1J�%�ߜw�v��"O�XHb���L	V�y6�Z:���`v�	
�ȟ�]��A1�f���!ˠ��a��Op�$�Ov	��ʎgVz���O��d�O����O.<��(D�/^@�(ݙW�tq���+�H��"�%e!���g� �'��'�iz�NG�+s�$�'��9��=�D�Լ �tD��$C�z���o�!��id� ��I<�%
C*��pScwΠ�"dKb~����?���hOv��f�n�% ]c!�ㄔ�e@BC��*YA��XҊ�6`��e݁ b��r�����'��	�;��D���]��64����L�&1���Sş��	ӟP�Iwy���̀�u|<xf�@�E�	Iin���G�W��+�jʒ{%��t *<O���G�kJ*��u�J3r��{�d�7����i2|v�"��$<O�����'$�����ǭ/���#U3C�v�V�'�ў`F|�k2#�:���A�	�̉!�y���7p<8Rk8/t\���0���Ҧ��	[y��Ί��6��O���|>���
L84���v�rp�Qc��O�i��On���O,����v��u�D��#�� �ug��a7صӧ�ө&Xz�IA��OJ� L��v���)+&���O�+�T�95&��VC`3��¤z�$HѽZ#=Y�ȓ�����G��+��C�Et6\��^"6����	��?E�t�$h���G?a�.�YrH�A� �@�>H�I�.�hy���M1�@T�`J�20�$��?)��?��4���ӥ�D���Z0�� Ҕ5�ׁ$OУ=!Gg��|(0hr��iR��pDRC��w��%���~ڑD��A�~���Gn�D-��hS}~r������,}*��$^$m���e��	]��ԁ$]�Z�&'=?94�>	G�WR�d�K�S}�|á$Ó��I�%Z��b�Q�}��L�0��<�r�[�\QԘȶN��+���	Ҹ9�O Y�Ov]Q��>q[?-�6�]/`�E �/Ӭ1����+�O��
F�>)],"�zW�mh�(�Y
q��Ţ5���?��u�dt��d��F̛vIƮI$��ӗp�R���j���D�O��Nj�?�Ĥ6#N2g��!`�t��n#�~BH�����|�k����'�J�!�c�9'dFrî��8>	p�#b8�; ��l�	���p�i���|��Y�J̍b�`�L�U;���ɟL۴�OjX����<ц�QE?釈&@��C�f��OQƐ��K��r�'=�l�����@�B���/�.m���'�t��U�ZG@�E��'`����ߴ�?�)O4��|�S�l�I˟�х��.J�X)�v�*N���
�N�����O^��hO�S�K�$)�4�I�&�Hk�I�W��C�	�]���7b�2Ŋd@�&��C䉖jq��P�ܔSI����L�#��C䉪�=�aƍO�:ٔK�nC䉲z��@Rb�˃v��요�C) (jC�I-5�:��$͐%.~�Q�k �w>C�I[�|���u�\���;Z��B�	�aRDl�QF](C�*5�PJ�K�B�	*!wN �6�R[X�0թظ+�B�I�F��i�EQ
~$R�0�ɷ�lB�I�d��H���'H@(G�GJʖC��qt5ض��w�`H6 �7`�dC�	3��b�Ď%��Q�q`I�4(pb��QrJ�r��R�茰5�xCgL�/���ᦏ*z
<�����b��V�J�Y��t�`%�a�0hȖ�Rg�D�/A
0"���5���V�����E�e�:���#�U����S�V�r�Tl@W�|x�):3�ޯ7BE���#K���4'�>� -�p&]�v�[�&Z4J
!poq�ZLխn��P�J"h�����Uҟ\��/)dd���h�S�,O��PS����	a�V� ��!r��x��5�O���3Bڮv/�tw���1*%Y��x2�L5�?a����'�ħr��1eJ̾n���9�
�=(3*=�=Y����<�T/�v>"���@���Uؗ��U8�s���5U�J	��#tWr�#�/P���d�Or��D_�٘��~*|k0��"�!���<��!�S�L�)&�W�!��ݏVC����̀+WҮ��7���m!�$���Ԫ��0 �ݢ]!�Ӻ�ࠚq�C�z��+��Ͱ�!��#ж�H�-�r�L���
9!�䋌ac�5Rc���.Sԁj�-C�S1!�� 0�`�DAz>�j���jל]�"O:i�0&�6X��C�W�4�&���"ORaf^tռ���.h��aS"Oыp�72���	"�����1�q"O��I6��	z��3��2"O�-)aj �[s$7�:m��0"O\%�u�H��ZH���Ƨl�V��"O��j�?dM����H@����1"OB :��F�2P�1'L<�V`�t"Of���-r��j��J2U��rb"Ob$��A��7�v$��g�^�=)�"O���8 p�$�]�*�S�"O��S�>⸴(F��l<��"OJ̚���]P�@��A�'���"OH�ؠiٝ۠k�	�,-��XQ�"O�4J��:�J| ��\�����"O�I	� ^t���%�V�8�qJ�"O���Ċ o6��C�v�f0�"O� 0�鞖U����"�Y�J<�b"O��[��߁g�L�!�
}��"O�$�eo�E��%h��ݨ�ąsr"OޘQS���>��Hr��!3@`2S"O�\���	#8��X�=A��@�"O�}b�C�)p�br�5P.JYV"O�)��@�]�L�	 �ۤ5�����"O��r"�J�<���Ԣ8�� �@"O,�PgF49�=�$m�������"O�-��8P|���잽��Ի�"O��&EM5?l>��lǴA�00"Of�C&Mx� @*�
E�VT�U"O�1y��8y�n�ÇI\�b,�5"O�y`*ܲx($�0�n����	�"O�ԑ+�:b�$m���"�s""O^2��6G"�@�G��	�@"O^y�'/��J��0J�D���"O��t�/S����Hӎ>�8��"O>%�'���~�����͡F�2F"O��!vҎjN���cm
B%�a�Q"Oj���L�ț�!���Tq� "O>���>
�����P$	%�"OV ��E�*;���dL�a��d�`"O\�Q�Zv�>􀕢y[�	��"OB�����*R�E	��E��|I�"O�Й� �������� "\�$��"O�0�D.��-n$�2 �zYі"O�q#bD*j�X����$�>��"O����a�.'����S ^�S��]�V"OpS�E�$�� чB�py�Q"OJmx$��D1:�.էC���"O*�z�U%�f��q�	�+V�ɛ0"O$1�s�r�֤k�Kn���"O|u���3�L`� ǒ�q;���"O���兤��!���+V3���P"O(t[�� m�����}.H��"O|��'L)~a7�H�Z��a"O�qg��࣏#tt�6d�9�y��>��c�l��9PMr�����y�ʏR� ���˞�.ʹ؃�h#�y������D�,�6]a�J�5�y�,�gt�27!Z� ��p�Ö�y"��u<$+2�G�����3��y�Kмm2l�(E.n<�A���yB�#s���3V�'~+8�ZV���yh�V�t(��I�y)HH������y
� �qR�KT-� 	�Ǉ��v. �"Ova�r�@?Vb<�4-ӯ	8��6"O|9�$@)zj`A��K��L}j���"O$ ��ڢR��L�3���Rd�m��"O]1w������]2��8T"O$9k$H�@E�sdFγ\uh� S"O�y;e��0Oov#���N�H�"O�%ʀ�$@V�;&��88=
c"O�yX����L���շ8�}!�$�b����k͇_S����:-W!�D�9x��1 �K><��[�J�~M!�=wPف	�~3�da$e �}�!��M�FJ�UZ���')�فtd]:�!�$�<a'�0�e��w�`���{8!�ā
b��1�f�94 m��-3�!�D�*H� �q�R;\Ձ�BT�4�!�D�3+nH�8P�ڼ`�N�X5/M�_�!�ރH^���*$?��,`WNM$P�!�Dg�nܻ0���:hl!HH�P�!�Ğ�w�.��'&>²P:Vh��u�!�$:>��u�T*�Ҁ��-Y�!�$ݺU{��CBI�}
ޭ��G���!�4��Y�GM��R�L`���6�!�Ĉ"Q�r����X�0Ly6�յ"�!�W86[Bȣwf}����[�)�!���/2�p��,�$r�=M˷3�!�?l	8��R����Te�|�!��.H�B\��ҝ2�B�9�CǗ|�!��V��J�I�&�3$l۶�ҫ4f!�d�;S����҉��V��[3,��b!�dā5�:IP2�Jl���ٜ/�!�$�#yn�#�mَ4��0 �i�x���d�P���H���9SQ��#��	:�y�j@�3���#g�"���Em��yr����ǫ ln|�6��,�y2��3��!�&��L2S
���y�j_���I�o�� @&�УG-�y�"I��*� �u�.%��+/�y�Ūv���`G+�l%��ʢ���yR��2
_ځZFҏi��Ű��[�<�!KK'UnlP��M��!�8�kz�<91�D�	�:}����*J�uL�p�<9$,�J#�%B��éB%<��n�r�<��g� 56�����(\����w�r�<у��'�`�nJ�f�m#�d��y�+�����0A=]*��t���y��ʅ
�(w�R�8 |z��Ť�yb�ɣ5��@p�J�|��]`��@��y
��̓FZ<oH�T
��y҅�[�݂�J��N^ز�׮�yb�-d7*�zf�M$P-�r�R'�Py⤇,G��%��-%p5��S`�<QBoy�|U񤨃s��jT�ET�<1���2�ro�
<q�KP�<Ad��[�H�C�����`��]G�<Q3�S/s�`3f�K*�n�c���M�<��Ӕb�ؤJb��K����寁K�<����J".Ti���B�@�c�bJE�<�g� 37a�=&�R>�hiC`gx�<�V)Ã7��r���^�F5⩔L�<!��Heb����fz"A %�H�<�Ό;~g��H�b��~�!H���C�<���X�bO"�P�m]0R�:�ȄCIX�<I,�e�n0�')�+1}�iȐ��z�<� �@11jΝO��Hӊbz�y�"O,dbŠ��7�h���F^T^��"Or9��G�x �4����B^LAT"OdX4��(e��PTfţ���"O8Ipք���2f�'D�2�b�"O�E�eM(U+|t�ʂ�&��U��"OTpa�J\���%[ 	����"O�l�gF�'���a[�B���S"O,DAqGϹ3S�ȫ���.m�Req�"O�����E",1�u&��-�멋q�<�&��=F7<DJ�.�V�(��w�Bw�<��CO�O#�I(�a�|Ą�H�>m���һ?P^�y�3?��ȓP��Jui�5�Ĥ��*ߕg�84��yD���eO*O�$��C�D��ȓ>�<�� ^|AJ�.��R8�p�ȓ����c�"B����	�P���ȓ$LpP�@���؁�k"Y���ȓN���`uk��Fy�4�����9�a��Hq:��d�ƞS�� �ȓN��ŨB#�CL\p���Ʋ|�0�ȓ��yec�9+����!�
�xc�=��*��H�c)�:�|���D�Ǯ��ȓO�����@jΰ�A ��DS�d�ȓbX���僕Y7�5	1nO
/����xLM#hK��Q��(�\.�\��E��A�& F�b�da�g�L���ȓ�f�ba�
�gg��T��-� �ȓ;�֠9�.W���܀@K_�^�jU��-"�\�/�;0S�t���% n 5��5t��h��I�_�N�iU�5%�q�ȓJ�YP1m�#Vr�A����3\�ҩ����tcd@�'�Hp9&d�3;;�H�ȓT�����D�R���F-a��\��)���br��;3 i�ŊX,$�Ȇȓ!���d'I�^�d؀�E�IV�ȓl ]��'�<����ɜ�>���P��q��jd����N �D�ȓt0�]+�I�6`;�c��8<�ȓ9z|�R�L�U����iœw�����[(���5`G6k�L�r���g ؉�ȓ4�x՘��3>�Z�S�F��?����t��E��#�Su�A�o�>G�Ե�ȓ"�{�f�*�|
c@Y=1��L$������e��dR�7 )�ȓkI�]5g!x��Y�h�%�d��ȓ;	`�X�Ι)�<���P
o{z���{�t$��V�+n��g
BU�B��`J��W%��U�h	<:(����d�zC$Z�^�zbκp�:�ȓJ�\-p��6E��NI�s����ȓ_LX*��ڊ+odБ#e�2H��X�ȓ<�B�0v�)ՠMAb
2jv-�ȓt����*ӭ5M,0Q��M,Z���ȓ�`�f� �h�ꌫ1��i��@ж%?m�iK�iQ"8*p���$}��������"KU.x��LW����'΄	bJPAB��+�Hą�B�`��T�U&R�d}��E y~hp�ȓ	8����kz \8�d��\���B� W��h��<����?�&��K`�LI�N�r�$ȓe?{���ȓ&Y���)cK��¢5w���[�e�58���3��ƙl*Qr�����'C
l(�M)�C#s�$���S�? ��i��p��`ӺO�L�P�"OR�
a�Ңwȼl�����"O=�ɇ�J>�M�q��j����"O�Hq&h�q�$��r1�`ZS"OB\�c�(5~ܑ��[?e�HPa�"O�X���L/0�a�h�\%��e"O�л�f�_4\�s���u�q�D"O1��,�#a �P��$���1�"Ob��S*��%3ء0OʱP��0ʇ"O0a�G��e��<
�o�S���f"O�A��LG&Dl,���.Ǎ7�2�p�"O��c�d��G@�! "�Ȥ��T�4"O^	x���z�A�BZz�z$"O�ڀ*��L���rD�UI�"O:�BU�	�Z��`�ʔ�&KV�St"O��Ӵ�{��ͩ0)M�(�U�"O�q�.C
EƐa҆�"a{�� "O&Y�cFȂd{���1�J;z���"O�(����')'�	��>O�M��"Or!����� � ��I�+mY40��"O�m�T.ˎWю��u�]�pP�D"O�Ux�%��h ���ϻ5T�M+R"O����ˎu�� j-E�D�T���"O��K���{�j��Ti.I�H��"OxTR3�¹!����v�� *��]Jf"O�1��)�)Ja���%�~�f"O���&m�DoTu���"}O����"O���S�M�'��9�V��"q"OB ��QV.r��Ph�x-�K�"O��vG��n����,,�H�#F"O�	��I�*KT"�2�eL�(�^�2"O�ٺ�˸H?x��E%T�'��8�"O��H7�ݜ6>M+��dV�,�"Od���E�"+�V	b��Z9M��Y��"O4�2ရF�~�Z �ɀZ��A��"O���FNd`�!�՜o�0��"OT��o]7lA�xXv�6O¨�!"O^��e4+봔���T Fl�@�"O(�֌�4?��2ᆀ�hk��8c"O��b�n�:l|�}��L$�\��F"O"L��@l"�Kg��e�"O�!�+�1FTz�kt��/zbT��"O"}�D�&r�Niڣ��3[��	�"O�0*�����*���O(<��"O���g(��.�.�p��3d�ؔk�"O�X��w�YtO�)P5iQ�"O�|ti;[)�ŻA�C�v�,#E"O����a��[X��F�-��	�"O�B��d�`�<莀a�"Oԭ��oD�x�bUXq�X Qz�i�%"On���9s��0�5�H5s��*�"O���G�Ȼo��l��D ;���s"O� !���c�E��E�Q���Sw"O�P���zŀd��"&���"O���A�N(n�4��B�&)u��"O���R�� K�6a��}`�CF"O��d�[pptE�dΊ.6_�X@ "O2�8'��=i��%�N&m���cb"O2�9W���0�Ь!#Y�ҽy#"O&�`���Iq�����:ۤ��"O��C�놓Rɪq8F
�/4�:��"O\Rp��;l;,uiU�	?��s�"OUrM\:<��C�" 	�"OƐ�#&\h�Q�77���"O� ��c +���80��:4"O�l���m�����
�+֤��"O��S�7Ξ�!�h�@�!�"O�"�BF=>Dp������D���"O"@x��C?3�Y�QN��%�0�y�o��s��� ��r$�p2M�'�y��Du���u�ՙx�����CT��yr$���,����BX1�i��y�Ac�"�Y�I�	݄�h�A]��y"��#S|�����Q�\Jŋ�y̕{ʬ!E�Q'~�� �E�yr@�&i�1�CEZ�}+9p%.W��y"H��.y��ʅ�Vq�Z��4�%�yBK��h1@#E{�`\R�g���yRJ^$#v���g��	�	=c�B�9BFʕ�D��Y���2Słe�^B�*f�ਃ#	I� ���Q��>N�4B�Ʉ!�r]���C��#��){�C�/7�cwg�rl0�#i�_h�C�ɝEKj�A�� ��q"�ʇU0�C�ɡ"�J�#�JՔQ�eS5�I�r	|B�ɀ@����p�D�6�� '�� p�pB��:s�1S�'Q�j��p�NN�4"8B�I7�rdIUƒ��%"AO�H_�C�IDyx�����,P�珟;C�C�ɟ.�~�26KC���L0G)M	?̐C�1dE"�@]l���$�$r�bB�ɂW�6�h�f٪R̀���ٌ�yr���Vz*�)��X�z	��ڦ�y�iϨV�ZuJD�0Qt^,c���y�C��2�;s��u#�tJ�_'�y��W�|��裮T�f�̑�#F>�y��@.$����G8c[��"��7�y�̊%S�9�'n,n����*�-�yr�ս8`��+
�b�J�S��yRƬc���`ee�t#�Z��ybI@�tĝ��
E00�.-��oN��yrL���Df (\�a�@���y2@^�w���'<��ɡH¾�y��#by�-P5�Y� 9���4�y���*b�
��YtD���G�BC�	<&cr�#�Q/��#i�{�fB�ɕe�>�i��+z�y#�G �C�IE{��1u�9�t��g̨e�X���U(��ٕ-�R��-� �H�Is�4�W�7D��P�#ML� `���"�8�eN#�E����.��O�P�Y��S�U:�� ΍��=�
�'nK���H s���=H��bȟX��w��؁0Qy���Z�|ie����K�6>.pB�	�E���qa]���	���J�9�N˓5�vM #H�k���9	ÓoJr��Fʪx;�����3_X����+GN�}c�㋲�=b�!��$�&)��[+-J0a�F�(��I�r��㗀GMk�bEˑ=H�<YԋT�2� ᓈW$��`I|z*Y�3���%ڛ<
�(A�h�L�<A
!1��8c"��I��L�'d ��E�f��� �؄8B`�D��'�:Mۗ�'xg�-���W�}.4�3	�'���+��_��V�����2���Y��˟B:�d��eU�[�p8)�"K������/gآ�uDF�;����G�(vp�{�'ʞ�Ԉ`�'Xz��֥V���ڽy[l҂�׈-�j�'� �I�l��a�l���)O=xɑ��D�<8 ޥq����X���G����v"��"O�|�
ق4"�2�y��Ҧ.c�<�4k�y��I�q����Ìq��D	#	�%:\����^	�f�����
SX0Hl�;?:!��ע"rś�*̉a� e"&J�%X�~,(&�iR�;5D�DD(� c�~Fz
�  �3���#��{��N3$�s�'+�52GI��pw �1���un��� ���N� ��g�'ߺ�X�.LO�a~r�;,h� @S�i�^��B�	��O=#6�J;6��q�.�tS��@I?�k���&TS��7a݂<9$1D�@�v���R��|{']#����4-W
�(��ޗ7r�TR4J˸)[ #~��i�*� k��A;3i��C~Q�ȓ1l� �0,
�0Є�
$�Vdq����'C��
E� rh�C�{F{��2�j��pʑ�}BW�_��p>q�M�>�h��DX�b��:7u6�8%��Ґd�B�X���\D���U눼y�ʌ����	[x�D{�+1*�~�8&g��r#1��qaeɨi���y�(E��ȼѧ"O$Q�B��y��)���/ .>%@6�'��6�J%3���ȵ<E�D`C*��0cu
Y!J����`?	^!򤈻3�@�*ܕ>0ī��KZS�k�`9�S����<1f�U�M���*P��h"��T��L3b�����0��#%�t�z`J1@�ІȓH�P���aH��<�C���^�p��K��؇��h�CF�VKz���yk �6j7��"s$[�'����ȓq�މ���ˇ%��!�����<��h꽲�
�6~�yJ0jX=<\`���w6�t2È��Ť͒�CY�hq$u�ȓ36
�#�̩H��dڄ
ev�������c	��L�w��W��d��D?�H:d-C,��)x��P�q����+��ɺ�'��VA*�a@oM;Ģ���H��q酤R Dh�p5����ȓ�����ڳI����El��+J���ȓ��0�F��-D �@���J�l�<ya�O>��i�JÁ
�Д��k�<����Uk&h1�$�+�0!����k�<���_�D͌Mk�؄X���%?T���7�It��řS�A-#	ı 4D���D_%!.�`�&d��1܂�KA!7D�Ta�C�g���P�$./~$�f5D��R�B�(�� i��N2�
����5D�b��2 L��`M>x���$O3D�h`+0eXx9P%�������-D�@���ʠz����ǐEnm�Ԅ,D��i��޺Yr/F��>��L=D�@Y2�7S��H�oE�-_���<D�DhեX�Z5ʩ� ʁ�*��K��:D�� $O�F���D��q���W�,D��3V��Sm�u�kN.L�̉��%+D�쁂�H��	��]����ժ-D����@�F���ڡӆ��B *D�,ې�ޫTT�Se͟�R���,D��#Įώ4��ACKM�>�$l5D��ӈD6�\���a�<9 �N3D�hh�3V2����
?k�8�Z�!�D�5T4ҏZ�Z�<���O�s�!�d�#��PI^()��q��.0�!�$,�tb���g�N�����(Q=!��P�ϸ[��	<5f�ӳ��&9!�ՐC����*%�h�a�QE!�$�K�Irץʛ1(�'�!�^�BB̹�s��!���q���{�!�Ăv2p�u�� 
l"��U.ߒQ�!�d�$P ���Ǭ͞e�@A�'Ch�!�D����vΜ m�L���`΅u�!�DZA���*ߟDäA6�ҥ3�!�DS:?9c���&87<���!	�!�dS�&	���D�F���E�����H�!�Dє,t}0��!E�8\���R<I�!�� ��;b�˭?wiA0�_E6�P��"O
4(ЉW�Ov�4�Q�L41+�"O�Ր��MLE9#Ȟ�jT9a`W)xZD!�`Y��l9�dE=<OBab���5"fH��L؋^H�Ÿ&"Oڜ���%�0�`�h�Y���"O�|�P�
)���K�%}R�|�"Or=�G���J�F�ށ�"kU"OHi�%�Ñ;��Mj��E3��8p"O�a�C N-\NA��C�)�%"Ona!�?<�|$	�엿
��Y��"O����	�i�a�L �~(9@�"O�� K�;l����EG�s����"O,�"��M��Bݘ�5��L�g"O<�3e�[-W���� L�
�h4#�"OE#�cE�:r�;A�үU��JA"O�A��
t��m�7�ϳˤ@K'"O�Q����x�j\"��vY��+5"Ov��e��O��Y+��˘U�u"O�����M"gE�M
@LM�HB@�"O�T;D��&n� TQ3�
2-B����"O@x�@A;9�R�%Ǜ2k8xP!�"Oj���G��x��j�%Τ9��(r�"O���Q K�,%ہC�W�2"O��a�C֙#|�0��L*�"O+�g�<�=�Զ�+$lzC��  p����2~�!Ѕ�[�B� J�Z�Cf`B13H��� �IS`C�ɁDP>���X���v㟵4�B䉦*>�=:sB7s|���s'�a�B�	�0 yA��8WgxU���Q/�B�IX�t���C$�
8�tfPvs"B�	�Az�$�V��C����v? dB䉋fb��T�71�������Y�C䉜nJ��Ё7��XG㜈|�tC�ɥ0�b��b����(�f4p��C��$h&�9u�B�J
 )���I�MK�C�ɻ]K���H�A��ș�뇄nd�C�I73>�}ʠ�J�x�ZLK ,��>:TC䉁#�.蘲"�[v��q�BzgfB�	2+�@ZA�̯n�%�$�<,iLB䉹R7F]� ᪝�g�N.�C�I�yH��Xb��50�x�;Ң� �C�	"�X��A-G�@�X����DW�C�	�x.��FiA�'����W<j��C�	%g�rBe��{1�	�?}O�C�	OE@Hb��`���r�"�C�	6C+���	�L��@���ç{��B�	�<#Ԉ+`g��|��@��땑1�B��+���q��;~�б��Fo��B�	)�NP�S���yṳ0�	��x�B䉯Qj��9%,�4aɆm+�gˮm��C�*�,ak�Y��R��c�Ȃ��C�I�/"���I��&D��F.��]�C�I�e0�Cq뚺O(Q#��F�n�C�I�kf�}ْh	�vLmiE�H?C��2;=�	Z#o��VJlTp'�ō(�B�/J
h���"J�N�R �,F&�C�ɦU��A��� X�8��#�ߠb��C�	&Q5r�"­�9�p���L?e�C�ɬoAj��d!הh����)A��C�I0ς�т�ã�,�JT��	��C�I5Lʀ�׭ԪJX1��^"#6B�	NiÀ�ʕ[J%1GJ��J��C��I��,['&��?��ئh%�rC�)� ��jO
&��j3h�m��H�"O���ւ�2: IG'��e��L9�"O$=��L��v�P��,7b�XC"O(�`�\?���&��_�� �5"O(="E
P�� Jޅb�<ٳ�"O|���NҴ=��H
'�Ź=�k�"Ot� �))wUh�Ȑy�$<CQ"Oи�����L���B
����
"OXp��c\�`��0�N��z��l҃"O:Qx!/:/���RN��`;�x�G"Onx�`�X�t�kq�4o d �"O�5�5�G�j�n��f�\�<�T�w"O��"�,E:Un�tq2J�&K	ri�"O�Q�%�W�J��!i��[<L� u�"Oֈ��.!������%:$4���"OF �
�R�Uѕ-:�$��"OJ��T�0f�#�Thpt"O� X@CQ�~~Xy���\��K"OZ���덢B�^�Q!�)_? �yS"OD`��,�
G.�Y�	c n��B"OXL��I0*���ƀ���i��"O�PJ�E��n�Ջ�+С��I�"O�L�وu���:���!���g"O8,Jg���L���� hȖ ��:G"O���Ϟ(�DqWlA,�F���"O(X1�'T�<؁g-��.Ę�"O�����q(>ay�J:p�\��r"O޽�r/V�*�L��v�J�[0Jt�e"O*THf��f���B���62�az"OЁy��0J��b�ɱb��"O"-H��l�����ą/��8� "O�9�C&܊`� $	��Q"<��q"O�����%;Y	� Q<v&<c�"O)���˅c@=�g`�4\:�L�"O�e�gA�<��XRr
~'�u"On$ �H��ph�ٵ���nF֨z`"O^0��FC�$����7�L9���3�"O�=P�ƍ��Ҩ��m@�~�>LY`"O�$���+'�j�h��{��TYb"Ot��(M�o��E{�;`�:�{�"Of��g*N�f�0�!5��D�0��"Oҵ��%;r)���.|�I�"O0G�֛ d��q&_�Ch���"Ob������Y&�娧%�`���V"O�3�܄�H|3u��Km�X��"Oԩ�r�["!X����-qe���f"O��S���w�x��UۘOVX�1T"O��J/EZ��QP�K1GvJ1��"O����3f�DdI6NǶx�N5�"O��s�Ҭd0�҇l�Yg���"O��X"n�~�DD,��k\,kp"O�,�I�odȲ�H(]pށ�"OT��ai�c��F�m�Ƹ*d�$D���S���n�Ҳ	��*��k!D�XZt � ֌�"��Z�v��t˳+$D�{�)َ{a�A�%%�حr��!D�l0��#fB�)w��4A���2c�1D��削^[�	(vE�>�X�{!�=D�4r��=�\@b6b 7M 4��(D�tI��%E&��J��^����%D��"��9-���+B���j�ܡ�3�&D���,:*L;1�ځD@y��(D��y"O,1J�=����j(��O*D��P�/f9<9Tpʁ�2Cax��)� �T�D���f�d$��i����$�"O�L�C�"��s���7dJ���"O@�H��9*�5*�/��$�3�y��4s� �u��i4�}"�A��y��S�coT1�gȝk����ȃ�yRn:^�ā�VL�pEd� 1���y2d��i]�8�ܻ27 ]��K��y�.�x~����
�.�^��WO#�yi�;c�M�����
~@hb���y⍈�_�֜kJO�nR0�(��yr��!�lס�"RQPR��yr.R)��yh�
�}bt��+�y�o3wE�T����m�4 �A�y��Θ"��M@�Ԅ65���,��yr�Y[��<c��ǎ,����^�y��q��0Gˇ)Wy��80�E��y�V'p�ܫ6���R'. �bH���y"������;�ֈ���[���'O0����t��D	H�	�X�'�`7$P�%N:l��C�d�ț�'��1A�#���J �Nrɘ�a�'T� KQ"A#R�չ��FB

�
�'C�%S�!� �xذ���r���b	�'��Dsn�8b�X\���6W�f�#	�'�LYۖ�:ix��;� S�S���'*\��G!�wi,ջ��6PC(�Z�'�*<�˛�Z��x{��ݞ��0x�'�$�Q��L	E��vOE����R�'/�y�BAX�z���*�@��;�1K�'`x��T,�|qZu�ʿ!BP-[�'%|廅/��0i<�����FTh�'*�%�S&	��+��K��n��'M��i߾<f��e�8;��ܠ�'�&�K�$�e�.�9��Z� �U��'Z�Ũq�ī n�*�d�T���'���QN�w�ĭs��H!Rݑ�'Į��v�Nu7�1��l�H�'!j�Y�	�w�`I�����&gj��'�x�
��D�1�2Y�'˖n���
�'�2�hď�!,>X8rm�EI�#
�'~���f��9^xq��hD1@��
�'A��4���U�3�|ܫ�'�8Iؗiʋ#� ��m��Yt��R�'5f�ȗ�W�'�� 	s&ĘS"�}2�'�p�aqK7i��y�N�7Şp��'/��P���)�\ݡ���0+[���'*>,���[�Bg�x
�I�7w����'(*i��'�;K r�0`�^�.�x�q�'� X�/ްf��qV-4��'��"q�,3.�,�%��-��R�'4�	k�g;)f<y��0#bt�i�'�����$���S��Z�1�'H�����#_�Z#e�@�����'��xtϑ&k#�kRmҌf�5��'X�iä�Drp�YJ̷K7�
�'�Zm�RK�'?N��PQ�H�Ze
	�'~b�YW�X4t�X�b�:BT���'�l�j��K�AGp ����:1
D9
�'��A�W��%Wڐ#%�V�0$V���'OL���
|���ȓDۍ5����'�:I�!�����F�|��\�'��]:LˤH�y�Ӏҟa�0�
�'!: �E�'hf0U8#a
uk(PI
�'c}"�8�8�y�J�rF��	��� .L�!��]A䀠LX�~ό��"OL��peFb%4�ru�7.�ֱI�"OΈ�BFHZ����J�HV��kC"O�,� ⋌'jh��I�r�d�%"O~�A�Ǟ�9(]��һab4���"O�e��!_��s���\m��IW"O�pŦĆW���cq�Y8{[�0��"O>娲�֦0�yf�=절�s"O(��E����2��Է=�9���ݎc��{��(%��P�Ĉ��y2���_��)T@F�NPE��D���y��D�0g�ATA#�Z\��̎�y�O 8\*�XAꙪ"�z�O��y�h�9*"�# ��2`�NԨ ɩ�y�%É`B��2i��qх(��yb.�?i'F���� c�N`i�e�	�y�cԴ������A�XH�1!�BC��yR�Ȧq���C�~��ڣ�F=�yRGE�3sݢѥEJӞ5SA���y��|P�����?�Z�c�'��y�BA�<��Aˀ"��>tZ����M��y�
B��a%kҨj�F=3�L���y��uz�	y�GYS�r�JR�Y��y�B�2d��! �[�Fq����%�y���l�r(���!f2��Qd�?�y�eD�(��E��@.08}�#-Խ�yr�C0/J@�C#N�20�Re@�y���j��l�$�åx�F�*q���yb��,�h�i"s��J%���y*ߤ�4�妀�d"<���̧�yB���oxTD ��=S<�Z�+��y���0S<�CV��x���O@��y����HX`�L�n�n9I왗�yV;N���PbG�;4�������y2��w�|��X�d��E�Teϰ�yR� }?|�2��(f�<��,�y���0Q�6l�$A#3&����y#��v�Řd�(t�[����y2�B3G�Н(�8~�&�����8�y���1��<�S
M� ڢR왪�y"��V�h���b״$1��dZ)�yAR�U"�ȋr�˙o�@�(ˋ=�y)O�DI|����T�p�"\�����y�%��*(r�I��3��2�����y�Ƙ �F�	�ɇ8w֔"��4�yb�=X9�wGE,8�F�h�Ο�y�%�&�A���@��t�0�n8�y�͙�<6�����- ��-�E�%�y��5L����T�V��JU��y�hĸ+ �As�ñx��0���T$�yBdܐH��	.��w9� �w�׃�y���$a`ѱ��ܱӰ�27C!�y�H/]<���D�l>�#W�V�y �l�G��y���x�I���y�.��<d��8\��قuk��yb��l8PÐ� 2��W��y�fF�}��Bé�.����B����y�-Q�<!��`	N�j�q�a��y�ER.a�%��/@6vJe�a ۀ�yR��;L-z|p���3��!5�y���
/޶�ꡡ�W7b��`/��y	ZB ��IIF�1J�	Q�yҬ�Q��A�����v��` )P��y�.��SR���$�ߌp���2$f�:�y
� ���ECmR``�0�>/a��"OZ��,M�T8z�E�%�B�
P"ObE���	v{��x�F��B�yȐ"O6`��/� 4����\@�"O
��t �YgT<(�* �p�Q"OT]bqM[�l����x��0�B"Onٙ�ܢx�P���D�>}��Ő"O�01�O1G��[&��In�I��"O T����1B0)�%�S�X:EC�"O�����8c�C��{*�1�"O��ZG��|�,1)f��5*��j�"Ot:��	g��,@��Q)8��2"O�D�'��ؤљ%�_22���t"O����<}����0m�'yR���"O��@�L_ Um�Bc�5c\v9k�"O� �4�܋f
�E��f�،��"O��F��L��SG�K"0��D��"O������g��%���:G��8��"Ob�PA��N��b/�[ɂTqD"O��􈈵�젃�m]����a"OZ�r��-^�d��b���v��c"O����A�1��{��?�P0u"O�hP��	{�9�@B�W@ޠYU"O>|9f��� i4��#6� :C"O ��Lh��y���#|��� 7"O������NϜ$�D.ޗN�ĥ�V"O�u�4"�6��-��,�)�ƴb�"O��⧎�(��e�f�Zs�@�"O�T�c�#}��(���6���@""OT�"΁ ;�M��jɛ�X�)�"O*@�G��<b'( �S�6�iD"O�Qiu��(x�"���_	(���"O���%���f�,Qd�U��q"OfA��3	F��s�aL� ��8:"Oؐ�K��F9×m͚[ङ�"O�!�%��9uZ�`��iQ��v"O6�� �.1ȁ��*���"O�b��m��Ð&� ?�VD�R"O�1֍Q.��Yh�$C6:
�q+�"O��`V���c�E�6�x���"O��27B��Lг���j��5��"O~X*$j�e�*=�׭��L����"Oeʢ��3c�\���8"�����'�N�� b�KsPt�U�r�D���'�V�ɁHʮ|-t<��Z(5 ����'�0�o :
zdt���E�+���'g*�J�΍%)pڙ*��Ml���'�FXQ�J'8���2V�F�dN�=k
�'�v��.��D�&�K�x� 
�'�`H�B�;XU\QІ�Ov��i�
�'R���Alͷa:n��@b\�g3@;�'�j����Ԣ<G|�	p�ϴ`.P��'Qޝ	`���B�
��GL�_�V���'4<�l�[@ҍ�ck��m����'9(�"�G��:���"�z�(�	�'IZ娷�܁y:PI�Í.(|ʈ� <O ����V���胄�%�}(A"O�����9D:����G>%��zw"O�1z��?B6d8p��b��-�4"O6��@��%rʶX�t�� UvZ�ZD"O��E��2K�B�iR�q��"O|���_�t4�e�6TLE`�'g:0��JO����0����p��',҅��NG��^0�!����Y��� V̱�L�N�f��"c�������"O���¸^*d���J1 �����"OڹK���$m8�bK0x��᪡"O�T� �'�<�aKW=[َ帀"O �kb�̒q%v)Hd�W�쌴Q"O�m�����A��[%	�l��v"O`4��\�LTd� ���ZD�"O��@ִׄ �9P������B�M�<��³&"��W�w� ��¦G�<��U<#|�)4�U�F�@Y@#�YA�<I�d�%0QI���x�$��2J@�<�5Ł�<��qJQ*m��p1��z�<)tM�7��\0��&>\�x���_�<1��+^I��2�F!8K`���e�\�<9���xUʵn�6�^����M�<�׬-�|0�%fX����eJ�<1r'- fb�UnQ̅!�.�^�<�`�ְ+u&��UD� ��t�)�X�<��2E�����ʛ4Q��:�`EK�<9�CH2���h���n�t�rLP�<y���:�Ȧ	$U�x���g�<��C=�:Xy�+\p� f��b�<AqIɻ~|���Η�<�^͐�VW�<��	M�Y~�J��L�\ًF�I�<�u�Y33>�@�G�B�6j~�0�JQ{�<�%i�YO"�ѓ��I>��`_�<a��܆Q��0҂ ��.X�ЄK]�<Ib�Z�X=� �0&K;jG={���\�<J	0��!u�41�0d�d��d�<�5.�5; ѶE��z	�p��A�c�<�Bj�}����-��y�2%"֋�W�<!b.Խ ~�8h���A\����V�<Q�Ȍ ҜP�&$�P�YP��~�<Y7Y2���ba�+}���q��C�<1��ɪ�vm�pDīL��0���}�<qQ��
���£.�9)M�@I�v�<�&�I���)Ce��{6��"�Hr�<��=$����#�m3���Y�<��.�%$�<8���5&\�D�3�U�<I���R X�K�杜V�l�G�O�<aǅ�	#`<���F� �h��JOG�<q��7(�dy��Ww�4q3�d
h�<96�шY�^ ����4Q���#SF�b�<�	[9(��8;�◇Ec����A5D����H��G�$4�'Z�0����0D�d��J����6|'B}C@M.D�<�`i�YN���O�&	1s�*D�\�7�B-���V@��+%�<���%D���"m��e!(���*L2Z0�d+��/D�h"�i���T�,�,ʑ&0D�����Iu9��ÇBіi�s((D��u#�Au2Il�<BA�}5&t�<!�ĉ	 ��3�6��$�D�ȓ���R���@��k�"Ǝx��܆ȓ0����#R��̕�֢��d&��ȓ*L(��C��)C�4e�&Q)�=�ȓ5�Zez#�P(;�"T8��G���p�ȓK5ڕ���ÞBS��B�� gBR��@�3C�V�lJ>�4��eo�X��lV�%`�8O��q���;�͇� �z�� L��9��I��ȓ@��XA��P:J)bQ�\�D�2x��qha2rg�#��R��ǊM��>�n�@�e�7��,���P ��х�S�? R�xu��?0ܐY�i��X ttj"OV�qw�F?u�t<�T�޸y8���"O<ɓ�Ξ�J�25��ņ�'� 7"O4A�#��SDb����(p���$"Oi��D���De'~���ӳ"O��uH�r�����f�%7����"O4@e��2IfX�!Š�>�:=R�"O ���jN?hl�@XC������"OlHb"�]/c�V�3�G�,?��a�"O�8)�͠q r�P�K3.R]1"ODdC��ڠ�=�c�MM��;���O��B`�M��O?�IT��!��[�'��`҇�a^H�*Q�k�`)y#�A>D��8�b�E�`��>����ްh5��)E�
݈q�G���D�i��衦�ظBF1�	L?B��p�ҪOa�c?�؜&ٶ�Q�őF5�U2ԯˏ�b6M[�6���'����?�D�ܴ�]:��J}Q�U�7CA�
��?����	3oX�ip�(ˤ})F�Y$�F�<�5�i��6�!�����m\7(t�i� <W�ƽjTD�!��IZ��Z�4��<Qǫ� _@ce�[�Ȑ�R��Aӄ��q��2a�r�������ޱS��O^��Fx��˨C96�����r���`'���R(�Ls�%]62c&�:ǎD��8X��t5h@/�`�:�zuj%�^!(�ZT��jzha�c�'U6��u�'��7/��Y���	T}H5A��Y��ƯE�**��(�y�&~�H�*�씂-�����G��! �n3�M#-O�d�o�J���<�PE��u���2���4��<��b��B�$�20�ϭ��<��B��$�s�K=E(�,���GޮP� IՂr\�T���R��p�9+'�h������&�bQ�*�=F;X��3Aށ~#le;c U��d����=}䉉t��$#�^�dӄ}�QL�*t&tS0��	�,�`IX��MS����$�O��ʧd{h�āމi���:�`��6P�T��3>̒&��7��RW�
�]�����N���mj�Z˓b#d�T�i���'��ӡ�^EHQ�иo�
!Q�ힹ"�:�'K�?y���?��l9�M�aeԩU�ޥA.�=I<ڱ�'h�d؈႖�P�����n�vFz�F].LW,�yrmL�uj��c
*]T�AK�E
"�@��F(["ym^ͩS��f��"=�w�̟L�	�M�����鉿Ж��d&)� ԰��,X�x�	`�S��?9��2Zz���7,cH�QK�#�ў�&���42[��C
;����K6{Ո�{嵭gG<��435��`�_�ԕ'����O�'#�t�K vʼP���%FI�1���q���r��_�h�9�\=Wh�r����Ͽ�tON noȄ�7�����`�˙񦅰3��@�j�iEF&̤�2�n��7� (��\c�"$lG2RSś�,R	]��5޴C����IП�4�?Q���i���	��z���T'�,� ���',��d%ғD�Dpӆ	k�� ϐ���Fy2&hӘ�l�~��")�ծ;Q<�l�,Ghh��aPZs��'�rOQ[�����'5��'��a�~*�47�Ą9Ў�V�̌��Y�@'"M; �@�9��mx�n�y�\%I&�/7����Q]�'����kӍ�D�Rѫ�:.���8�JvӒ�[ /_Zn�m[�Z')��O��`S�y�>p�B��ă4:~���lP�T�H�$E�;@����O�0J���	�'�����A�	���J	��QÌ�8,O�����";�K����-�P�1�h��Mc%�i��'����O��'��&�O |  ��   4  �  0  %  f*  �5  ?A  {L  �V  �_  Zi  Yr  �x  �~  M�  ��  ӑ  �  `�  ֤  :�  ��  �  !�  d�  ��  ��  (�  ��  ��  ��  ��  ��  < �
 � X �! ,( o. �/  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h����z�"��h���J���y�Α� &�n@y#Ov݃�*J?N�Z��5
	�~Rdd�Dٌ��s�����&@X�fD?C(rap��'>qO�Uc �G7x�ֹ��,�TI�"O���#^4�H��Ǣ�X�#"�$8��?u�	�͈e��i�p,�`�3�tq ��#D���B�]�Tjh@�$�a�)y�,���>)�7#�)1i�$�6&f����$�>D�a+�YQ���ō�yɄ�Q�'lO�� ��FiL�ZP�N7/j��h D�01u�M5*��JA��H7���� ���<!A��&H�u���0�X��<Y����&/F�{W����0���Ɉ ��C���4�$.W*�zM�V�H�2r��>ь����T
��!�� ^��p����"�!������E掄1J��;�`��{���M��H��H�V�:�� �	G���0"O
P0��z�h `g9�6A��$5�S�I� _����#�6b.u�-ŔKR!�D
<k	l�{�#�"k��͑M�s>!�d��:+d�2P�0'�D�[��$!�Z'=N�(fرK� ���O>d��'�X��<�����S	�A0ԫ�U�)�#���E{��iĀ=+�o��hX�0�Ƙ�O�!��Y�x*1;�*�J�=P�X�-���>��B�->�B$�Εgh�CN�q�<2�;6Uڕ�n֜��(��!�w�<1`˄�SO�����w?��&* r�<q�h��*t{Wh<�:��s�<��B�3��A�*ڽM�,l:$��q��&���¡Z.�H�5?j�����6D�TPd��������f]��� d�'D�8��d�8�RT0CꚥY� �'D�� ���_!!��X��q�T��7"O���&jޤ`�249!��'�"xg"O�����DY0V�o�,�14O���D�G�B���=���6 �)Ba|"�|§��)8r���'����"=�y�-� �.%ȓY?$��d8�.թ�yR��\l���F>�6$I�#0�yR�Wx�����$X1,��뗏6�y"��/A��i���T2"��ɢ�ɣ�y�e����1� @�r�Ҋ�y�E�/d��iǔ�f(���,ؘ�yrE#@����m�P�2$R�EÊ�y�L��x���E\�C������4�y��ڊ�XEҒ��6eƭ1��<�yb�ۯ�4�T�Y5*n
(���
�yBI�$qظ�T��)�!��(M#�y�$�+��xJ���?H���J�?��'0���h �D��Q	�F��91
�'	���I�&X��:1)G�C�(�H
�'MB%鳠�q�,�WmP�8���
�'�X9�a䊂D͢b����U��'�xґJ��~�|б�z��3�'Kў"~:Q�K�w� qa�.}�l�Z�<q`%Ǜ-� #� #_�c�L�^�<��C�\� ]�b� +$hʳ��X�<��9U�΁��N;t�Ȍ��T�<�4-�u"%���7��R@��>%�	���<X�%%@�l��}��a��+p�9h6Z���j�@�2ّ��}:�.h�@j��(���Z��\w�<���ȸD�v`�+	�Z�)��J�<�����A����W� ''�Pᡖ�Gq�<�d�@�Uj�I�Oե,�ԭY���q�<A��)$V��'͓C�0pI�l�<	 ��Fj.ĉ�"N`}{�Bb�<���x:�@�:S_����BY�i���Iv�����P��	��
��8_a@�w`�8�yb��0�ޥ�ւ@�b�4�D3�y�j�% [�H�7��7U���q�[:�yr^%\�v�X�P�L+:��K��y�N�d��p�Pb��yF��qn��yR���G�Ё��O+=Na���ՠ�y�F���UI�NА��ʍ�+���$,�S�OG�P��5	O��ґ�ET� ��"O�x�S�N0���)e�P/o[�{�"O��1ekͤU@2A�W���`�.m��"O���J��UZ�p�@D�Q�(@�a"O*m"wD��&x0���_�]�@�@���O����x�vǜ)C�:(�SH�7Z����D"OJ\�І]{�(�5�Θ���R�l8��Ô�U��I��l��� E9D���EA�b	��1VE�q���d�*D�\��� (:�T�1�ϖ#e|��(|O*c�ػ���R�� �IV�S�\k !D���P!��l\N���o��t�+q�4D�0(�o��D�Y`GΧ_� +4@1D�����]5՘�+���5=��l�@�/D�p��׺X��$�%"R�F���u�0D�p)�#ܻ'��,9`�P.>in8`r�_h<��eS�#p��ɗ23^�C1��YX�xGybH��a/t�õ`ͮ.����D��y"H�#Gl򉓠$�8=�e��o����e��ٴ��S�O� ��F�ßV�H��W;!�9�+OTXi����.��=k!M��p��8q�	
�d@�O�1Q���M;�S�? H9�Ԡ��:cT�q��+����Ǘ��l�����L�0m�*(����͆/e�D�3j�8=�B�?�iA��Y^QnX*��]0P b��o�s�'��'fdܲ�,T>zd�C�ݤn�4����'��#LS�av��#���`->���'O2�З*�5":��&H
�BY���*�S�t��<ݬ��
ƺ	��U�
��y"�H
o��Cge��p���#P�߀��IU���O��	�u+F) ���ƥ��v,P�	�':�h:2i�=e��9$ٺx���'%j	��kD�.چ�c�Өwt8��
���~���>;&����ƐA+>j4I��y-�(*|� ��͵#��h��M��yra�d��j�i�*�	G ��y2��B��H��c���j���y"O�	PRTZE
*A�P�����yb�й;��2�A;���s%�=�~��'Y����ϒ���"����"�R������W�Ia<�pa �J%s-08�q�Ҩq�jB䉾S��yQr�K9u�2��N��"0�B�'s�pP��%*$��VCP�#PB�ɿ;V}B������׈Q'F�C��6VA˦ ��L{D�*Nj\C��'���
P��/I����%N�iJPC�	$	��Ź�"��6E24/͕M5�C䉿=����T�g�\T�@2�TC䉱l~���=/\@���HB�J B�I<\�^yZri�	_4���-�9+1C�ɘrf�aŋ��x��!O�EC�"$)�-�3+Ȳw!�Ā��I^WC䉨q�|�CO߷VrTX �O��=B�	-t3,×��+E�h��	=;N�C�I>��xŨ�Y�f���	�9�|C�ae����J4I�2k�iL�9x\C��"[6ʵP ǚ.D���_�B��C�(&pPԥ©�&I�uޙ_�B�I�U���H���T8噢 W�
߲B�	�x��i"�� 9xbd�P�T�D��B�	 @��"����ZI ���&ƸB�Im_3�!�78p��3(@�^�\B�ɢl6�!Y1,�&"'`��^+Q�B�3z	�3Ev\���j
$#FC��*pq �h��z�A3w�ZH�FC�I�zR�����+�81䃓`�>C�ɖD�����Ǆ�rAk�
CkC�I!�< c`�*ZYA�a���yh�B��@� ��P�ٻW�B}3R-K5�TB�I� �.=`����6A�&N7rBB�	z�)Pŉ�P��{�fZB䉪d8�0�b����adj\#9`�C�I�tp�pT�O�/����#@,J*�C�I�K���&FBxĘ;�D=�B�ɁC&��ʄ9v����ϗI�C�	8��É��s�ݓ�N�<�C�I3O�b��c��.d� ͕ �NC�	���E�ʡv�x �W=Y54C�I�|�B�r�4���J>1�C�ɞ?�R�J@(ה�<r�D�G�:C䉿^��͡7"Z<ߺ����|�B��B\�{�M�	%�,aW��8q�4C�I<(e�Y�"���sY����Y[�RC䉉o������w��Ÿ�B�;�C䉈["��ԧZ:5$�	�5��9K��B�	0{�V`1ǍI;[�҅Z�NF�n��B�)� d��5��"W4��q�N�j�!�"O���?(��)��"]{p�0"OF��#D(8�%33G6mL � "O��DHGq0�� ALQ\���"OP����\8b����7��hR`1��'�'��'���'�2�'Jb�'�)����2����4A^���R��'��'B�'�R�'��'���'��`,W�i��+P��pP���?���?����?���?���?I��?I��7W~(�hģ�49�N��Ї���?y���?����?����?���?Y���?9'j {��l���ͤ0�8i�!Eܐ�?���?���?���?9��?1���?��#\1;è�t��'�8:���?1��?����?����?)��?q��m� ����K��a���۸5�
(c���?q��?���?����?I���?q��`���X���Xhv�* �*h�|+���?���?����?���?����?���<�2��!�[@�])��'*ò Z���?Y��?���?!��?���?	��7�@�r0�����J� �<������?���?���?����?����?������!�"T>+��/�q���?���?Q��?)��?����?��,��ڵO' VX=�� �3a�0`��?����?9���?	��?��?Q�U�QسC�&����r�6T~<����?)��?i���?	��?Qg�ih��'ƾ����(7­K����O���ȇϻ<���󙟬c�4 cx᫢)\�U[��jtK�$%�@�2�[~~�!r�n��s�@��"\�"Iv�% �T%���Q#�)��៬`bf�ɦ��'��iH�?y���ix3H\�q��si^�s��a�D�Oʓ�h��� ��ߔFpz�X3遢pe\ ��Hܦ��..�I\��^%��w�"�iC�B��S�X�<����'��;O��Ş"bm�޴�y�dǍ2.ٚ�@^�a!�DSG�^��y�1O���	4u�ў�ӟp{�"]"d���G�F���	w� �'5�'� 7�܌�1OZ��*B�`89�K��npr�`�,������O����\�'$�0��P.,��̱ŏؼs
��O��䀐Id�x�����?qѣ�O`�R�k�wd&���O�OO��"�<�,O
��s��)be�x(��@$s�$!U��<A��iR���OmZb��|�УP�c�\I�&i�e�����<9��?�����Rٴ��dz>-��'B� 8�lH�a`�h�ūW�>�1b/"���<ͧ�?��?9��?!��B�J�lj��@.#�\X�����$[��)���ҟx�	ʟ�'?q��/^N�x�q톋f
H=�&����ЬO����OD�O1��<�FGO�<9�88�����~���a�H�6�8?��By�l�I_�	}y�T�h�<˲	�S��t;�ǘ#$1���ן�iyr)fӬ�h�D�O�(��E��YZT�h	9�Ȓ%��O�n�K�+�����	ޟl�S�ƺK�4{�)�7"�!ȅ�� !��`o�Y~� *~O���t�'��$@ݝ/���R-��3� ��<����?����?����?9����޸6����'��e��XBǫ[����'.�le����1�R�$�Ħ'����^�`��p��rP����_R�����i>�;�Cަ1�'@.��� 15���A��R� }��HF�E+ �I���'.�i>E���\��(l��A�(ą3a��O,|I�(�I���'�`7MO�L�����O���|Z���)W�P�# ����&Af~rɮ>����?1M>�O�h@�0�IC~iXC�Rc$!pd�pF�qf����4��������O�a+f��+fL��!׊�!�" O�AnZ���`����8L�4A�0&�4z*� g�Kgy�lfӶ�p��Oz�䛶d�\�i6��z~T�1�K�jJ����O��Ad�gӎ�|"t*�?ɗ'˰�X$w�tLأAlO
�ə''��Ɵ�����8�������Y���&C����X�'&Vo�� N.6��#D�d�O��.�9O+��y'ɂ5���9$��2& �K5�@<e2��'�ɧ�O��F�i6�dN�*���*�iP?%j��&)ˬ��$ήH�����o���O��|��\xI�E@�f�^  P)�=�:����?Q���?�*O8Ll�0{��ןL�	#	Z���n�I����N ;�0��?� U�0����,'�\ك
͌a� A)�L�]�<P*3�9?�Rl��F,���P&�L�'@-��d��?9v'��Z���SccE=��툰a��?����?!��?y��9�|EّLׯ>K��+��Ī$,��P�j�O�oY2���'-�6�1�i޵J �D�7�q{bALx �d��eq�$�	ߟl�	e��oZv~ZwZ�4���OHJ�F�Q�J�B)F�N.?� ddPs��Ly��'��'R�'�ҍ <P��Ag�a�>5�m�-q��	��M�����?���?�K~��IS|��.������I^< ��\�����O���(��� ���%*_�c���`��0<��9�M�\^���a(h�{��'���'���'�$�+2�څP�<�S�Mw�|j��'r�'9�����P�4x�4]������U���H�OC?D�@)�kҡ-�X5R�ݛ����~}R�'���'�DM���]#+Mp��!./T��
�"�o�����X�/L�Q��t����� n$"e"��I�z*Y޼u:O��d�O��$�O(���O\�?Y�P�n��iC� ?�:���.uyb�'=l6-��V��I�O�mM�Il2��o�3Քa�$��
�''��O��4�F���~�l�.xd��Mq"�%�!�6#��;�("!���^�����4�����O2�D�e���a�M�`�\%:�m\�T�6�$�O�ʓk9�6-��Y��I韔�O���2`ܷ(���c	3�2�Oj��'�R��?Yy�`�h��`��<y��H�֕'ʘ"�D\ ��얧����ӟ�#�|�T�];w�ת ����n�!�xB�e�$=��JK6�Έq��A�Dƴe�Mٔ�����O"�n�u����ڟp� ȏ')b�8r��o�4�����p���l@�o�Y~Zwsb�(�O�4ѕ'
��DL�r����`g�P����'g��ݟ��	ϟ(���h��o��"�2,�R�RS���8�B�:�6�݁@+��d�O@�$�9O~Qnz����ȉX,�� DTzb��� ݟ���y�)�7v��l��<�e"8YT��(DlEh2e��<ِE�/{���	A�	}yR�'���7Yv����\T�0��7��B.b�'uR�'�剘�M��L��?����?!Gd�$��y@KK�J�μ��o����'���?y����	0�,1�[ 	.r�aw���	��a�'\���ư?SvE#������l#3�'X�p��R܌�aTCI�I#����'�b�'��'%�>�"p���$���栮=��\pb�'�v7M�<HrT���O2oZf�Ӽ��o�5^�(�!d�KiDФ�)��<���?��.蘁�4���ih"��,�\Ayd��~H@��+.b�82�5�ġ<ͧ�?���?���?)��	E$�1QC�� a&���%I���DBߦ���^Wy��'"�OXrB�j��aUg�W{Z�*w��G����?�����Şw촤W��z �P���$
�a�Q%�P���'4��v�
ߟ|!B�|RR�� eJ�u�脻T��z�hJ��Ɵ0�	���I��yy¤w�zTz�K�Ov9���
�%�\�&GP�@�
�O��m�y�|\�	П ��s���
�D8� �*G�|�"�떫�tl�l~"��[��}� 'Y�O�G+H�v�����&�,!�ă�y��'<��'p��'��i9Oؙ����_/E0v$���^�$�O���W֦�Yb��Jyr�h�t�O��x�&E�g�ġ�ϗSfr��k8��O��4���4�r���Ӻ�ݴI�)��Qr���"rɋ4�'��%�̗'}�'�2�'����!U%u�;���� d�']�U�P��49K ����?!���I߮)`Ȼ��4( �A;2o�*x������d�Ot�d!��?9��+	*0�fC�O�1P�d
�bփ~���h#o����$�M|?!M>a�
΄&ޠ���s�:T(b�?�?a���?���?�|�/O�o Q�踋�`\�T͠�@vIߜG��2������-�MËB�>�R�~!�g"@ZR�� �D�8^��#��?����M��O�������O?�(0g[��(��A2��"�}�<�'1r�'��'oB�'�� UlM��N�5y/&آ��XT�Q@ش�p���?�����<Yq��ywV�F�����	�:}b�+`�Z�w���'�ɧ�OU�]���i��5�x� m�&~�p8'�5:����%�r`���t��O~ʓ�?���O�R�&�K�<��l�!I`+���?��?Q,O�ilڒ
�y�I�$��;H���uS-dt�5�W3Q��?T���I��d'��I�`D�L��S�D�hO�c�0?y��g���6�^�'l~�����?��J0��LäA�>!Ɣ�G�c�<��II-x@H�fýf���!�A��?QU�iqh0���'G�{�L��$~�!A��-�>z/��������ϟ����N��u7(�;{(����i^ʉ�$��Bɘf�Fh�$�Д'<��'a��'�'�Z1[u��1W�l1���(|�6Y�<cڴ+OF@���?�����?�6�����9�.N����S�_	 �������k�)�S�l�j�H�h�Tm�6��/X�m+ BD�t�n�a_,cF��O��I>y.Ox��&@ܾp�N�B�Aɏk��8+�`�O���O����O�i�<Is�i�c��'v8�Pӫo-�u;��@� �!�'�|7�%�I����O2���O�Y�mTDC Lr欚.dj���OV��7�7?yb��?vD��R�S��}�$�ӳ2G�1	c�=;�z��0q�8�	H�������⟤��C�V z�.yf���}��da�U��?����?1��i��I"$W�pٴ��|�$���ʔ�B�Pp#D���U�O>Q���?ͧSb<�ݴ����6��`r � ��$C�$fF�ÁoL�?Q �-�D�<ͧ�?i���?�Q)��K�|����7���V`ո�?A���]ӦU3�f��p�	ٟL�O�|,뒯gpT�*#�\0�����O�1�'���'�ɧ��ɓ�X�o�7�RI�C�u�<i��	�x˚6*?ͧ"���	j��,G	8�sd�;\���8�	Kp��������ҟp�i>���#d��'�7N�ڰzu�̔=���kbň*8��7�`q5�'�R�j�f�O�Q}2�'d����{qhqpb�:!c*=���'�,=��;O���^������vBV�S�? �1���A�D�}a��ɋG
�<�37Oʓ�?���?Q���?Y���IL�5I����pŢhi�O#&Ӭ�n��`\�I՟���Y�s��R���#V��NH�-�0��4��'E�3�?����ŞVf�5��4�y"�5L無�"�[*?�@|���ybN�1,��������?�Bbe
�6}ؔ O�Pfn8��O"O @mڑc^�t�I����9[�4@WIP>T�=�d�@�L���?��[���I�4'��`�6	}��c�y��ȘA&!?!�Lۭ$�0 5�M���'/�>��L=�?�������Zr%��bfT��-ܽ�?���?��?�����O�a&���6���#��L#S��<ɰ#�O�n)%���Iߟ�4���y�`H?I�$ç �7˨�����y��'���'_�in�	2*���I�ן$=�%K]I��c�"� ���+�b;��<���?���?���?�"m݊ �����
i+i�d�G�����y��n䟈��̟�'?��I�g}���V'�� �.��6�W,v�*8J�O����Or�O1���9p�@ (r��8�FÓi (���6�1?�`���{�L~rʄ�>2�DXB`�<u"R�BB��?���?���?ͧ���ڦ10������Z�*|�<ZA�]�A�V�x3�}���޴��'����?!���?qu���{S�)��J3 ��P���ޟ8=�ez�4��dҲZt���Oj�O�gN�'Z����pf
L�DyĮ	��y�'�v1��Ӧ+��q���":6��8R�'�r�'a�7�*6F�S��MkK>��$]9$ z<��d\;~={����?y��|�&����M��O�nV9v��)�w���G�1hй�׉�O$�AK>�/O����Oh���O����rm$�bt��^Pڶ!�O��d�<���i����'!2�'&��|�V�sE�˜7���9�FU�(D�pI�I�l�?�OP�šaJ�*�֬"�hІH.�����F���i�+|��i>1��'��5&����!��f��2�/�!�
�@C[�|�	�h����b>��'��6mӠ͉^un����mٜ.� ;�
�4�?���5��F��v}r�'tʁ���ǜa[r��ee��9{(�KE_���A�Φ=�']~eW�?��3S��8�a]	'b�#ÇS*���&,~�ܕ'pB�'�'�r�'��Ӵɪ
 
L�y\hh�S'^2�K�4�ƅY���?�����O47=�Dґ�Q�	�dy��a�,�$)���O^��6��	�4��6~���.˅\��zd�SV��p���b�T�� -G��OMg�ly�O(�Ȑ�ϖ(q�Z�GW� f4x�2�'���'\�ɹ�M�FC���?����?���>fN��=��������'k���?�����>U.�I��PԲhr0dԜxH��'��%�4*m����Pٟ����'�&A��.ߚYZ� y$m�{�A���'�2�'�"�'��>�I��^��� Q�hl>5�D́�
���I��M+ㅧ�?�����4����(j����)ףdb��4O��D�Oz�$	\�7�??��(ӁR���) t���̊$="1�scD��<%IO>�+O���O��D�O8���Of�C��]V���C�)	'�2H+b��<iw�i9�=��'�2�'��O����8�>T�E/��J<h�����Kb��?����S�'��Ly��M!�n�I%$$a4���R��M+�P�$	�� .��d(���<�B�ZP�SI:p'l��[��?����?����?�'����ۦŚ5���䐔h\�&�,5��i�h�d���{��[�4��'m���?����?	��M�U���	f|����j7
p� �i�I0<��˰�OGq���N$v(%�f��+K(��� �Q�}����O��d�O��d�O��S�']3���qmT�fĔP���������?I�.����0����'��6�+��%$G���W��#d1qaAЂ> �O��D�O�3YE�7�;?iD	��2HN��BN�/?��٠FѧA.ě�d��X$�ĕ'��'72�'(� ���
�
�3I�}�4H�'��_� 3�4JU��k���?����I�6L6����θ^.��g��9aq�I�����O��$3��?�cD!d��x`B�}���!"��0|@ЛBꂛ����D.��X`��|�!]��uk4��q#����阝$P��'yb�'��O
��SL�j剋�M��MP�h�i�d˻_�|�R��
o,d! ��?�ѼiZ�'�B˻>���r�(���&H�D��o�8DI�)���?1��7�M��'�2�[,M��1���q��vU��a��Ҳvb�����61�E���|�]��UT�v�C�a_	["� 6�׸b$2 ��8	��P����4f��+$i�j|�a��~�Vh0�X|��P87���l�����È^:�&�D�zXh��˼��H!��y.$�Fx#��q�ĆB=J�8��A�n8d���é/�\	��L���A�IN=M��Z2�˒~t� aD)B��s�ƣ;?��I�P��P�DJK7Y�B��uE�.Ci ��%�`���E�b? �;�krӎ���O*�����@�'��y�ѓ$���~4 �ǰhV�9�4W�����䓵�OE�D�/�źB��%.��!��SWl7M�O��$�Ottjb�Sm}R^���	o?�a��ƈ�v�� К0�
��'�����|��'��'���Jrk�&kK
5���JW�:�h��h�d�d�9.5v˓�?���?�L>��x�x�B�M�_�썂ԥӞ����'?|ٚW�|��'��'��	�� �h����3ΈR��D%i�h���&~#��kyb�'��'�r�'aV���)j�&\%�]#!vrȖ�X�L�'F��'t�Z���[������+0{t	�Ȉ� � ��Q�_=�M[-Of�$3�d�Od�dN�4���ɇF�6H��!�; �I��A�L��?���?Q(O��pp�{���'�6d#p�_	2ؼ�� ���PZ2\qc����d?���O����*<*l��A)K�g���.GlR�RaԜA���'�U��.����O��$�he�FOZ�>NX�Fm�bdB��&b�K�ԟ��ə2M�?A�O�����!J�ٱ��n�L(�ݴ��$A=-Ʀ���۟��I�?�OkL7x��yjF�4U��b��Y�`���'�"fA�W��OR�>�1�)өf� ��Շ�	�.������ǌ��9�I����	�?Q�O�˓ևB�O����J\�V�d�i!����M�E"��?9I>Q����'>�*�Oқ	�T�S'��I���(�,~Ӷ���O����2��'��埀��w�~iPSȈ�Z��BΎ#)���>yϚ����?i��?�I�wh0
��D��Mږ��/l���'���m1�4�0���O��w����n���S(Bs�6�<�����O����O^�7�P��I1~ݮ@��Ƈ�=�T5�4�A[x�'R�'��_���	uB��o������8{��������Iu����	uy��_�����^�A�!C��L(.��`������D�O��d#�d�<�'�?�7"zq:)ze��)F:&T��aP����럈��Ο�'�ܵ1E&'�^?:�X;я����@���6t�n���|$�(���t�'��ZJT��9[��9�f���aJmn�ݟH�'�ҭڰ$���L�I�?�X�8q�%ʈ~�p�1��r*O��D�<Y3f�Q��uG�Ѝ[�B�*�).E�(<S!�ɗ��$�O��WA�O����OZ�����ӺC�Ǽo��A���9���#�Hߦ���uyRǚ��O�O�x�R��1X���v�ܨ� �+ڴh��|���?����?I�'��?�R���O�=*CI��v����\�����5��b>��	O��P�JV�F�l�%���$�H6��O��$�O������I�i>���M?��I�9��Лt�B��(Bg�YȦ���S򉸐������w?�K�&,����+�$�p#F}��X�t���xy��d<%��.2Ad�	�jW�-^�$�4��A*�����'|bA�T��pW�yu�Hw�[�a�AZgUay"�'��d�O��ɄI��4�uA_� �!ܩV�7M�.D��ğ`�	ԟX�'�cUeq>ٰ���'�M3p@P7M?�����>!��?������O��'�?��.�F���Z2M�L�33��f��������ޟ0�'s%B&'�~"�.��L�!��p���C'Ğ�㔹ia"_���I矀��p��N�ܴ˒��U7Ԉa�:n�t�n�����Zy�$e!z꧱?�����^wZq�wO��]T��0�5=�Z��'��'�r�]�y�|�ҟ�x 6�U�1��Usc�Лq��`�d�i��	�|����4�?q��?���f��i��0oϱq�ڜ�ՋRj�*h)Љu���D�O"̫�>O*��O������5�� 0�l-%���O�r����� 0�7��O<���Od�	Yr}bQ�Lѥn��P~��kv&���x����<�M��eg~�U�4�Z�9��08�����<;�!({f�:�i�r�'F⭊_�������O��	p3\�S1��D���R��&5$6M�O��d8��S�$�'��ҟ�@����<*dl4�1�وf� 騴�i��g�ʠ����O���?�1t�t�9%c��j�F)	�X78� �'�2ٛ�'���'2�'��s���qھ�
�:��: K
�A!$�M��ЩO�˓�?�(O���O���˞"��7ً(.Ȩa"� ����7�~���	̟��	��0��JyB�
>=
��S$O�\��e��EZd��Av!�7;<!�����On���O�� V<O���
��Vʚ�f�O%�|Cv v}B�'B2�'��I�N\R����$��&��D�PiZ�"i��(���&�n�ş��'h"�'������Y� �(X�����U�ܰ���v�����Opʓ㸄�5U?��I���S(��H��,[���JU�T5fd��Oh���O����3W�$&�D�?��'�DS�7�ރU8�� ��m���	���b״i���'R��O��Ӻ�EJ�k���Eㇴ&Z�  )�ܦ-��۟�@$�a�p����'�!4D�QGL�%%��z�*Č'�6�E/�$DnZџ��I��T��:��d�<�!Jӗ�܍�s�R&3IF�:�!C�v@�l^1�O4�?Q��	VThs��G���xACO�v�j!��4�?��?i�K-88�	jy��'c�d�,0D8���JN��@�5���'�剔&(�)j��?i�,0,(x�$ër�l3��̻Qh���i���m����O��?�17��)H�*�`��5�4e��A^��'����'���'�R�'��]��b,��*�9[5L��7�d������ ,��O�˓�?�,O��$�O��dE�ML�-� �,%�T���6��A t0O����Ol���O��ľ<9��F/��;K6����䉡jR�ɦ�i]��Y����ry��'R�'wY:�'�l�5��C������b|C�D�>A��?���$��9�OB"�)� v�ZC�&2f0�Bc�,�5��i
rW�d�I��,��7e�b��~�l�t!��kǏB��m[��+�M[��?A*O�	'O�z�4�'�b�O
��R�ɛ�c��:%�?:ԓ���>Q��?��|<����$�?����	[�l��(��P�r�!+qӰ�~&����i��'ZB�O�r�Ӻo�����;q����W�}�	��DQW-��$���}�1͏�z0m����V�ڀ&Hܦ=(�*F�M+���?���J�Y���'Fd����ү[�t��e&�I�1�l�2��<OȒO:�?]�ɓK�\��h��E��E
��L���ߴ�?q��?Q�LJ5���Yy��'�$��|����Q�i醹�wH�?����|��Ҁ�yʟ����Oz�Ӏ5���i7���D����+E&s�6M�O�m؁hOy}�W�(�	Zy���5�@әk��ݙ��ڱl*��5�P��Ms�H����?����?����?y*O��h��I�Q�()�.�2-,�ղ��0�l9�'��ן��'���'_"ǎ��(�Vz#�ic5��[�6i��'(�'�b�'��R�l�7�V���E�o��0 Ȇj��ٺ��<�MK+OF���<A���?�"���7�F�����7�J� �m�NVT[��i�b�' 2�'��ɉ_|j�뮟���_n��Sc�Մ_��9�amV8t���lZ��'�R�'��i��yb[>7���q1����	�s��Y�'�վ���'�b^��T������O������h��T3b����@T�
v�����Yp}"�'�B�'�x����Ĺ?e*reE|�ޑ{ �X9�d��(vӬ�!:����i���'���O�d�Ӻ��i�9%N%*eo#e�"(�w�T馩����qq�0?Y/O �>�8u*īp��IC�ϧ5���6�o���8
����'"�'��Į>�ɨ� �ّ�.Fhҳ��[�2�{�4'�d(Γ�䓽�O�e�5f�2="��@��� 1��|p�oӜ�d�O��ͳ-O$�%���I��L��B�ҫH�zUyw��`�&�mI�I�t�I�K|���?��>H`�E�!:�t�p�<)n�f�'*�;�.'��ҟ�'��ث\F��zF��%@$�XC�$X�=�DEb����d�O��d(���dDE�,Ν9.B��L��x��9RF�t��?YJ>����?��놧K�epc�JL�j���Gxt�����$�O����O��^���P0�D���&��TH���x�U�!D�~}��'��|��'��a�$�­�b���&�9M4!Q�	L3)[�듷?i���?�*OD���Tf�Ӈ�=��-����ȱ�B�$��P��4�?�/Ox���O^�$��]W��'}rD�4:�d��
�oN(	��U�M����?	(O���0B�]���,��0:L�ks��D)X��2b��8�J<Y���?y��D�<�I>y�O �$�$^-�]��l]!Y����4��$�)O��n������O��)�l~r�^6&�LxV!Q9f� h!5�O��M���?�Q��<iH>!��ԃ�D��06"ɦt޲XB	_��M��rś��'B�'����8�ɺ�v�����!�@F��ew�X�4Z��܁��	�O�q2����:E�Ӥ������4�ަ��I��T�ɑd¤�ۋ}b�'��d�e3<u��F۞1��5z���^��|���e��T�'n��'�f��g�	�?X��t*���<��jvӄ�]#\���%��I�8%�֘"��i���<.���
�.��V��,=XM>)��?�����DL����/�m�����=���2I�}�	�����n�I����ɓ,���zA��[0p`���y��M�Ǩ�ퟔ�'k��'�BV���E����$�ޓi�Y3"D��iU���g��>����Ov�=�)Ot�Dδ\_p�[���#Iȵ��T+�8��'�"�'��Q�x24	�ħ\��\�A��a��%K�o2�����iў��'5�~��"��B	�a�dD	;e�P��.�̦M�	��,�Iܟ�u��j��T���S.Q=8��#�������z���H<!����ȡ>0�֝�rzxd�PX8.��I��FO�1TN6m�<y��@�^y���~����*���h��\)l0���C���!j'N$��b{�㟨�3�.2�ڼ�&f9 ����+�	�����W���'^�'E�t�'_�U>�(�G����!zT"��Lu���IБ���m>�b>���hF��Č%&��$�󤗅wȨ�4�?���?q!)�eV�'���'��$( _���砓0�������R`�O�-�T��O����O|�dE�k��8a��#/��wWԦ��I�~�a�}�'sɧ5vL�F�̤�5�=NDa�'�A��� �i1O���O��$�O��đ���H�֯N�~5���7O��h�I�<����?�����?��'L`��$��`1��츳�4}�''r�'�"W��p�玁����ְ��]�u��\��TN_�M����?����?���'f��R�Pԁ�d�>�l����I�|��ʟ��	蟐�V��A�4�'� �S�ź|�r��C��zD��bӈ��-�d�O��;��H'����V8�$�
�'��#et���b����O����O^z4h�|����?���\��-�'���e��1�d�u@����xb�'�剂^�#<�;mT��8�22_�M�܌���o�syB��h-`6M�O��d�O����L}Z� �%�#d��K��E�� Z�E���x��'�ў(�Oj�(�FjX���cm�|8��P�i��1�p�'+��'��O��	~��� m�*t�Ǭ�gF�Iz`)_�0�:r�Dx������|o����
~��i���K%)�kIH8�iqq�4S�a}BaۛpC|4k$�Y��\u�ʘ6�p?I��̅oj�	���>e���PG�(�>Di��'wh��3���!�iCiD�l�F�0y�f`��B�<�n䩕��1[0T��c�<�(1"AJ\�njr�0�@�#*�0�r(���
g�P9~h�ss��#�F�j�HY�zB"� ���Mw"$
��6.��1�� 
3��! PN[某�I���	�i�!�	����'�T��5G��s��eqF�I�%���J�'�&c�~a��%PE��*��C7��X��,^���+# �<^~���a"��3���h�L�;\�q��'�+
@V���)ڶ�D��P�"�'
>x!+��q�&���#�B�����	N�'�J�Y�K����҉e��9��' ��2�I��e҉��`D�o�ļ��'eZ���d�?IgȰnZƟ���~�dMP�J��9�aU�^����JIl�&q�t�'���'� ���_�s�|���.Yj�T>�11LN��\��U�x�	V'-�A Pb
@�+&.������ħ.\IS��� E�uM�- �YEy�?�����'�?Q�h�A�X�k�n�!}��Ppb��?����9O�t�.��ބ9��͞*�DҦ�'�O���`�}x<����מ-t:�7OX����h}2�'c哏M�Ұ�Iן��I�'��!U��9���2C��������R(f��p��_6 3�S����'�*}I�dZz�^���$�=(���ɡ��#xM�,ɕ{- h�a��O?�DV�O�l�`�
�"Ԫ��ԃ��Md�����O���,?%?Y%�)���(z0�f��6[j<���=D����&-��`4�BF,`X3�:s����'F�J�h�o�:MA^� ��	2_�0���?�A/��c����?i��?	������O�B@��|��@��
�O�رbe�O>\�5�w?����HXs8���eC�t<"�k�ԯt,%x'����R�8@��=�M��p<Q�Āt��`ʡ�&+�  #��`?�w�ǟ��	l�'��I�D�����79���UF�=��B��'{�\�:g��
'>�|p�b�1��I���?͔���A��6GXw�L��M0Ƙ��!P�x�P���Op�d�O"IKp.�O>�{>ٸ�_�3Ǯ,���q��*6���K��^DR9�R&�d�6��1T�X59ԮǰP �D��a��8x��S��t�a{bg��?���Z&@��&���SQ����9���0�Y$¼����%oq�1�ւj�܆ȓDHxy�7/S�86U� 	�8ւdΓ �IBy���m 6M�O@�$�|�dbD�
�<`0K�7h[h���7��(���?���X
�̢�Lߐ%}ɧ�i���с�Z�xF�(A!�<?�Q����+���D�D�C:9<n�(�-8�� %ʻ�(O���%�'XR�'bU>!���:J�(��
L�L26��џ��?E��'�N�֌����]���C��
� ˉ'�<S����g�:�A�ǰ' �9��')Hș���>q����	�F(\�D�O,�j/ΡڢI��0|���e$�2D`!ص�ѱ��
��W6kf�YP�|Z���>���A:.l��
S�DD\���Ġ+�\Aؐ�F' ��E V�p��?�R�J����y�y�Z�X'	�+r��I����z�r4�!ǾU��["�!e����`��x7g��l1��GN��DGx2F"�S���;XxZ��S�6&��r� 
�q��'GN����SW��'r�'���ß���dčچ+&=��P��*Q�}��(Ly���d��>Oh���
ٚk��	1N ͠t��,.����땍)��D��ڟў��٘N�@��ճP몽j�챟d�B�O���%�d�O����<��!Sb�a�tj�
Fda�'��J�<9����
�����0k�áFD	Y��']ɧ�D�'o�I�Jhx��4N��@Ԅ̀1O�q��ݳIJ�����?���?�[�?Q�����.+TrrM�d
�n%�\��۔3#VA�b-|hH�$ǈXXH��D��k����D54Rd8�(�I�I����X;�D �ɝ9�$��I&p�����O���9Ķ�Y�����F�(E�2���OV��0�)�C�)ɰ�˥�O�C>� p��I�<i�$(R���0�_7qH�[�O��<٢T���',j�C�ei�2��O0�'x2|�� D}�(I��J=N��P@�I޷�?���?a�ʁ���T>��#CR2DF�@�r,-1����  �`o�0����Z=n���G��o����S�Q��3���OV��O���|b��4lE���\��f�N8�?����9O��kX�H��d�!�R�	�~��'h�O� z�� -rz�T3�%܎#)��g<ONI�D'����	ܟ(�O������'*��'�,Că� Ҷ1"Cҩ��$��*uN�	���W�-s"��O��t�矐�@�>���!c�M�0�PA��8�|������ه.��?E��{l�� ���e�gd�|z�צ���?����?������G��1 !�89�h�"4ϋ��yR�'��}�˸M��H�� ��D��W֑ �"<���U�T����=:��Ќ_>�2�P/+�r�'��	Qt�/-���'���'?�'�?���\�,�Z�b��u�~ ,������'��y�R�˟B�> ��@�SF{�
��8��̦'NM:�*�8/�`����28lzC'ج�p8���hO`X�M��B��Ey�R�fɼͻ-�O�l"�o�Ot���O�Y���IVy�hX#u ��cŚz�r$�Jڏ�y����Z�u�C�4A���YF#=Y/���O���{s�yJD�ؓm�nu�F��3:�!�d�
}d� R�_�[��K��_c�!�d�"D��a�d����^�p��"O$����ˢJL�d�Ǯ�w����"O@P���R�vL�@�l	�.]v��`"O2E�Kː	�l�H�l݌VX���"O��bg�|%�Г�ň�[�0xE"O\��-�$I�z���t�� YF"O�8�w��(-:6�рf[��9J�"O��x�� {���$@I2o��M�B"O�|���}�~�S#
�
D�Ҥ"O��%$ܓ�d��-7�=�"O�y �Jwt	v�U�^�F!��"O�	�W�$����I�21p�"O؀ag��;>N5��"P�V�T�K�"O~,
��VjN���QD����H�"OFlzD�l��0r�	[-n9��"O���#�^=I^��;��T}�@b"O��6�G�>0�T�N�b�����"OH����F̾U"e���lul͈"O�u��$�UR��VI{X�UcB"O�Q�� �(�}�@�ZD�zL�6"O��+Շ@*�.��6g�#sq�je"O\MibΥ!���&5^� a"O����ĝO+D�i1�Ҁ&��١�"O����ᖧQ�ޱ�b���z2"O�\ ����V�d��%㌶o����"O�`ѧ� wA45 WD��T����"O�}����=P�퓲��AN�\26�ȗ)}~@���i 8�8�#���էY8k�ǔ��0A�	�	��$H&���$X�9z���BS4���P �$x�џ�c��
(Q0�'���O0>�$@���R8B���Tj� !razb�<a��u(�G�0yZ���!W0Z�$bn�),F��u�ޱ����e',�&�<���^r��#�"�B���2�\!���N��i	�"��^l1O�h�*���(�*���������䘟E+�L�f��b�~��灖�}d�ɺa���'G�-XUl�x�'��M��'N(]WRi���GZ��qbʤX���q-�������ɻLѰ�;q�;7dA)z0�ɰh-�ȱ��M��0=�1
O8dP4"��M�� ;�#�͐��ƓLm�`0&�J�0,>��/�#l��|�˓r�X}%N�X����]3LF�Y�,�p��)��ECBl���'�(��(�Bm�����I.�W�M�`uX��R�
��I��x�T1z����"̥s`*���a0�<�c�P:?r���� X%�� ��C# Ykۓ|�
��)7#F�h6D�,!rhݠ�Z%>t(:f�&����PT�)�;��D�<���(��',R�g'��5bߌ1���3�:B"zrJ�����*��5&͙>��E� ��Db��R*+R�(�7�O��~/�URX�}&��Z�$]�g
�)u��e�R��sF^LX��W�$qK��P���<A���)!`)��BU���I�7��3d���
��l�T�Fy��E �H�3��Ӽ{ϛ�QSZ�#d�B�#���a�HZ<yǋ�(����:�2}HgF��&�|J+O��0C@z\���H?�I�I/�8��V&`��T�<P����=52 !c���"/����'�XaRe
g��4�
�.�Ti�'�6�rB�Y3~*�����'�Du�4@��@y�D*�(�G�Zp��O��PFA"s(��M����3��#� �svᐵ�v�S���2���%!4��pR�H6z"@I��U�z�*���)�(gŎe�,O�p���>��>��!k�i+�g�������+h6�ad�5$��[e���U��ԡ��D`��bŃ�9K����I~(�aJ �>�5"E�~|P�>7MJ4�d-�7n�6u&�r�B �ayRg� Z��m�a����$��._k��D��a�e�/��I4�|%����m��y"oς�\iR��-c�t0�vf���ēNn�"���i���|b@�� a��[�K�C��q%�8��T���4.yB�	.1&Ly�!⊍bXU�F��>.)�P�ʅ���9�B�!Δ	o�D]�M��:�wdH���ed�xL��gH�Q��tI�'���!e�Q<<,�B�8F��̢ڴ$�9ŉ��e Vӧ���E���K?2t��+��N6�83�&D�dJ�E�G����ӥC�4��%��K�>����n�J�#"&!<O�Y���ھ�D!�(�).�T4���'��j&��kTpm�ӈ�:Pڭ8�o�*�~��&L�Vh<Q5Eʋ�	S�̟(p�� ��m�'�n��&�U#;
������@�x�A��2����0$t�<�� Y%:�T
���VGJ�M���%	�L�
���֒>E�ܴD�l0T�3A%��(��$�LE�ȓQҭӴ ۖ R ӯM%@�i�'Y���
ȸ>��)��I�C��c��Оl��}��� W"��dL��E��i��Eav�#B-���Q���ͣ��X�'�:� gX!�<Z6(59��l��d�(�	�7� '��O�l���aI�7/�1��� '��L)�'���4"E�'�,H��S8#:���ݴF���L�%	��ҧ����G2͔09��3�� �I��y2F���`�kv�L�O���ao����֞&��e��I
=_v&���hO
�*��̀=������)�@CE�'�P �6��
�(���?f���r�G�K7��%�ɋX��a�ǘ�p?���E�4P��_�oJ�D��0�q�ċ�h�2):��ß_�ݥ����	 �lawʆ%�¥�"OX�p�51 r�
��ҴUs��)ֆU+'1.Q(� (,LY1�ݾ"��>�	.?�P"f�8%���!C��:b��C�
NX���k�!�ڜ�Q��o�¨�@��->�F��9_��h�2&|�QF}�+O~i��A��m���!$ʝ��=����C��E��G�v|�`ዝ\�p9냃Q�Y��� ���Q>��	�� �T��Qh�"���0J�(8�=-C!I����������n���Oh4��n��m{Aa^=F"�D��'QB8h��R"'J�		�)��q�F��-��	($p�̊� 2��i�Q>���'�ɀ�W�M��0�Ł$b����$��E�#�2�,򶼃D�
`�H�(ҡ���\�&g��`�T�b�|�6)�E6��R1cG��nիf�&,a�[�#�);�O��%77�T�u
�p��,����xTN<h&d�h���:��˙¼!�C�ԣ&��~�����������>A��9]'�~b`�/a��lX�c1�t0����ZX��!����?���cS�B]�,�mJp(��p�')Ё@S� ������VC�#|L ��+*���A�(�T�3Ư�O^#|�"��$)D%�2���R���()�6p9e�8ʓW�i��	��T@�K�@76��ё��h*���t� ua'�>]	Zኢ
����Oح0�l�811r� d+ٔ��i���'�f��d�.?F�H��f�1$nf�91E�Z~�0��Me2��2�n�Sӄ���	��p]��b�+i��%�>L�c���!�~̦ph�Ǖn����N�O�;��[WHJ
-bU�T��Q���/qh�`�J�	��U�G��9Y6  ����Hf���GJ5=��	R�O2lA��l�f���!_Ҥh�7��]��FN@�R5�O�m����8O�f�������b�11@���a��@">�A� 8" ��8R�b��MO�+�9X�	�!zў�#5����Fe�W�Z���j����1��9U�Lrl2�����G�I�?��"I��F���0Y��\�v�A�2����fH�.(ZLb���b@�h�L	�A$�-��)�@�O�8e,d޹�ĉNxa��D�JhAH���?��ƅ'_���f捰@�d�K��
 �\y ���-��		`@�O�"|��L��|���a��q��0�~���%�%(�(9YN��P�gJn�g����� �=)��T�;T�"���A �ё��^%P@�Aq��ƈOt4�D$*��PѠ(�=�e ]1k@�a�b�^�HO�jT+Lh�0���`r�����O���2\pB�\�],�����_�ՈO�VЃF�K�O� @��u��[R�����v�"w���B�d���ōfܐ��}N8�n�C��O�	�E�0v����|�E�2r�Ăd�W�O$v�AȟT��9z�e<^d��b�4`�� ����ϼӧ����D��O*�t#j�v����<zET��$[�p"��hC@\`��K~�O��0��g�L��C��j:5Y�AB�o��{��~���褮C�U�$���ќ�J�K��:Kg������Xy�%�Ž0DN��pN�Z�ɝp�>=a$�`��ĥH�	b*��Ua�s��\�V,�$q�ը��	i0V�KF�t|�Xc��58�6��>�B"	.�^l�K>�F*)nx��K��?I��Y�"ݐ`"�t�Ug��Y�N5��=扡N4���e��"�X7�V��-,���n�=�r����~ �����2r�%���	��r��Nׇ��)�� ��x}0*Pe�;Q"�(cum�Y\q����Bզ�!ʛWF��'�4����U
��ֳz~X�ȧHL5�JH��J�p�j<��ů<
�U�Ԧ4<O�a7 R�Q4x�$�G�
�@r [��� �J6	�b�"}�dЂ/XL��W@T�|�-������<�SHD�<q�,����{�,j5��"s��m�0Gd*%�����A �	�$D�2t��Y8$Y�0�赘CCAW�T]����*���3u��-b��c��1q��"�ds�C�%|:� u�l�N1�C��Ln���"";4�R�g�G�n�:aZ�L��!���I$��i ��f�'�h����0a4�N����p�F�\P
\�Q�!o�)��'�/W�����5P��5��s�|����@�u�W���D�+ �DIu^����T�`Z^ �!�'VhU:D�XM���;BլL6��Bg�N�#D���MB�3a���f�'�hT8@�X(��9J�~�h���:V�yjR�m_8e�:�
�=a���d�	*4�P)C�C?Dz�pc��6��ؠ��O��Bv�_�k�vyj�ÿmj�"=QǎZ9R���B>L������]��d���$ە��c)��I�Ξ���\9��,�4�_
|�Rچ�Y�$Y!�dS<,Y�L��U���s��T���-�	`�tS���4�@1���F��M#�.ȩe�ڄ+P��ٚ,O|�<��[N^���m9�D�m��/�^�����\��L�v
�3ғXl�Ӕ/�? ,�pS�[�n
\|��I�.�\}��F�p��r�-�4�i@�C5`Y�KGZ���ɺD\��{T��9���GOI
&�b#>Y�60:�|ړڽDn쨂-*C�	��l�k�<����D�����+U.�Ɲ�<I�CN;~�ȑ�<E�4�Ur���gL��c����a䙠�y�
`LĨ�揟�p�M�����Y��%��'�Aˢ��uF4��&�&�, �����)�K�$'b�;�
�d\x�� ��I�$���|�ya�@�+C
\�9CB�uG|��k�);��i�`g�p����81��Ę;hq!�D�) �$e�:���-B�`a���V`S����	U�D��O�'}�>��gK,s�B�I.(�h=X��,.,ܑ�e��{�B�`�Ly����T����Ԣ^�2��bM87>@��`,�OhZ�`�0VRH5b�Gћg
�M���lx�
�'�D�A�L�w瞁�rO+}5�l�����c�v�G�T�J �U	���(�XM�&��y2Y�H2tL��k�p  ���G!�yrX찔B�/|:q�UE+�yi�%�D��5�m%f���y"NB�a��I9F#�;+�*�(ԅ��yR�q{�#`�6u:����yB�
8i����j������y����-�6��aA�!]l�1�B��yB�X�&K���i%@j}rq�E�y��M���A���v�b��/׉�y�j	's���%�q�X�A�m@-�yr20
D҄�
bI�рA���y2_`�9*d��0W@���E���y��I(i�D��fÍ: �s��4�yRaߢX�`���#�?*� I@LK��y"��>/ЌAiX%�"A��y�FGi��ˁ"\�O��H��F��yb�72ͪ����M��!Pa��yn�F2T�aV��D����Tl��y���'���� W�$R$-ؓհ�y
� x�[֎v�j���#A D\����"Opջ�&�`�>� Ӂ[ yWd@�b"O~�pFK�Yf��� Y�7r�̓�"O4�t$�= �J@�aEՖSg�� "O�ـc�4t0=8q#�8L-� "O������5$�Y�P"8��T"O����0]��Y) ,�)��Z"O����cЍY��}R�L�H5�`c"O��[Pȍ�7|lU�CKP.*D�K"Oj��-j�n]	6�I�� �ɴ"O�"A*�Ep�#1�I
n�p�3�"OX$B�
�0�X(���F�Z��"Od�{w/W�O$�CF�V�?�h-H�"O�����͗(�I�!h$�@���"O�w^3N"�+vE���l��"O�(�⇚2g��|Rũק�y "O<͊�l-(!��2����?tZ�#	�'�M�d���%~ 9�n��ef�-`�'T�		���:]�u(ËQ��b�	�'c�\�Wo""z큲+.}���9�' 0ȥ��>p�,p��F�t�pm!	�'P���&Ô2Ċ��kS�Bp0	�'�֠�DlSp���k�+y��i+�'a����jI3eX|Z�昆p��p��'�L5r�#�3{<���� o��EQ�' �]�H؉m�v��e��S��}��'e�ź���~8�}�W#[P�hа�'�����3P�5��DW�v�R��'��L� �:jH��r�gؗl�2�	�'�ĜH��^(>ȑ�0,���p��'�@�r���K�Y�T��P�p8�'�n�s�	P�G�a�ΗJ*���	�'<r�R���0�(��F�z
�'>�ȑ�舚��T��Ĉ�7�~ ��'t���r�D/CN� �1IS�D����
�'�ԝ8u��*A�:1�͂:���	�'D(�i嫆�)�V �C��<����'�L#j�-~���b	Ékz%Y�'�yjBhȺ[��i��fν|_���'���Pf4|�\���*ץ`s`���'<~LfC�2:�"BeN�O��3�'���L��!���
\U4�r�'�x�3�F�"#�����$��5��'a,�z�&��,���Qn�����"O:��돃4j��֏<M��1"OXl�u��>P�Iїm�b���3"O�E���Y�!��	����tYQ�"O8�POڶvΡqc
ߚg4Q W"OTT�D���,P�QI� ]j�+"O"�0�c2{�2`R���3u!��"O�e8�"���!:ƮJ2�-j0"O �S���(W<�e��;��X��"OK^�*���ҌTJ������y�AӺq6�1����9�1玲�y�[1<*����lU/C��0�r�;�yR`E�z�N���H9�|�����y�%� yâe�qF˃ �q�qˇ��y��4��%�+�49���y�](t���g�D�v��h��eӏ�yr@�M���ȶ휬���k��(�y��Y�8�r�������1C�_ �yb� Cn�K�.Ѷ
=�xe�7�y�"�8mO�y�6+�9�XM�!�5�y�.Z�CC�`qF	�~���a����y
� $0�'��8�h��Ez�"O��h"��to(pLہ5�r�id"O�ay��()����ȓ�v�����"O
Փ�B��XU̠8q�]�o�U����-ړ��v�1���gh��1&��cMHA��� i�Q.ЍE�$r&;M͖Շ�cF�k�"C�L$x8�E�� }�b��__���.ţE��:� X/�؆�%�,�9Q��\/Эٰc֧fz�H��ov8:�^$l 8���O?Y�-�ȓ9i�=�d�� ������]%*��ȓ	����S#}��M;���	S��d��U'nM�6d�%i��J@���TC���ȓ0͘2�� ��tҧ���	���ȓ!�>�{�Γ4ttp����0�Ć������l�n�H�J�[����ȓO`$�Y�e��]���Af,̥r���ȓ��8�d�;Sv�� � 0����r�da�I��C]J	�HX[�$h�ȓP0��('̭O�$�C(�
h����ȓ���@%Z�m��m�n]�3"U�ȓ��py��R.T��T��IN_m�؅ȓ/���VD�Y��D����|�T��A@b�[�E\H+���9S�4���G���5 ��(f���~쬼��J����V�j�m�'x�楹��-V�ɱ�9D�X�Oш�Ti`X9-%lRe6D�ѴE��ʮ�'`A�PDI��K:D�4�ɘ�6�RF�@0�*=��H9D����AH���9�`o�E���q�7D��!F�W=�@KG#[�$|[��:D�hU�N�"�-��h�)�~<"�9D�X�t@ʴtj,!���V��G	"D�8ѥHG�W�Z�b�X7_N���e,D�`��k����@�R�I��t��)D�h��?�=Җ��
�)A!"D�ܨ����`����*O���`:D�`Bcc ;���"�̈�}v�o<��s��`���I�|�H���!�1A�^���+ D�Dk��5r`�0�C�_7a��v�;D���U$Ng��ѥ��P�0���5D�t��-[)F%�Ѫ�� |X ���>D� 8�I7 !�h�MAu�7D��ʓ�	l���4JӹP��)��3D�d���pn5�����e��d�&D���0gK;���Ι.Y��)[a2D����"]	�P�W������Ũ#D�����L�]@  $/��=Щ�f� D��j�g_h�RI���EN���b"�È��pzS��7v������ڔ�9&�|��)�S�kۆ�y"Hm��Ոŉ�K��C�ɬX�:\c2e�(P`P�!0�W���B�	3t�0��
e�]���[�AB�ɿL�uZ@��+�u�Y�v��C�	:�ơYO�	�~ɸ�*�~=�C�	�h���q�΄�8fj�)s��3C�vC�	�AL��b��MuQ.��"K�NLC�	2
��V�U# ���F��A��C�I0	�Dc7➺4`䴡��Z7y"�C�	�j>`���\�q(���3;�C�	2$0D��w�4{2�A�<O8lC�	�g,���G�%8x��'���B��7!�����k�.{�`�D���D.}��I�\��q���rU���ڒ�y
� ��r
T
�䑆OX-*l2�"O|@��
�>��ӈ�'�Ҝ�B"O����m�z}
	rA��v]�%34"O"��g�l5�E����@v�)a"O��cwF�%B�4�#�O�hj��"ODa��A�+V��D�!ܣ|b��e"O(S�'�������J�>'-��G"O��HӬH��b���I�}!����"O>K��ȮV���4��k-��h�"OF��ԧ�0U`�h�&Z���#"O�@ o�|���z� E$/iʥb�"O��p���_�0��1��aG��"O�A�D��$(z�� ;&�֨h�"OR��J�#bY��b�L � ����"Oz=B�E��B��\��;V+K�u�!�d=��� �ˮF�,y���͠o�!�$�2h����醇I�j��-�� ړ�hO��HPm�_N�!3��k�H�J�"O$���$�<\!P3�Ety����"O�%�6�^����r%���jp���'�ў��
`�(D: �a`�xK�+D��W�A������,$Ҋ��/7D���&�['W٢A��N5�Xɺ'!7D���f���|A0)�0��10 �]�� 5D�(j
Q�x���f�V)B��R�3D��j'��,0�+W�� k{h�a�0D�Ժ��J=_�<�G��fS4��h9D���B�I�&��U{�߬��5��<D��ha&K�vL�"`JR,&��f�<D�l�R(�0HI�|a�H�F�
AZr�$D�L�T�M(gF�q�cƞnpF�{��>D�$	t�G+u���n��=3r��n=D����S�o����eǟ9���P�n<D����"�<���f��<{�H�be:OR�=��L�r�P"��CNAٳ��F�<񑂙�  <�҅
��F�NY����L}r�)�'9�N�2�%ް#��9��)h���j7Dk` W4,8A���R.8tĘ��]
ʴ�Ee�&N&T��۩b# ؄ȓ0�F\2����!h(�c�("�
��fS�}����?WT�(���N!b�@q�ȓc.$�"��ʝni��#iV  آQ�ȓ(��`��kE#i�2�t$�}E2���d{()�"�^�jL�L�4��w�|�ȓ.��I`S��D ̠�_?A;��x_�̱7&��u4�T�W��q�<��6��2  �c����7�@�i� Єȓ �0��%O2VX�ր��e#(�ȓ��(D/���H�'9y}�5����5ô��x�`�4' 8��-�ȓj�BD R�
�8,8Umς}�ȓ-�<SVCK�c��A��
>��\�ȓ
��q&���0��uڦ�K�����1�F �'B�F�ڝ86l?+H�h��Z����'!&��!IA�C�f�ȓR,�(�씨p*�Ď;{�x<�ȓL����4��Ɉ�ό4?����J����0˵J��d�Š�8v5�ȓ.m��e�W�u)��©p���9|��+W*�.�L�g� �N$�ȓ[�j�j�A�7:�|!�=f�lD�ȓ	���G�D�D��F����ȓ��� !�n�XE��Z;v�݇�-g�u9�к0��Q�ЭC������S�? @`�q�@ ���#���#&5�5"Oj0����S5l����[�>�9�"O�1�+�P�<��7dW
F�,��c"O�(�am8b�jXZ��V�3����!"O�Mp�C>S�R��d±qS��z�"OΈ��F�$���r�R$+L�Q{�"O��:a��y耀:�KK�v[b�i�"O ��L!f-2yh"h�4S.�WL�<9��]Yppl+���R�8���)�\�<��	X�˳�Hd_�m�4��`�<�4��F��f�>,��Y8�.�U�<!��@�rk$e��1[�hგe�L�<���.V��{��ͰzܜH@-�K�<�C҇!��w��6B� VjK�<�A�Էs ^u� l�+*�����DJ�<�r����9�g�'&>V�F	JH�<�g`��,sd�h���,ex<�	�D�<	�h i�T�8ce��$=�q��h�<�/Ú���c�S�P"�g�<9F	:yC2a���D�`	�f�<y��
���4)�ܦ%.�����a�<Y oE;mZ�[�F��"������s�<A4�-iH.��퇟[C0�j�/Xp�<If.M4u��,b&Əqtz�㏟m�<q4���PNP�A*�S�-�ĭ�B�<��m�8l�bA#qX�P(�!bW@�<�X"	b�t�g�ԍ�h�
�z�<y��P�B&��eBn|�Ҵ�Cv�<1�%OD~Ճ��X�Fr�<�a ��9��T*�\���)Kk�<�A%*��@E��9AN���7�i�<qd�_n��)C�`C��h�K�}�<�Тˇ  ���-��`r��eI�v�<كM� k� x�ے�����\u�<�cm��PV���[el��w$�j�<��L�\�ZQ�d��XW����\e�<�&��59�������b�ha���^�<1aO	B��:V^�$�0i��^o�<�d �?��e�%G�{Q�I�v�<IKW?O�����+�l5x��%�Kp�<��"�3�*1�@AĂF��A�ho�<	�*P�D�1��C��W���ia��h�<����1t��5��'��TuI�B[�<���d�\,JA T&��#� }�<�piHV ��7,�
R�l�S�<9�&��	����ϙ�uw��T�KZ�<)Fb@��jHpG�K�< .���a�<��Y|^�m�G�ׄqb��_�<�㯑�+��Z��Y�"@U�R��\�<��l�.!�qD�Z�1�nBB��Q�<Y� W���RF��.x��$�Q�<p+^�^9�w9O�<ai�h�<I
�B�t���I*X�0��.�e�<�7��A!���P V}���b�<��O(��§�D�P�r$��%�I�<!!$\3����b�En�C��\\�<C��m�t�ˇ ۄat@�{�'c�<1b��A7�c�
�&�����)]\�<��g^�8-�Ċ���_V\�զ�Y�<!R�� c� ���͍?��x�͑U�<�d�Ȧ@2 Ӆ\��d��#X�<� +�2�(��ꘜN� 0�DNU�<92��G�V�P�J���XT�\J�<QGP\���R C�6��Q�\K�<� .���+�	X�"��;�}�"O4;Q�N}�|tk�Hu@�ab"O�qk�-P*E�"92ō�"uR��e"O��)��-��ػ��+��DB#"O"%� � �α1q�H!z��""O�y���&!� ����ruZ�G"O�%	3�8���� �
�z\Ja��"O���PJ-y�X�Rc�ʘVnF�!�"O~P#��W M�T�"đXt�Z"O���5pl��x���1 M�Ik�"O�m�&+Z�W�p����$b�b�"O�U��!ܨ,�����&��#"O41�R�H�;�i���X�0r�"O��ip����r�8L+��A�<�W�רҜ��f®J���3����<�u-��I�ZȂ�4Q�"xs�L�v�<��.Al�>I�4������t�<!'��Xh�}@u!�������l�<Q�Mݛ>��"��؅.LĬ�H�M�<y�Í�~6d��Ac��L:S�RB�<Q���,������ -��I��A�<q0�Bx�Bc�Z�ej �9�x�<$�����Z�˃m�`b�J��ȓ\���%[$_q4�q��"����j�:�P�#�_d )�ũ�.��3���w�C�A�pm�bI��^��ȓ.y����FԤx�i��j_�Z�f(�ȓ�钶���g�����\#@hY��5	t��9%˄@�E֜5ށ��BP~HJ�!�2���C�Z*> ��ȓ|	uB����8d@��z=��S���f��;x�ge%�ࠄȓY�R��bM?L�L�T`��ט����"�*�AK=@����d �<>�V,�ȓ@|"�P���7�p���A6G��e��g<�))��z2I�rhܪr��ņȓi[�����tbjE�|^<<�� �.�3�e>~��$D�(��ȓ
Ć𠦣Шo�TP0��<V`a��B�t����7�MH����&"V��ȓ:��M�n�4/O������4_��t�ȓ<Yΐy #�����F�A�h���ȓl�M��JeJA����d����c��W  ��b��g��	�ȓ�ʭ�'`T}6HH!i;>�̈́ȓH��l�t��0M�ԣ�� U����F"���֬�i�\�\I�:�� "O���$(��[t��u��h��"O4K5�0I��������y�"O�,I�y�N��#U��DT��"ON�І�λ3�Pq�Ӈ/1��H��"OH)���!=�M+a��4<�&"Ol�����60��ń�_`1ӕ"O.�� F	)K�ڈڀ%F�A�@P�"O���A�;P�8Qrģܡ��S�"O� 1�b?H�+b$�8w.ۢ"O��K0�ϧ��X�!��J�B�"O��H���L�x	y�����Y�p"O��t��k P� AG0~z�H��"Oh�V���( ����a���br"O�p��C %)�Zyi�Є*z08(�"O��P��P�(m�7)Y�;|p�it"O^�#��[>M)�K�g�8v��a�Q"O
ģ,�/u����?�����"O� FTq�-�������͙���
�"Oh @�<{��lKVMFG�P�"O�MZ�Ğ ���*�̈́�k��T�#"OD�"��H�����x�6"ON�裯Q�!�X���V��j���"Ot(y�fZ�?$HQ5�"y�bh��"O���i�2#x����;:�)�"OBT)����v��,�I��&��\�"O^M8�G��d�Ps&�ڽg����R"OR!����5�a[��v��q"O�]r1�G%i�U���g�d�zQ"O��xÄЈf�^h{�ai9|�B�"O�T!�ʙh�i��R�h�$�#"O�ɠG�W��
pJ�mR�"O�(�Rh��(\ҭ���Ks^���"O�c�"�	j��Ec��Xm��ٳ"O���C�h��}�wÜ�e�I�t"O�h�ã�e�0]i��?\D���0"Or����� 3)PA�'Z0���"O�1�
�]�$0z�≐x�\I�"O���G�xz�MFD�%���� "O<uxb�	�lUȔ�! F�< �v"O����?2�+ª�z����yRي,b|�/[�b̌A���yBNY�(UVm� T.�+R�ݝ�y���'k�f��r�à2��`��Q=�y"l�}�>��%o��M8Tk��y�さu��l#A��3ڬuT��yr���>7<�tk�2�bQ�K��yR͔�N�5� �R�3�J��3�yR.�9g�4R�cP�S�3�k#�y��X6t����Y�
L���ꂤ�y���*$W(S�}�X�r0"���y򦖨)��LK��	(�|���&�y��Y>3G��Ʒ&�^<Ip���y�ra�Ŋ�8��x��,\���'�����9�@0��j� 1�����'-��)A+.D�8��Ah�0�`x��'#UZ0��ʸ�S�(�{w�l��'�Dd�JОT�:�{$%��o1���'2��&�Ϯ{`����bVU�	�'�t���H6s��t��
ø�"Q�	�'~��J娅O��0���:�qR	�'�4�0�~��#�"y����y�h\�&vlRCUN7����P��y��Xv�䉲gCU�HHp�{�FZ:�y"��/b�2l˦�]W�`(�B�E��y�]�u:`3� l�(�G�Ւ�y2��@����L=B�X���A֘�y�K;[T@�u�I�>f��ё�N�y��û"oT�q�BO+5\0uC�Қ�yR�̦9%�u��$C���#�ԃ�y2�ŇO�b���S=fu�,C�iX�yRa[�k��0��U_u(�"��W�y�Ţ3٪T�pꜾF��G1�yjS�p<Ѐ5'�%;8<�t���y�h$VZ���`�ÎC�~������yb��N��@'7߶lh�B]��:
͢b���
*�4ϛ�}�tT��2��|�#	$#��z&ˆ0<��0�ȓQIZ<jW�N0����g�7C��A�ȓJ�\��nzi h𧪜��x@�ȓF HY��ۦ0�l�r2�Ҭ~2@��{��%���ц]*�M���T!U�T��S�? �T�6�*=uv��G&^
B�FE�g"O�}ӤoҠT��3&^&.����"Or���M�� ~<Mb��G/��q�"O���`��& �2�˚i=��t"O(�pc鏈3*�͌-0$�!�v"O���,J"$Er"��U8ȩ"�"O�d��ʝ1���`,l�b|4"O�(�V���\���REظ6�J�?�y�É�?z\ٵ�Yiʶ_7�y�b4n��r�	}���HV�O9�y�B�(w������_��4�f���y��'w̠�ʆ�YFu���Ո���yҨ�`�f�a5c��DW�8˲	�����hOq���
�T�t��m�Cn��z��-k�<��_ 8*��(B2}�I1	f�<�ģJ�y�*t��ǁ1]�����i�<�D���lu	��j��`�r�0�i�<� ��m��t@�eZ0yZ`�P& d�<�Í��}��5P�H�$��𒅂
]�<�B��L����E�ܤd�")˧k�~�<�n֨H٦]I���$U�L�*�j�t�<T�y_��#0kxxU�O\�<�B_�g~��c��%*���˲�Y�<Qv��
 	6���Ɣ�])�x�� o�<q�b01M*���&��L����7
�h�<i*YJ@��r�Ji�F�(pg�e�<y�Ɍ�8���Q`�ѶM%:�;��i�<1�-��ic`��6.V���]�<QW+�4!�1�,$b��,�V�<���Tn��
`LT�
f,%�BfM{�<����:]q���;���Vdx�<w�W�YHD����U�\r21:f��v�<Y�H�-Gc��x�ݬ0Q��"#o�< �ҙ~Dxaz��H���!�Dkyb�D.�'C`<���+O))�,�'��B��܇ȓ[,V�#�� L�@ə��d�f��
t$R͏�3$a��)Î�*A�ȓ+k�(Ѧ��6\"<�@�@#�f���# ��r��#R�0�?|�1�� G�]*��E�\FP��Q=MN����m��Li''�~5�����wd|���Kp��8iD�%JFO\F��ȓO�TYUK��W�]H ȉ�=�<����AR�JY2gL����#C�$Ƭ��� �DAfivUtYR.�9���ȓ:�<��-
5d
"�9��G4:F��D��<�%)��3H��0��P�rE��FDcC�o�2��A�'1���r������4a�M��	T8�BԄȓ���yŤ݋,U.�3oE�b掔��M�5���'ai��#6�T���qY�#���j��ءeiV/T9X%��`mͲum���.@�#�d��K�h]��I	dR� ��N%9��0�ȓ�6��)2Le
`� o\Z%v���]ڼ%A3�\gb�u�Ġ�D(>I��Q��Q����g*�a���r=�ȓ�� ��O�7�����+�����[��}zlN D<�OO	�݅�N��I�K�`��p�Iшas��ȓ��0O��x�ppp��@�
����Ɠ#�6aPZ�d��؀U��.V��Q�'�1i��A�Nk�![�a�����'�B�F�f�,l+�G�Y<2R��� �L;�0��IP'2u>�T��"O���̩�p�R��)n�&��"O�p���Qp"��a����e"O�8��^�u�b@���I�t����"O��k��ɫdJv퓐�ݜ��c��|��'�ў�O���B"y��� ��?Oxl��'-��4�Ƙ,�����n�4�����'�n�`�@ 0(U�fFɜ%����'ZBq.�u�Dt�ebP�\�pi�'��;0+4�|
�$�Bh�I�'�X���)�=�p%���աk�Yi	ߓ��'�X1��F�u���0��58FX��'�L�����D�C n��(�t��d4�'$�xU�V́!zh���Z�0���?����j_H�m��DN�ar����a��[:m�F�|�p�ȓ?k8�'�_�f�.ǂm-�����mK��]/�r ��i�O&�ĄȓP�[�,��4��|06o�Gt�|�ȓd��Y�ע��1_�%�BF��4�i���Ɂ(�y5Lp���0E�za��	��,����J��DL/^��U��]�Xp�&�2�Yb�Q+u�0��dA6Ȅ�]�"[�	JDL�I��ч��T�`f��'k�`Uɰ(�|�d0�ȓN)���[>J���s�%��Ѕ�ږ5)�,�0������M�l?4���	R~���C�$i'L�U�v9�˔����?�
ӓ8%B(�gI
�c��U˴L]�_���}��a
Lr�&!s��9Qg����Bh��,�(g�F̢�j��p�f�ȓ^T @�������/1Z���^8T��p�#�XC�4
P���@�u�F�/ɬ�"%E����b��G{�����4��LY�)!�XCbF�y��J/t)d�	���C���y�oS��$P�'.�9i�pe�H׵�y��M�'�����)P}�`*Ō]�y�R9J�9Ǭ��^9y%����yf��:o�Y񥖘 ������<��͵
�(��BgW VQRF(�
����3X��ɩ1ǔ7X�Bm������0?	�ć8f��
��])Tɬ݉uJTZ�<1��^X�<X"�ӊ,�2E�]�<�"BF�L�����V
e��`s!�`�<�w���U������D�3&��F b�<�'��4�i�%g�O2��	7Qߟ��'ў�>��e.�&U�ܤiPj� D����O,��2�S�'@ ��Ғ&:v���YZ>��Rui7D�$@p$|�@�%J�C��HFo9D�4ʵ�I=?��3!��M�����A2D�8"@�Cݖ)�ސ:���S/D���_�(0h�eJ^P�
$��+D�����ۭ
��]��c^7#[��� �5��刟rqȱq m�E�rFx�{��|2[���
`$�-�cV�"��#��-�&C��'&`:,0EL�~Q�hRq�� �C�ɽ}4�I##ҼO�����M �B�I�>j]�@晩P�RA1�a��~��B�I&?T�!cqɏ�
R ��!���,D��:�G:���U�θ)EA�g;D�����֒,S
�3��K�vV�����4D�t�&�MlF`���#Y�U)6c1D�4���
Y����SI˪i���F0D�� ��{��������;�`i�"O�����2KH�bD�� <�&��"O��JL-Q��DJWJ��3����e"Od\#T���9�pК���|���q"Oи�u�IvzБ�I�zn���P"O�)���	?p�Z`.��&w���#"ORA���(����3�eY�Œ�"ODT�A*?9~��VN�XH���"O�X�6�	.�TY=iDe��"O��J� �<<��P�K^�}�"OάqB�6F���5��!c�} 6"O�͹�� �*�u�ũ͜iU��"O�=:�ヿf^��G�7Wb��F"O6�p`_	�PR1_N�A�"O�аG��v���ڕF�%{��!RB"O���5�� @�D�2��.�ع��"OF�{���"�ޠ ��
b�`��O��X�-M{�*y[��N�S%8D�dS�ZN��F���W�࠳#"2D� Z��P8.�TA���"��;��5��N����*<8��v��
 /�Cd�!;
B�ɞN��e0�����x{.���B�	yw�=��*(�j��N�S+�B�N�6Z-*7��X�$H�ܔ�� ?�g�m����d�A�T�P��Q�<ѳi��PB�ǅNqڇ�K���̓߄0:�Zby@}q��K�l{�I�ȓ�z��&��j�����T"W��E�hT(�I��qTrpӗH�(r�y��=��T+�)�4�1�6��D�ح��R؄#��:�8�ӱJ��[� ���������.$�|5�W+E�	��uۡ��(�B�	�23��G�W�HĤE�`��6�C�I�-�j�(gO;~�1��+��㟈G{J?=aB�^|v��EU18f��jU1D��*D��(m�Ĺg��/[!�(��/D��q�)̀:��ٕC��`nnز�.D�x�e㉐�"XbgOʖ u|԰�/'D��A����5�2��"L�r&D��9�ؾc̶���� o���%�$D��q���54�q��(��R:A��E D�(�t�G�y���x�L�}۰�=D���eÂ5>}r���)F�����k.D�<¥��i>���� 6rؠ��h-D��cn�`xN��$�]5R9�\Y�7��Z���ӎH�Eb3

1��5X�(ىr[2C�	�X4���G��nI�gd 
C�I�t�B1��&E���QC�4b}2C�	�\�����x,�DIA�<JB�	�ܥcwad�P4³f��B��]|E�%��iqVI�kZ�T��C�I�X����%k�@�"�x0FM'kJ�$7�S�O�����D��q:�Y��(A)FL�`�"O�� 	o$l��ğ-DV�M��"O��!��ڡ-�aذ��;K��#�"O�(�

al�ݢ�jA�C�2]� "O,��UY)Ӫ@I��!̪���"Oh��v��r3<�вgB�Ä�8C"OP$ɤK��,D2p��%�z�V"O2\Q�Q�lj�o��� ��"ON�`IL�<8Is���=c$��P"O�;`��zA���ѿsVn���"O�i �ٴR�(AJF,&C�	e"Op8�b�̵8G�aKc'�8/8m8�"O� Nձ�FWnnx�G�Ha��ȴ"O`�,�5{zH��5�ȳOX�i�"ODA
�α�mI�n�J�rU"O�]@�#�9@��A��2<��hv"O���P��(K�P��"P�;��5�@"OD��aڭ�� ��b<}����"O�	1���U2�a�^���"v"OT��,�<�E��"�'���`"O�l{B�d���Ёa�(������w>}��.s'�8���6S�ݩ3C1D��J��-B`ɪJ%�xQɒ�.D�dH����9�B	�Lꚍa���Od�=E��'V�%�,�â%����h�4��7K&!�$|!�\�ff�8_���%Ɋ%3!��W&.8���D�"6/�y���� !�$�	^�<�X �/]u2���&U�>!���r�T�����-o��s��W <o!�D�$�¤�"�P�k���x!�7U!���-'�<�x�(�Ov��z��� �!�DV�A*�SU�B3fE��P�㗩\�!�Sf:�q3�ʄp�д�@C�=�!��S�Z7��pU��T�Ĺd���}�!��
/'��B�
=2��hSa/S�2�i>MExrj�<uP��Z����:�,�Hi��y�D *�$�� �4�\� 1�޳�yr�@!*͔i�q�-3�`�̳�y��#�0�J�f	�#�<HG����y፼�F�Y��M	'�x-�iڈ�y�dS���ZD�وP��5����y�(�/�tA�"�#V�=�"g����)�S�O�V� 1�"q2�,+w�ژ���'�$��p/{�Pq�@9�8��'D��{�]��Id�6��X�'�,F�ǣ;�8�� z���'� �ە�M5S�䴀�
��
5�'* T#�%c����4R �t�)�'�6\a��=
�����h��	�
�'�^� ��y�p�3�ԩ]�Q
�'m���4fI`������>l!�8��'��dzb(��uG~*�BӒeZ���'�t��ǀ�N ���5C�\ �'�J��7 �Cr����e�*�i�'����6�Z|c�����k�.
�'����Ô�pkb�y���a���	�'�݁g��6ܙ���'*����'p��6fѹk6�P���(h"��'j�d
�J#p6��7�"/�9��'h�9�
,�@����"
:D��'\�m��,L����g���20�'(�Ͳ�ʫU����&�ZJ�uy�'o~��s�(0�T��FL�xm�
�'�h�A�'Z�6(h؊�(H�8֠��'����Ӆf�ҍ#t`��7�7"O�=B$�W%7p�'�3i.)х"O�Hqphܦ~9��B�X� hV!q�"O���Զ?m�A:�8q>N�j�"O\�2��7d ��L=W��"O�����������?`���/D��R�!<����% ͚:���";D��3�#r�%
�I�@���8D��(֦�!k���3ƚBY��aa�6D��֦�y_�pAEЕҮ��4D����\�����E��/P���0�7D�D1��&D)`IiR-�&:����q)D�� �e��O���l�)�Z�:2"O�X�s@�h-4QzR���;��Hs"O����q0@q)D+͕|⒉ �"O�Y��Ϗ6t(���'ʬm���'�!��&B��!AbC�Q��q�uA� �!�C#8rB�"ǭ��00��"G!�䀏]�Q�!J�+�"�Rf �x)!���a�~���O�y�1�  B
!���|�^@Y�ĕm�B�U�/�!򤙿8R9��&�2|bm��Ü�!�D\�@G>�j�M�L�N*ԍ�A�!�$	�-тTS��ƥ����0.�!�D�*nb�i�f���P)�3mw!�d��� � B):�����M A!��-}O>�r��+:��e3s��9џ�D���))��e�Uf�1
�P"9�yRā�#��`;Tɟ�kwb�(P"
��yB�ֆj{Y� ��c1b�#0'�.�y	�< 6mOW��E�'�̴�y�lR�M|��9PL��Crxx�蓶�y��H�+||��WN�:�RA�雼�y��<� ��R�?���s����y��h�rN7�P)d �y�f�7w1���
�<����CEȣ�y�M�w��y����
�DiS됀�y�ꏽm|�r�,V�Qֲ}K@K��y��
1�J)s0*ίEb�����y�Kޔ����6�ȳ>P �R�/���y��� ���FU�lZ.�(g+֤���hOPc���A$�݊uCX� ����H#D����I5�8����T�r�����?4����hƎ}�^�AP���TT�<!pI�[�Z|��ś8�"����SN�<�A獺m�V��e� 5x�X�Хm�e�<����e��Y2N7`��w�<���ƆF��y'/�0N�Ӑiu�<q�0;�2)�I����3�MZf�<�N�'D$��*<Ě��d�<a��X�� ��0@�;OC��S�U�<���D�����ĺ.z��Pơ�S�<i���stM\�a�&"�e�<abgò8��K��5�8� C�h�<���ԩ>�`@�Ő<��F��O�<q��6E&1�6��` �tR��q�<ٷ���RѴ(x$*Z�J�q�ɋR�<	qoB/P����%�|��!!��f�<�����D����I�]t>�@N�a�<��N�o�J�*�� �]���^�<9u!I\!`w\e��頶��]�<�F�3��,�rX3�R �q�P�<�A*:H{�)�*)pt��
^N�<��Z8�:���&J.��@��\Q�<a�ۋ�v� ��"w��!G�S�<�@�٠^.���&ɴWIX-����s�<�F�� `t���@���j��Yt�<Q�./�4$���(D�Hq�<��C��<m��g����9Z� [W�<�ga@�-�>���g?������GR�<�1NΌ/�*�	�`E�S��Q�Vr�<i�����l�"�G�o�ry�k�n�<ᶣ�.$�$8a�)C"7��a��
�_�<�� 7"�=�W)N_��,��q�<	05ߠ��J�=��l��y")F!8�I�B�:�Ui����y
� ��A�CdD��q��#F")�"Oxu8`/�"��5p��	O�D�2�"O�����~h֮7*�@�"O&<�2@,E��E)��9K��[�"O\�2%�P����QwB��i.a�"O��c$CE�K���0�.X��"O-hӠ�   ��B7@Q.i�N$��"O&L���v�Zģ��AK�U�`"OV�aP�S�m�L�@�:<����"O����A_�s���3^�uҦ"OH�r�o;/,�H�&�����$"O$H0l8H"*R�N�D��`�%"O�TQ����,U�UGf�4��A"O 2YG���8p���T�thY"OA�FP0wS�����%���"OnI�ī�g�4���ދXr��
�'�b�w!�e!J��C�{;�R�'о�v"N(@*83����B�d��'&@Q�,��J[���=�T}C�'��5�a��5T���둅�:��Lb�'h.��sH�'_�69���9�pls�'��-{�E�2u��h��g��$z�0J�'� "�E�	\/pa�ǤY2!_H��'��=;�'��\r8�ċ�p�ȅc�'���š�C� �W"4x��'�*X	�Œ/vp��ƪ͔@��=�
�'�l�Qv�ҹE6�)f �=����'���ar�Z��||����&7��	Q�'��mw�� &ѳ��<�m9�'_���t+{�q @
 ��d"�'���0G�!''hh�.��A{����'��Tm�)�4��cl�!g�4�B�'1laR(V$L���3�H,d$���'��up�K/'��=6��;KFb,
�'�Z���l~u�	�RlT0�x}b�'`V-���J�H��1	R��@[�'0����l�0~�����H(C�����'VU�'I%V�����%T�Q����'�d���/ڧe$l��%�ܹ�	H�'i���:2\yD���T�8�'C�@�q	�=&�3����'��$[�!�>f�nc��H3e/T��'2�@�aͦ�6̡"��'I&@}��'�V}�6o҃OC���1cމ��L`�'Ʉ؈�"%q�b���O�b��i��'r����煈"�:us R'a�^P�'6���'' ��9B��?i@q��'Wt(�oP�ѱ،g�0�'T�y{�B:Zћ�l��d��'�P@!�O׸\!�<��E?X����'d@y��g4�@�`/[�?�$�
�'�J����/���G�O�<%���
�'Cb4�@(��bgX�:��DA
�'K��ЋH�dshݱ��6	`��vH=	��0j*A� %�������%����J�_JP(�����ʓF�\ժq
۱$(��oZ$7��C�	�l�4�����I�U2iRC�	�<��ʳ��
p�	b"��t�NC�~��-#�លs�¹���N4�C�,n:��ʱn�>_6�1� [��B�I�Uta+v�A';\��C,�rC�	�٤����َtaV雵�U�
0|C䉈�:sDْU�ژj�H3 �B�)� XX{emF�]xh��́@�Q�d"Ot�(��)�
��"�*`"��"O���BX��]3F!]8%�Ve�W"O��(@!T g�
��#�;�tl��"O��r���'r��9�g/��!a���Q"O�5s��8�<�@�/�RS����"O�0���?4戜Q��[5@=K"O�����"(�|�S�Tl �y��"O��Ks�+^n��yblU�O� rD"O�����; YhA�Jф*iz���"OZ�
qK�!� �Qj�#Z��;�"O�$��hϊ������(?�]BF"O�yK,��B�\
_�
�AѡեR�!���	v�������c����4	8I!�  Ԩ�P肅_v������U!�K`��1��E�nV��1`�/�!���*w�c �X���� @H
�!�D�6�@P��y�eU/�Py2GMed�Gi�0H��}㢁��yRe䝑#�ф0ެ:�k���y��*#��3 d�'��X���<�y�Fd�n)�4	��!*:�!�#�y����<��Ⱥ�� m�l��DW�y���p
�u�t�A	q����y�m� #Q�-Q%��^��Q(���1�y�f��9��+S�X9Y�&�8���y��PE�X8;7D�Gn:D8p�A��y��1k����*��CSn]��L�<�y⌏�CzXid�
!��H�yr�H�CƄ$��G�]q��eF�y	�%L�A�P�\g��;'��yD]�M���В�=3̝�aǗ0�y��͗���DOt�~�@�����yr�L!�L:e��$i��eA���yR,��//�T��ʣ\rHR�ၔ�y�ؽl���R���*gw�@���"�y�� Nr�0����\j`�K��Ж�y¤�*:@>l���
�'-B����9�y�H��5v  �l�2�4�hV�y��ч`BI�u�
>��3�ѵ�yR҅L:X�b!g.��1� �yL(�`#��3<S�pRQ"۷�y��t��A��ߞ`2�@�X��y�	7T�Ի"g��Sx=�0쓗�y���w3���K�}Ev@p!m���y��6s̢��I�!#�ir�$
��yB+�>s�@��W�$1����G�	��y�F'~.:r���'��y`L��y" Ћ\`�A�v� /�\�����y��q��`�Ĺ�Ȱ�G�Y��yҎ�o���s=P�׮���y�+�7j���l��w��%��>�y��
AdP*�.Ŕ��ō�y�CJ�� 
%�a�l�[�yBPrl��A�FWj.h�T�0�y�&ыbJ�da3˟274���B�B"�y�"B5H>L�15Gř=ft��R@Ԡ�y�*֕Dj�`& �;ǌ����y��=��Lہ�_�15�y��b���y"�R"U1�9��*�1y�k3�T:�y�J�>���BLܘ4���Q���+�y��TṈp�A_(*���� �y��T�.��g�!�0�cs.���y�`ۉh�|�b����E��j��^��y
� �h��-H�����CJ@�x0��"Oށۦ��$
:��S�Ʉ<~zt��"O䵢(B�S��PA�	���S%"O�͹E�Bd�srA÷-���@�"O(i �m�zQ�� �O @ 
�"O�a���j������hu9�"O���&��(	<vm@'+K(>f4yC"O���raZ��@�I��_x8z�')`��p�Ŵ�Dx�nR�����'�X���ƾb�~��,B>$.���'�:3h�<+��<��&��FU��'��18���)O��;T�ȧOy��1�'A��%İ:7��BV�C6F��
�'،P��!¨X�Fx�p��+F묐�
�'	"�	���9V�As��,t*���
�'�΀�aN0k(�Q�R��Cw&�c�'M��Q���)\a�l�$�ln89�'j��2B�DP(<�a�@�,����	�'E�}gB�U���6%v2�0	�'!�d�iŦ��P!U	&I�y�'2*����0m���ڄu�4���'�����:#u`4G�ȿr� �'������<�<h���_�( ��'G�e��Z�� ���'M1f�r�'�ش���_�+G��Z� L)P�2�'����V��8��lB��F��P��'��MIa�G�l/ ��vAW�UP�S�'�h����G+�P���m��V�6iq�'�ȕ0�Рv�����)\!A�'�m����H�b�� ��9yZ���'K � �����P���!|�E�'��͸։L:*�$��c���m�'g�!��Ȕu~�p�ČH�^�"���'�d����x�&y��A�3'�����'I�ݻ"�YyV񡐌ƈYP��'� 1�b�����l�	�@�'e����%�l$tcULW<�\#�'�J����U�.H@���#�<>"���
�'�$����R=em����B)6m�	�'a`���
��D���O8G,j�;	�'��X��O�9�Јi[�F]����'3�@0�*�3HN����fK6Ix,��
�';R��4�*��մnBH���M��y��տOC=!E牁�5KX�}�	�'u�@r�gT"w�$:��� �`�b	�'���AH�'���@g��"�~��'���B�jԛ[u:�!@��v��8�'�����\�N�{�lG+�"�H
�'p��ZѤkC�	[�G!/L��j6"OBЉ�I�>�^q��jɗf4E�"OR��֌V�`�b�J$j'D�J�"O ��F�)�~x2/�&
���R�"O�y*%c$6�f/5ªDA�"O*!C��78n<}H��92�B��S"O������.@�}2�Æ�y��"O�$밦�g��������"O4X�R,\�v�:a8��U8f�y#�"O>��냣P� ��E��A�!"O$�@�dǵ�����,�riXT"O Ś@ �#D��M _d����"OF�$�5.@nТ��M���be"OV�b�!4�-��.>	�h�"O�ֆ�}�<Y4�y���"OF�`p
J;��Q�My(�2B"O� , ��o��s@�c�]�r�l0B"Ov�p �/W�v89�v�"&"O�E��l�w*�\��j۝H�,e��"Oȕ��kԆ|t�ɹ���XfFA#g"O�� �U�S:SD'D2�eX"O�!��D'�| �]�`8����"O���N�������7��� "O~�awN�*q�UH�D]:���
�"O�Q�G��5K�9�dT"h�%"O���
�L9F\c�bV6)BޘZ�"Op��A͏s�<)qcB�a��S`"Ol�R2��+q����∪�0m@ "O6� Ä�Lgν2AS ��)��"O�L1F��!iꙐ�o�\�R��0"O��OA2n����A/J:k���s�"O� C��Z�Y�L����N���1"O�is�m��_g�y�&-�4o�IC"O�-RG�Uߢ� �־��l��"OfTy�3�$�JV��+a㬄��"O���'���0%�t��q$4M�"O�JȚ91�~��u#�.v���"O�髶��,!2$��a�8�l=��"OvTc�%ՑJ������t�f�%D�\��A�aLy#aʇH�*}���(D�D:6k0�&|k���.�	�a'D���b"�m���bS�C _��sVj*D���g��92M�i�Bn��M�B��#(D��#��[6w�D���/x�tyD+&D�`cɅ/D{�(`���j�,�b��&D���6�?f�U�n��(:,ܓ�!D�PR�/Z�O�����G�V��]1R�=D���� �70��12�őf��}"q&D�����v�p�vȞB2�Q*��'D�`�v���H��xs5�ں���3(+D�Pq"#	�W� ��m� `�e,X:C�I�$�8a�2K� X��C�v�"C�I�~W0T	���"X����曊#z�B�	^�tR%���&
�]�7�֑e?�B��,;ƺy �d�*}�-�����+�B�IR����!��"�����		Wҡ�$�	���[#*Ѣ(�j��t��<A#!򄞌5�,I��\�ڂQ�����.!�C� � p�3 �#`�H,�b!��pe!�L��1�һt~��NQ�Z!��&Zm
�)�,����v��[h!�Ę�6)�YiB�L�8�ԝ�^+4�!�<��4{��NnI�׀W#'�!�$���(�(e��_��j�@B�<�!�DGm�-P�o��,�V��k�!�d��z�I垛W'Rj5�W!�d�+�@���g�	>VpB��_�R!�d� %��,�n��c ؤ�Ǫ�!3�!�X� �B��J
@�6�W�c�!�	
�IH�c'u h�AE�9yx!�DſJ�b��o\�T��S��C=Pv!�DH[�T��t��G�Dq�+N<cy!�*�D@�K�����ɂ�3�!�^"r�&��1���(��I�D�!�9DTQ��B���pZ5�A��!��$t���d�Z�n}{�IK!9k!�ć�d��	h��L2w��cS!�d�?"58
�c�_mcA��YG!���/���3�kʍ�nᷨ�-4!��`�<|Z�FԴC��d�㧎~�!�� 
8��ڞr"�rS�܌|�캲"O��i�G�L��-:&��)�|a�"OZ���!�g.��f\�$��9;e"OСb�j]�f�������Sњ�s�"O8��U�C���ps�ʮkY��"�"O��z#%��B��[�aBMR"���"OU`N����	`��3�pyr"O*�5)D4
��Y�[�f@p�"Oz,s��5T1F��\6g�b���"O���bn̜C�t;���<�3"O��+�!�P���G &'X0k�"Oh}�C�N�ęQ�N1c2�9W"O��ҭ��a��H��P�)n,ʐ"O�Dʗ�
�G:,����=Cݴ��"O\�'g�������I���G"Od|b1�Æk�42�d����h!�"O��CGO�/�S6��Y9���"O�Q��-|�����zl��"O ���K)z�<B��ݦQ��9Y�"O�,�cl��j/���Q
,�& ��"O�����K�9.\���	gx���"OR��S�'M�X�˵^svF� "O8|K![�
�:%�&��
Ndڡ	a"OY#e�tӜ�[�G�FP�AH�"O8��w�[&`�u�f�ۋ ���3D"OP ��Gҝ!QP�� ["�9��"O�Xh��	�3O�c��U4wj����"OPH��@,5V�\�#
r.@�"O� ��-�%t ����i�p�	��)D��!��.:�"	SЬ�x�!x4D��6��	bۢ�+VA�8;~�/&D�x2���0RDT�(�l��U�d}kb/9D�H:%ɇ�n���Ka���d$�x�e�<D����O�Sod2A
N����q�:D����G�>�h� ��Ivִ���4D���$�U,����@F�c|ܱQ��>D���e��7v��l�se�*NU�Չ��<D�$�`���z����=�0���F:D��9N
��2r�ȕ$�����9D� P��Ex�$�D�E�""�!Ȁ�8D����*��ut����A�0c�A	&G1D�@�j\q}\b�Y���y��9D�����f	��m��Α
V m�<�t�Y�{B]:�6U��jtvO�q��P�B���[ M>8��]�"Ob���͘7m�dq��A��%{w"O
��	7k7�����Ʉ�|0�"Ot�C� ѸV#�(0�ފZ���"O���P�D���W�܍����"O�!���ˣN��($+��\�b���"O�)X%Ƌ"��ܓc	#GP�5"OP��sn�;��"鋆Q�|�Q�"O��j!�)	<(���qۨų�"O����Z���f�+ir�`��"O�h	`�\�t��Y`'�	���pG"O�y(��J�.A�V�arhH��"OH"���a�r����XU`iw"Oj4x�Iӆ.W`8�h�
3:���"O�٨�Ǜd0r��tC|Q�s"O:�1�@ɀk�\��G�[>x� �W"OHCM��%ն�����?ST��ȗ"OR�DP�/���yg�����b"O�MQ�	�cm����
���j�"OXEb���+n��}�դ;ȵh�"O� hd�aм9�ik��F�:�^YY�"O�ű�#U>2�����bK&�TH[$"On���̺y�LcG#�q�p�
�"ORd�RF��h.j0���C���Q�"O�A)���(w�ڌ�B��?ID��%�i�铉�)��d]d�,�kD���t�if$\��a~�Z���uL�HZ0�B�Z!zT�5J�>	��R�z�ѸRF�뗡P�@q���"OL�sզٮl*Q�f㚬9iƱ)""O��d�	�,����!�$g����x��'B<�"�B/p��J`FK�6�H�	���~�cO-d�"����7r�L9�RjF	�yB�2%N @�@�M+VRl���R��y�)9,���)RO��SΆ< B��y���-��ͱc���L�'��y�gU��y���3G��&)�.�y"�G!0��23m��>���f����O�~ʖ"�"�u-�
l�1T������cg�TPhM���VD.D����@K(8��0��7+�`�B�L6D��A�bO #��P ��k�rXX�H`Ө��IyGqO�">yWb�",(1兓3�`��Tq؞tnZ����c����/�%R1�p1���9�|C�I������X�H�Њ[�v��b��Cő�ʧj@`�4)Z>q��D�f�\!���,~ �d��4��УG�ݵ1�P{�Ŝ��Q�\��j$fQ!G��<$�LpBKK:<��"�	=
3܈� '��4`�[f*E�!��7-���?)e�Q�����$�Y����x��4����<<4	��B̉b�d$�s�N*�JB�I�3��k2�&r�Sr�L�e��E{��9O����f�|���3��<[v�	Z�"O��SmFrZ~�h�-�.b;b9�:O�b�h��43�M T���P<��0��":��C�9l���03�Ҷ@���� �˒M�C䉀�zT�冑�5"����A�-��C�I+p����Th��ʍI���I��C�I�삵�b)	�^�L�%F��gH|C��.#Ct�z���X�A�Ӎ�"@<C�	� O�m�U*+e��8Ql�@��B�6PK� `�03�.=�B4w�tC�ɘ\wN�V��[�ͩCj�M�@C�	�~�01�MX"�8�ń?.�C��"0 �G���,��I�_Vv�I�'B- a�J�*8��*��_�{�4�hO?7��9�� ���%SӰ�ؒj��_�!�$K�B8&јQJ�0�r�$�ǑI���HG����&7s<�p�@� M�6�4aF�ybI���2@Z�'S�4F�ԡe����~29�S�Ow��@ �#_��8Z�*^�M���
�'Ҩ�2�NĮy(X�2L!F/,�kJ<�}6sѠ�k�����9�"�Fx��T]���)�Q��А6Ƅi<�l�!�Q�!��Sr���/L�d%"��T�t�Zi�<��Op�E{Zwp1f�)A�^1��E����lÉ�$>�S��@���S L\�0�
0Z�LX
�y��9�= �o��^5�6G�~ˎ�=�S�8�?9�3���dC��cC�m�'�ax�bǢ0���a����Q��ԧ��=Y�y�DNq�֍�3����E��yrd�Q�L�BD�3in=;�JI��'G�z��
i"���#+>$:fe��x��5 �9��5����-��֦C�ɼ6�.u`�X�s�p���N-+�zC�)� �EPG��<\�T��f��"`v��`�"O�eCe�./Apy�5��Yt:E�"O�0����^HqZ�(ɦ2�h��HRH<6�C�s(QH�̗4Ք|
�l�H����>�U��)r���"��N�fd���G�<���)G`(S�H�y��иs	V?��{"�O8"=yRɏ�w�h��Z�H�t@`�lHg8��&���e��#� I8�iDIkX�2D$}��'�V� �Z|��䍆M�x��d7�S�d#�&�*-ғ��"�0C�-�
�y��@�v�HR! �n��O�۴DEz���'V��EHI���1�ԭKM�i�'o��s����~3�EaaO���q�O����K9N�T�ٸ�n-�ՈQ�.���V�O�2�胑j���c s���"O
�ɔ%�f���"����_��(O�=��r~�%�r�V$Z�����kꜰ��n� l�a F�`Z���/dC��ȓi�L-����
#
|Yg�A�R
���_/>X��а7�ư8����d��ͅ�cEtx`s)�`OV-²i۠[�d�ȓ,�X=t`J�]�x�E�G��,�ȓ\Q�$�G!��K7r�Q��Y�m��+�~x#di.��-�RI߂����=�tpw�D�3�&�k�cPdc�	�ȓK�(|)c�8uQ������;xl��ȓ\�N�7b�o��y�s��55�-�ȓk���#�%A��rh)0�����Un@�%%��h�@�.v�� ��m@�ď�>G#Z���	I�����ȓY����Z5/.�h � C(` ̵��r�J�����| iP����^���;���ڣ�+q6DD��>B2��ȓb��HB��?��E���H�V���ȓD��"���;y)�h����.���>����?m��$Z�������^�X!�^�<1k	�'=���@��,V��@0�)xD�ӈ}R�Q�Q�P�'O��!�͞�{�!8`.��)�'#�-C&��9h�x�XǠ�.E��'�ι��D���#�jJ���(��'�����A9��!�uKE��>e�'��@�&��9t��J�gخvW�H
�'�L@��2�^��&[�oK$��'��4!�˘A���x�噠c�`,��'H���3��5�1IE�P&�h�'��IJ�I҆����/ t��'Ԧؚe��������Պ(�Y ˓�(O� "3hf���a�Q�=)9X�"O\ũvj�,5N�((�!�22�
��	T����=�q�Q���h�P�P�ޖ�!�D�"	�PȠ�f:(\zL �#ѐOk!��	id���h�`?�u��Et���Di�&�8"��)�cV��b��ؒ�"O� �!��N�$�xRG� W��E{�"OjuP�gäY����e�K4��"Od���]oPTG��*�Id�O�=E��(�n�~)æ�T!6o��5�ރ�yb#�.#���bN�,�d\�u͙ ���BX���f��1\5ƌI 	!��H���?�OR�+?�)�� �t%OH�V�$�ȓ@t{Ee߭_nĐD�Ǉh���,��J�>yŀ,��
UN2�����0�%O����i�ࠊmY$Q��9�앰1�.�,M$���}��4��S�? ������,:�^����41\lM�"O0�(҉
	��J�N9
�`��"O��(G"Z#-�Rlb��@���2�"O���� ��$�	�R,xT"O�CUf�+���j�EǾh�\@�7"On$�g'�4r�ȥ�Q#Q��j|"O^IiDa�6�����W�ܖ�$"O�pX2�C�.������v9��"O��Y����*^��0���Z�""O�MpTj�=}�I`�/�2�-�"O愨��L�>�$x�,Z��Q�Q"O6I�Tk�!5��\�Q�J'����"OK�Am L���.��1�&�y�ȅ�&��cl@
WA*�pe��yb�\����M]�@��|Z�,�yB�t��S�OX�=А�He��yd�mH�"+L�%D�ȓ֯���y�BW�S;�+Vg&��r�,��y�OT��<Õh�8'����MF��yb�4�`��E����f8p�Y�y"�?3�V ��nK(/�n]�R��-�y��9�Q�č�+��(Q1
 �yr�T�n&�$C��G��<,�S��,�y2�Y�B��$��\!c�pc�0�y�BH�G�r0Z񄍬&��L�"��6�y"� 6hZV�����$־-����yr�9J�b�Sbf��j��E#+�yb&��<�\�z���8�b��*�5�yBfF,%|�9�Ͼr���y�*�&a��I͆!w�eza"Q�y�hP�1Čȇg��.�4]� �R��y�iј!�0���gΎ"	� C G5�y�%pz!qC�� ��a�����y�h߿yi M�@b_�
R�(���V��y��_VC������-s���eL���yR�^%�D\��eT���$�G��y�AICyl=�ga��LO�Ԩ�a(�y���.5opmi�K�jI ��ӆ�y���
�dJ���[찈PMУ�y"@��^E��IA#jԬ!��V"�0?!��P�}"�Z3@>v�>��%�ֹm|8���Y�<AV�6d���*%��9J���"v�0T����K�3ʄSD$�=+z��<D�<�S˗bu���U�\�>G�H]!��,:��ӊ�Rg��<Z^ʍ�"OLU@o����vM]�3�u0�"O�5�'���n2�Qc�=M�а 0"O�u(%�ʷ(d,$�lD�G�K�*O:��u�w������i�����'��\�.�����"X���8�'+��s e^c��� ���,T�� y	�'�ܡ�C�#m�8)�o�Yd29��'4��I@�/F}��R%ͦec�'9IY��f�h�ѣ�
�x��'���ˤgޣmlh�
�JY��'�h����^9���6^�w
�X�'��yvc[\�sf!���n�r�'�8��&���9���{�'4���/ŏj\�ď�V�Ei�'��Ș� 7<~h�yc�L<K�A�
�'j�:���#=�b�zS#_#<q0 �'G�a����\�dMysEϨ4'^��	�'*��`���Wт�qB��!�^�Q	�'��m�i΀B�<U�$9!�hi���� ^aR���"�Zɀ0H�:Ф�SF"O�tXu��nB� X���X���0"Ob"V%�$h8�8tF+{�\�e"O�Ԛpa��k5N� ��{w�iSU"Op2��Ϫ=쬰2 k\�P}��!�"On�'bƌ;�b���;cj,4*�'����烶��U"$�6{��e��'yp�E��%o��RM�z�$z�'?��уO�3�t��W�BKV P�'���Zĉ
(Î%#�oK��	�'���[�K�x�� �w��8<��`�'<1�f�m�v��@�L�pH 
�'0L|�%N�q�\Qp�F0`z�j
�'��3�ŏ���pу�x�r��'�$k���lW\mP��h��x+�'F
@;�e){B�1{6��Zs��<��I�=�(d�s�Ȯid}��b�<��j�31�Z�ʠe��f �:��@A�<9E� �X���q�%��r �]�4��B�<Ɂ�ԯ1�R�KRǛ�K�pQ�CM\[�<	P*N�x�lQ�V�X�cH1SAF�I�<��H.P�([5b�<p�L�SN�|�<�'G(x���0�Ð/��+v��=jsv�&�;V�}�g�䎛O,b�bv����[�!�ēL:I�CͱK�L5 ��S- f�Ӑӥ{4���J��}�����#��d� ��b����I�W��T��¥�6��'�)�ĸ4��Š7";wPM��'\,��@	=E4ep�DP<aR��L�`�H�}Ȱ�QE�O����!D�S���y�aIt�fQ�'4��Xd�2)N ���=���c�vDB�1��p�G:�3�d�,U^�$
���g����D$�@��֫,��mS�HH�)Q�I���4i��M2�J5��l�B�>�O ��j�&�ԇ�	y�����'L�8b��Q@+���[�T�c/B�F����䍦r��ҧi1D��"ů
_��Qb� ϼKPνi�K3}�D��}���+s('P��?�)���, �5�@͌f$����+.D��[%�hP�0�fi�Q֎��ǐ86Vh4�.ODQ2/������-��'eN��V�*l�Nh�ēD����r#P��h�Fi�^0s�Ύ�.2(�	!e,�O�(; "u�0L�e�ض`�\�e�'�4D�E�X�a�(�$���Ҙ?ǖx¢�6��C�	 g,"�Avf�Co�(���Y\�lB�I�SF��R���F��a4�V�sBB䉄uΪ!7iF�4�8=��-h8B���ƭ���]eZ'DOv-B�I'5�6Y�r!�8-��x��G^9
��C�I�~)*�*T�ܼ�����(YB�I�|�`	����=��@ЪV��C䉖����!o�k�������"������#��a��46��Z�AR8@VD��eU�=����x�.�0�+�j�V�A�Ę1���Ez���NR������ �J"��ɚթ��~�������)AP�˒���S�ݱ��[�b��F*��3[%��h)�i�M� `��O�Up��X��x�ĄS)S+���$�ɴj�Ty@��-��t&?����WN�� &�H�Π�� ���R��5#p]*V�'���JP�[��j1C@�85<)�I�`�I��iֲ2��C�O�O�ؓC�I���b�M/G�õ`��F�f� %-K�<ـ�:��"a�Kư�)�����`�tbE�#�bD tN�]j�':���;��	Y�νwZ*��@Oֆi8� ��Ik?��P*��N����皵2�E��+[&i��(��m�0t�i{n�t�d��b:��?�m�N8:v_
Ry8é T8ў���,��-�W��C�O���, 	Z���N��;KR|��'�P���<rԤՅ�I�'haIU���z�����d�e����VW���w.��KEhi@��'MMleh���% j��#�����p�Z]h���1D�� R�:�	�,���!��}�|\q�Eo?q�eت���E���9-t����V�Ɋ�ywF������� .�P�+W��>YՋב0`���!Ƙ�Q~�+v=�� rt��/3e��8Ձ�c�2㞘��哩���A�:`o��QI�.^ �E|�!_�[%B�zWL=�O�&���ٻDW��r�O�7����'?���3h\YA.4�wX>;�p�'���R��B��ݥO�>A����C�`tR��alj1H�?D�,؃��c3V|颢H����A$�<D���w��1Ndh!��p�i:E?�O�a*5�/�M�!#(01�0��^�YM^�:�HCz�<1���( 0�h�n#o��ZAD�;b�'��Ja$�;a�ɠ""3����e͚� �&���a�h�xe+�w<�EM�4FE���H:&������7L ks�T8��Sr)Lq�Ă)
~�~�I�d�d��FK�alt���:{���?9�Ϛ.z���E������ƃv�
 -T�x�x��ެj��D	k�^��S�*�0=�#Ō
�j�j�D7j[�au�A\y+aּEY��T�sq��cjـ>(t�� ���H���4X����a	��y"�T8T��l8���_N2@a	J$D�S-Oz-�P'/L�`H�?%��'\�ͻuZ��Sc��J�/�	�^=��Iw]�(�$��.e�>�Q�撦-	2!*ѫ�N>�RV��`o$a�Oh�,�����?)�B��,��P�Ng�(�!GJLO�'(�h($�C�<e�u�@�?i�a�j>�i¥���	VI���p���+��-x�'Z扠զ�4�%aD�{*��a$ZyB�S���=�TO�jq�\��#��7\셰5mU�!8�3(�*d��_�r���O��b�ŗgR�K�'[�l� ��뀼/��ɟm`��;����Z�e�����V�|��U��]H�,F~��SL3a�^C�I�T��	;��: ���K�
"�n-17 �1p�2�;"����8��ҟ�K�;!q��d�	ia�ia6����]a�j�q��x��Y�k`
�g�x���#�$�9BEԧ-<~��B�S��/R�!QHe���9}&� ����L(�W
I��j|Aq��oK���t�n3؆4�t�Hz��Zc�1[�~�(cKH�.��`�w�ۡ4���իǉ3�a{.ݝ,٘QE����xIR`���'K�
w�\8?S��j��"~���$��p�ʭ��e§n���A�	�jT��"�W#3�!�dȫ	�fm�s�#WQ@���`J�ya��� k�4=��"��(:��g�*
�jy�c��$olމ򅇂�2#<\�Bi�IK�as�-D���E�7
|�Y�Qʙ�Q��	(ʑ{X.H� g����zuX������"�I���+�'��h	b/����ԛ�FO�Y"�\3
�zP��Q�E�mK�e���592�Chѭ?V �!�@�?��hã��횣E�0az�䏴6M�h��G�6L��j���	��'��=�:��qc�[)�:%Z&H]0d( �s��S"D蕣8T[8E��c��h 
B�I �bEX��u2�蠣'Ae$)�+� #zd9�я
=�`
��zm`�B&����[�d��~,�:P��{7*��.�j�<����%�H=C�Ax��	����m4�9
U�tZy���m1�ɬ;Os��u,��T\1O��W�'��f턍~׬��p�'¨����7��Iҏ��Hs�4₨T�"�5 ���s�ɳTg�#/�@�rQ"ق�����&G�Х�D�D�+���#�&ω)��O��aEI�����ˈRj=�WdMVbm�􈛐f��`k��!, �3�k�>B�	,7���c���6=�]	�cΩC6Z�jh�eW�H�c�QB=��2�6���k���2�j@@C5��d	e ��>o<�+"OĈd. �<�9UN{��3�J�O lɁ㚑P��쀗G�?A��?i��& ���H�.R�ze�(AR�f�'	0=v&S@yB$L�5���OD�`�O�$� �(({�a�� �
0����Uܘ9�@L��[x�`!P�>�x�-�2�6˓HG��j�6d�.ô�6���{�,9QbGŶEy��J�'�;Az��ȓ}���q$��150����A�c������F��sC#�."��?����憘\F�Oڀb�/�"ou��:U����HC�'� |�f�kH9���[�/��Y6k�Ojx�q��=��.1������'�h�Waϩ����C���U��1
����E<�0O���(�H�Z�*Ƙ|����Qfa[��՚1"O�(�g�+h�R�h1F��axlʣy�0��"`V-��)��<�󆁧W�X�4NTR̀�qL�r�<�(CD2�lP,�8��m�p���<QtH��+@�?\O����: 䱫3�)��\94�'�B%8�ˢD^A��o��������9>���7�y
� ����"Y.e���0�/�BTjC��"Aj����3^�Q>�8��&Ҍ��2��<FO.D�HC�*6w���!�`�(�0TI4v�H#wn���S��y���h6���̻X2�TI����y��`k���"+��D�TX�bg���y���(�l�z$	�e�����?�X��&JO�r�|(��)�O���e ;$'F7-�,n�HP��էa��!i�X!��)l�>pz֢��{�� !��ދ/0��x�a���q�>�;�$G#xb��󊑞<�$D�t�&D�����+��0�K�3eN�4�$D�Ы�*y�4������lL� D��z2*��c�hHbPE�E`I�A!D�P�䪛�N��I��+#r�S�A?D�0����hd)Q���B�`DЋ?D����ě:�����!��I�^A�M=D����fJ:���a�� (�h�R��=D�p"�*$x-�p	�t����G�8D���蜁b��H�����(,�I4D�lC�˄";%��;`)��m:p�5o(D�9���u�nH���I�1�<��&D�\9U�A'W(8ɠ-8 ,��p"%D���S��qP�pj��_��� c/D�4#P����3FEޚV=ָ�ӄ0D��bq'R��4�j A��1�����.D���R�]�4<�	qKP+EMF�I��,D���@�L�Z$,i�&��\�4�K*D�dHd眩.����HM:qYڴX�2D��zs��'�6�yiL�̭�*D�x+��D�"�X��P"��9�(D�ı4���;�L$ �3�C#D��(�:���MK8e�@|Y@�2D�آ�E��T��"�I)E|���0T��2�'�~��ī�W+"���;�"O�Ļ@)֍-.�9�֢ߢ?��5Ap"OF�ɣ�=� 	V�Ţ'piؓ"O$�����qj����D�i�%�"O<0p� -��|��4vF��f 0D����B�� 	t
2%^�9�5��L.D�����T�NS��HDk�/ux1G�/D�1uč�-n� fĂ'l��+d&+D��[F���$�4p
�d.E�IS�(D���(D-HY^����'٫�$=D�@�@�]:$n�}�Kω��1�%D��Q�̛+�^4�W��c��ɸ��"D��Se�?U��|�SG�2��°�>D��@��/)�d	�+\&��9p/?D�d�SƏ��|E1�Ț
�fC�B=D�����I�_��|!�c۬=�Bx�&
?D��"�� �J��֡
��!!u,(D��8�I8b�.�S@�����b�y"�Ƕf
�=��@E� �\peN��yB�ұ	�l���$�h�,��y��3�BY���̂�Nb$�8�yb���*�[�d�۠9�t���yB&�:"Iw�UK���d�M<�yr)�> 5c4AL��s��	�yr�P�t`���1,� 8ӬPR3����y2��O.�se΁0����"K��yR�=KS�u�)�*-�5
����y�ӄB�]B�I�g�D;Ņ��yb뛭8��c��Ņe����W��yr��$��c���%��Rtc�y�[�mLf�Ȗ�~��)�b�Ҩ�y��ۆ8��)�J٤k�Z��%-�?�y
� ����Lj9�(igf�!�B�1f"O&�
ֈ�:�
$y�c� 7n�aA"O��i����@�x� L�<�t�q"OJt��cXXsvO�9#���"Of�+��nqy�/Z :b��b"O�	Ca%�"f�
9;�N�c�B�6"OY�P�@�On��s�K<!�^�8�"O�Q�r��"B�^ 20K�,@�A�"O���L�T`(�*�Y���D"Ov̈ �)C�U�wJ�$�"O" ���A���Y�`=4 0#"O�ɠ���-h)"���n�7+)���"O�����ƙ��q;,�"!ʀ:�"O� '#�8	�,9S�l��CΉ��"O��"D����Y�3�
�p��"O؁J��ʟ,�����d`�b�"O&D0C $q�����bD�*۴`�"O0i0�'G�Pj0��!@�a�b@R@"Ol��T`ATʰ-������E"7|!�Y�**�SR/�M�x�E�J56!�Y�/�t�S˙K�D�0�,2J!�$ުD@��� 	�41���;t-˲K�!�䞿W��\Ȑ�T���5� ��5z�!���;��`j$#�+<�p󵄊�>�!򄃾I㪹�2����ԃE�N5]!�D��E�7%ң�a{R âq<!���"�9�`˙G�`4ó�]����1�|��B�\���rRhz@l�6jb����"-D<�ēZ�08B���[�MJ���~�H��sJA!a��U�9�O�8)3�C/)4d�F픧M������'��ĠՊ�4P�:��Z�P���ܙ��|8��M�-���B��=D����ʛ nT)�I�'?� �F'}r&K*j`@���_x�?�YT�P;	�j=�$!�N�v��G�'D�Թ1@�XO�J��"{R�V�_�	��-O�p��Z�����g��I��i�)ha�asoH?:�xi�Uڪ�ɕ&��#I��ۄ���X��1Ȅ�̛Zf��Z2���̰>)p�SMbp��PfĬQsV��k[8����B��^�	5�l}r/�57��#��N�]&Z�`��!�y2-[���y�9 z �aC���p������mG��e��RI1�R�04�+�bć�y�ՖE�R-
�F!h涍Z�&ΉTuq��<��E; 8�>�O�=����A�
]�ӭӱ<."�ѱO�9@CP
R�85B��ȅh=�} ��]<&5�%	ӣ��>!�ȐY����	�C�L���k�Vx����I B�H��'�b!ص�C�L�� ���L1H�0	�'���4B�9��3 FT�W�jQ��'�L�" �u|:)S /ۀ@��
�'��0��-��|����+V<���'o��Cr�6�z$�O��V&�0�'�JA�8�����@0��$:�'��`��d ^� ����}K&��
�'�N 䂌=i�F��#��@S�$)
�'�zx�L�QעIS`��=e*p	�=g.x!�g��Q�E��x�~�9sG�z��� �"O���� "���-E>v��9鉱qÌ�)�.PQ�O���Gn�'($�rV��>C�`�	��-�v��._�$Չ4j�-�@�2A��A,lXQ��K����(4}���d��?94��8��a #f��A�4�[@�'���JAԳe��D��������0�-�8>��i��
��~�e 0h;������k���Z�����L����0H,2n�rK�[V(��&��%�"��Sⓤ�2�&3\��m� *
�s��j�G�0r�6�"O���@�Ĺi:T�\��5J�,}�����m�ҠϪT��Q�#e4/�Y�H����7�l�ա��������I!�%��'#�9��FW�T�Y���r׾�1���&z\k�XvYA��Z�-�<�Ҋ��S�? &�+���� �`��F�.f����K��Q� ��q������$��9uN}3���i 3e���~Rjp��eCpfi��<�@�E0���;�eZ�����`�OX��n\�V��a���~J|����	�$�`�	7:X���[�E����!�Q�C\C��\�L�"Q#ƗXx�hRq���`|�<��'3�܂��b-���A�|#n��I>��7�p!)pĉ�m������Ԑ;�Z�*�'�^�`�ד@2҆�J2,�D8Å�;LH�H�Ń!n��(Ӳ�AܓFT��|jt'E!�$��u��2'`\��j��O�� �1��rF�$��		/G��`��6PS���Qh!�$W�t0߅tJ��`<!k�D��8�*��sBĿ��)�'v��:�*Q�W�	�]!���cRFUˢLF3}����S<A4
̈́ȓw&̠�i�� ���ܻW��(����V�� hw�i5DM�r�b�|r�ύmCZ��
�'��H�ĩ� ���2�8С�(��
0�4���N�^�$�0��w�r�)#�� %�� jò ��(�	�'�vVʎ��-B�LԠ�y��iD!(�lH*\�(<�$����U��M@���(R���(�$bdda����5n�RXD"S�g�����O�b��Ӈ69FT"W�yN*0�n�2���)r�b�#��(u!az��I�hT�S���|4��;�FK?������0F��.���>9���x�n%A2-އ�|fДR��)�"�)�!��6z*0q`(��&���,}��H�W�䳠�S�4��=�7b��K�Ox�C�w5�+�@�m����&����@�E0�=K��G�$9��E��;ayu��&�� Wd\��<V^��N���VdF4~�q��&J�":9Ƞ(ˍR�Vܘ�����O��@D���*;Ruc!#>��
��7�0�k�cF�.�1+E��y?i�A^�9V-@��9LO�y���d�n���-3ox`��]���U(ǦF�ؔ���Rw�'[d���B	�-6ڔ�$��	HZ5�w;��b�6D��k#�N�!}�QsA�N-U������84��ʓ:�L�&�J�U����%_�	��yg�߾b�,"�C?]�|ҥaP �xr��?`|�XTmۼ]|Ј3�a՘S���X���GӶ���'-h��#|r�.>5��1@IW.5Mr�ie���p<9F��%\��<�M<9�i;,�<��[eı�qf�@�<��nQ�����1G��V�)$�@�<�v��J�n�Q%�
0�&�POCyr�*� ��I�O�%1�iǙQ
L���0���$;b;p��	� P5����F�t�ڴ�q����e�r���;.��cn
dg�$Eyb�f�|��ՠ]G�O6�*��^*E���@/ҁ\-xQz�'<Q)�
T��d���P�v��q��q�T= Q�I���)�矌�GLϻS�����NO-�Ni��&%D�X�"��}ĝiV��#]��3�Ǡ��sP�M�t:
���'y,zPΟ�=���Zr�֥W1���[�P���ҜH�(�ԋޭ::����Z3q- ��v/D��rWbʀp* [Ҋ�0�.a{'�1ʓv����Ks/$#|J���K��*fn��h��7���ybHC!f�jq*RU�s�x(�c 9�0R뗥'\�)O�"~�Ɏm�����6Fƌ�ȄoM:U��B�	�~���"unVF��U��c��O���I�r��,��l�>Raz�!�	��ڳ��>#�&��ѯ�9ܰ>A#�q�0�3A�@� 䀧� /,��ò%>x�!�D�K����ڼ'} 3rў�Y��"p�o�`��aH�|����hب"E�B�	h1�ܑR�g�r�Z$ԁKX�B䉅OvR]�u�!��]j� R9�#=i �B':�,�}��/� �'�0T,j�n�Y�<	@�
� ���!��E$ \@�`�� %��#�iCNɧ���BX�=������Տ|����n��yZy��M�h��9S����NQ�$R 牔<��U�[�@�r�m|@1R�nͥ`�Ne[�\�X�l(��I�g���C7<�=�JV5f�4Cd��{�`�S%�#D��Ӡ�ҿB��ɸD`DfV�	��<�@�ب�g�'|���|2�˵	V����)��EM�y�<a���e��������b��S>�r	:��
+}�ӧ���� �)JS
&�ʡA�d0N1Ba"OJ�����?BhH�E�q9p3P=O��C���V��
ד��5镄!z��<QN�#����	
r�R(���	o����7o��*z�/�.B��)-D�P�l��3�0	� �T&q���!�/�~�֨X�rb>�|*��d��Qa�wl��X��C�<�0�_�
 F<sC��8��ѣ�9����"�140^ӧ���d�0�n�sҦ��b�}���Ϝ@{!�DA-6p����j�;kh�qf�(��$HK��}��&V��p=9p�PF���2������H�e8�ڳ�أc�
l7'x	����ol��X��ۼ�*B�I�^�ً�]��,Q�i��$�B#=�4j̯y��}"c�<R���p���kB��H�,�h�<�"��}����SB�U���E �e�<)@F��.��3�ܝ�d�ۢ��z�<�4�P�<�|�`�(rM��a�|�<q�l�D$��r��-5���j�E�<��h�.న��HD��ȉ��K�<y�
X#YgL�(5K���`J�KY�<1R�Ϭ�!�@�ku��9��Y�<A��P�H5	5$�~�Vd��	�<!�L�|�z�˘�m9 ��.��<�5�M>j��S�	w��+��x�<ё�V�~II�"ǆAB&�˱#Vy�<�0m�"t=��^�#�̼�3�]w�<qb��Ҵ��oł1�ʔ���X�<1�IA l[GL�y^`��fMZ�<�у�I�.�'�W�f�����(WR�<!�Tg�j�H�-خ]-h(
G�J�<YO�G2��A��¨	��!a�͏o�<�� \�"�u���]˘%��)�n�<Q��N�dᜫ�v΁����'��q�m_|�vdѫ XpQ�'�X����F����+�U�ru�
�'�B�����'�����.�e�d}��fʈj��t�(-�w�>y����ȓ[��"�>J��Q�?�d�ȓ%��=!A#��l�@A�B�2t�}�ȓ/�>�s�>1�D5��;�b��ȓ9GR%F�E�/t�8LV�.CrԄ��ڱEy��AP�g�]�n���c�X�SP�NzH`��Q�g�|���&�x�����YM�,���C�P�,���#�"E�G�W�Jl� �E�o{�I�ȓ-&� {f��B֨�2f�st �ȓ����`H>3����-ْN�&���J���[%ˈ���08��bl,��ȓ^����@�y�tC��X�^"E�����>ŃR��0Px��6 2jE`��͌i��$��w��AB�<�>!���>E��aXT��d�!Q�&
�<Y�jZE$�O?����A��"�%�p�]�G�\=B��I��������蟌�K�S
N�nq��+Ȥb�����~~"eIĸ�&�g�!Ñ	E�{��c?��6���ޔ�Q��`��y��gD-�?A!�	D�&K�'N~D���q;��9wo
�*r��(Q[
x�F�3��IaCe>$�e�S�O�ҥ��E�%$��D̀�XeV5·	�~]qO�ᓰe^�X��::���ա�<Y��=�@j^,�a�4�W4|:|pAC��:R̚!�ĸ��I�(t�(�%c�	q>a��M��=�$�
�:8��D��~� A�P1��q�e�T���z@�Bt�ٕ�Ԑh��ܷ_���DY�D��Y!�n-}�����(�TG�?IS�E:�gP@�f�G�HtF��$��ȸ5�:�$<��<b�s3�Չ���*�l�#j��	+4��;E�9�X�CӢK
��ap����9�真�#���iz5z��9�T���[�O�8S+�{�r��<O�a��� 3�`-��\��D���O�V=:��G VL)9��̘`9�pbŃ�^xh-O�ӧzpj��|d��3� �@9A��!]�d���ɂ����;Q���
2���]�>-�0�%�Z����  vp���Ւ��Xb���8�}��J��Z�*���aJ%��Dؒ�0|Z�Ӯ#��d8`ʗ�M���3%/0�2"]�\j���Tua�t�&1T�ZA(ˊ@T�XZ����/V�l�cU(��^a��#�&�ԀXV�Nh���������'�0Q���Ol&T��v�v�z�#Y=O�e8I>q������Ou��#�E!ch�Qs I T�p{-O���1g-�O�T`d\�D�XS����'�AXt"O`eq�O܊K������ L�pı6"O�՘������D�#'=w�
J"Ov)���Ry훱kԥtH�*q"OR������[!Z��D��9rr��"O���Eܼ\$���Uv[��W"O���d����%3����F:[6!�ɂ7î,th�)J h�k(��~!��X$a��a��f�˦�޷e!�d�&u�u��oA�v2��#e��X!�d��d��#��yf�qQDϧH!��>��9�aΈ7� y�i�/U!�2(2@ر�t���cSH�zA!�Ĉ1U�`IJ4�5�����5z>!�$G�\��l�8��a6��!��5MY�l*�C��b7����!��B	���[ǀ�.�0Q��"Zh!�W�)В\�eN��r��Vc��y!��Y�}je�Bf��y��P�a@)'q!���E� !��KK�6��׊M9�!���:/DeRr';}����#�!�� 1,����
:A�Ѐ4Ψ+!�� 2p��7b
�.���E��Y"!�}jС$F�*ء����/7!!�D��-�ީ��À�Z~���퐜\�!�XP�
dI���(Ђ��!�G�zq!+]�m�����a�(�!��p$(a�b�È8�(�Ca�*Dr!�B�l���[c	��f�(,��>gT!�I����8�g�7�K��w��t��'cD=y�MK :Â�Fd�-vAd@�ʓlL�%���r�~M��Q>��l�ȓ7^>��r̃��ԡr�l��J[&���9�@�Ais�1S��
���'L�9{�� z�ְ�/E+l=r	�'x&�@ǥK-Sp q�pn��'4��R#�U��DTypHŎn]i��'t�;��Do��$!ܡk:��(�'D�[2͗�"m~X����O4:�8�'��,#j���	��ID��H�'����K�F����Q���9�"O�)i@�2Z��ң_�/ah�H�"O��mY� h�b, N�ecF"O�T�� �r��(ᄬ�<H&l$;�"O�Ma� �?r11��P�{�ZxJ�"O�Y���}�41�C��w�|8�6"O�$r�BA�bHc�B�qԨ��"O*����;Lva��F�/\i@%"O��A����2���)p��"O��[��wf>p)�I�)ϜZ�"O�@��>�jx �8F�� "O�s��%�iap�^T���{�"Oȱ��+�����X�>X5��"O ��cE�oF$�D]�J���t"O J�	��<q�d&>e.�F"Oz�s��K�f��cɜ<\�`8�"O� Vd
%%�"t��e�#��;�d�9F"O�O��z��ap��b����"O�b�ɎeB.H�Dю$���c�"O��;���."�*!���@1q���*7"O���r�ށ�n�
��\�q||��"O�43քV=$���Q��( 0��E"O�A�D=`��l�@<ر"Oppb��ЀC����e�Y�(њG"O�г�N��fZ�M���C�D�`P"O���v����`�s��y�$3 "O��2g�ׄ2��*���4ed,j�"O<��D!ՠJ V0�D��`d�T"O��(���<��y��CJ�`>���f"On<2���s�N�D�
2>�г"O@	�͆�q�>�j�(�=n��Xf"O����-�"r?N��H�1eA�"O��ǌV*3X$�p��|O�@��"O�ł��\�V3@Y��[bA���w"O�Љ"��'�0cD�=|'����"OU!��պZ����s"_&=ֱ�u"Ol��#��
<��6c�%�k"O���A��) ��{6�ԩ���t"O�٢Aޮ,�2��B�� ޞ���"O�`���ft�Jǁӥ
{:�"O�̲!�"V�cEV�L��"ODP�q�Hp@�IH3AY�/�.zt"O�с0U�vv\H95�WXq�"O�4	r�"�@�@�D�WJ�h%"O�\�d�����v��:R�Ȉ%"OF,
� [��Q�N d�aa"O,a���ۧwq$(�sV2B^��`�"O�U�B.N�mg������3lC�y"O�mZ�@n�����%J7|A��"OB�����N�;�گv*�A��"O橂Ĉ8�̄2e�?��[ "O�)��=o����%�*GjZ�A�"O� X�eR�}�����ы+r69�"O� �ԩ\�|�vD�sV�][�"O��UF^4N%�AA�o��L@�m��"O��� �E�����":.��"OTc fU� !`�b@�$�c� �$�yr��f��r�[�օ#B��
�'jLa�S�~���!���3_&0��'� �H�M.]w�U��o�1�����'�Xɓe�I%,��)�u�X0#� ���'~�1S���\ b]�@��!d����'�bX"��R�sa��� �M#~Bh�'��:wnF+�\�a�DQ���<��'�A���؞ #'c�� `- �'^n `�
ig�0���zp`Y��'|�1����ht�]����J�NA�	�'��@�i�9Z�R!���Bs����'�X1�	�_/�U���6ܔ��'i|x��N<:{Ƙ�B����b�"D���#�D=A�����Ӟ~9�e��,D����KҰI��`X�hQ�"n�kR�+D��#��F���H��I#\"�h)�)D��F.�p^`�`t�L�s���ҩ%D�$AD������U�s�<9a� D���%�B<:�
8���8����V�!�/3 $����(�0�u���!�$ךN�����Q*���Į�d_!��T�&�i�H��@�<�|q�"O.�y��ݘ}�΄���@��@�V"O� �a{ -F$~;Z��7,�q8C"Op\3 �/T9V��$ʐ"@�[P"Oʔ�c끌F$���Ϋr�1�u"Oj�H���V>��ڵ"5Ԭ�`B"O,��A�U�M`� �f� �1�"O|@��M�2���4�K�k�`��"OZ4�$�y�)2�D*,�c"O�  ���9�j��ԣ��ڜq�"O�\�d�Z}uPA��ВA�N��r"O �dkC.&a��;B�[�[ߪq"O0|J4 ]�p�!��$j����"OXɃ�G��m�n �᠘;3!hMQ�"O�����x�-��l�Y4"ONp� %(�.	�d�É$�R$"O`�ف�(q�r��
Mp�X��"O����ۗ5%|0"�/	#���	"O�Ŋ���?7��+�P�*�� ��"O�)��)�%+C1Y����Q"O
�iFn��;�p�թ	%L��4 �"O�({�j iD�����ˈ8�f�x�"O(Ț�@inܜ�F	8t� T"O�M���ۖ>��@i�j�
Ah��Q"O�D��ۻvBp䑁�!+Lp�9�"O��Ħ�tq�W�֘]Cm��"Of=xՈ��a�t�aDmRP�=��"Od��E�� ���t��X�ҍ��"OFX��AG��^�K
Ժ\ǌpá"OP����A�i��9�i)s����r"O@:F�^(�@k!Iw���T"O܄Ib���Gำ���#� ���"O�u���]��lA�iک^��=(�"O�A2o�2p���SN�9U�^,Y�"O.e��eP(�]���Wb�e�`"O&9h��ͷz��̈��O-6*��"O�������S��L�S�^�e$p�
�"O�A��89fA�1>�����"OD��J
j�02�N=I;�}j�"O!���L�I^b�P2�Y�f�aE"O�<ZC,A�g�2ayu����r�"O����d��)،M�׈Y:i��Pi�"O^��ņ^�=�B=�&څ�:��U"O�ũ4l�[�͹�f[",y��C"Olq�Ӧ��[Im��f��s�� 5"O�z!��I�lh���!Bn�p��"O�=�*�FhH�cʼ]Z�`7"O�˷jz�3�Eòh���*6"O�`�ė%*�)�ď_�\�	�"O�H��)��`�:%�� 8ߌ<*�"O��7��9/Kx�#7�-d��9Y&"Oxu	`���v%`�U1����r"O�j�&G�dqH�eN�h��"Ox���܃v#"Q���ÿ��h �"Oґ��(�B�����a�Б""O��QÁe���KgN��Z�B�"O@t{g�L�8�qڔ�˻?kz �"OZ,��#�� ��I�Z��h4��"O�)
�� ig}s��^�j����"Oh�3��J�|�*��-{��p"O:	�p!��q�ڨ8���>~s�,��"O�q�%�;"�����_���j�*O��Ŋ�+VZ��.@k0	R�'�H��Z�3�~�  !A�&�)�'�����GH����2�]�% ��8�'�@-�F�Y	���3򨞜$i�u��� ��O@�?�\mZ���t<B�a�"Oȭ�ټ]���BO®>�Xձ7"O�yj�B/u�H�"���)����"O��L*OMԢ���9�Z� �"OE��范;�L�K�(K�E��� W"O�SC�Ue�� h�K� ��"Op����+b��I�G��N��B"O��R��Є'��x��&;����"O
=SP��I@J��`%T=L���"O@x���K�b|�*qiT':�����"O2,��爯��x�Q�r��`""O�m@��� n�yx�R3%Vp[7"O�hC�x ��M�>�� "O��   ��   �  w  �  �  *  P5  �@  �K  W  �b  m  �u  P|  9�  �  c�  ��  �  O�  ��  �  <�  ��  �  {�  ��  6�  ��  ��  (�  x�  ^�  ��  X � � � <' ". �5 �; B �G  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����iX���XVp���#��I�� @L*D�<�ޠ�B�"�ͷ^���1<D�<;Uc��*�"bi_OLa�'y1Oz��#�~����{���"O�@��_4#.]dᎺ)�8��"Ob���/�k2��Y��A��(zR"O\���1?��1E^�n����E"O&�2A�
��1��kI5��A[�"O��p"��kpRur�/�8�����'�!�ĞeH����d� 9���g[�l�!�Ā�iޤ<)�eϫY�f��D�	lq!�Ta�dZFÅ;;�T{�mI)�<F{ʟ&%����a���qa�(��s"Oڌ(3��Q,I��iH56�pp`"Od� 6���#� 	P�9x�C&"O��kE Z1Px8� �B��$A�"Ö��?b� �E	�7|�(��"OV�" ՞����/@�����"O4���U� ���ȁo��	�a�IU�O��̊����v	$<p���G����	�'�$`)&`*G+��K���A� 0��O4Dz���W8}�M9����
�"�Y�)Ϊ/!���T�|�&GҚ#i��ч�̑|!��vr����e�()�����*_�Q�<�'�Q>]��F<`���Qr�A	h"�G<D�X@ǋ@�^����c
M��5"�>�N>	�O'����Q�g  Q��_6��h�	�'���h�IR(b�� �N"��q*OF��e؞h��hܐ!���ӆ(�Ľ�H&�pn�/?z����
�0�m�"_;I`R�	K��d�Tˊ$�N$�-O�Mj1�p� ��J�F#}���P�0�����ɴQG�zQd�~�<�	��)�Ĺ��c^��Z�#}�<T�=�`0ȃ8(�ɗ�UO�<��*[��p�[�&P�N�^iQ�M�<���j��D�G���L0K�<9U�q D�����C����#��S�!�$_6w)�l�'�j9���ɑ�7�!�DB8N�:0� ��+
��h�4�\�&�!�����-���Ѝq|j���Ȧ!�dNT��)¦pc�$�팪b�!�dփ?�5`���$GV��8��Mhf�F{���'��%��cK���\�↙����2�'[����d��5��b'�_��	��O���¾U�r�S�`��ޕ
��R�>!�;n�r�)�g�:��鰂f\�#!�"18�5��8hY�m�D��W.!�DG�OQ�I;v.ӏJ¤bs#�6!���
,5$����V�UI2�㖂��o�!�G ��Y��C�H�i���W�A�!�d�y�]+/��k>��B��~!�$���,+�d�%*�A1��8	i!�$��d&Z��߰qX�t�	��!�d[�lQ
}�S��^�8�Q�jU��!�D'Q�(�:C��>A�%1�(�Y�!�D·���C��q��y�%ک<ڑ����)� F)�ő�<<B�2�-?�uP�"O�L1���;j��P�T)l��бi~C�I�F5&aP��e2̼x��{�@C䉥 L�Z�ʇjT�`����4�:C��;�.գ%�N�zv�ђ�3�(C�	;cDDT�*	�"9��K��57�C�6X����B���ؒ��cUbC�Ij�&�JRh�\�^���h���B�	�#WX�
uOT4(Sf�z��טU%$B�	�3���t	K1o$q
.?��B�	_�A�d�8y�T�6���_�B�I�k�੉a@�Xa:ѻ!��2ND�B�	�~��Q#��}8!�A�a��B�I�	ɖ�Kt�-D��0d�IT��B�	򒴲Q�n�i��I!l�
9��"O t3�CO�,0N�!́	-��PG"O�"1�֝6���R�l9"�|LU"O�pǬ�.��H 7���]^n��W"O4A�פÉA�, �5埶/����"O<���eh��aCY�f�2̑�"O��4�Y*���RN8n�l�""O�1��H)bt�\��a�ԆT��"OƜ��&S�}y���a˄x�\R"O�غD�	�m���3$ΚV�
�P"O��P��k$��"�F�$L�"O.=w	�'?�N��o��n�8Q��"Oj�a�*&��-:�
��0�"O����E�TU�i�R=Oߔ��"O���K*!.LṦ*�YmBy�s"O^��k�.6�FIBrOߪ2l�աc"O`5b�̢O������u�x�[�<���/1��)`k���M��A�W�<�G�wJ3cD�
���9C�G�<��^�6=jW
ߎi�vY�.�@�<Ѵ �)�j��e���ky�<�H�'e�D[�!�
G}��0�t�<���ۅ-�P�bA�������d�<�&/�9Gt`��0��(��yǤ�\�<�2�A���*�@��+/P����Z�<�b'�	Q���P�4v�zy�3m�m�<&���:��Қr�����f�<� @B��4�K��"�F�XQ,HH�<)�	�pX� ����P�<�dO�l�<q��ɡ73����I,$�4���C�d�<�����0�2��t��'+�����b�<���ϡ�������[۴���HZ�<���A�:� � �c,B:y��a�{�<�6*ւm71�iC�8^4�
x�<��%2Q"�1%�ͫ7�he�F��\�<1�d[�j���G�L0v~M�&JHC�<����?(�5�`gE�[��m;�/NY�<�'�A��zuG8y����hW\�<aEB:���q���
|���Qm�<y���;ith�@#�G�����\g�<A�!ץ;A^uC��Q�4�B$i�<��G�8n�H�I���i)�H�HL�<�f�"Y'��15F T(�t8�#�L�<�7LH�Z���S$@]�*6��X$�JF�<I�n�@y"Y�BNv��8��B�<����oc�(�af×f��s��@�<�fcן9�Dpv��2Tƹ��E��<�����a��}�D+k�P"�O@�<��$��m�tɣ@��N\�hr�XW�<q�L��P��P�K��z�ㆃS�<� �xڐ��h�%��IWdV����"Opt�˙�dy��X8��A�q"O��;�CĨy��V(Ӎq�48Y`"Oؘ�lU0K��Ma�S�~88��'"OJ�!���nD&m�G%��Q$�qBW�'�r�' ��'bb�'%��'.��'����(�0�l��\90�d��'�b�'�R�'��'��':B�'�ȂS*	�vN�|S��ǚ
��I �'���'���'���'��'���'ဌ��/0D	x��^�<z���'b��'���'Fr�'xb�'6r�'lRi�D�1I\��E(�2��iu�'K��'�r�'��'"�'�2�'E��B��KNy��`#[۞X���'@B�'���'X2�'h2�'���'+�H��	�!��9�g ?=��ep�'��'f��'>b�'���'���'ǰA�aCB%4<�(x�+bJ �Ѵ�'R�'��'u��'B�'��'AVI�C���6B��H��[��24�'���'u��'$��'���'���'� 0����)k�Ua���:���*��'#b�'B��'
b�'}��'�r�'-��Y�H���:S �_���C�'���'>��'B�'�2�'���������89�I�k�p����ǟ���ԟ��Iߟl�	ٟ`��ȟ���ş��C	˾s[*պ��PN�P}�vm۟�	���柬�I��,����M����?1"�����е�ѭLT$p1�.c�4�����E禡�6���}kfYR���	)�Tt�El4V'\�{Y���4���O��"��،G���(QD���sJ�O����THH7�;?��O4H��$����:�&e��S�Ϩ���$˘'��_�F���L�ZL@�t���`�JO,7��?@�1O��?������H7
�ر�[�Z[��Jr ���?���y�U�b>�qW�Ѧ1�w���$ȗ�D��Iv�V�9�͓�yR�Onu҉�4����גefT�u�W���r��>
�d�<9L>	Ӽi�x��y�A_���	�f�=2u��H0�OB4�'P��'(��>T�ƎJ���Q�lu�Ju��A~2�'&2�(��?�O&0��I?j�2Jܸl��p��E��Cj��	py�󧈟�� $k�h����a��p;aF�%����r�0?1��i%�O�	�=L�����0b~���f��4/��D�O����O�y��.j�<�����21�FfQ�Zǌ cD�I�U�V`�"�������4�"��O�D�O��D R�A�A�e]��G� rֆ�#)�6���JXb�'ib���'��]B�n����"Jǟ;�~�6¼>)��?)M>�|��lL�Vr���c��kX<i���L�fM��4w��	\��4�w�Of�O˓y::7��Ӣ-Q7lO9R��=S���?���?���|�/On-nړY���	%�ƙ�A�jg|��Њ��e�R����M����>y��?���^L��1�gì8ܒi�CS��]��k��M�O<x`u!U�������w$4L"��= ����� �2t��'��'}��'"�''�b	{����zOYk��=��� 1M�OV�D�OH�m�h)��Sʟ\�޴��_����weM�UM�����GP>ѺM>���?�'nڙ�ݴ���W"2�n	��ݒ4U~ �1��rd�UJ�I��?S�'��<�'�?	���?�2�
�0l��8�b�v��<9V�T��?!���Q˦ek���џ$�	���OP4;u`I.�:��T�������O>X�'�r�'ɧ�)@	@��ՁkF�)z��5ĝk� ��ݴbj��5?ͧ`���d
*��H�FM�A�C��8:�&�4}7tT"���?q���?��S�'��d�e��4~�ɉ���Ze�E�E�=1��ܟ�{�4��'#ꓨ?I�҃IKP��6m#2�P��V䄳�?��p�T�ش����<�I��'��S�/GT��"Ǖ=|��;�
Ga���Xyb�'?��'t2�'��P>����O�C���5��}�Y@�;�M�&V?�?����?	M~���cC��w �Ge��NA��:�=��e#E�'42�|������-��f7O�wC��f�d$�㈱Bh,��7O��4M��?y��;�Ĥ<���?Y��i%��y�M�
(R��)e(�u������IޟD�'��6�Џl*����O �dY�'Z|�(ŎJ�H#�X���M�.����2�O����O�O�(�p�̵S�*��3!��a~��+M�\WbB� ͢��
QO���R
ݟ\�g+�RG^��!��$wp���vo�ӟ��IΟ@�	ΟPD�d�'�:@!ҽP皱�w�Y�h��]ٕ�']�7�V5P���
���4��h
���-�Ū�m�&Z��,aG;O��D�O2��˖L�*6%?�����3J���/@�@���1m�	Q��T 	VM$��'��'c��'��'��Ǣ*a�����N@�	��_��:�4�:p���?����O�x1Yw'�&4�~��5�M K��>����?AH>�|�bI�$Q��PPƖ3nkր�b�]";��u��~~��Dd�����}�'b�,{�B&��2
L2�a�6`x\���@���P�i>	�'��7�բ=`��0@X�8Bv�β�(QQe�58��T���?��X�8��Ɵ��c|��qϊ$e����C�kn��݅d�����L���ڒf������� �����%��m�� ��!�h;Or���O@�D�OL���OB�?a�Ģ�#8֦=� @ak�@����֟,��ПHP�4zL��'�?��i�'��C��e>�h�w�A'��J"�|r�'z�O�F�&�i&��>r �x�����}�@��* ������Wbo�w�Oy�O�r�'��Z�%XLH��N�k��ȧ�%>\�(;kO�	��Mc�����B���?�,��u��1e������1?ڀ踄<O���_}}�'	�O�	�O�e�p��M�D(�Y�:�^,�E	\&�Z��1LB@X ˓�"�N�O
aIN>i�!֖`�.�肆ŉ*@���ڞ�?����?��?�|�(O�Mm�2	l�3"��@9�	(Eڰ	��������"�M���>a��M;*�j��- �A�C�]�>�`����?��k��M��O�$�E�:�O�౪�H�yP��hOh��'��I����I�����۟��	\���i�k"i%L�LC �� /�@6-�XL �$�O���7�	�OB9mz�)0�W�BJ�}"�Dʱl�4���+��D��f�)擞j<�m��<'
4H���0Z��d�lip��I�Jܠ��O��N>�*O�I�O��b	F�%����E߂ �����O �d�O����<Q��i��'[B�'{.AJ�A;�r���v\��4��Q}��'9R�|B-�,�����Y�$A�g㌯��d �r%*����Z1�
��_���*2���mJ�r*X�;B��}���d�O����O���>��[���M�|�0�Ɔ�3٪PZ�ş!�?���i�91�'	��hӢ�杢	��<Q#�a#�(換#���˟��I˟����ꦱ�u�㏞$�D�3xw����I�	q��Z�k�!��&���'���'r�'��'����AN����v�D�1q��\�P�ٴE�l��+O��D:�)�Ot<�CN�7Z[�x�`��[��]QdA}��'5��|����J�Aj(t/����Ã�V6��M@"H(\�X��@/�1 ��M�p�Iqyr.��V?�����Cb�Az�A�����'���'[�O�I)�M��J�
�?1Ƨ��7� �U$�'�ņ� ,��I-�M[�B&�>����?y��h�����˝ao����E9�1#��ћ�M+�O�H�̛��(�����Wh��ec�?%a���d��!��7m�O����OZ���OT�?���dĦC2ȳ�/��o[��CAU��d������ܴ?00�B/OF�my�	km���żhHh�!��<.��$������>�\o�Y~R�Z�z)n��U̓+b;~ k��+�����i?�K>�)O��$�O����O�liA.2�0$�e	�R7,���O���<Ⴒil�� �'!B�'哞䀣rƃ<N�Tt@MƧ8����ϟh�	z�)�sLˤC�!�4�ұKm�d�bD?��L�R�ݔ[�<U������P�`�|҅]HdH���رS�t�"
�3fR�'���'����_�\ ݴ{���Ȥ��+��D� ��,�ޙٵ���?I��d;���L}��'z	2����v\0����y���Y�УdLڦ��'�pigE��?��S�;W��~��ѭ���*�8"i}�T�'�r�'�R�'M��'�SvRR��c�ؔ�
ښ��o�yy�����h�	�$?M�Ƀ�M�;|� $ISE 	<�U A�]�	�,����?�H>�|Zs�[2�M��'�>I���0 ��
 U�S�
�'�,i�
Q�l;՞|�Z������z��B�Yr�@����XH~�٠�埬������Pyjӄ|
���O��D�O�!�� I!.dy����[�%�'$9�	���O��$>�$��`��=:VOI��*	�>[��	�vc��w`�|�Lb>E�'�'�L��i-Y�S�ע(���b��יK>��5�'�2�'#��'k�>睨Iln�itiɳl�5	ҍQ�>P��	��M�@톺�?�0���|���y��Cv�3t�W�fV�i�c ��y��'B�'� x ��iU�i��#a��?�:Tm�+`a�y��Q:`���0�E�+��'��I矀�	ş���ݟp�I2H�X�`,�E? ���M�+5�섗'�7�!h�T��?)J~R�_������<[ʶ���O�-!֘y�C_����͟ %�b>mb�%מ>H�a �MޕQ|@*0�1l��l���DP�)��e��'�'�削H�}C���R���*P�@�f�������؟�i>u�')x7m�D2\�$�p�j-R���k�5*��72��D�&���	����O@�4�X�B�M?��<+\4)P,0�\��Êe�
�98tå�� \�I~j�;r�4� �.*T�)�v�)̊$͓��?� �q�j��%Hb�\T3�@��D�O�o��"X�'Q��|Bg��u�ܜ!�i	�v�H3V�F v�'�R�����y������$d0wCHTZ&��F��NV3R/�]{w�O�O���?����?��#~|UfD�TK�h��ަx��$q��?1,Ov�o�.����	�����~�Ԅ��P�u0�Ϭɴ4*�����$�\}�'�|ʟp�Sr#�E��i�s�E�Ru<�P�$�827N@6�}�*��|Ji���$���#P"Dxbh���ş{��`s�ń��`���|�I�b>1�'��7�J F��Ҧ^��ċ<!�e�q��<�s�iU�OF��'��%�4~�L���(0vJ��O^!9"�'Wr)ײi���4n }BCܟp�S�? ��H2�@6f6���K�2,[�6Oʓ�?Q���?����?�����F���	aF��x�R��� J��m�OL"���ܟ$�Im�ܟP+����`ѣx�H�e)ު��q鎹�?�����S�'s�TL��4�y��CD>��:�H7ɶ�y4i��y��N�s"���	�G��'$�i>Y�I#J�,�c� �S�t�,�-���I���ϟ��'�H6D��z���O��āT�(��A�u�Zi����i��T�O����OR�Oޜ��ELs=�La�iӮUTl�r��ؙ�o��{dx�� �6��{a���۟<ӂ�/U��Շ[�~�T�da���0����h�I��G���'(��S�f�|1���7Fs��AG�' 6-̹0���D�O�o�I�Ӽ�dTVn�)��N�<�x@�h��<a���?���r��Sݴ��d�7>P:�O����2�L><N�<3gwm�#TY|�IIy�'���' �'��b��M+~�ao�#m���N �di�	��M FƇ�?q��?�O~b��{aL�8���5�\Y�Ҡ� 5��2�V���Iş�%�b>�ꆮ�3+��u�%t�Qk��I(�j�oZA~R�ʹ'�n������D��=�8�(�C�A��bX
73����Ov�D�O��4��lX�FE� ��"��X�!�ҼI�p ��D:[-2�dӂ�Hb�O���<�U@�&�4�kO$R˸�tHT�W��}��4��$�!J�|���O2Ғ�l���˰��0IZ�A-��ه�T�w��$�O����O���O��D1�S�T8����Y�0�rE�@�3OV���ʟD�	��M�H��|B�&j���|�f�*(�Reb# I�^ �%(��G*|g�'�������6�������	J�5�(�y��Y~�=����6PS��'���%�����'���'up�&m�UwXM�,ԗk˰�H#�'�R���4_[�l{.O��$�|���K	?��x���<��=Wb�S~)�>��?�K>�O9J���::����a��QS��D0^�0���i��i>]ˤ�O��O��2��Z&Aڠ��k�#hXҨP��O����OR��O1�
˓Oꛆ�O������Əi�a��B�_�6��',q�0�4;�O���"V���#�
8���b�����d�O:dZC�i���=p�H��f.��a���N�}ʂ�ߧ#K���ny��'�b�'�r�'��Z>}{�O�I��Bv�\�A���H��M��C�?����?�N~���x���w@j�H� �\?"x�c��l���y�'Or�|��D�B�o���?O8p���`�)E���r�;O>|p'/ۢ�~R�|�]��ן��D��FDA�Q.$"����S�	ޟH�IJy��x���H��<)�"_�u����(R�.��3������9J>���y���ş���_�	+*�ʵ��X7Bx�G
Qa�n���a	��M�F��t�_?i�� �,b��LO�*̠�DǸ^�p����?!��?9���h���d��b�6١�C�ȉ%N�:� ���Ϧ���@��������M���w���I�C�4u���0���	!�����'~R�'�r�$	������j�@-:3�);�����
�D�*���D�T�@�O,��|���?Q��?��腁�w���F�._��Ss�H;��æ��c,_ZyB�'��O����'s�z`3"��&���+8F���?�����Ş,��l�6F@:q��d�.ux�8慘!�MK�O�ԑP#ٗ�~Ҙ|�\�t��E )5��-H�/�dث5NB�l�	��	��iy��b���z7�O�$�DC��;�DQ��M	U#�@��O�nZC���I˟,�i�E��8���&��i�̥KŎ�Y.4aoI~�.+.E���'��'���E��%�a���?3&��  �<Y��?Q��?Q���?�����e!�����y?@��c卲Vr�'��}���0�:�J�D�ܦ�%�|��$G-9	t]� �]35g�T �>�I˟Ԕ'���;��i=��78x뎂+%�� �f��q��*େ1z�,��	P$�'��Iɟx��某�ɵH�(�d�>H2�Qhw��u��I�	͟��'0D7MX��b���O0��|��C��h�1D�C-pT���Yx~r�>����?�I>�Oc
ua�UG�1r�B=w�a�&�P'6�P��i����|
a覟�$��vkD"Axb��D�ł�U�ʟ �I����	��b>��'M67M�1/���a
�5<B���J:M�T�R2L�O��d�ɦa�?Q�R���	�1�h��'KB���Q�LzR�����@�Gæu�'Ӭ�s7�EܧAB����f�z��A���dΓ��D�Oj���OB�d�O��į|�Ul	�(�~�Y�LM�l�,: R"x��/�,2���'"����'�V6=��|+�aT+5Y��H"�8Im��`(�O��(���>e�7mj�����
Nc�}sԬ���Q��n�T�4"߳G���!�d�<y��?a"d��m6fT�w��� "��CÍ �?���?a���ߦ��c
ʟ���۟X��I�Q�	to�V�1�T͘G����	���z�	/;�J}�3aK�'z�\�5,P�F*�O@��En��R�@X�O~e��OTX��︵ DЛ9�|��A腗!2dX:��?���?A��h��NY����@�T�-�ƁQ%��s-��dT��*we�������M��w�V�@u��FD`5aW4X��1�'���'��O� �����@���!k�� .ZrK�R2��
D�~��+���<����?y��?A��?A�a��D	r�ۣ
�LY�d���\䦅�@�[yB�'��O?b�C� '�Q[eV�o��Աe�w�*��?���T��6+"5��E ��d�h9�4ua�&"8�剢y�tH�'��('�\�'�0�#C�^>�U95�/M��f�'3��'�����dP�r�43(�]��pw`Ѐ��e��(�gO�Z�H�
�5����d�o}R�'u�|FJi1g�4���A)�7:�̲Q(H����'��@@��?�������w,`Ÿ��
�a37wݬ���{�h�	ʟ��	��I����*��đYD�jj�pR�4�A��>�?���?I��i���ӟO��iu�T�Ox�Z����+�5 �\�4���+��&��O��4���gsӒ��J���U?s�Fi�Ã-"����d���Z��]�IKy�O`��'	rl�L�r�z�N�	WE�1' X�[��'��	��MKԪ��?����?9(����%i���´t��%x��a�B���2�O��D�OV�O��c�@�J�3zD)B��;X *�8v��H��(�'.?ͧp�r����[>6�Ajj�lm�ą-ED`�����?����?a�Ş��ݦI��#U&2#]//0L�4EG�0
8�AU�'�nbӾ�O��DF}��'9�ิ�!6G�ik�̑-ڠ��'9j�E�����֝76S�u�S�e�
IeT����6A"
��
*M�t�]yr�'��'i�'�"_>-X��"ղ� W&A,-��!;5EV��MC�%6���O�?e`���37�D�j	C���=����(�?����S�'SW!��4�y+QU�XQ��,o�z�xUł��y2��^>~�������O^����D��/��4z0�!V*��hv��O���O\�Y�v(�=�������v����O�'3�rS�KO��=e�	ߟ���f��mTЁu��7^��Y8g@�&�6�n�4�i�%�|2��O�%��I'����1\X�p#��u�����?���?Q��h��N\��� ����oE��7%�8({��$�y�U�H��`�	�M+H>��Ӽ�C��2���#�>}j$���<!���?��	�(\0�4�����$Y# �Ni�&�8tH'fY�}`��Ή�������O����O����O���ɸ0XR8�%9G%�0Ӱ�D�p�ʓu��fFE-"�'$r��$�'N|�ʁ��c���٠�\��4���>1��?�N>�|��C(�Ձca�'u�b�Sj 4��b���)���,x�T���g��O�ʓY�.��D�$V	(�#qB�H�8 ��?Q���?���|
,O��m�+V���Vz�@pa�j�ؕb�O��&�-�I��M����>)��?���Č(r���[�����'Â��N��M��O����7�z����w8�R+
=�2Ak�v�u��'�b�'���'��'B��`��ԶDG��g-J"�P�P��OL���O��o��xN��'T囖�|BBN�}�>U+�!%6\���p�
&�'�r����;zQ�曟�݃}C`�R�?(�qH�]S���PEFП���|rU���I̟���ݟ�g
�YW�q�$؏TM���ˉџT�IFy2�j�lı#��O0�d�OZ�'~��B`�U�c��J���0b�i�'��ꓐ?����S�$&@&G��#��
�7<���gN c�rW2����O��G��?��k#�$Q�$Z��q�ۿN���H$œ$�$�O��D�O���I�<V�i������
&w�x��C�\�Z,y���_m��'��7�+�	���d�O�Ps2`�*5�g�z!V!Xu�O����Md�7m>?A'�Ȅ@����xyB�Ϸt����D�3��4�`(J��yRW���I䟄��؟P�	��O�<�*�GJ�lDP���&/��a���j��(ɇ-�<A���Ou�7=�N� e�B�{���#�*A�}@f��O��d?��iȧK7�~�D۷�)a����ŵ#����GN`�\�B��=���/�$�<���?�@�Ư0�K�mЃ,�.�0ti�?�?��?����Dަ9�!�П���ΟS$ ^ 8'�M���j�b�å�p���Iȟ���]������q�N�c��=Q��2��p��=R�$�|��O0Z��,k`�u/�l�8E)�?ޘ���?����?���h���$�-�ݒ Ӹ\�f�	��^�)>��D���!Y��S̟��	&�M;��w.^��&��v+&��J�
��E�'���'�2a�E�F���ҩ�2u����Z7/�0\H��]�_w�Ab�͇h�pp'����D�'�b�'H��'���i�f-��A�&�ǥ.�ZAQ�[����4A'6q���?����?	����c*�/1�i��ɐZ��A��O~�D�O��O1�h�`F��p�\зf�5R=�2�`��=��6m�My�ΐ���������&;TlP̒�4  `��˧a|�iӌ�`@�O\�(gb<�$�*Fm�+���Z 0O��oE�����ܟ|�	�( �M�|���(�G�%]<�9#��7B�J�l�g~"������'�����4�K�D	�-�J��<	��?��?A��?و�̛�Jb0��MA�	���h��-V��'�".v�p�:�:�"�DA���'���ՁȞnIB��k�F#�t2LU^����t�i>]���R̦��'l5!
� Ru+��[H�(��P#�( E�X��7�?�D�2���<�|�i��5`��|$�Ȩ0�!&��MFxb |Ӕ��� �<���� �� (�#��+.�Ԩ@ǈ��I����O��D ��?5#����3�X��X-S�$I��3b����Ə ֦U�/O�	W6�~B�|BD�:6����@N�p�й�x�@o�n�*����h��8��B�76��7�E�D��d>���$CM}��'��	�#�u�H芁�.��X��'@��֗/��&���iݾ��ɬ<i���ls�q�I?N͊dHG��<�.O:���O����O��D�O��';Jr�Pg}������_�(��!�i�tp��'W2�'p�OU��}���RM�����'LYi3/ؔ%����Ol�O1�~�P�r���		poP��v�>}m<���m��I �	(lc0�ۗ�'�f]$�ԗ���'ށӗkľB&x�7O�P�,H���'���'�[��[�4m��/O��$��|�����6%pX��(�s��㟀y�O���Ot�O��A%Nێ �p��N�)g-�)斟��Ý$<t��l/��By���ܟD!�Ꙍ\nyX�o��a���ʵ�ݟ,��Ο\�I⟠E�$�'h�c�b��R���\�#Z7�'mv7��U�:�$�Or�mY�Ӽ��aG:6p1a�O�O1�D��<���?��K[x�{ڴ�����M��П6hՆ� �|i!T���a��� I#��<ͧ�?���?���?a�J�%E�`��T� �0��D��&��D���� ��(�	П�%?!���\xД�X�T�M�4$еNI*-R�O��d�O��O1���ۄ�2�%+��!�p�Kf�VjXt7m'?��^d��Iq�	nyBᕣ'�Pف�Q
��2� �5r�'/��'?�O��I��M�&�L�?����<6|]r���":�vE�w��?q׳im�O~��'�rQ�,�.�t���;��sڰyU��� s�Tm�j~�ԄA>��ӷ<��OH��	mv�qQO:6	t$֏��y��'�2�'�r�'M��i0���-�$�q�� 	�bВ��O��$�O� mZ�kF|�Sޟ�4��Vh����w�hГo[iE��H>���?�')nl��4��d��ƽ��ˈ5�\��Ν>c��������~�|�^�b>�I9�b=���R�o�m��	J!�"<y�i�.I���'4b�'��'��A̐$1Pe�W�Ճ;1^�!���x�Ij�)�g��a�\eYWE9.<��y ~NY�ЇD�MU�ؠ(O�����?�b�+��ݑ^�lqPB'ٛZ�V}�U,�����?����?I�Ş���æ�q1!����p�P�̳"�Q{WH%@$��ןT��4��'�����n�,�-���8gm�ԛ�O�	$����П�ZSO�ꦁ�'BlX���[�'A��h�4)����ŏjT��ϓ����O��D�Of���O����|�ጌ'E|b���H��L)��V;?��F�Ao2�'����'th7=�F��7	�	@��u:Ja�m�O0�%��Z/uO�7M`�4���H�r�Bs�-�2$Z�"y�H�d-G�4�+b��my�O\rNU�P/���A�7w���ʟK���'@r�'��	��MV�ջ��d�O�q`膡|o^�0g�<y�x1�2)8�I�����O���'�$�0K��R�ةB��"�a�����S����ɰ%�b>�۵�'�����t���kX�_�R�@$ĉ�����ݟX�IΟ���n�O��O��1Hh�0�˖Ѕ^��sC�'�7K-���d�OR$n�@�Ӽӣ��,M]��  �h�X�@��<���?���A��l�ش���Z+~,��B���.��F$�@	E�$u0�"���<�'�?����?i���?	U�
�y�eeq�Z�G� ��ĞǦ���yy�'��O�2Oſ	6֐x0�\ & (h�r/ۼ"Bꓙ?���d�
�&z��2�㝰]���3�e�#xA��-Zv�I�}�D�a�'�h�$�H�'��ũ$�I79�bq��h3R!rW�'x��'�r���T��ڴ]�8���);�$R�w��(�7Cͮ�����v�$x}b�'w��'/�!j&CA�}���S���N�������[Q��������j�Q>��]�x��T1�e����u�M�t��	՟X��ɟ���џ��Ii��Ruf� ���'M�u���An�3��?�hi�&o���ɓѦa'�l9pG�)l&@{���0H<��`�T�ʟ<�i>M�#	���'Z���s��D&O7I�5H�
�.,�I�Ae�'��)�s��ٶ'��'�vA�����3�0$YD�>ÛFg� ���<�OV�fA$K"�;e�_�;#pYz�O��'cb�'ɧ�Iޢ1���S��#0A��S��+��-a+ϡ9 �6m�Cy�Ol����c���`�M��V �HO.̾ą��FW�V��gᔅ�@���8I�MSa�ӯ.=�yF^�PR�4��'E�듮?�d�U�'8���2ft�2����T��?i��/lxh)ܴ���	�]k��y�Oq剁?�.=25ŷO�] ��y
�Ibyb�'u��'�2�'�P>uJ�ɕ�T�H<y����W�$$��ܵ�M3�Z��?1���?�L~:��w��y3+��0��9zP�E$z�|����'���|���ۆF[�60O� ��[�]K�~�ؓ/z���:O�u0�j����9�Ϟ6`��ץМUǀa�ɚ�M��9�̅+kq�ف4�T9�
H3䍇�s'�����F�b�1s-�/u����4%V�QXy��Hމ�� ��h'Uk��D��d�`i� I�~�@��ڶL���cR�@�#��i�`����^T�dȲ�ݚ3Faz�s����gL�L�f%K3)�"�����n�.j.-+��U�>��L@�lG2 � aaݯx߶Ŋ�.��^T�Bh��M�6�^�VB��%+V�7(Q�� ��?�����G-U����%)b{.�R0Ed`�$��M�
X&�n��ɑdV��K��G��v��T`X �ze�ٴ�?qL>���?�`�L6߸'���H�$�ea�U�d��9 {�M�ߴ�?I���d؏f¾��O�b�'#�t!M�2�$�&oݜJ�
�+��"O"�$�O�<@�!?��E*��L�z\�P�4+E�=���2�&�⦕�'y�1�t*w�L�$�O��$���֧5f'�l��l3e���ꡓ2$Š�M���?��'��?�N>I��d��#�V���Y.�zQ���ީ�M��픪-t�v�'b�'?�4�>�(O|q�T�UE��1*��:�I!$���xJt���OqB(I$���A��.� t�`)�
N�7-�O4�D�O���2�p}�Q���Ii?)�&\=T 
@�ߨNS�`[�JYS�8�D!sN>a��?q�p�^�{��Z����qB�'f�t=���iN�%_�H����O��Ok�W	Y}h-GA�"J(�9��ʌ3F ��$9�]&��	ޟ��gy"��8T@nѻ�n�__~�yt�T�{PJ���>�*O�d5���O
��*9R���&��Bu��wm�iA%��O����O`�a0���5�&!1o�K�~Q�3�Ц�y�A�i!����$�X�����r�D�>i0�� �� 	�H G�
HS���M}�'$b�'��	�D���������8<"Iz�X{�a�I֩bcP<lğ�'���IğH�e*F\�H��a�GО(�JMaꝧV��o���P�	iy�F�$��'�?q������x�q���X�.)Lq#�荝Mى'\R�'~ڙP"��?=����y�RB��tR��,x�`ʓ:�J����i�B�'R�OyR���,��QH����F	pn����.X女�	ӟ�`Ɍx����O�=�����
T�dEn�)ݴ�9�ųi���'a��O~����O7Q�Tf��V�pM�ׇH�S�"un�5&V0�?a��4�'� iCˏ��hQCR-�
����Jr�\�$�O��d�H=�D&�����7�D# ��z��X����!�nZݟ`&�����d�Op���O�D��#\�WWh��G�֫n�sa�Fܦ��	��
taM<�'�?�J>��I %B�Kx����TJŀq� �%�X�I@y�'v��' �	�[&I�$��> ֔x�ʇ5�2�;wG�>�ē�?���������Xf�VC��ۦ&Ѕ��i�rX�<����4��ay�O�!0غ瓀x�Z�2��B��@|�6F�5x���?������4����]�[����FOS�J� �dJ?<s\h�'{��'~�R�(;�,Z��ħ,+Q5�ͱW�X�Ӆ��TmH�i�|�\��埴��dX��&�#&��c� �J}��3 �i"V�P��4�ؔO6b�'F�\cEx�id$�4M0�Q�U�Jbμ�L<����$��\~�֝^�Qsp��chH	����?vH��?����=�?1��?i��*O�.��~̢*�;�@� g-�kc�v�'U�Ɇ��#<%>�Ha �9��KW+�2yЙK��j�<<c���O6���Ol�����S�t ЁOkܗ�d�6	����ќ�+wY��pA�'�S�OY����N��I��8k��Z�0�U2�/pӼ���O^�$ݳI��S���>Q+U�>�F��#NܳK�E"�ҡN������'Y��S�c+^���gm:���.}K�V�'�Ȑ�\��[����[qj�� вmŅL������tft�<�����O��Q3��
�L(!`��Q4Dԉe�F>6r,˓�?����'1r�O�@����,X��� Tw9Z��°i�L-k�y��'���ǟػ�jV�p��59�:`jtg�4�U1�c�����IƟ(�?�����ux�v�ħ2# h#�Ψ��=�ҏ] �ē�?�+O<�D��stD˧�?QT&��~�J�8���Ot�r�̺X�����Oz�m���&����E �n���%�j��Je���d�O�˓��Ē���'��\c��\�oR&�Lc�O�<ŀ�Ob�D�<����?�H~�Ӻۃ(����t	�`8c��YRG����a�'��*��r�N��OL�O�,�vr����LO����q��n�ޟ|��ܟ��I>���<�.���b��w�|Uy�b<YVQ	����M���/�?���?����(O�ӛw����A9G�F* ̞�1fx��O4ġ��)����5oE�)�̉HcaW�-Z@y�Á��M{���?y���<0'�x�OnR�O԰x�C�vO �ю��k��!�Ĳi�|���~��?A���?q�"K��"�� IF�Xu�2�@;���'�~��@?�4���<��������+%�8��n�<��B�x��'��������<�'J�5BУT�Ó���*��a��޸�,O&�d�O��O$�Ӻn�5qy�����+}˔ݻ��Ҧ��	Zy�'���'i�6#1z�H�O��x���v*���׼o��d�޴���O���?����?!T��<�v� �Ce딛}���j�/K1�����i�"�'D2�'���($i�)Z��z���v�[2$�<>[:0ҁ�ғ$�L}ـ�i*�V� ��Ɵ��	� �$�ҟ`��4�z�k�˜$e��ڃ�[Vi �o���	y��~U��'�?����j���v�	�֣��h����R@�=��	��@�	ԟ�ke�i�D��y�ן���s��	W(a��h�${��y��ir�<]J&��4�?����?Q�'`��i݁s�)V�ka0���D�T��a�t�c�:��O�*A��p�'Oq��dR���./:J�e'_�(��e�r�i+���5)g�
�$�O��d�����'Q�,miX��Q� �T���q𧟽[�0�4j4�̓�?�/O��?E���$<����(�\m `�A�V��<S�4�?���?��Ք��	fy��'$�DC�\ �
�d�7.��G뒛;d���'��	�Y&��)*���?��\ �H+��;�T�p�#K�p��`B#�i��vx�����O�ʓ�?�13w6A���L��`�%K�3�P�'l��ћ'Z��(�Işl�'ʑhi��Z!R	�c)�0^�`	�-SFi����$�O�ʓ�?���?a���2��܀��cψA�@J��z�Γ�?)���?)���?�+O�EZ�F�|���Ykh�p����z���5��ݦ�'d�^���П���+/��G�� �1��<'E�an��mZ�H��џ��IRy��k��'�?!��iV�8jբ�f���V���<Z�6�'�������������l�\��M�A�V��l�r���v�dxE-�馩��ٟP�'�.L(�~����?��'L�z���Y�rո�oJ]�ੳ�S����՟��I}@��ʟP����T�'@�Д ѪQ	Z�䅓d䏮+��lZZy2�ڦ#�r7��O����OV���n}Zw��=x���[e`uP&�S&P�J���4�?I��g⾵Γ�?a(O<�>����!VL��S�'� ��W%}�b(�`ʦe���P�I�?MX�Of�T�	� ř*u-\0���X������i�@U��'V��'��	�Od@ap�]�bLqj��(/9��r�o�i�I럴��%��e�r}bZ���	r?��\��n}�fI�,8rŹ7����ퟄ�ɑr���)����?��s����VA�Ě�
�@�j�X��i��-�R9���d�OTʓ�?�1h ��Y&���m��h�$�K�<�4m���%�x�X�'���'CrU�V�H�KH��XT怾g��|z���)"�����O���?�+O����O���E�U�A�痄����g���_fĜ�7Ov��O��D�O��D�<�2��E$�P�Jy`��&�^����O��O���Y�p��sy��'���'.n�I�'��X:��I �*$֮ϒ �1@�,w��D�O��d�O�˓= �+�W?�i���@L܄�0%n�WV�U�,s����<����?	�9hx���i��h!˙2�˰Id݊)��4�?����d�C@d��O���'���	*��JQDE�6-@��D(��[�~��?a���?����J~�R�\�'����C+w ����qu(Im�`y��=UP6�O�d�O��	�A}Zw6�(c�k�(q{��"�bƙ	U���ܴ�?��rTp�͓�?I.O^�>9�&NM� D�}���А!�Z��q���`����	ȟ���?�9O<A�sjb�@�&߽ب
���ư��c�i��p[�'c�'	����OL&p�솉PrP8��F�u5�nɟ��	�<����ē�?Y���~���Y�p|�2%Y�-~����,�M�I>aU�I�<�O���'��C�>"+���v@,#��O��0�4�yB�@�ǉ'#"�'"ɧ5V��r6d̑���bO@%�GN\.��dţ^'�d�<����?I����~8&YF��N#,����9~\���cMU�I�x��^�	�|�I}�t��%�
��ŋw��f��|3�?�I�H������'����s�p>�0��z�ѱc�I�M�8��5�>����?�.O�$�O��D#A�$���HAZ� P�%:��H���+�x�'���'V��ädG��'֥���=�6)3!�7�"�P�l��M����䓧?��]8�����I�2n@�W�޹:t��&�ø!�N7��O�d�<��{4�O�B�OnL��NĴ{�,��,��d.`bf�7��O^���%����<��?�f'�:kC���*FHm޹�� q��ʓ� D�ži"�'�?i��"��	f��4�r�2�DxG��0�"7M�O,�߂?����=��3� #jna���g`�f�����En�z9/�V9oZ͟$�	֟�Ӕ�ē�?!Q#<-������8��AĂ�g�&g��yr�|����O�hCp�@�2�֗��xt���	���'��N<����?��'��H�3R���ggL��ݴ��@Gz�+����'���'��{�.��G=L5�c�[#([pxI5%i����XJr<|�>!�����Ks���u�RmARjϪ*

1��oe}���rz�'*"�'6BX�ԡ0'��O�AB��ĿK�vX�gO= ��L<����?9I>���?�W�(W�1���K�~QZ���kf������O����O6ʓi���Q6�������	�tK֌�O��Şx��'��'��'^1C�'�x�P'(��u�\��2阕��%#��>Q��?����aU�'>�$�$;�hSq�
]��9w���M����䓯?��bFf ����	QwP��a���q���#��M�	ڟ��'�,�i5�I�O����U�����)A�����J]_���&������Ԙ�f���'�4�g�? ^,��֟f*R�zt$��`
Bɺ�iu剪��H�4 �����S;���I�0���Ӵ�A|0�j` \���fy�'��O�O\f�A1+�E{�ͻ �֏ol�0ߴ$~��K��i���':��O�O�	�9�j�3�IW<���۸,����'U��i�O� "�5.P�h@w�VV�J�L�֦���ڟ��	i�I�J<ͧ��'34�T�06��؛��X�Ն6�/�����'�?����~�5)�����ǔ�|��uI޷�M���n���*O���O��|rMʿi����1�{�1�o��0;@K�x�m ����O"���O��B
���(qa�x�0!�"0|C��@:]��O��D5���O��Is�x� 2��7'*Ti��b���	� ��L�ĆÇ_�)������Z՞��$D�b��?�����?���V��h�'Y����⍴H��0�҇D�n��Ѩ�O����OP���<�f-�2\�Ob��	'�J?-��y��͇�������q���:���O�D��}�O^��FcR��vP)�c��
��%Xr�i�B�'�Ic	`ܸ�����O"��D{���&��L0LDRMS8d`�|�'�r�'�2�F���Ĥ<��O�4�B�� ���q7aV�x�*���4���6���oZ���I��`�������"��O 1��x��Q=�V�S��i�2�'�$�3�'L��<a��e�1l�J�O�2	4���u�ߘ�M�3�ƍ8����'l"�'	��(�>9+OЈ1�mLQ>蔘4�
N�H���h�Ԧ=J�b�@�IIy�)�O�4	�I۝7F�8p�:��lN�)�	�����Hŀ-2�OF˓�?��'p��zb�
�~S$����(y�ёߴ�?)O����>O��՟��II�s�G"2j����ȴ�ץ�����I�f��8�O*��?�(O(��Ƽ�5č�p�0:�L@K��,T�	�G=���ȟ���(��]��';��`�4n�qYGϔ2>����q,D-Z� �����O�˓�?Y���?�fA
�(�*���=v�rmA?������O~��(��G�X,�ϧ8�6�����"[��9�tM���4oDy�'Y�Iğ|�	� �-m�HpC�0q"�q�R�� <Ș�ȕ&�����E68�Ģ���nU.����Q��H�t)�#d�h�Zh¥r��!0T*O<iaf┨\t�#�тU�TP�'�F�z��P�:��� >��x�1�֫"6�I�B�u,h���돺��m�0kS]�nɀU�K�\N=x!n۳ ��n�b�@+�ޞ-�n�j�l\a��i�ֈF�h�]��k�%@1���)�f@ʵ-ׁaS~p�T"z�P���F�8e��ő�	SYxH���W̢�K�������lZ��O�/d���i��y�l��\4m� ��Xе�$q_�#dG�����wϘ��&�� 8�z��ፇ�u��h��C3T{t��Z�0س��#87���H�G�P�f����܇��E�$i� �h��'nR�����O�aB�<J�l!�d�
#�X;"O�ik�+[�+S��C'÷r���I��HO��|��S��)���3�� �������T�!J�8M�	Ο<�I��3^wB��'#v����s��}H&l�X�&�q҄�O�ݚD/W�t�jX�wKN������ҡZU�q��.W�<-�s�
=����	f�bQf-^+/?bTR�ޟўtqr$D�*��M-4��
���A�����S�����O*�=�(O ��roڄM:����F�3�h�bc"O�ۖ�׾A�<	�S�Љu���&��@���ɰ<��ɏ�E���@Y�V�M&�!�ʍ��/ǯ b�'���'�~ �OK28�l	�cKk���۝:�����Ȇ_$�)`��:8�|���/m�Ɍ��"f�~�� sW`�4-p����9\��'�X<h��$R�zx0#hT���-bQ�'aRY�D�	R�S�db�x$�d�ݓ"Y���p��ybo��"��z�̂00��w����y�L�>�+O����H}R�'��S�>��3`��/D�Q%�J�)�x�T��O��d�O����v��%s��#�T>����N Y�������k�>)3�/�r.l�lB}�}�l$�*"��d�%%�lX��,�9�<��c��Ă�4ڱ�ց�t��>1�؄��`��W$����6O���-�O�A'dP�t�\Шt��"wҔAd�'�rO��
XNd�w��:'_��>O�@�$A�U��ş�O���E�'(��'G4l��H��W,u3t�̤%��%;w��~�b�T>#<��G�tJ�t!Q�k`!�E�>8��`����O~�8VO |��!��C��[Є��q�G�a�\��9�)��(1�)�;0"��h&�Ft��L6D����.ަIY���&�"��A�7�-Ƒ��Z:�P��ܔ1VbbM�[��I��?�UC�5w�\����?Q��?qr��x�4�dL��$V����
��/�~2Ą���>�u*G�OJ�\��M,%gfh��B�^?i�b�Ix����V�U�Ճ�h�A�2�+򭬟p�2/�O����7#��=��h�D؄��/��fG!�� �`Z���"j�|�C��D�L-���Y������4'LƦ]��ŕ"~�P�XB"��o�|Y�՟���ğ����,.�u�	���'L�I�	ןd!�o��@��\��L@B�(D�:�O��(�V��,�'\͊=+r��5
E��/9�O&a�'"mE(I��0�7L�cҜ��*���y�)̩UWе���S;L����Ԑ�y�&��L�C(�SD�@��dШ�y�"+��9`z��޴�?������U���A�dQ����#����O�$�O -�bg�O�c��'c{��[Tc�x�T�Yd�)TF��Dy�����=z�Oq���p�E\�Lw�@�� v ��d.�'\��(Wod0�s5,�!>*��)\�q�`^be��T�/���񉪗ēux�y	H5�PԢ��Eo���D�QCp�i�2�'t哪ghy�I��d���4�,�!�G�a�T˄/��v�$��E�˟��<��OlB�L3��	P���54U�E��@�C "<E���+���Q"J=���ٗ�9jJ��B���?��y���'-zY�5��
��H##@� Ƽ�' ��#F,U�]�H�AG��ɂ��DBI����L�tA�r�N"_h�@fI�N]����O� ؆�҃C�����O����OlЮ;�?ͻd���!8 %����e�$F�L��,�����:Ynx�u/��[���(@`ҫ%����=L����׌D��9�¡�
C�� �h$��$��'g\��`M8:���H �̸DeN�S�'�,����Y�LeIW�H�:��E#-�S�O�n��A�b�r2P�.�ptAs�V�1y����O^���OJ�D�:f���O��6<�D�O�4P!8p:��,\��g�'3���-O��"���qϾ0C_""la�k��p>�������;�*��-�2#Ů|����T�HC�=W��Y�a��"�Pd���/\-\C�I !2�z�E
?�v���a]mp���'Һ8��'j����O�ʧ/x.a�C)����0;���36���xV
��?����?�cm�?��y*��X�3�+XF���K];�BEp�	�BT�3E�hIR��57�*խLB�'��$���?	��?i-���"WN��P�F�
�JP��:t�vf�OD�"~ΓJ�6Ś�����r倰��p�,0�O�&��$��{��i����:6�8�Ci�RDI��M���?A.�T�q��OF���O(!Q�	��U+��	���P`DB�%���D?�|FxҨ^�=��\��E؂(Vpa��Z#�d9���)����p��8a3�����/���i ��C*����S��?yB�x){��! b����E�<Y��aBA���M7p7��v�O]�'>#=�O��]b��׌q�V�	�C�u[���'�BCڵ*4Sw�'���'$�c�~�;?�i�D��cF����K62����z�a�'R���w�ˮvo��p��^�]��,k�'�)B��)�O
}C���`�*���N�	���OՉ1n�O6�D�O�Y�p��vy� \��8"쟷a�8��)-�y�g�~��Y ����S���i��("=�O8�	�B�Q�40]I����+&52a�Q�
 .5��?���?�+�?!���$'�?Y��0�*�pd��p��QjV��3d<���Ih�ZRTJЀ^0��&�5Sp�݇�I=
�D���O	�6/G�:H�H���S("��L�"O���hDF�1�� v-#"OB)��S.����7���i!���2O��>��gş2Ǜ��'�bX>�xG�+��]���V�;�De�FL#*����Iǟt�I"L����i�S��� E���SȎ�>��% O��(O��pS�� -��@sb'WPdk���m��<����hG����71j0x�ʟ�<����$�y�:%TT�%�h[�H���0>A��xb)�=c0�!DėC�n��*�y��T�	N�8����3�\�C����y"E� ��jW%�`[�i�䣋?�y��	OZ|�B�T�UQ�zWϕ�y�2Z0��F��!Pm��2�OF6�y�G�V�dm�@[�CP�	��Y��y
� 8M #řOz~8HR�F+Z���"OX��ѪJ�y�:�ʖ'�(���Q"OT%��$��N
�"G���1��ʗ"O��׏GL2<���7l��0�"O��"�+وz�.}�)�2�ԑ��"O�T��K_�+�z���'�����$_y�<q�B�􊠃�_WZ�%�e�I>>!�D֒y�9�UBȭC���iC�S��!�d��X2RhSׄ��D�;�(��d�!��ȍW!��r�P�Em dq���]!�-_%��(���9��EјY�!򄜯s���� DǤvP *@��?_�!�� �ArX[*ƈ��1+�V�!�^{��`p�e�W$����9�!�[i�(@ƅ+Zi|�*1�	�!�d��AJ������yb`pB��M	\3!���D����BQ&�#�W!�dX�;���G��[1��s��z�!�d�N�@�_�:���P͒��!�d�'6޲�i!�3O$B�
T* 8r�!�����MݽA�=��HY�!�E�H��� O��z�ȸ+@��4�!�D� o�Dj��`�Mx��!�$P&f�p�W�φn�)�N�$!�ٕ��P��X8]��sN�%!����8�;�&*���65!��� l�f��.�� ��81!���gL�-���7�� S\�!O!���]�z4�K�	����!��aK!�$X�| �}�B!X4ADp�
�(!�D��D�`��vDSzފ�Z��ة5�!�$[w���$��s�hG�S�`�!����Ld� '�@ּ`6Ƌ�\�!�đ3Ta��ӗjްR$l��3��!�D��R�*I�	�m�(��"J��!!���o���A��s���%h�\�!�D�����K��l�t��K�!��  Kt�d���G�9xpq��>�!�$B'&�� ��G�}��z!��0|/!�dȄV�h���;r@	�F�
~!��D1t��� &W[�]�Qn�=�!��-E@B�L�<��8�� r!��]+p艅e2PAs�JE,v�!�D!!�&!y���/J����#*�)�!��#`$:h�ë�5Cj�E+�H�7o!�d��1<�(#`��-����"i�~~!򤊍s$H����K�\�E�U�!�ݳ|�����ift��E�5K�!�$YI��� �hb��;��  �!��@>�2x��?iW&�dG��!�ě�$�.�7��#,rQ�p�αF�!�DC(pq�̢d �-}�}J�.@2[�!��Rê�PjOp�؁"-�,!�ݘ ,�P2U 2�ˀ�W���>Peh��$1!�*�Hqj	6�\��
�f��}R
�b��/]�@pK�W�J�#5�ޟ
B!�$D�[ �{Rɇ^Q����ў�J��F�O�ɫb��(�q8 G�;R�|��'���1+�E�@�ʀ�JOڸt[��B0�>��O֌�(�d�+t�/ ��%9	G=�)���!D��T`Zv1Xa��،���Ea�tc���:@$����HFqO<Z�L�����D18,y�A�'0<Y����ᦹkR��#���B��S�leRpk�D2?�� ч*Y���D�b�!Gn�=`��:�� \ўP �YgL�'56�H��� �]�V���P���Af�
�9;^�"ON)� �Mv�z\"��	\ 4`���'Z�� ���g��	E�����ᓔ?�T�9��u�qy2�DE�`�ȓlP���m֮  I����(���}]f̈��K����b�d�i�,Ё���E/I'<RE��I%8Z e��i�H�V���\����G��n���O¸�_0�*	ד,7���e��l��x�g�@�t��D|��f0�O�pB+�- �p���|��`W ��
��)�"O���RǶa|ph�%>
�!����'EE�\�gOηb���
�Sn��� ��n��x�h��I��R�E &"O�q��_�w�5J"���<N�u��$0��zs!@�d�Z���'�>��f�Od� ��2g�3Gnlc|�Y�"O�)s'��A����j����2��'�|�� �;.&8�UB
S��(q���/K`�[��&�K#
�T�azBe!HD�$��^
~X T����)Ar�vMZ�����.��� �r���Q0@ɖs\�aR]�.��1*���i�B�"h"}r�ܯ�)�l;�~Zí�W�P P�� Q^�����^�<���("<<������9�NعC18�� ��3�	Q��ޒB��U9e��~BF =�j�p0F^onͩ�̇��>��ė"Y�tҗ�F1B��y���"��6�|��^�9`��&��(vO}��VQ�'�>}聥�6I�F�7m��mX0Q�����8>��Ve��%#f���N�l����w��8��[�_���� �/?�^Hx#�Q�C:�~2�f��%���ǣf� }C�h�8�M��ϖ$���z���/(�j�q�S�\c��P����+}����pKO�I�N���'� ,�0 �Em)�ĐN���ТK��O`�j��9�V*P�a8��'��C�.҂1M���+6<�q��P�����eƟGz����(ѕB���2�X	Ω���O\+���#!,��茊������	���컑��	}Q�L�g!��<y*�Mz����Z�|S�\zy,թ6�l����o�zD���<AR�h7�_��|j�L�	.p�p���"�<)sIݧv �e��
('��(*�Ó�r�|�>�ϿV����� �õN�0��L�<I0��ge֬x�D��snd5k���DC� z�}�џʭ[���67g��h���}?����<L�`H��f�u�*%Q�F�EX�TH�"�KV�q��k;ah�Q��э:�]�r�S$�?�n@95��:���%k�>Dp�c[�'锡����j5n#5 ֊r��A��D�4J�EP�G�Z7��cU1��^#���@L�Iy�8��5F(�8�1��M��~�N�q�����U,5V�2��ֵ�?�G�AJ\�Pgh�
3il\ɁFO�S�4����K�n6��S�o�����"O�Y�A�Z9d_���Ԓd�,d�c�5\$��A�y[>}���˒������0�g#^�M�ܛՋ�!��+3�O�	둁�[qb=�c�@�M���w�U( q�A�b�'���Ș�=�X� o
h�b<���P�x���c��1�ŨOW�az̈ <bՃ�#� ���sI�3 ���jL�m� IV*�$8t�J���sVj�db
 r��\$���+#�2�$���#'%J"�@!`�8��~ڶj�a���Y�&G�z~y��f�E�<I�lž>,�*R�'�-0G�ٛ$NV��W��bu|p`$��⟼G�d�HS?AR�ƙ2G�� FdQ':���+M{�<�pÕ�KHp�7O�G^���M��K7\�Z���>s�P�u�U�]�(�p��,i�@kGN�<	���"�%F +g��&�
���=�vN�!-��a��kA�r��	����(
;P٩@��Fx�(�D��*��M�T\j���E:�+�- �N9dA�=�� M��M�PBՅ6X.��ӞeNv��ԁx��!��J#El��O��aR�Ka�S��0#3��b'���\�E�@l��AW:ݛ��J馑��㐛�qO?�k'���V��{���	:��l�(�x�0��	��OǸ�{w��UDf�(��)ulHQ��#{X��d�O��0Tϖ4�p=����	�%7��г��Y�Dj"c������?��W��h���k�C36���)bd͓J�$P�*D�L�fF�B�!
������Z�'���?$P���4.��(�I�?�c��H����!uXɻ#�O��0
#�y���=
��G�T�Kxtl����5�ؠV&к1�H���O�&kq���L<AG*�cMb��ڠ<�Jט�d!�$�w�|�����a t�āl�8�aإ*�(��V�& gN�|��Xzre��zi�h+T X  �\X�'���Q#�Q�d��'K��H%JC�b� �����,�� #_����a��H�Ԁ)�NZjh<� �t@'@�4��xbqk�UE��r�+}���0ib�c ��n�`j�n���5@��&zlK�wy0v��nJ�M��Ҝ/���*��vqK��@<T������L�ZHAgʑ VU�� ��U�;�h�P��$f�cS�A>P��g��ɐ`��ʧ,t��3���
�Т?�W,��𙳞x�h̥o���Ȓ�C5.�锫�p�F]���F�LɾU�t�X�9az��[�B{�L�Q�F8�2�V�����ӏ8xE�Z�)�Q�����7[����0IA=]�Yҁ�L!��ʑ��!�(�S��zQ��n�<	�(�qO?�D �cX�x�,^�7L\M�"-��!�$N;Y��q0��f�(0@ ��qf����w�c�1.��qLJ�n��<�梃�[S���
�~mI�8OE��'O�h��ˎ.�n4��"O��Fb:,�PD�6�� 
�B��	kJic��)��Cr*� ����t��"� �!��B*&�Y�aZ�A���⦦4U�!��ݻ w����*�&2�©�`@�2:�!���5o:0Ċ�DG���QB*2X�!�d�21�<�S��Y�S���&�H�+�!�D�{����ҡ�7(;�8�\6�!�$�o���a�E)G�.M���.[!�$Ɩ!�Y���u�p���)Q�;!�$��b4YpkկZ��<p��1
�!�$�0�`���$��uǰ(�̈0!�d�F6���ꟙĶ ���ϴH�!�D׷l��(�@��������2�!��
N��17mG/P��15�B�!�d�\���i�o���*�Έ<!�$�Xk�I�ca�>8 ��y`��/�!�D b�Pą��b����*?�!�$��rY<]ÔąR�01c�C�Y@!�đ�|H� h������刾-!��^*IL�%
��D9erd�e�!45!�-me��ys��md<�G�N2`!�$�P�P�	�]��	�3m�!�D����A�6#v��`0ȝ<[�!���5�|py��J41�D�t��!��1�D,3h���v���Ę$e!�T'-B��Zf�ׇ$�h�τ�,O!�	=����;5�J�붨��s�!�䑰4�"F�( �t8��U�!򤅆6����A/H� �L=�"���!�d�)c�J�h_�]���0e�!�$;�>��E��ͼP[$h��<�!�$ɑ��5K��-��M�d�V��!�dW�Tz��ׅ�J����eӸT�!򤋞o_�m;�K�
'�,����D�Ey!�$ؕI��\�0o�+Q�%�6�Ɖ9�!�dܮY�Xq*V�RI�� ��N;W�!�8$�Nt)�b� gc�J��R��!�d��u���� ���	Ac!�ܿ���DHD�d��(�!��"&�Z5چ� ;.�Myu�U=�!��f[����Ӓ�Z �d��6�!�$_�"��L�a$H�ph��$� e�!���vTH���|��Y�Mɔ7:!��7�Y����Ф��՘e!��F� }Rek�jy���{^� D��J��M=Rp��U&X�&R.�XRI2D��"@o� #i�X�t�B��
���C.D��H��;�)� ӤB��z��(D�K����Zv��%Ï-���� %D�Ѐl�(l��tcҠΈCU� W #D���DO�=#l��	�j�P�
@# D��!�N�)�A�5mC�#e>�T�:D�� �ę�`�1Xcᦔ�d�tГ�"O��Dl���PFE̤f��)"O(�Xr�!_l$�6$5B����"O�`���Q�TG"T �DƯ ���"Opѩ��#P.���"�Y�E"O ���|����D�m��1v"O�lZ���� �ӣI�S�X�"O�)5	�:Z^�IS��v���:c"O�t���\�*K��� �����v"O�L�!��m��š���b���:�"O܍�E�g��L�2��$
�P"O���n�C�X|��NP�V�J�k$"O�m�@_#Lbz �1��9��yG"O̡'��9[�hf���Zt4"O�|9��ӤTd|�vBU�m���IS"O0�:�*���+���)nDR��"O�SgiLj�$uk����E0� �"O���&m�.��T��`��o�L�7"O  z�)K���'��"Ip� �"O�,g�D=\�h���9&#���"O�0CQ�_�h`З���7eP���"Oz�*�$	Pp�A��_�2��{"O:��u�A��Ȍ�{�JA�en��y�c��}b��C(ԇqd�5:dc>�y�I�?�`�	�ʷ~ST�ڒ�	�yB�.�PͲ��f�0�s��C��y"N�<c�Q��"�b��M[��ɤ�y���U�$���'��n�a��$�5�yb'�|�9��.`檝p��C�y�(�|*ƍ�T��4%L���CD��yBn��?��Pp��'�� [����y�C����PC*L����ZTƃ��y�ſKrp���n���4�C�ʎ�y���bh�,�1�ɹM8(Q���yb	A�H���
'�h��g��yb�ЧH�hX`	F�q�H��.��y��7g4E�7���c}l�H�����y���Tl��K�1^*��
4H��y"-L9�fT�S\�P�H��f?�yr�C����3ƪ�0 ¬�y�M_��p�kƢ@�0+�<�r����y�h<!�p1�L��33�:�y�+@�4�Zh���G�4�����y�ϛ�5D�S���H�I���۟�y�%������@�J:����!���y�B�r��y9���7.�:-x����yr�s/^XА�� \�#U��yB��&��ipU'�2l��{$��yR�(�8� ���&�!�MG��y�E��w��M{'�J��� KA$_���'�ў�p$)f�9=0�i�" _�+|t0�"O�D����FP�=R"�:E%����"O�1y0Hɷ �4��N�v�D���"OL��(�*���-۩���b"O.��p�&Y�Ɛ{4cLm���"O*�
�Y�{X8�{�Q]@pi0"OH��R��ln��#��Vr|�S"ORa�E�	Bg���t#��r9�<��"O�9֫Y�$����!6�p��"O.��%Ӽ��yzĊզ-� "O���cM�4��Y!aiήP
����"O6-�a)�*tr�I�/9h(��"O�bA��_Xza��!5)6`B"O� 1���ujX�Aa�n>*�	&"O� hX��昍+p��kg`Hs���"O��$O,aFd�Y��(*�A�"Ojp�c�	�VH`�E��/�,�)4"O���ъ8m:�QC������u"O�"�}���i7[�b�ޔ�w"OrxK��ݓ1��-��% vX��"O���D�4,�ΠI�F�(g^�B"O�)����n�X�P�EuMJT""O���$�H�ĭf�׺)E�E��"O���Π�>��Ȇ	�^! �"O(aW�U�.��b�K��5�Bs "O|ѐ�MQ<l���*�\�ޝ2D"O��z��ѥ_�T\�ъ�m_Z邰"O���3��do|�k��6J�r r"Of+w*������@N<9y��u"O̬��'G|S�aN�0���1"O�	Z5�H=?j��0���'u,��3"O>�ɡgT<�����+��Qd�T�"O�1�N�l�H���L�?Ґ�r"O���uO^>`�a��=!�Mks"OF|! J=lZE�u��J1�"Oz�x��M7b���3(B:U��9"O^=y�C��h2di�&p��ͩ7"OH�W��H�ܔSU��qjFe(�"O�jbj�OŖ� E(S�	O<�'"Ot%�!�D?B�Ɲc�L��?� R"O�ЊcbϱY�����
;3�exR"O��j��ޜ{Q��Ä�M<8\mط"Oh�B`��!d���j7�ʴ �ґ@c"O�H:� ��|��g�a��Dе"Oh��3�ʑ"�GG��5��"Oa���	".0���6��D�Xa3v"O 0��/�1���EڧW�>�%"O��q�ê#��!Ã�4vo���"OYQE�B����ᗔzU�B�"O����26���%���8�ҡ��"Od�.42��tO�
�F��b�M�r�!��K�R��Wd�KM��Zł̕B@!��z�[�"�.$<nP�v/�'*!�ȟE��H�\�nۢA��N�!�DP���	bd`S�7�j��"�;�!�Dׇ6^|���������⦢�48�!�$��t5Z��q��(Ɍ8�d���V�!�$Ƹ}��x�fˋye����!7/!��ԢD�G�a6��1�$T���ik�@��kͯ ��02�MeF\�ȓ1n4���O0h�0��b"�"}��Ň��X)#�It���$��PGvЅȓ>��x8Ԯ��@�0��ךc)��	[�'�T��f��a0�y� ��&��5�J<����iĹ[P�L1�nH�lu�e�nJL!�ė�Ef�JQ��a���R��d^!��ذ]�yJ�KQ�l���IuKA��!�dHM��0Ӓ,�$l�@����ʀ"�az��D\�w[�k��x:��6cC�}�!�ѷVgz��)Լc(�O+!��	aЦ4���N~={�FՂ�!�D�/O�<�e�Dd0~�",U&Qm!�ě6s��) �X(x%�M+!�V�HV!�Ӣ=��x���l9�(�㤋�GH!��>3��e逡d1�<�A
��A!�ŬSǒ��"�����u?!��+R����
V �f�g:!��X
���Q K��eeN�.�!�� ��v�@:6�H����� ]4�W"O�9��c��:G2ٚ�L��?��`�'"O�T��N$��APkO&O�����x"�)���V�Z����7w!fM��ӈ%LXB�[f)��	ݠQ�R��IX�jc�`S��X��x$��D��r���R���g5��?�U#E�D' �"�օ5̱I1�^ V�����|(<�`e��8�R��sn٤��h�<1P�E�4��a�/����|�<�����b�p�#�]�t���!�z�<�$vqNǄ�b��y�<��판.�$1HDC� P��L�c��s�<YgK��Ia��T�E���� H�<��'��5�&OPBX���SG�<��jZ	Z!8�.V%2H�|�o�m�<1s$ٚ"���������Zb�i�<��V-",�5e[#|��}J@i�<��aD7j4Xp`&�'����7J^h�<���a$����)�"l�m��&�O�<a,� �!�!ŎrS~��P�MU�<I�I�4\~��'�Ō1s��91�Gy�<�����j��@  I<>䪷�o�<���T\T�8u	��`�̹�w�p�<�c��?,����	4H��ljI@x�<�ч[b��C��$+�rdrE�M_�<���L�(�Z0�&'
�~L��M�f�<�T�Ə�b,�Ē�w98�I�!|�<���M�����B�OO�����w�<�qI�sj	Q
��-�qD�Bq�<A�j8wS�I�G�n2P���i�<���T��Yڀ�Ķ��u�G�F^�<�wȜ������(����4�Q�<�!�_�{<X �Ʈݗa.�(ʱ��I�<@��#&U�t*�NE)���RL�F�<a�M��H��S6���y�<�G�/n����٘�Di�m�<Yu��7!�.x宏*K&�H�f�m�<��Һ6�r��rl�������l�<�G��S�|0J �P>�XG�L�<acG�DL	`֒*f�Pa`�K�<Ѡ��${s��R压�A�8L�E�l�<C*�1�b��0l-� y�%��S�<�$n��}T�$�M6m{a�O�<�o��A��X��Ȼ���0�ˉH�<1 aE+x��H�4.��~|���B��I�<!�� �6 H��5G�t�
��MG�<af��v,�1]�}ϸy�vaOW�<����Zܠ�0m�<���
U�<�t'�e�0���&וj�|��IU�<��'�7e���۴����y�͒L�<�"�΃f�B��	D)H�Ң�n�<�Ký8�Xkb��u2�3�A\S�<�u�I�Vd��{�J�
A��E�U�<т���At��� �dP�er��U�<����r�	P��O�B��4-V�<���Yߴr�d�,�"�y��N�<!����H��ɳ��;r���L�<1���13�ڰ� ܀G�EY"�Kr�<�c-O�'^��D�<.�z�;4��o�<ѡ���o$}��8U�L#R��m�<a��[�$@��U�<�t[�`�d�<y� 	�����t-׬�����Oc�<� �4hya�@�)w"ɒ.�_�<Q��E�x](My����B���`�<� xyRG��}�$i	��8�z��"O���GE<l<�3EǱj���"OB��J��1�᠆�ђa���"O�U���� k�8jdcM/_o��"O��� ��>%>P"S"]��>e	&"O�`�u�>_v��뎼iB���f"O�����
	VČ��ai��?j�J�"O�q��iƚO��Dˁ�Т,<8��"O�r��ň�����M�)��HP"O�i���
�K�T�e���'"O�(�5c�~�@ɠ�C�aq� p�"O8ySs��8\�R�ɵ��HSH���"O��z��I�<���q��33`���"O���
��l[Δ�w�ǈ9/�j�"O8��ʞ6v"�j	�$�� "O��Ҡ�*W���T �(�"O�T�HY ?�b��Ճ�p���"Ol�X�+Ƕ�)e"O/-cx�R "O�� O�d3�q�aA�����"Ol�r�*V�.����{�v9§"Oɳ��`��c�Z���+�"O��v �?�&��2f��v dA��"O���&���˥��b��3�"O��RAG	U6\�����7F�̂"O��e��p�n��R⅞r@�8��"O@�[aߺ$�����A�3]�Z�s"O�����[�R�(]0#�0�Uz!"OV�R����L��� S����%"Oz�bb�<��p0����F�\h`"O�DkD�ъ"T
�ٰ�!�n��Q"O�髷�ߛq�>�CE��g���*O.�K�۾;te҆�/rn��	�'�P���ǔZ���6!�r>�Q	�'��i���)4�T��`͊v�V���'t��ׇ\8��TZ�I�-gY�dz�'A~��'�Ųt2u�$�܅\�4Ȑ�'N�}����kȨ�TBY>Ɯ���''\ �"�ەo�L�Z�_�e�*���'��4���M�Ӡ�QCmU3P�4��'),��i?�N`X��ī={�� �'�H�2�a^�u�x���92'�S�'�}�W�V hs�T@��*�����'Wdi�DK-`�\��J�yq�r�'u��cT���Iq�B.#Bĸ�'^�Psp��%sV!+�b�-��H�'6Լz��FrOFM�GI�8!D�
�'�d�h6�Z;D�m*���/��$�	�'t�@�5&�!����e�Py�1z�'���9��X�v���	 5����'��`�YD���9@)K A��U��'&~t��hOZm|��g@4�2eR�'�f��3���ʼ*G-�0)Uҙ��=�T���Ж!��P#���b���ȓj~�,���ŏ@��)[%A�Zk�d��PJ�-�F� j�JT�3�Αc�����v��$ꃂ���4�`D�#�q�ȓa��U�qW	�^��	��/�1���dQ�%��U:ZшߗUc&(�ȓn~=�ЇǸ#�~XA�f^�+���ȓ��Ya
O�}>�$	 �F�V�.���GnD�)�ר
O�`뗋\�p�^���w���D�3.�SG	l �����T�b��%	l;"�P
1��ȓ;�a�z	:u� J���S�? H)q�Dݡ.�4ұ���Dj~���"O40ٷ��k�ajt)�@��,�""O� ��K�1&pk)H��̩�"O��#����
�@�;��C�j�2�"O��4΁��4���M�w
$��"O��QFV�+��l�,�-b�a""Ot,"���uE�PQ�
�K�s�"Oz� �N B�r�K,<w����"O�Q�v���t���݂X_����"O|E+�l��E�8!����%]$�I!"O�qbF��b/� �7��s����"O��Xb� �$Q��̜�+�(Qi�"O��k<=�e�)��1��l�F"O����D�7I�����\w���"O�4�Ŏ�(F8��`��&i�j�"O��"��)p���	!�cШ�`"O*��ѥ��J��e�`�!	[z��v"OH����E1j$��RO@�C�a#�"O�1�"%�
�I����+��ن"O�S�C�=k>�hj1ț8% �BF"O�����ܱVQyǨͷE:0;�"O�����X�3�(�Ĩ&I�<<9!�$^;�H�7�Q(�,��%h�4 !���`G��W)Ӽr�8 �WD��P�!�$�"ܶ����B)�"Aa�@�!�d � �����P!#��uAqA>9�!��Ƴ%-�@
�	(7�&E�� /�Pyr��nv$̻��f��$gĒ�y�$�3e��x[�H�?lBHSĨ��y�$�3~���h�B��B���=�y�J�hR�a�e�ڕ���7���yb��5�L=�P'���ˆ-E+�yr��`jXU�p�0�>؃P��y���+D�X��cH� !�K�y�i؎	<�� F�ô�2x��N���y"nS!4�JL��뉲]@(j5 �2�yR	�x�\�f�[�t��5��%�y�`�L47nMj�����y2-�0G��I�*�$dozk��5�yB�
[��
�@[R&�����y�*�'ONșWMD��8����y҂K�7PaS�ѳ���xG�a�<A`��#d��Ijg�j�8�r��N�<QF�z#h}�@��X�C��UT�<�C#K&R�P���U&��ӳ
�L�<� A�Tn�pL}�eʢ�y"l��e�mr�& �І�u
���yW;x�T����D?^I����y�DŢ8��805N
�~�sk"�yE��T�@�`,_)(J4H����yb��*4��hs��9|z s˙��y�)K0sˆ�)t�X����AM%�y��I"�����U.Ib��y��X�#O̰�gx���b�]*�y�+�7�<�*��<]Jx��"�+�y� F�Y���Ņ�W�D��hͦ�y��K��!w`��Gfx����Y<�yR"�]�8��*�̋t
���y�[�!r"�$8�}�W��yB�д��˱�U�JϺ̘D�Q�y�GY
2��P�@g�%B���hAm��y��24'�!�����Ї�/����gs�m"�d�<�h�Ũ�pSB��ȓ��%	���8��Q�Z�u��S�? �IST�G�2��w[�R'��j�"O��+Bo��]ʦ`�B�p�`�S"O�a�Fn�+; (�cN�lHX2�'�ў"~"��^h��n������k��y�&��g������*I��Q%�yEAF��$;BL��c��(�&�8�y�aI(�d��Z�X6�8���>�y�`����y��Lt�)ja�֪�y2c �1��9s�A����@��B���>q�O��ZC�D�ڴ�P�!p�rph��y�d��,��x���Z� ���y�
q�*�iC�@!z�����g���y�"�)RF0m�v���Z��<�u�݀�y�(&'�A��M^�M�r��yb� ��|$h�c�1v�|��"���y�ǉ;U�,��d@�� .�#����y���,b!���98,!T��(�y�뚤�2�H���~E�x�G�&�y��>0~؃�[l�A@�K��yb唥~�n����<]���rl0�ybɎ C'h�Y��ҋ)6�t��N��y��Ȗ�n\!g�'��=��MV?�y��Q�	7~���G�I2� <�y�DLbx��\�6�V�J��?�����e�][����C��5	ӆ.T
���w"���h�
w���OM)�P�ȓz
n���X(X�`S'қr�&���M�i��ţr0��`ѝ_HD�ȓ=eXX�eI�%DR�[,"�b/D�A���N9X��/N9I�B�I�7��lyWN���t�@EJ���D(�S�OyQ�7O6V�V�_���R"O�$(C)��J�ъ@�A���Q���I�<��`ͣX�uw�S}4���e�H�<q#▕9�>r���M�a�� H�<)��&A}h=h��V:*F$�T��E�<Yf�4>.�ݰ��G�}����y�� ��z-_5I��듨�-���䓫hO 0ЗM�RY��RN? ��$!��.D�ȣ�A.]�yx��+V=���s9D��1U��""��H� P�$=TEJ�"D��0Q $j~��25��n|4ux�?D�0�6�V�ҦX��̌N�I�$�>D���0��2���y�ꞷ5�A�� D���@"��,�z��5����i?D���SaO��|���\/j�0c�8D�\�`� {�tI�HN�E$���!D�����aЧ��b���a4C>D��b&E�D{�����C�9�m<D��*$j &I��| " [��1�p�8D�`[U�:M��D>A/��c �4D���N͔Vr����QW�H0	'D��k0H�5"�5��N�	+� !�0D�dQ��{ܔ�b�b��mD,�b"-D��@�W�I��1���3`0`[r�+D����MS�X���T)ՃW |r�?D���h�!x��b�#P��}��=D�,:��N�x�`���P�#
e��9D�pQ�GL����R�΃�r���*5D����jU(��TXr�TT�D��j4D��Y���
�����-mL�ՠ��3D����a7i!T�`"��ظ��p�&D��P�BĻ;�vx����'u�-�#D���"�
�4�RvFJꖉЂ�#D�� p� g#GBF�!�K�m��R6"OX���o��7�z�1����c�:0�'��8×��'z��0˝�Y�p ��0D�p9��K�[�`����ٕK�H!��)D�xH�IµLw��o˧l����g5D�d{s�Ԋf�$YX�	�%4@1�1D�XA�!D
M<|��g��s����=D�xsr�_�/���էN?KQ@��%D��Hf��,f�R�X�h^ξ"�o0D��aB��"�5BuТ1.ԍb�F<D�H�$	6	dё �$u�M�wI8D�xh@	�2�p9����q��e1�e"D��2��έ+���AtF��J�Pً��#D���v
�nf��5T�Z%
-�4D��p��J>"�h�L�
k截v�5D���I�&�ع�S�ըO۪�1ҏ0D��qe��D릙A�S�o��;�B9D��U�_��ˠ	�IGR�y2��O�C�I�UPD���@46�L��A�5^B�I�4�ƌ��5X� h��8�*B�Ɋ1|�zW��<TP\�`'"ٰ1��B�	�=;�, !���V��U�K�0��B�	6(Jl��.�M�d4"�t�C��쐃r�c`�Sf@T9jC�I���:��6��!(Ŏ�VC䉰r�e���cP�a�2S��B�p����+ϗ+2Ny�c�K9B�>[ �V@�N�҉�E!1g��C䉳WjF�bӢ1y����b�vu�C�I3mԾ�!�XdV��{/�B�ɬiX�cW I����[+�^B��0X鰨�Lz4���X��B�I�E@*����,i�8Mw��'�C�	�w�T��,�r�V�@$�НP�C�	.-�jxZ�U���Ɛ�C�rC���T��40n,{�R|��C�1CU�p+%.� Poh�2eNR�
ubC��(�P!�1cxp����2�(�/O����B�>���ٖ���S�EH�!�$�6w*�"oY�C�T�0Ϟ+L�!�dݏZ�.U@�,SJ�\�kR�Y��!�$ϫP����0��D�1�:x�!��G�o$d\ff.�����\ @�!��&C�0L�O�/BwнKw/ٞL;��2O�	Xc@�X�XŠ��`� )�W"Oj���GI��~�YbD�0D�	��"O*�ʃZ�6H`�!�D+c�>��"O"��,��d���d�X�]�4���"O�x���K�]|}yr/Ю#���IS"O<E"���P7ָs}4��D"OD�Z�"�.�847.֫j^A�"O�[��9M]��p��9�ֈ�A"O�yv�	&r<9F,�q�Jأ�'�!��#y�C�	DH��	����K\!��Yzh �aN�N߼��u�ީ0R!�DG�O��q��C�0"��e8���uG!�DE0Bh�u��șzV�H��3E!�D
�����G='������Q�&@!���o���3�:8�'KYEP!�Dɧ|V�����	;Ҙ8z�� G!��R�\�ZCj��m�x��/V�5!��FA����G�C�.���.�!��1hE��e�'-����7"Կ-�!�ċǪ+�K�A�|���R|�T���G~
� ����
�*a��PB�"\%^�3t�'�!��3���#�!��� ��JU��)�'
����a��`�% ����	�'��D��B_1CJ��`$�(~b�%Q�'�n�K��8�,�*Y	E`�,�'�����e*�t����:�4�{�'�6���-w�0���*N�I�'y�@�@�C���9��-�$#��QJ
�'��薊V�n����#�="�
�1�'�$�deX�\�|�{v.�?QIZDb
�'�!X�%ԐmjF	� kM̞��	�'�h�� C-Y��Zp#ќ\\^\�'�@��)�+8��B���_��8��'�$����MN�!��dݦQ�dP����)�V ˃�o��)�Oغ:�N�S$�'��	�4P�� ���o�*��=9e�ʓ�hOQ>�{v-g}�{���,v+!C�����O��"��SVt�)�C&R2I�r��-H�B�ɴrH�U)����YY�Up�ȕY@B�0ю9� � ��U#��U�t2B�	�: ��3l�,z��{��S�F����+�	�:�e���ɯJ�Lq���r9Ԣ=i�$}:�%�]���X�,!��m�ȓe��F��)2��$Z�^qʔ�'�ў�|�ŉ�.Ln�U!��=f)&��Р�n�<�Ra�#�`H�D �``8��Ņ�D�<��A�r�r�Iܱ��$iqG�}�<1��<hU&͚p⒄�zQJ�y���Γm���"�LK�������:����IB̓9*LQ*��+o���f[�D����332Q�f�<�t���F�E�'7��'?ɧ(�����,D*CaH�AV�\�yMQf"OƑj�"A�8�r�@�ċ_n�� "O
���C'A����-��<��}�"O��c�DK*bJ�@5�b�p���<�Va�;t,({'$�(W���	�Bx���'H�P�w��K�����;Z�I���:������0��E(�g�3eM��-�yB�Z#.E�S�o�2<���
��!�$��"E�IK�#�6d�����D�!�R���K!B͗G�����`�2}�!��,B�T��lN�\��9�Tj�%F�!�"3N����	1
�T���/o�!���z��v��S�PI��7k!�d�C���D�[X��%(ŕ�!�>#},4,RJ}1�\�`�!��3Lވ;ecX;O�X8�&A4�!�d�%�n����E�u���p�eQ��!�$\/�ʼ�E�Q�f��Px�C��!�S�l.��1��P�2�U��`~!�D�-H��3�ӦC����w	�4c!�$��H؝��N'=�R��7(�=0R!�d��Ow�x�@���zd���g�!��Oh�hɅ�2-��%`i!�Z�EF,=� �|�3��!\!��M���2���=���`�9_,!�Z�S���am	� �`�vOK�5 !��%�3К �Z�G�g !�$
�&���5W4�H
aK�k�!�āu����_��zVE��!��#:^�H�l�\CN��!$ȴ.�!�DK<�V"��SCJqA̒D!�d�	bqɲ��	@�:��&�̿%!�C7���r�&Ƀm�ű�.ӕ!�!�� @�slJ-Z�2΀P�J�"O�܂��ƧS�b�5�H!��"O��$eЅ?��p8���W���r"ON8�r�VS�A�G�"*�Ѐ�T"ON�� �N�S�b[ե^���"O�ձ  _!���BM wP&�1p"O�Y��ba�B!�l�ф@�4!�DқR�" c��.g�l������OZ���-9�P�	K��R5B���!�S� O:��@�I�r�,Q�3��9B�!�����*��_���(�Jp!�d��u�X��%�L/�ԸyV��^!�d?}v)�R��(���q ��!�R|t�X�u�2mbS`�.�	m��\����@
�H�-��j����F-D�8p�W�-�����®0av��v.(D�`S��@ܔ1kF(�m�#U'D���d�{H���$��wK\|Iri&D���f�Ң]�*��.:gy��!)&D��d�_9���)W��!���AD�#D���S#שs���Q���6�~	��!D���a��*�4!)��+��{$E$D��i�)�9T��p�$n����O(�=E�h�00s&���ȜH�v�6� G�!�ɕ3CJ=��f]�M�.tu X�!�(h�j!K�h��c���Ec�A6!�$�.�B��Aa��
e�� [9X�!���2}�@�aTg�?Yx.���*��!�d�:h����Ӂ!wd�R�)/C�!�D�����s��N��\�T+P,d����dqr#AX�f���A� +hkRB!D�L{��;<u �˓5��U��E=D�D����p��s%���!a��:D���ڷm��Ec��΁MZz1�q�7D������I2<跭��;:�	s"�<�
�sV<A$��m�jt�3) 'JF)�ȓus<�	�`^�.R�Q���p^�ȓea���5��pD>�qfIݵ�J���f��F�yO���G�D���P�ȓY��J��w�l���*0Ot��w���$�D3:� @��Qv�ԅȓ6��\���������2�L0�ȓ��=��QF� �R(�xt����<�Ʃ
%l�D�6��E2L�FϒN��O� tǉY|N��r�X�\��"�#D�x��FN<�v����ثl|���?D��p$E�,e�l�a�c�;`�Qk�"D��zE*��I��G��3�	�9�!�d+rd���$ �})�P���H��IX��(����������$���J���I~��I��
�|�����C&Y��b3D����U8w�jL����/��	��/D���pY�<Zp<�R.]#!����� 0D�<r�Olq�P9�`� K	8�d3D��°ʛ�Y7�}�DB̝A��\ڂ!,D��Xb(�R��,!�m�S��L��*D���B6Q����`���\��<�G�:��V���ꅦյ@,�#�	� j`�+D�P@�È�jB������
��Y�3D�P�A���WD�qږ�\=<��r�(<D�Љ���r\�\�@����G�6D���`Ֆ}��B����5�O:D�xiD�	4=: Xpk�1��ٻ�.7D�tqp�_�un�Y)����P�@���'D�� |\q6MZ
{��-�*U*
���3�"OX��� �%�����RpJ	�C"O�
%KYy�T��v�Z�oQ��AQ"O �+��R.�|��U�A�fc����"O���h�  2�`c�gF+jQĈ�"O`M��苬C�F�H�бh�6�rԓ|��)�9Y�ahR��5S�9���H
�rB䉽�j�Pa�	i�I��']�n⟜��ɟtDv,[���r���C4��!F�C�	#yHh]!���AllkQ���ܐC�?�V��@j�UC0�ц�U�H�rC䉢D3�u!r
��cM� �H�\^C�I�}=��:7�C�W�!B!E!��O�=�}��E�T�q�h�:\��6]W�<	�bF<�΍�ՌֶW%>�9��TI�<�C��! ��zp
�3I�j-��\o�<�C��)�ʱ���!���󅅄U�<� �9��%�K��@c.�� X�<1��J>���x�R��Y�"�Mo�<A���y�Q�W͓w�캥�ex�`Fx2$�>����F�^:���d��yↀ[ �����sD� 5�D�yR,��n~F�h��8I�]���:�yR@�}~<�v��6FZ��hac�ybW��9Ҩ��:tR��03�yLÂa��qF+K�0���'E͗�y"C�7�x}��∱�Y�q�7���O�⟢|R����W�(�ȗ�R�d����{�<�d� �N�q�ɒ�lo�!���A�<q`jRC�}X��[�А��X�<%a��X>(� I�sB�%�c��{�<)�.�4 R`Y2�Y dպ1:Ad�R�<�D�}H��.xe^��Ni�<q��+>����@<@��C��c�<y�KI�yJ�c������a��S�<��/M�[_���(��i���K�<QF���^{�Tr�� ?'f�����G�<��a�H����U�R�`��%��H�<��d՜.�dE�7�
B��9�0��_�<�g.�;V4!w��; �|!0�U�<�6�T	lY����Y�m��p�iV�<�LbC��BjM%� �"o�M�<!��Ώ w8�q�	F�-b�{��`�<QĂR�z 0��d%ݾtI���r�<ׇU�Ef<AN�;E�cw�Dx�<'��q^�x��^>x�<��s�<i�D/;ʱ�2�<k��<p��p�<i ���ƭ�2��Q�l��G&�Bh<�eɫ&+��`A܃s8��fJ#�y�)��r�%g`�!r>ΌR�k��yb� u���b�	L:|eI��X!�y"9"�Ð�,?�$��L1�yRa�RH⳩G&iJ�c�o�0�yʆ^�p�a��#M�I���y�DD��e�0��'QMf�t	�y�)�4v���BQ�U(�Ы�Ų�yΈ)h(��[S�J�"��@J���y"LH�G��Y �*�>!�v@�B���y�eK&����`�ʴ��#�Z��y�䓯=��tj�)S�aQ�F��y��ժf��U���B�u�(�@NF��y"�Z���)Y�}�~���ܽ��=q-On�� by�M5&�6*l�|AC� ��B��1{Sjp13a�a���:D`s�B�)� �0�q'�mY��²/g�L��"OR1d�S�2g����"��h0"O��`.L:�x
p,ç;�,��"O"��ц�l{�9��YKk�u�"O�d�`�w�F��U�ܠqM:-�'=�ā�w�&K���4���I��Y~!��P�H�* "P�]���as�"��!�D�7tt^��̆�2��tQ��ף&!�d��f���p�N�,����!�d�[^4 ���y�@����К&!�L�9N �"�6��
"�N�[�!�$қLN��eh�\$�h"Wl:!�DL!�>@��N1>?d���� ��)�Uc~�k��U�aL~陑�W'T� �'O@1g$Q�z�*���c�=TD*���'��r�
�1öE��NԧKND��'���z�!&rD�` ��E5d��'�l�Cn^h��9��Ӯ=�$ ��'7�{�-[�J߆R�I62c�}�'�>=�6`t�BP��\	6̌��
�'�a	���b��x�Đ�'���2�'d�C#�ߏWc���ǀ'!���'����Ak�,<�;��"�x�2�'���[�GW�q�U��.?����'�x�[��_-^�
�%�w��A���yB� I��1`O_	�e��M5�y��)A�ne�s�ѾXy��<�y��L�<YJ̰��4l���9#�[�y��6��X�o�`ArZs�J��y�ߑ2eT���R�J�����&�yR�̦i{Vs�P7J�M��,�0�y�ͪ�\AH3���Q���ѱ�G	�yBFú�q���*M�rL�s����$(�Ƙ'$��+�#��� A	 6踚�'��	�G�#F��)  d.o5X��'�� 2��U���Pz��	m�$���'��OU�6��Y*B�ٙR>�a��'D��b��������6CX���'�x�ao�vh��0f�_�HP6�q���d�3��i�a�3"_��f
L�|��	۟|D{��4
Ѧ>����� âK%F��y�^�d��Q�r���*&����P��yr/J>qw�M e/�x��E3��Q��y��Ə~��	�������5�����y"h� =�Eg
�n��mⵤ��y"��J��}�T2��A���\��y�×�@��CD�ץ7��A�#!N6�yn��#j�*6+��?"~� ��  �y�K�2�p��ˋ-��QA�,�p�<�R�W"7AT�Rp�)Znn�Cs+�P�<�J^�L'��!��t���#QT�<q���Hidp�mV�Y�xw��S�<1�^C��P�2�R�+)෭�N�<qu)��q�<0"�F�4q�Vx��FxR,Q(:���d�)�0�R��"�yB�I�-��,�ț�O=N�`Wk���y2��6
R���@T<��W6�y2�	����,��b�D�����y����"���g�6/(za#F��y��F�)�|���$C4Q:r��<�y�JЋl�Dy�g-ݳ~YD�:g����4�S�O�����IV�^��
��	%��Z	�'��� �תb	4�IN��=��T��'@V�p�N��������;�:�{��� �lI�N��L�-�5�S�]بJ�"Ol����Ӆ,���Rdb�1bp"OL9�U�G�Xg8��B�p�ȼ�"O�p��mRgT���AP�@��Ի5"O����(d>����5�6���"O��xМ �X(�`FR�CH<�pQ"O�$��;e��l1�k?�Ȼ�"O6�pC
c���ZS-F�3L�S�"O �"V$�:���J9hI�"O�,�"C�/LΘYPɘ�M-���"OLЫ%	�>�B��Q'�,﨩a"Oh��ľk02�isŎ'.�ܕa�"OH�HL�C�=��d��|�K�"O@82�* H������z�)q"O��a���%ߘ�X�I���
��g"O���wk�(]�������.�ҰA"O�1*1��p��Q3�+
=TB�B�"O�(�7�YKl|q#�E�VI�Iҥ"O轱ՄG�Q2�h�tˊ�zG~�Y��'@�'��O�����3�b��3��?K6!�>�(�6E�Ysp�(�텱 {!�Dɤ2����8U��S��"!���"0[���j�$GJl �-�!���� [���]2�Y� �[n�!�G�?J�թWi�w%�%���^"X�џ<E�4*ѧ5���s��wĠ����x�A7���V>Z���0��aO!�d�T��1C�,<�6���K�=>!�D�Bz,��!k�(~�v�hRu"!�D�Y1D��'	Z�gj��I��)
!��q)�,G�Jd.���C6(�!�S3�T�H�8D1�f�.n�!��$o��4	JM!�$C�k�!�$T3Fd�)e!��m�~�SN6[�!��nF�����h�������Nq!��D���t/�HZ��nK\GB�I�8���v���l=�K�F�0C�I�R�*�*E�� �4��펑]�C�	�3��@��	rjiC����2o C�I�D�&��V����e3֭��-��C䉰;=� C��>N��*�-�7��C��?��,���#N6�#���x۸C�ɬW�m��*�_��\�d�A)Zd�C�ɨ6~�Ո�� `�^�qeGݩW��C䉢N6� ���v���rV �q$LC�	�@ՠ̙V��2��$+��B���.�X�Q��ω$����A9xq�H������%A� 5+s�Ր(����|n �EAtI���qv����L�ٰFѣBHNLk!�[�����/��"���{)v,C烐�bc�Y�ȓ&�XS3(Gk�̰Z�	�l��ԇ�81�i�1��*mV�9��K ������K��^�����n��n��(�s'0D� ���C�sTDk �9(�Z��1n.D�죥B�-�T%x#o])$J�|�'#:D��H�.�7/�4;��'δ�R�K8D���$� Z�cP���P���&c4D��ceNڼl��Ѓ��:�p���e5D��y1�0���2�D��:A�3D��:�$���`��T�H7+���Å$�O�ʓ��S�Obp�G�¥e>��A%i^y�"OF��ѠM]V�p4�M-a�$q�"OE��Z�|
���}�Ԫs"O� (9�@jF<f�P�:T��\Ά�SA"O�Ͳ3�O'}F<����9G�&A��"OT@ۤĀ6=�h�M��O��a0F"O I�e^�Pc������-����FQ�\��Ii���QC�M	:h@�alƔ6�NB�'~ƭ���k�N�	��n6B�ɗQ�(b��m�HwJ�c�"B�ɲ���2pI$awn}@G���TB�&87�p�R)
�wN�˖��>*�fC�I-�X�I�����iXW�*zB�	�R�B���
�	��@�d�ݛrB��C(D��'Ӗ�HI�E_|�XB�$z�1���1#�ɡ0JX�a,B�ɻ?v�ɠ��V�4��y���[=�B��:Tl�L���_�@}�=��aY6t� B��
`-�iJ7�9f��9�'O>�JB�	��|@�a�=jq���7b�q�0B�$�!2RKS�	�qKY�쭘 "O�Ix�ƳGA ��l��/��e4"O���Gc�~yR�3D��K2fu�0"O�M�A��#�� �Td��8��b"O�a�C�1C�\��-�M����"O�x!�c²�NlJ����i	�"O:�9��T0$Q�c
Ppʾ2�	~�O���j'�Ӽ5��9�
OI׶��
�'}^�J2m�P�`���/U�>��
�'i��{�h�&ݔ�eB2^����'��Y�ra�XH�aQ?W)�Q"�'���Za*�Q��h$D�(S�����'	b��A�*q#
�����z	�'ʂh�Qo�)�,%ʱ�~��iA��D!ړ(�-{F�J�N��Ih�T�r�=��'�4u���c�yq*r&���'?
`��{<�4��gG�d�!	�'�@Y�또s��q�o��x��'��EC��/hx��*�!�+�d���'�,	S�L�9uo�����ā�'�
qC��8> �8s��)CO>)+O
�O���yrjV?�tlHF�2N<�Pr� ́�y2��S;z!e8D�:��ɱ�y�#\�������e0� ��G:�yr��4K=���\	���W��y���#�D��D�H5qL�}r�a�y2!A��\�J�	�c�<c�������?��I�6cX�؁LZ�N�N�Ġ�V��'�ў�>u��'�._~ �����%e�$yЄ<D�8��Њe�|3�a��A� a�8D���3E $w�=��C��
h�P�P�8D���V$�_8H����'۲��6D��P�i^�.r|)��S��\�҈6D��TeS�28�ÀFN�h�c 1D�rg^����\2/d|���.D�pD
T���ի�Gu4Hqa?D��s'��!���h�j�_�&\�"F=D���&��t�֢̟[��-��<D��c��THt���M"���`�:D�\j!͋~^�$�aaLO��P�K8D��!HPNT�L���5#Z`����2D�3SBW0)s�m+1*��F&$�0d�OΣ=E����0B��yQ ���c���0G)Q8!�D�J�A$$��V�`��J
!�dB�r�F 	ҦL7&�1	�eS�!����D  � ΋$�t�'B�0!�1T��i��ɢFՈXY�'�3!�� F1ّK�'J�̫���mKt��"O�xY�KGrd�!�L� ��XX�"O�q�󦙓&:���#&D�~���"O���%�V���I2D�^�T��"On��$̞�⭘�oލRT�hӄ"O�8�#�L���3�I�B휤�"O�u#��^/t����L=G.�$"Ol���	icF�2��"���R"ODX³.h&)C�K͇I�`���"O֝b��W��pi:]��MC�"OTЛUO>b\(��h�/SW�9��"O:HPsA�;g&(J�œCU�]Sq"O��+��,N���qT'ژIL�@T"Oz�
F�#p$��F�>P3��3�"O2DJ�E�S���$��R �|��"O0�P��%7��Y�fH�b'�v�<�s*ŗ>��qqG��D�ɶ�p�<�r�
�(J!��(�m��$Kk�<��a�8�`�� M�s&�h�<IC��>L�x$����8̣��L�<)"��8Z�!H!��� �qb�H�<�q�E�.��S
�>�H�xS�z�<1!�=}����A�:bk�P�S`�<т�d�P�C��>A��=`���Y�<������)w�F8I��x nY�<�a
�<h�:L��ʴF>D��E�X�<Y@�PVAB��d�[X�X3�Q�<)à�zx^�qAj��C�@(��
U�<�G�0:��J��۫Ժ�TF@O�<�R�[�B4v��=
a�����v�<���� �t�*��ȅz"�a��p�<9�+�KlF��� U��֭j�<a�L�,Cu���S��L� $b�\d�<ga�:��ԍ`&p�yc�f�<A�`�	^h
QeR��Hp�l c�<�Bg@J�4�:w�ȅ77|�q��Eb�<���S�-ص�&:Ir��%�y�<�$�����0"I
�
�a�Au�<�Gb��u��'�4X6�15��w�<)G�ͥWVZ,)�B��`�Y@�C}�<!!�ʍyEbE	s M�D�Pi9�%�t�<�잺3ظ��E��R��I��.�v�<�1 ��~E�|���C1�d�[�<���;rX61Z ,��8�|=��%I\�<�cˀ �L�J2'Qf����ì�T�<��X�Z�$����2FN�<���I���[P��k5�(���[L�<i�Ύ$�j1���	�
ap��HG�<����*�x���� �Ȉ�&a�{�<y��K5#�B	j�'�nL~��3�E`�<a�k	N��W�?3���� (�Z�<�T�)(D=3BٻN �(Ig��|�<���ކ��� ����e�`@�<)��?h��Q�oW�2���@y�<����"@�>�3��>7����l�~�<Q�K��h3ٸG�8>{�s�H��<�Q�3�,��B���8I��U�x�<1��A
54�q�󤝻��f��[�<1�e0uŸt����V]���2�FX�<	��Vn��S�!$v��QCLT�<���A����ՠQ:�����z�<��OM���`�ߙ&� ��N�<�fξGEz��6��]�	�6SL�<���	#K� �)T�J}��s�N]a�<� ����^RC�99u�G�w�@�C�"O9�� ��I��j�mXY�T\�"O�,����T3ʅ
����"O�PI��fSF��w��P
�"OL����ՆizZ�"�EGu�I�"ODiѣ���k�9�3�:GU���W"O�0�D
͏g�غ��t��@�"O����WPa���׊rǬY@1"O4	K���K�^3��ѵ5ɈܑA"O�͡��	={p��d��=��\Qf"OpU�tmV=s?2uz��nVQ��"O4���؉1�u�E����*c"O8P�-�T�}:�D�
�&Qq�"O������$!s$�����"O6��%<��5*gl��z�)�"OY�a�bێQ�^	e�=X�"On�i���9|xs�H-l@� �"O���Ӎ��x���K4��;,_�8q"OTL��敐H?��E��a��2s"Oʹ��g+��E��"��`��ܺ�"O�Րd�ġk�ș�����c����@"Ov��(��U�B�	E@�(���"Oh-��M�0c'i����"O�5ʕ���j%Y `'íC�T��"O��(��2à�h��'.�Y�"O�)�
���]��b$^>�t �"OH��A�\@C�: ,Z�	�"O��h�)�%>�"��ޯ{�A��"OBa"	J�z�͙-C� �"O�)���j�%c��C*0:�*u"O �#�[�}�9qaR+Wz�є"O�S�lX7j�BL�F %]���˗"Ozx�uZ15���BU�w�H��"O��_&>�p��FQ�$ߐ`�"O��)rlOq�8$`a`�V��y�A"O�!0pl���6ْ�-��-R�"O���7�M3��ঌ�#A\�Æ"Ol����fk�,�K�O�`�v"O�a�?M���!��@�g�� �"OH�j掤��Հv���a�lQ�r"O���5G6p� )��;R >̂"O8X���3j���J�tXy"7"O���'��I�����-l��`�"O<�K����ʲ��7Ơ�v"O|0!ƅ�� b T��R�"O��	u⇎XBU+Ů!ؖ`�"O�Q��/ÒR
R�: lB�$vN��"O�qpGj�0#tl��LŞD���"OJ����\�}�ڵ�M��)3�"O����&IVĬ��J_�CD|R�"O�	�ĈE�*��e	�&���$"OX��tO��"�~��]4W#r$#q"O��HD�'�~��"�ؚ#D3�"O �H�`P�:����5^a�"O8s��-J���A0j�6SE"O�q����C?�-��$ǵ�4��"O�����cb���i'�x�W"O(Uh�@���fk	%^����"Oz���D,	i���B*Ō|����"O�P�#�UX�Ԣ1�S�f��h��"Olz�Iҩ ���th�[��h�"O����\�S���7��o��z�"O��[�+]��8P���!���5"O�� �>y�JD�mE#�Ip�"O� t�����SM���O�_��2"O|%���HK��0k�	+Ͱ&"O����ҕx%�U��ߣA*б"O����ӊeu�8�ʏ:%:���"O�]��߹ +D��I�v2���"O64(E�ӣ"-��O(
�~)k�"O@�9t��: [`����Nٖ�"O��1̒���m��$��ic"OB���`��={��Q��0m�.�q"OX�C�E�r~������1�P� �"O"L!w`�p���kf�~����g"O,�&��RHB������"O L��>M�!b@,O)$��2�"O44	i�.͘ ����MؽYG"ORܸ6�˞	&�yF#��]�:X G"Ozݺ"kM�}�$R4�K�.��E*P"OX���Tc�аD�J5�x\0�"O6i#�.я4�
��֯g�>��"O.Q��[� ���>0�`d�R"O�=�6�ռ5I�X��
���"O�M����'+�ԉ��V��*Du"O~is���=���Q��1r��*b"O��5��"s�qbH�;��`"O`��V�Ǩn`(!�;`�<�g"O*�+�c >0S6��E��� ���f"O �`��� O>�`���#PE��"O�)(���*4�h�fC�3r2v!"O�Y�j��������'tt�� "O�yCU윏p��Xa��O�,|����"O��J3l��x� �&Jt]��"Op�׈����hԪF��@�У"Oޱ�sB]����8T�j�9r�"O�� �N�u�jlZ	_X��5"ON5��Nyq=z��X�Nm:�"OT�*����w��C�Ɩ&�^�`"O6�q#
?_%�;�ûzt�$�u"O�A@u&ˣ�$I��׃7�V��G"O��Q�����KR�	�|V(��"O��چ X�AB�]�^��!"Ob6f�_*�"�+ݛvUН:g�'D��MHd:h��v�ǋ5̙�'�%D��n�,'.�jӥǝ8����'D�؂T*ת)�܌���b�D����7D�̛%�\�`8����ID�rv�"�L"D�h*7ؒ)-�52��h��˄a"D��KdZ��Z5� �ܔup����>D�,�cA�~��	
�;ۚIa�h>D���b��g���烌�H���yS�:D�p0�×�ht��
v�J�+��(c�L4D�H����l�'	$��,�E3D�@�.�0!ym�Y،$(V�>D��d�d�� r'�ˊ`�� x�a=D�\����fmP<"�nK'[-|hq N/D�$��#R]!���.\�H�@:� �ɀS2��W�
�R��4Z4��C�ɬ=Ơd��ي��QQ�A��v#?y�,�'�h��B� <���A��H�ȓ7�\�s���X�a����Eu�'bў"}Z#�%���"��1ɼ��� �h�<��Ĵ#PH��G7a��� h�<i1+Q(6
5Z�nX�-cp1PT�e�<���X�sP��C���|T�d�q�e�<�����e$���o�x�x�"�|�<I釚�4�����g����aQw�<� ���g'�.�@h��_rx2Т�]�PF{��),�R9 g@0t�����ƳK�!��@�/�(
6��n����j��h�!�[�:��Ӵ
K6A`ⴸt*ǎg�!��ћ2��Z�'��+,���(C6O�!�ć�a��:2H�C?�T���[�!��ěs�p@jR ��{��ߟy�!�E�Q���s�ۊ�5!!��.8!��@�gn2�i���Ij�����<!�"�~�*g*� �`qQ\��'Pa|���7��xs�-��u�d�C� ��y2
V)k2`�Fɜj����3���y2K��7Q��&C�cU���aS-�y�-��S6�Q -|`�ђ����y���;i��ڷ�H!Z7F� rlɩ�y�)\j��q�2O�Rja��NJ�y�$	�$� 3`�%:��� ���HO2�=�ON�X��04�}���_6�0�'$})�M�	|��HaE[��l�ANL�<9�#̀VhppS��e.�jRi�KX�P����5$���OL�n�nE��IO�H,���>Q��U(aD���ưR����
W,�',��'�I��O�Ĥ �ԪR�\t� KX�@j�(:
�'�T@�WC�X��8�i��^A��0����X������y� ��E�~��e�M�*�����,�2�p?��O�(	2�A.TdT�`f̖r�&��"O�`1C��XP�u��eҽlF����'��a+��YF��_:��n_.�N	�O���d�'Ĵ8��������$	CE�y�቎Ejl(�cO0i��zVbɖp�.C�	,;������l����nG�)vHB�	�
l=P�'d�d!�O��:B�	V����@^8�1K�aɆ,� "?I��)��@t�5�p��+`�Ԉ*7�A���E{ʟ�(��S�Xd�T�?k(��� _��F{��)S(`M�p��Gqv���E/
��ay�E�*�qOj����y����5��0�v����$|O��C���r�h��c�p��"O����,�N,��u��������"O����-v�4T�3����!�6�i?��E�)nZk�(m�̋�Y}��=X�ٚz�hC��1Yæ���!˾p�R%�g�[s�bC�ɇ6�R�+7�>U�N�P�X�Ɣ���.}⏔���m�:z��qP�dO��y⇙'�8��ѽB iFN7���򤔻���O����� �����sL˿f�q�'�Yr��V�x�(-�4j["���J�4l>���3�~FxR��:�R|�$,ۮJ.� �c���Oz�E��@�JĀp���U����/�b�,��p?V�8��cdc�7[�8�VHX}��7�S�D�|�@��872�5JSVg��kY+�HO����).��|�A��0�FA#aKߗ9�<����Oq�2��<��J^�b@�,Y�l��|c
h�UaCK����>�ʟ�Tlr��p/��;~��#��C�<��o29��u��#�dy؈3�z��0�'KL�ڐ��4o�m�J�y�x5j�'3�+2��,�N���! %���'�PW�� 8�J|JIۋO��y��'t�As�D�3t\x�4읊LX 	�'sў"~R�CZ�2H@s�$��s�
$�c�c�<���	tJ�X�4��M
�M�b�<���ȜxV��7g��e���I_�<4$�"��aڕ뎞\�V1AHI]ܓ�hO�Od���Ί�k��)ycC�J�v��O�O0��� D���>N"��9�Ȝ�B����Q��SX�t1� ��2�"�rD΅-�l`v�8�O�OP��eA��05X!&ˣ!5��Z�"O`�2�9ZNb5"�D*c�0e�x���_�Km��	�d�@A����d	O!�DG���� -�Y��y��M��9L!���9�4�����"e�|(�E��_Q�p��ɚO�"TyR����=�""�8�f�Є�I,
��l�$>bq*��W){�rB�Ij��i��W�Hd9���fB�ɚ�
q��I"W,���������$7�S�O�t�n�F:.<�oZX�i��"O"X!Tm��t�X�%��4{�� "O��i���N8��gL�bT:�*v"O4�g�>������s:dx�w"Oz��!/�R�8Y��V� ۣ�$]<���D�	;R֘I���)G�@y��@ E_��oӸ%��M΋;?���f'��,lHrS�HD{���Ҡ`��lW����$�/>�=�ȓ>��=��h\�#l|1�&Շz�x��ȓ-��i�'ƪ|ڴ�Ч&��\����o�y^���͹jI��(��ĭl���ȓ�>��V�1J:�y �W'� �ȓ�
aa5�	\4aP'�Y&t�zцȓ\r<90n^,'��) Dg@�\���>	����D�c ���nL��R��F���y��B𰴊e�Ҧ"F �ӑe�/�y���.��8	�a��l����V�$��>��Oh�n;+P80�ҫ�n#p�e"OUr�IN*ba�mJ�
ǎ8��2C�u���?���wRF=�N� :ؤR#b�9}�M��'� ���e�4t�f,h�D�@�۴⑞"~nZ�l�V(���N;5QD,�'�1C�	�)�%�&�Y�lt`�uG�,��	:�MC�1�`٫�f)m�(I+3�ӆ���'�x��)�� B�A!A�Y>�� s�_�(B��&n�=A��[�]�)�#��_��7=��I s�T��~&��ƈ*]�1�E ���.<Oң=��F�+S*�H�F�,/P�I6�p}��'��\��".`(��eH4��Q�
�'�PB��]����T�J
�'

[q*�2��e�E���J�'2"�<`���$�t����!Iq�<�S��ؐE�T+�Yf�,7Ȅi�<��#�%e A񭌒&�`�`!G�K�<�G,P"��f �/r��ìLF�<�#
� p���Gc	�˜ap�=D�TC&��(/�aT�$�R��9D��9&��N{d��qvPT���:D�z��6Y�$��ǮG�6p���:D�T2g?i�ГЅ��D`rC6j7D��Ç�,$E���(�'$~��e8D��a���-JM��'�@9!TΩ���2D�����ϊo2@���^7Y���9v�1D�@A�� 2l�lD�p� de!+0D�H�eB3�b����[?�BA`�,D� �A�öU��q�aM� u9Ґ�#=D�6$�l5�T�s� ?$h����O;D����+,/^,��Q.ۼ3� 8D���sh��x��]�!�3��=��+D�H(V�O�)�19�Gf�:�'D���" 'z�8�%��K���#N&D�ܘ� 
�/kl�pf�G�UJ�� #D�d�C�T�L�hR���g�$���"D�� ���>R�¦��(j��Qc"O8=�0k�������s?�"OF���h��B''ޔa  ��B"O�ݫ���:*	��)W�.hܔ)�"O���FL�*BL��8��@�S�n�I�"O���2��(G�l���p��`�G"O��O�ۦ�2#H^�3��]�P"O�	�̱%�zL� ���%̶ňU"O S����lB���VGODaJ��E"O�tk`�.U��#�\�e��"O��6��+5f9;YHDaGN_*b!�$@�n��h&���W�2Yqb͇�g!�DɏWQ0��o��|{�˅1,�!�䖤.�ERЩ��@�ke�!C�!�T86ňT�����Bm
�!��?V���g��>ko�����<t	!�dTl��9�N��pg���-�8{�!�ӍG�i�ˀ,TO"@!����}�!�B�B�y�9Jd��+f'�!!�D�7>扺��(4QN,(�`ٛ`�!�<V?��р�U�n^T��F���i:!�$R9-�l�:NU*<[w�02!�Ď/	\2��:4�2�̑�E0�$ĢT�6��Q�R�4��"�#O���F'U+3H�����7��}�'L"D�,Z F��\�2���) \F���l&D�Ĺf��bQ��� bV�h�g;D�H��%Jml0���oT6��`b-D�\g�ޡg�`��@l�
kL�̣��-D�ly�>?#d�yV�wg*�(B�*D�$�&�@�,��D[Q��[:�(�F?D�H��'�1RcV���L�>e����!D�(�Rd�N�"�a��cHp�<�`�T�@���(­Z�4T��O�p�<!��r�>���Ӎ4}r��t�<IG���c"4m 1�
	Z��s�nOH�<�g�5Ȭ]�1O�l<�����F�<y�/�6aƴ�@KI�^�Hl��A�<!�5Y�{�f��uC�hJY�<�5'V8����hM:��D�AfZ�<�!�X E\L��/��Uv��D7D���D�B�\9�1��A>1��a�E4D�`����;Ҋ�G/KI���� �>D���Ơ�<���2���1y"�jfM8D�� ⅊�B�2 �$cǡ,'�D�-9D��c%�5^Hz��ӕ3@43M(D�D�cӜV��9��2�x8PJ)D�к�I53?���R#�:@�X$"R�)D�L"�� E�PŘP.ݭo+��#D�����+V@����)/����4!D���"��j/\ +g�ɸ�����!D�$�D�^>c�薬���F?D�8;w	�"2��-)��/*r��rǋ D�d�� �8j&<4��F_6\j�H<D��zm�9HNU[G�a�Z�4k1D���SB�+Y���(��1# ���//D�P*����n�hgEB<H�"�1D��"'W#8�	9EGݽpG�1�4�:D���dM,s�HU��/�^4��vM"D�� e�Ν~.�i*�CGB^j�:u�<D��I�h�9)F��#�Z�v�"u�$D��d�#�l�de׮(�p�e#D��`��
�]�����4�qh!D� *1O�{x ˴�G/ $�S�!D����G	V@r3�}���kV+>D�� Dp!�Ȭǎ��CC�=Plqp�"O� q����}����&]��x7"OL CT��3#���n�;c�\�"OL�k5�ܕ�DlB� W�(�P"O�� 'F0n�`���X�EI@=�"O\8���M�a�@�^JAX�"O$Tqt�\g�]�ץ�, ,8L�"O"`�Mŵ# İ�0��yp�/�y�&\��<��Ϡ޼��e�7�yb�ץ	��H��8�b�J��y��OI�}Q�	E�9>�K���y"bȮŊQ��&(��bӧ��y��ݲ)�"|S�m�+.a�d�3@߈�yBH�5T���!(��49�&���y���[S.5Rt�L/_�,D��"�&�y<X�ִ�2�	�{ְc��y���	R��3%��1z	�a�E)�yH(��(a�Y�X�Z}�D��y�lJ�:!x� ��Ҥ�Xe���@��>��C��'���Թs���
�N��`�Y��� kS!��X�9tF�K�@��k���4�T�EZQ��I�E<;pB�G���O���}S�	0Q)�
�y�ό3g�	7@U�r�~������|&��sP��O?�I�q��,�rϞ5������Z�y�&C�I�ik>�cፊ e�qb�7�2��9ظ ��&4��z2��<^{&�ӳL�U�QB�A��0>!�h�	h�#�$�^���j#��C�x��3�͏y���ȓ|:tHȓ�Cf0@`S�l�BGx�힉g�j�����_�O"�=�SeK)j'`��@��P����'�4��j�p�@�I
l�
���/g�� ��I��	!Tӧ����Y�t�Z��AΓ ��p5�Mi����٣u�2�����	2�i0�	� ��}�l�@���c��
��H<RAG<H	b�4�l�
ml��.VM!#�g^|��SE]x)�B�� x6�C�,y��P'��p���(�����:����Etx�!���7(x�m�^�µI2D�O,ij�"W�-ܸѥ��&A�	�d�&���7L��2n�$Y(b�aW^.u]*i��N� Ȍ��bw������|��5ۂO���.�Ac�:�>��'(_�,�$��*2>�1�#풚���ς;�(5ۡc^ӦU�;7[��I��׹J��]┏A�V�B���	>�V�2���ge��k5�3E����ĉDp&��pe��ꥇ�!F��X!xh�C	�rg���gY#@��d�L~�%�C�EjU P�T��S�ʺ�(O�������y
���V�@ș�/ʻ���B�5��s��?O��s	ʣC! 1k��A?��Փ� �>��j,�Q������ J�K������7M +� i� �B#���qL߿x��,��� ��<}��4�"M��>udUaӎ�('��3ʞ8������W0�Ɯb
�!ޜ,3�J�;~�`�U)�6%�>dC"-ȱV��d�#%_��E¯B4#،k%�M<u�`�5)��#�*L�;=Jx��۪�.��sI��f����	??�d;�n	8Mv��ve��q"̨��O���rt�jP�p[wa\�(H�
^*AK<@�&�I�t:��� �C�S��Z��'oN=t<�+�.9�4!�?�eG�$!\�(e��
~�H��֌Xz�yR�OB���t�ʦN9:Q�G�J)N�ȨI���K��6�'(�"D	�	�1��3�p��	��X����]I�VuP�J9�U+2򤰁��H�\m  �9���>	�WE�tt�|�@� ��ASGBυ�r�)�+6#�@��YtX���&�A(�$�ȳK��-#R�˂ɔl'�j��C�:�J��"�'�H����0����Ś/&V��'��D�d�?3J��;�@0�l�ߓB:�@��O�O��6��0j��B�ĂN�$�)��Գ��F,6H ��
�4w\!���>Q��4&�<5DI�3�]1q��D����'���"�'͆}b�F���+�nY�V�iH��C�͊9P	�J�����q��'���	I�uRF.O���� SkN8\ވ�D�1}�s���E�7��Z�:^?����K�& Ψ1���0?	�″c�@��6�/S׾�ʐ���<16��>hv��:�yZw��/,���E4?ygc��V}�]R��p�t�w8�xC��S�:��d�,�D8h"��6��ɡ�W�U��'n�=h㣃.h�����SD0���f2Q���8�K�!�d�#$1�	��eB��8Dn�+o��4JJ>1d�ߪm����'Z`�LO 44
�z��ˣP��s�'<D�CQ� �2�l8: ��;�6�#��;'T��)� �����sP�y��T�|�<�8�"O|��SC�I��uS�Z4;x�=�0"O8 �!�<v�ԙ�N�4e`*���"O�U;��Ҋ Hy���ʗ	�%�%O��ӫ_�C�:Tp�P�qϪh���1��1��sfa�`�a_x0C0�R9��I�41�q�%@F�	'tX��S�P�R�Z�Ɵ�B䉒NyRxZ�	G�d�$M�B֖Q�(ʓ��=�tZ_@)���3�'oLɈ��l&2H�$T+lM����3�XX
�S"�Zl�ԭF��@8sE%#>��E�I�bPҐ��r�3�����=z�@�X$��5,��-+���DE;!^�˦M�~IҊ�-QN��b�ĳo�����O�#�z��D�./��ւ�j5��!h�6�ў��g��d¢���[�t}Lz���|2�e��u�\�����u����o�<ck�4#��q�۸h*�ӕ�	�&Ă3:�l['B�'z���TF��H�k̓iP4�p��()�6nW�K�!�DJV�4i�瀨#4#�,h>�d��M �B@��1F���Vӟ����P�>&��1ǜ�	������|�>Fz$CT�+�ҕA�O1/֝y�Q���\�a�� !����=I!�6=��8%�7���qd�y�'EL���58��x�"�1Թ�!�D9�R'���}�DP�����[���ѢEp�<AcnZ�'D�s�M^�U�4�xSH�/4䬩+��U>2��9e��1�p�z3�;���[4fEą�M��@N
�y2A7K�
��d#̎���M�H�\�N��8G^�Qb�	�K7�<��O�1�r�	�n<TM���T�\��p>1 �SvK�|8R�Za~^�!gֈ|,32�_�FQ��p&gTw/p�p���q���2#�K;{%~|1�O�5U'ԥȑ#.�;�
S)˺x-lTm@n�^�{�C������+T��3q�R�#6­c��X�<���']�^���)�5P�r@���e��뗪s0Y'��\���w�Ͷ�H�k,؛D8�5"Rj\
pgP$ ̛N�!��Cz��!�C��"�h�eF+z����G�=�i
�Ҋe]v���]>�DxrMۛI i��/܍R~�����?�e�75=
L����V������
N�lB�j �*|��C�N�!�p>�$�A%�|��FQr��X��^Z�'d�2�EC�6� ��ď�>��� 
@R, &b��6nH� ��lF!�T�$��H����.]�$�/֮L��	�Z�xyҌ�Z�4���`���A&��Mn�!@��P�^$�C�L�"�Z;Tm+��O�c�2E�T�!}B�E%��i�}&���qONH�`��s�X��h3@�<4��9q(�$t��H�Œ8푦� ��L�Q�'K��;i{<�a�� \�?��y��'���ⶦM�{G�<Zr�,?h��'[F����	\����a�% �4I�'�,�;���1��m�p��H*�%��'������W�%:�i�SP^��'��	{Ǯ�j�[O�9��I�'��r�%!v2u)��+�'��8��`�@��V�M�m��X�	�'���u��z�l�bG͔r�(	��'^��/Ub(@��H�(>� �#�'��=���� ?l����+����'���+�#LhK�*��E�#�����'��J �P���tR��<+���@�')`d�R�<#Q���&�\�"
�'wv�G-��0����ˌ�\R�'?@]P� ��4�ӭ�7} �`�'�l���a� `T)�b «h!	��'���H�G�#X�v�����P���'e�p�t��n�zI{�#ȴU��A@�'H�0��ȍ�W����A�Q�BĲ���'*sd�^62Z��9qHL�d]��'hՋů�FH���G��R���'��D�I�Qr��`�*�����'Ƅ����[� �ndZS,ĳ
����� �����#<\p��@�u8���"OZI��nb����:7N��&"O}7珿���31�,A�u)W"O�庄h�YL���Q�"�*�"O�ę&F�%���P�@5�$��$"O`�Wd�!$�P���t��.�!�$J(3�6��1�L:u�Փ��O�f>!�D��l�ro۾:�Y��ˏ:=$!�$K"Q���O�;��GlƿN&!�d�Q����e��/r� -����!�<zF��c˚7����gMزtx!�:m1�i�5o�r��=��]�~!�,&����WY��}Q���`!�$Ȫ4ռ�`��Z?8Z��;�LPo!�$�:`

	�ŌG�\8mp��%>A!�So�,�[���:J4�Qʊ�E�!�DEi�m��B0z'�%"ND�!�@�o������8���Sb��$x!�d�6pn��Ye�:�v����pT!����� ��և�"5=.!I5g̓RT!�J�o�!�&�B�MJ�	�0_!��B(L�%j�BP�l� '�$TO!�Θ`5�H����W��]@H˘ �!�H�b�84)S)~�%ch�r���b�<��F�=�Fx�v&�v�9`�	F_�<I5 j���3�X=欜�Ө�U�<q��=�~��e�κU�m�&��V�<i���M 	� L��c��#!�Pi�<��S���AT�W>1��WD�'�!���
f��:�����I�����!�$��}u"�R��E�a T�"�a �Bj!��ȑ�(����٤~�0X��U�^R!��ʐ�P��,�:����P��M�!�D�V���狑Cu`D����t�!�P)�p�K�#ŧLiP�R�R<D!�D	�g�X��KR 5�s�E�|!�d�?�����ꎜOj��@IQ/|!�D�7��ٱf�ED^p�A(�E!�$�_�¬fƜ�"���F�n�!�DS�������!� !���з:�!�dL3}����\ah�`v�Ѫ!��Ķ	$>$���U�a���ƍJo!�0`0!�7lX!S~��Gf�0zS!�d�)���o�r8F�ce�Ӳy�!�$�]����Ҷ?@�E*��1�!��;tѬ�@��իn\1研�6�!�$ǹ7���w�	%g�TLZ����b�!��Z�p{g�)7�Y0m���!���8=�´q�Q'�I�e픰M�!��(:$-�4�6 �R��3!��E�j�hc�	�l�xx��<4�!�D�3*���rg�0�B��攫�!�dQ3Z+h �MՃ_��D"uD�(�!�dM�v�^U2gO��M�
����Y�:�!���<v>�y'�>�v0�#"�-�!�Y/
^"X8F	U/i.����ߍ.B!�$_lK=#$�,�F�����n!�ĀHK*�"��A)T����ԋ��g!��?}�iHGoO?C�rMY�K'!�DO8����L�-E�,Yq_)@�!�I�37��!cΏ� `�}�t䂶x�!�D�z�L����,niժ�j�"G!��S�h����ɼw�iC��j>!�dÂ 찤��'F(Lx��Z�FU�)!�� ��s�I�%pV�!6��RSj��#"O�m{��=Om��5#WiH�8�C"O�h	Ջ���mGB[:,I��I"Op�X6�uyL�J�̡ E���'�����H�ݪ�Reh_��Q�'��:�+96Pl��.�7Gd���'6���U��L�ҩɵ!B8�(%r�'�~�4EA�a"��E��b)^���'*�L�ү�4I����X�[��%y�'fiz4j�wi�l�1�2f��M`
�'(�3�N�5-V�#6(Y(T��s
�'<���֊��\ ba�jzԠl[
�'/~Y��l�.LW��a�E�2|ZN)	
�'����ȝB��Q�-�<ga�1��'�l��Ԅ̋!���Q�!N�Y#�L9�'�i�� V	x���:��[�MH�'-�dZv��	[�*�b$+Ůl�B=��'@�X�s�Z>-`E�f���$��'�0��3GJ�Z��yv��x�.�K�'�� �˟w����(�t���C�'D8�:ǀ�Iz0�ktIY�E

�'�⠃v
�	J���ɣW#�r1	�'��ͫDB�/87x2�H�H|���t-���O�pa�K�I0�0B&<d�C"O�� �5aR<k�Cۣp��IT��S��u�O� �qc ��cak�q�
���'�H%��J��/|`��:�n��T��;���ۡ��w��s��&�:�H!�D5`]�(���-D��bf�L K�6P0��Bx���v���i��>�	��'Z2��d����+'�Z�BC"��`Ќ<z��A�.�Rp*t�M)�Zm!�8:Th����\�<1� ��=���
"5׬]���A�'r�k�. 3t|��E�D̂!b�,��� 2`�{�D�<�y2U�� :�e�Kˬ񨲆P0q�Z髷.	�6]LT�O?�ɴ>< @V��j0���I�r���$Z�?8�`��ԄJ�R��Dӝ$�z�� j�G^JE�ThT+D&�i��x�P�W(�H�<����\�v�9�.4��F�J�'̼���c� �z�)�d�qZ��ǌ�%�A�͘9�D�cw�:�s��d@G���<���S�L@�I�r�P�# ��)���w�ʌ��!?8�Qj�R	�'@z8h@��0�88ڦO������a�G\��Z��lX���	�f�
Ȉ���!��8���~��*���*�z������gᚫd���2�� ��4�A ���Mc�w}h)�E��n�� C��,AF)I�Uܸ!���\FrU����h/�!���=�M(Ḑ<� �&b��>�����cQF�t�sO�k(�9�3�+�I��Q倀Y�*��:�h :VB۵Xۺ�<��m��T96��<�pj�ڷ[߾�ӣd���92���#�Ғ}ߐ 99J�c�P.8"9�wM�|Fy�.Q�hn�a2A���0L�$���H�q�F�% �kc�N1n�x������'i�n��d��k]�9�.�%�U�#�՜`�ؔ:�E�u��(��?�O�eb�cJ�5�������(��A�Y�7�0X ���M���p�C�L�}"K 4���`	��2ܻ�4�|��(�>J��E�4��ja@�� �'��5�fFU* `����.&b��6BC�m��M�`%�i�&�ZBF[h(.Tæ��Z�1Ȇ�ү%e�!���4o��Oe,���H� f�y�!�<%e�Y�u��L>(�zqұ)��B�ڶ��|@�ԃB�v>M��E�Y��x(ƚ�oQ�:��ULV��ݴ��L����@����O-!�E�D��}�1��?l^��S*gLBt�Μ����Ӷ�λ=�91�)��R��+2��p�v<;2�\�,�f[�S��A8��G2!1*����ג��?F�T�sE���@˄k�81�d�T��TQ���I��:�I<C�X��E���	��}���0<�2a���C46��dSLP t��S�M�P�LV����F�4�X����p�/I-p�j(�D�Nׄ��O�c?M�p�l���r�# �R�2��$]̲���&|؎��H*���#�T�E�
G6�ȉ�>��k��t�>�O.�i.���^�7�wꐑ����e��	��o�D%�禕Av�$W�)S���Hw>�p���;;,pe�\��a~�"Z�O�)�m��9q��K��6�y�$� �Yo2�i��ƈ�<v�-�'�@��3�K!_���
J�lp��(�z���r�L��M�5/_��sa�O�Y
2,��K,}�V�y�xh���X>� ^�gH\.E��pF	)�~i�E"O�����X$:�b�e�#v�z�b C����v�r�Jp��x�D�c�vM��F��l%��RH��xb��'M�|m��A����}�f*Y�u�4��f؟H���	9�9��DV'x��(D�H��G�^���s	�j&����'D�(�L��R�D!g���I�(��I(D���&Y-mk�hJA��FҤ��E*O��L�!�&��s�Pu�a�P��y"���Zr<�#gU��&�
�*^�y���Q鮘�
^���2d>�y�߃%�a�K>�"�/�y���JRԑKT� �R�ċٴ�y��0s�1�j�-�L)h��8�y�D"Ѡ��N�7.C��GZ:�yBLظ*�
�Z�扚TƶU�2I ��y�
R����
Q��<�y[��Y��hO|��tb�!�H���Z7��7]��s���:H��3"O2���X������	�:|����i����S�Y:\ɧ���&#�4�`��� ��g����Ί�yr�ųj�B��f�\�z�J
�~��5p�&�҆�b�� �'M*c�0]���"I��P�"�O y�� � ��Y,ÚA�1A��W�8��q#d��%�yb��i��M���N�KM0�	M�(O��8�(�o��Y���N"��h�@a�8;\�{��{	��'��-�r��ec\Mr«�
QZ��橝#-���;^`XbJ�"~�	Y���CЏ�tے]�6�҈�4B�h�yp�FϟSbP	��*U�{���	�7}�rC
�$T�az����E����J�<�l�%�\7�p>Q�%��v�� .��p���*z9�<���
Oi�C�	�qn\{�F$���@%F�e�v�<Q�̗!v`DS�#&§5!�|��e�Ei����\�7�
Y�� Y����!v�ڈ���ܓ;8��o`3���n[�)��ѡ�'��p��{����&vHң�?D� Zc��b��ıE��[�q1�<3��1T��dJ�Ǻɧ֜J�a	 ��.�!�D�4�8��1�^�c
��Ԃь@�!�D���|��/���$������!�D� /V�9��7�XIzҬ�C�!�DA�:�~Y�҅�66�} ���=&!��>��\�3ȕ v�b���'�-l%!�D�+f�̳0B�.[�`� ��7s!�$$U�Z̀pN.|��\HK\'7U!�Y%�l�s��`�TG^!�dQ�E=����c�Uj�L04��3bY!�� �v&�9 )ԑ%jH��KL!��Ã=� �X��� IJd%��I�C�!���"*ry��d_�o��\��G�2�!�Ă�*���Q�‫E����`��K�!�d�[�(�c& �>k��S gQ��!�_'TT�*0%�E:H���l!�dW[���0r����3!�D�:)ve�fe�r#"����R!��<f��J��DJ� ㊙ZF!�$8?�����ǃ�4�=bqiA�yM!��ש*�0E����+6���*.L�!��3*�z�s��
O�`Q�&i��j�!�Dܓm�X!�Gfʿm���Q.L6T!�H�"ttu�t�k�N�[�-�/Ge!��ƌ,Ø}b$i%����+�)X�!�ă d�P�v����j�)�/d,!�䜥L �S���!>�dep����,!�D�Ζ��A�X%{�����6}!��9)uFt㦅J�xQjtAB����!�� �}��c��B!w���L5j]�"Ob]!�m��{��U�N�	*��Y�"O�}c�"�;{v����7?s���S"O���)�>|�e!�lF	��""O�᫡�T�N�>!�RkBl�z�b"O��9�.�?m��YJ�m�p���S"Oza� ��: �����`�X9�""O(��DE��Ԍ#f-��w"O6��U� bY�T�Jɸ0�1�P"OH�s�ǓC�J-�ȗ��t�;"O��p&J1D������A:M��ڧ"Ox�P�bޠI��yP�ΥzB��+�"Obچ�_�@��$s�iHiB���"O��F�^$*虒�J�+d�ar"O�8�
� �졑VJ@,;���b"O@��@�RG.AAR)� \��(�"O�p2Th�$���cÆƎ;Є��f"OR4k���*��u[5��ո�R�"O.��I��0��pn	�t��q�"O`��e�?7 >	��\le��"O~iEJH�
AB��tM3@��hG"O�My�I��|�����#z�,��"O��H���9M�P� �P|`�"Oj���$Gal0�[u��~.B��5"O�@���#F�dM� K� N��r�"OVye�U(�y�!
2��c"O°yw�ԏE�h�0�TEP�"Oȝ2�#K�O=$$�Gi��A���S�"O
y���(�Iw�O� E`��d"O8���@��5e���T(�z6T%�e"O֐�s��D5<��r�Χ(Q��<O�T8�#��-x�@�aѦX�ȬɃ�I >C��k�H�A(��8�bC�ɛS3�� %)$> 
�pQ��:8bC�I�g}�]���������+�N<C�I�T0�0��0vv�r�l�92VC䉤ꦴ�g'ԎGd�B�V5q<JC�I�s�q�j���Qb��6\Yp�O�Uj��!�)�1{X��[��_��U��`A8;l��~Dp�z���)�-/��1؁gI�;�P��ÎI�E��*[y�O>�Br��(�M�f��K�l��g#�@	�����h�<i�'�nD
5�Ou
��*W3<��(I�����xD�@��~Be	ڢ��>9�˧<��e*�$_8xh$*�� (R�+��'N�����""a�ڑ="N�?�qb  ��Ppq��"�,i�c(��R���M��*�"����M�F�O�z�S�^�Q/>�b���,@زĈǹe��1��ì�M��%�[�����O
`�E�Y�����Tk��ض A�[�h����`���C�&�	�0|��Iŷ
y�����-W_:��� E�m�Vxϓo�j�z�ӿ9R���?�}���6��A��5���T,�Cy&]�lG�8��o1<a����y$���X�����y�gx��I<�2��B�SV�H�Ӥ��}�T�#2�	HA�-�$�ѸM��O����ӲP�&L`��V@��g��~�v(EN�D��Z��.��M׀�+�n�Z�($�&xAt�O~��AM�$>c��A4E�?`���&)ys�h>D�H)E�)j�����;o7��v)0D��
�GF�4Ȳd9eG�#��	 O)D�(���
}�B��s۫]�Ze�Rd(D��Y�(���!�s<95H'D��ï�6:A䠓��E4k� ��#D�$��M�~��"��c����`"D�̭<\v�9��#&�H�I3떄�yA��f��%,%Cp��2%��yr�X���Ae�&^�m*����y��p�z�as��68uq�ٶ�yRf�"{ܩs�o�����h��'�y� C&D�=P�	��������y
� 87�P�9ꤓ�մ(�`+�"O@A��j��r�8�B�.U�Mk�"O\�$��:��2�K�NI�#$"OLq����g�bY)D�?HG��8�"O6��v`L-I�����6�ջ�"Oj��΁8?�բ���}�@I��y�!Bޤh����R<�}S�c���y��x��(�!�x�
`�g�yb᛽T���r�� %t�&N^
�yB�Q�_^ ��J��"�|MhѧS��y�\�o}���U�/J�L���y�-�R��`Z�<(p��w��yң�8a���z��D�+���q"��yҎN�(�FΚq�YC'�ݶ�y���7���F}�d#'�ԍ�y�G�^Pư�S�CA(�D���yrJ�
V.����
�2k~>�uF���y҈ �]*г��(Rz����V4�yB�P�EKd��$#I&�<
�M��y��A� U"�a��C�r���H�DN��y2g�]��#��(a��I ���6�y2��_ J�HOK�R��5+Q`��y2�`r���阸L���V��	�yB�(]{���dZ,q�F������y2BA8򰤲sF�n�l`5"� �y� �v8X��m�:R8���ǳ�yb�	��ᙖ&/	d5 ���yR��PQ8���Ό�2�Hِp)���yr˂�4��5�fa<'���Ҍ���y��O�x�Sag/$��� rKK��y��B>�Qc"�O�-��Q��-�ybh]�4ȸ �tg��{34���o���y���M��I���2MJ!$�8�y�ʫq�ƉC��NE8taiD��yRNK[��e�
u!]X��ٲ�y�����x�N��p�X,8%��&�y�(��kvp�*Ɇgb�$Y�+B��y��ӊAb%*�n�-���0�ω�y�Y�@
�E��(I<-/����O�yL�'b�����p���#���y�;�y16cI�`��������y��
|	$0�`I�6G�X�W��9�y���.MQ5Zj�FU�
ǥ���yb��T���`gV��y1I��y��q�R="V	[����)�y"mH�`�p�@ͮ�ȴC��D�y.R<tnА�*�2Ĉ։�9�yBi�I��HH�� �n�@�B��yBd�+JR�<�% S ��D#�����yB��jer�(nא���&�%�yrL�:9�~�c��&��ѨVV��y"��-��
��$m}腪*B�y���9*-�E{�҆fm"�5cK��y�C�`����Lذ��%]��y��\�w��q�Փwo��p7�6�yb- ]�^�6-��aD*(X'ŕ�yn^��1��@�"V�p�(0 ]9�y�g��ICK������ ���y���)��Q�:
i�y�gDC�y"��z���"�n4ɘ��C0�yr���G��ј�ぞ�MS�EN��y�D�R��1��&�+t�\|����y��B<�hZ�.�s֊�FHA��y�+KVš"��3l�`
��.�y
� ���E���CA����.?�@ A�"On%�����uՒ8Xd��<s�ޥQB"Oh�@�lY�z��`N;K. �Ф"O|4��!9�jX�sn�y� ��Q"O��xG�T����r̀7:�S�"O��Z���s#a+|1V���"O�ѨB!��B��[������"Or��e���T���6+����&"O����Z,Tؐ&��EwT��"Oȑ�Ń�4=M\��N��}�^9aV"O*�*��$l�D��uz)r"O��Ť�>:��!5�W�Ol޸2�"O4c4fD��$LC%=h�� &"On�ЩR�7`-V�=U�y# "O�p��ۃRw��KU�L}����B"OꌑŃ�F��# ���5C""O�S��	�D�a*\_넍�"O�;0a�9 -�͛"#@�.H�7"O�A���-c������	w)<��"O�i4��*p��UX��lG4�҇"O�̹Al;p8�B�Q�u4\�Y�"O�I� ��)Wfd93�S-  �"O8��L�O�2LF`�;x���)�"O�|�GGGJTp�ˆe��i�"O�ZF��1Py�xZ�*�/t��"O@�r/̾?<��`jF�}j�!S"O0��aN�<N��
�N�Dsl"O4�q1��0$[�<Y�Ρμu2�"OP��q�@� �B��W皬�DY�"O�}�E�FS�IƸQ�fE�C"Op���*1Qκx:B��-d4�"O��q�I"��@K�Lϡ$�P���"O����H�H�`%g��J�8re"Of=x�AF�$9�Ez�c���@	)�"O¥[��Ɛ �0%e$݋U�V1jW"O��:��j�x�!���:xZ���"O���2DՋc��x�A�><t�x 2"OZ� #%ύPk��)����v�6��P"Oi�(X�"�Ћ`J�  ���*O�@�Q�,$�iHt�y��}�
�'���lE(/�B�Uj�T�
�'"q�F��{̨��,W�u�x��
�'�B�x��<l��hr ��ef��
�']��s�����К�'V��
�'悵(�Y��$�3��%R��!�	�'�	h���Dz42èZ�H�ʑ�'�}����J�s#��)ZV�
�'d�dC'
Z�q���B�J�)vЅ1�'��]��Ĳ%*��ʵJ-R���'y@@��iB ���	q�k�'$҅:�%�=v�N�q2��:
�'n�@y�eI1�й�W��8i���
�'�fͩ���i��LC7	�9��,i
�'d��"P�G�s���+G�9|UT�+�'�Z��⣞�2�<i�Q�^�r���
�'wZ�S��F-_[��X@��,��B�'t-��� P5�B�D&fJ8�(�'�5�a�0X,@�Ы�XA����'e�1�&�׀���I�T���I�'�fM�q¨w5h91VdF�Z�j�'���[(Nϔ�+W��H:�((=D�t����?�4�T嗩&���O:D���D�F%ִ�sKS�&�h��f6D�� �/��HeE.#���-3D�� 2�y�D�) �X� !�S D�*�ye"O������P���T
�b�teA""O*��%�{�dA�H��H��I��"O��f���|�BHD#��)�d"O�a�"jF�rP��Aա�*��2"O�h��K�A��B#� ���"O��pdD��`4�7X�L�0�4"O��ꏱ`焄Ѡ`_# R�(c�"O��:cU��(�#���e�&���"O�d�g��t
���6��?��@�"O�$�3�� i��8j#(T�Y攰�"Ov���k�|��p��N��$
"OP�5��# hm�Fh�/��%"O�EsC ��~+�Ũv��$g��`"O|m�'��?q��А�R4f�,Q"O�𡰄�yVp"6h]	S��h�"O MC�jD����ƈ����&"O��;��vsΜ��V,} �i�"O2(�$@A	+�1��Az���"O�%`1l(����V �m�����"Od�8X���0���@�h٫4"O|��͔=g��8���O1aK"O�lIJZ
-���w��p��&"O���T��tv�	b�b�FFEK�"Oޱ��
��P�툵��" "OD�����,�����4T��T��"O@{"��6�.ɢ��~,-��"Ot}[��ت<�����$j.�`"O���5��Gh� #֢Y�c�+"_�<����Oe��h�oB�uA��q��[�<ф�H&l ���D�M;W�,�p��@M�<1�*k�&�r�j5ID��(�cGK�<�a�+�n=��
1�ӗ���<���x�4�:�۳u�*�s�I�g�<9@�F�V�`Q1�-�~�;��Q{�<�j@46/Z Q`��L���u�<Id�T�]�r=�C!�4=�x��G�z�<a���>/�I�U�#}��Q��z�<!�K�a
�Q[G��
J~��%y�<����E��%c������O�<iŇ5{(��0!ţ)f�aX�BA|�<���+}���7 
�)�`��&J]�<�#j�3h ;�!�rfި�Sg�S�<�"�,/R��Ì�I�N��4I�<)Β���P�1�C9"���2,�F�<�p��$ٺ��S?/z��BB�<QEEϫw]�uۂmG)"f�%��~�<�n�"/��ܐaA��*��8�u�{�<遌_���2��O���j�@z�<�ׁŝJ��A�K�o��:c$y�<QŇ�O�^�h��CP��F�|�<�'��D����`�8+�ēQ�<!U$q���إ�Љ
hRT��j�u�<��= )p��>p����v'_u�<S��(O��@�U��<CI�$��JPq�<�Ē,z�u��	\"@N��qw�<�bk#PR8�if��q�F�����q�<�VJ�	"�=:�j�=s��yH�U�<)6�Ǆ%	 �WD�:7���2�^H�<��o��;���:@�Ёh�d�c3��B�<�gE^   ���'�� �E�"�#����Lp��'vd�b��?;Tℑ�/	
G�T��'7P�e͑7d)�q�V�MR���'|6�����$ ��3}4�a��'���Z�
Ja�LF�y�4�
�'�q�����]��� ��jx`	�'y��1��hWfI����&[�z�'�*�"F�'@,����LG�&�<�@�'�}��FKF�A����U�
�'7�x�ĝ�q�h��a
'<L9��+<O�e���S�4��T�@ 9�t�A"Od��F� /��l
��:�b�B"OI9��P�k:�Ɔ�+/;�t��"O\��6H��n�;1�]�}2�	b"O����-O/k8&�Bs�C n~���"O�h���/}�P�ԫT�L1���'9��ps���R¬���F/~Qp���D�s�<�!�:'�~��6玟?.$�C�q�<!�iUv|y�2/��Ey��q��k�<�R��%��L��$UD@�
及k�<� ~�1ǋ>XA�8"�%�!�ހ# "O���(��,�DF�!r��q*C"O�
��2T�E�S+������"Or0YS�Y�s� qDA$8�� "O��gMK�l/�b�b���rl��"O��AB�Z�PT���lI�-��| "Ol�8%��{��2G�i� ��"O�ڢ�ץ@������#cv��q�"OFt��k{�Z�!!� {tΠ2�"OBE���S\U*�A�o����"O������9���ᄉ�%li,#B"O�qģ� � 8B��K�7T��!�"O�x��q��@���!�R���"O̜S�f��Vq��˟��u	�"O�(�(��7����-��I��"O|�����[�|�%�߄��`6"O�U/��q! `Sqb�%��S0"O"0b�d�!m��� �9^��h��"O��JV!*��U`2��".�����"On��vfJ�M��9y�fB�i��1"�"O�,3.%
��e�% �t�h�"On����|1J�d8g�v�9�"O��03�S���lQ�H�E�5�v"O��(+��rO�`�\N�^��"O�L:!싮{�r!)�٦�+&D�2dG�uB�ɵ�\���Y��h'D�l�A≽E�ꈁ�ޖCd�P��&D������2T'$}�0i���ĩ2�-?D�����/�Fq����4W��1ȅ�2D�(:���:Wo�����E�kŭ5D��XW&�lF.(q�B��j}f�-D���uBY44n�L3E��/;��@�H,D� *`/�!}=�5�ٛ'��=��*D��������A;w1f���#'D������)�8Lz�iϩ(�F��$D�0�&�0H��刢 �*���"D��2� }^bXz���h��ബ"D���TL�f��:$�Ǿ*��"4A D�����#�9x��ڟfg()k��"D���v凄W��I����[^D<p�#<D����.�G��T�7ED�Fw�p��%D��kē��>i��`B�
d����o D�\�f��'�Z��q/�f�Ny�b�9D�Dzq��?BiD����&:�BR�5D�hA�#���	�)�'�ƍ�Ud5D���/Ґ<Ւh@b�9u��	 �$4D�0QPC�v�8�*f�F�C��mz�M0D�Xb���NC�H��!L���8D�:D�����C;��d��E�+n��J'L+D�PI�a\<lܨ�B� v_p����'D��s�ȅb*b�ps&2'�J���#D�L	b��7&���Z
'D,��6J>D�@��l��s�a�#<����<D�`�I�s$��`�c�(Kc�<�'D���`	��mPX�����(�Z�a֌*D�8���ȕ9�H#�F��:V�<D����^�RQ�C K7�̡�=D�$��`��b�mIcd�5۞Ѫ�#/D�+��,n��k�GE>�b�	1D�,`Q�2A��:u��)(K|]c-D���eG'b�0땏QrB)��C/D� t�.^�H�2���J�6�+D��[��T-��II��~��9)�%+D��R�H�	�vm����d����(D�� :1���L�����J-]���j�"O���4gJ�g����F)f�H0��"O�䀄%�	N�"����%!��b�"O 9�P��J6�Ԡ�9� h�"O�͐���?Q4���i���:��"O�\��⓹r,@	<IAP �0"O.��FhڨV^u�@��w�L%��"O�t;䊖%���[���1c�����"O���/��P�H���I#��hw"O��`���L��_�f!��C"O$�lG#6%@̚�ƒ�Ru0}S�"OX�c���t���!��Qmd�r"O@Ź$��j�b@zĕt3T{2"ONp���*��8��%^up]��"OX$rSϚ&U ���� �u�ɪ"O��h�HÆ	�ݨ��]�Cd�%��"O2��J �6��X� �حj9J��"O�b#
_t�d�+J�n(jU"O%:%H �v^���/A�~gFQ!P"O�x�g�5����ͲPR� #"O�$��%�A=ՓSb�!M-.�bc"O������+���v!��#(�lx3"O���EX�<(T���F6uPM+�"O=ꒀإXr�`1SI]��{�"O�IR���4�����ʬ	����`"Oʘ{d�E�����U�H ��"OҔp!��" ����֟,7|j�"OV%@�B�5	�H(�Rl�7�@�"Oز��zZ����jF�E
l�b"O�p3���zM�1!��6|�Y&"O�h��T�Gez8�7e�g��5"O�iC�
>ʀ�C��$�DM�"O(LJV#�-I�:u��G�x�aw"O���8��X��Fr�����"Op4򇎛�6��Aˏ����"O,�y��S8V=���!D��P���"O�Q��A�3~�T}���1Gt�x(�"O U�UME��� �Q4��
�"O����׃up� �c�]��l���"O�쩕(H�i�z��E�ة�Q"O�P� T��#�D�ح��"O���R�9p7�a�TX�w�H��"O&m�gO�n��8��̡k���"Oб�&h��] �Ӣ�� ��D��"O����U!'��:��l�K�"O]��a�}�޽��@�"�(�S'"O}5�q@@�*`*ԅ�T�"O(�)B'��I�(� )�
�a�"O׏��Xu��C�-Ţ�I�"O�L �kJ_x=i6���Z
P�q�"OTLx�)S�(p3�,�ZT�"O��z�hJ9��H�*ǍL��0�"O����\�>�(�)[�t�P�"O�I��7u���8�Ɂ�i��%!�"O�͒cĈr�
]�w'E8g��Q�a"OL���C�sk�����	�����"O\���"V�T�UhY%�����"O2�F��BY��aW\��0+�"O�x;��_��p����itn�@w"O�p@D`��s�fpi6O1up� PG"O��r��O����ɉ�fU`�y0"O�)���'WN���$��O��D"O��:Uĉ�7��{3IǕG:n���"O�Y�a���@���?(���"O� L9�!L�-J X�g���Ta"O��ycN�FN�a󐄔�VJڍ�"O�l�o�mp|�0&��+\�@�"O�8�7Ƙ�L��*�b�.����"O`@wH�� �x�rp�Ɯ��"O�l��Oϯg]hKQ���e"OfM�#΍�AdX�0!g� ZG��4"O��0���Tm`yJD��"~M��"O\���.Qژ��$�(��ݙ�"O�M�2gM�.A&� %����U{ "Oj)��e�6v�|Cv�Ĩ֞�B"O$ds��+W-�P��@��f͙C"OhX�
ȟ_{r`p�@���2�!"O2���� L��ܨ�e�/a�V��"O��+D�sP�ٺw��i_��"OԜ�j��Uz
F��}ґ��#?!��ձ,{�qa%O�&���j�/¿�!��/&���:b�h)8�8#���!򄗎8D��*�Lׇ�9@T�F:C�!�dY��J$!�B�,j�]�K�ws!�DC,���s@cZ�+���� m'yc!�Ý6���׆��ы�(_!��bŚx���/���k\�0/!򄐖|ڜ͑��ޅP%�T��j�$m�!�A���9�2Ʉ4")��I0�!���D^ d�(>zdhX�刀�{!���I|*9�I�,bc�eb�NX~e!�$��� X���ґO!�+C�^!��C:lª`s�"=5�ѩI�?Y!��8PM*"�o$FYH�ʉ

�!�d�@tzu+"��#y!z���iȋi7!�䂣�Fȳ����=�E��8!�$îg���A��[�z�!�@j�&R%!򄎗MFd���Kצ�
��f�y#!�$k���a7*  ���խ"!�؄{���Z��U��ڵ�n!�����izEiۂ� x "ο*�!�$lh=�d���(��1��T!�	{B�cBK�G�>9�5��u�!�d;_�t"�J����,�		m�!�B��t�Ӄ\�'؆�вg��!�$@;J���Sf������4�!��zV��U�H)U�<�x d�%f�!��ߥ� �BcYg�dE*b��3K�!�$�-6*9�����E�^mJ���8�!�	�o/�����Z%Ɣ�be �"�!�̘�^��w�;2�p���o��l�!�d;��8rqL�4�j�a���0I!��L�h�y�)@��L�Տ(:Y!�dr��0��1+�:!X#��?!�:����w�̰�J ���Ĭn"!�[tݮdB&Nэ-@�pC�G�5!�ӶtT�!a�k�=�-�#Q�!�d��3>v��U�̸i�깃��� �!�D\�SP�
4�ʆX��p��a4�!��9I�@�׵9ΦqQo<�!�$����O&Ǆ�xnթR�!�D���N8��MR.%΀J� ��W"O���`��XxL1D�3�i��"O�I�te���D�B��$\����"Of1�f�"lNH�06��.�����"O�qR5ԢM�q#�O6�:��4�'	�ہOT=R����7	�;!�D#VyzP��%��LA+%(Y]�!�� ���b�UѴ1�ffȴV� �{w"O��J$�I:g?}S�/v%��""O`Z��̊W�~�Pt���PM`�"O�q{bo��"��Q�W�	:La�"O&���Ŋ3.t�с��hT���6"O�u*B��MrV ɠl(UI"Oz ��l a�ڔ.:�X[F"O|쑤�� |j��
�c��)�p�"O�ٳr��$�*�1���:^Pb"O�-���Z֚	�Ń��|ؑ�"O4t�L	{P��`���)�v1�"O��ÆO ��p��B�
�$��lp�"Oz�j��
\�P��DKՂRxD���"O"�ag�{��9��I�vu�hx"Of� �Y��(�*BH�"��0�"O��@��Y'D��=�����	"O���7�k�/�3jV� "O������V���Y�¿G����"OJ�8q�IG,iZ��Ɏ*N����"O��+Ҧ&^[|�8T�ҥ+�V��"O\���.si̤�4� !��<xV"OH5b�!��A�r�JP8�S"O(��,T=���K�"��"O�$Ka�9sp`�)���)S�@-a�"O�ةC+YQ����ON�V	JH%"OTx� NX_��@�r�t)"O����´{�-*r�	�Eb��q�"O@��e�<,4U�X(%!`G3G�!����e`�-aAC��`�!��^:l��R�6@���"�O�!�$��by
=@�����kM�c�!��K�����%�Z��3!�
!���?%k4H�� �˚�'yx&]��3�x��$�ʄ0T�{B� �t����R ��Ɉ�c���p"�m�d���J�
DH���n��͓�H"4��:O�%Q"T�H�*m��c�)�N5�ȓ*�tD�"F({� �� �
���ȓc�bH����R.詗��C�F@��ly���Ѯ�).�ppɂb�c����`�2hu���T�4PYP��'li��a%��e�R���h[V!� ^�H���2i���`�.; �[�D=St��ȓ#�,�V�]�x�t�$���RB�	�2��E�&GR|Q(��V툏?�B�ɪ+��Pf�{ب(��0��C��5B  �C#;�`��EV�4�:B�I�����S �dpD�TN�^C䉿1����mT�Xt`��s��
C�I�A#X���V�I�:h�jM�]��B�I�yz���WAзIj�H��g���B�I�&�}�M	���VJ��*LhB䉻!قƠ��m�r�r�~B�I�4�4�(��7�6���]h�C�(o㢩y�F X4P��3�+-U�C�I+Q�);�D�4 �ny���-��C�� �|y�D�� Y+G��7Cy&B䉳|´��׮]�w���ȓ{*LB�	�&D����nO�?>v�HuE��Hp�B�	�Zkb̂ S�F�*�I�4�����,?!��҅SPe1�n�o���@c�]�<�TB�5� 	��ι�x�⪌V�<	�h9x��E��2)B>0Ic&�M�<�GG�-�������/$O24�+�M�<� �2���nް`r�� ����"OF�2�_�D�ʳIW.N�f\	�"O���&#�%�Ve�$���;��IF"OH� pBO\0\�[�,S�$��D��F�O�rq)�.�/v�Jdc�H"�'�1H�W�)��(�`�W�
��!�'-���� �*&4TTk��̸ �ݨ�'�$��,ٽ\�T���	ue>�R
�'��y04č%�L��7�ž~,P(�	�'h��D�*F�R�`f� ���k
�'�z0�'��2i>(�E��H ��'�!��O7\�"���@'`	�'� ��DF�6'���Pc[y�P��'%\�'�@'RuP�v��h��'(�[wD�c����8T�Z!�@$D�k����*�aB�N�F�Z�"D�L�V�/f�"-SvE�_`��q,"�OR�b�J%���K� ��Z寙(Q��C�l��E7"L����%Rg )�ȓ\����aE8d�
�r3�
��m��$����Z�\N��� �T�GO����֭��f��@�R҆{Q���!Ir�s	4C������X�^݇ȓzy(Iy I�F��M�W��@&ft��	ӟXϓ*���&ѻp_��4�֮c��� �:��R*¯]ܪ�L�$nLXX��X��9�d-(3H��$� }<4�ȓQWEzkP�4t�]#�T�7*�I��G:fI�F��]�6Y���Ϳ#��d�ȓY[f�����./��{�Π~N��ȓؐ1��5q;&�8��%��3�� �!�M�:[�D7RV��ȓ=��s2��33�*����q-�ԅȓN�b��o|aQj o��t�$�\�<��Ӎ�� x1�g.���M�<�厓.���Y(W����fM�<��ǉf�P �rD�0:�x!�F�T�<є
�1I0�rXQ�İ�o�v�!�ę�p�f�éUfVk���+5�!�$D�$W��k���(X��c��o�!�L�9�<M(��Si�L��D3u�!�D��X�Z���坔e=\QH�'
0V�!��	��0���UV+���5G�!k�!��R>����%FƦu���Ȑ�1!�$��kV�d�	���iG�N� !�DX�:���(gKX>t�����A��OH��ڼĢ�RS�G�||ĥ!�"O<�����N�V�{GL�-7q~U �"O`���|�I���<j �:�"OzD�џi��P@%.R�<aT"O^�0�L@����!	�:�)Cw"O��
5�@' Lv�9�ə4��1�"O�%9,O�>S�Xs!(�>^�V-B"O��!���T�
�c�e��#zѡ"O2IY�VL�*���$<�,,R"O�	���^�$��ϊ%lJ�8�"O�P�7��9h��5+��F6m��C"Ov�����k��@�f[��<��$"Oޥ�LN�i><ey���� B�mk�"O��ɤDZ	5�0Fd��4
(�
"O���i�������W�μ&e6���Z�D���	&,�L8�sjH6hz�p�ȓF؜���	C�F�c`L2	ul�����k#LV�[2,�+n�
���S�? &0��M$&)>�3팇%�TLa�"On���A��n"(�#��|�P0"O�����Pj6q�!�#aĜ�Ч"O���pdË\;v �v�\�>��@�a"O��S�"]�Sh,�Y3/�@�f݀"O|����;��S�_�Zզ\��"OJ��*-���#%��X"O����S�R��S˘-eT�Q"O�X����89d��V� �b"O�	��!ߨ	B�ma���a�e���&LO�	��H�b�>$0Fנf�#�"O8�1��[�MU�6�φ@��CQ"O$��ʏ�?.D�&��H�DS�"OB�`.���`���"�<�*O�9tK��?��A &j���'�,���&4G �*�a��X�'���3��ەkZE Δ�Z xz�'IheQ���%f$Щ�&Kb�d�'6�IH�-�O}R�C7BG�I{�D�
�'�f�Q㊁�d�d�I�!k{ll�	�'��XAd�W�J����dy2��	�'�p)�1�1r�\�����3�l��
�'�n��B\�v�L�$��c���k	�'rLA
0��*s����d�d�E!I>��k j$gM��M���Y��r����������h�%kN
_����H74�t@�O��8W���@F%{�zрu�Ir���Z=5�����%�V�K3�2D����� ژi2��˿�6P�R�.D�T*a̘��D���.h����U�-D�$9��F� c�г�� P����l+D���Ŧ$;��-��\�u��ra�*D�XI�ˑV�|y'�Q{��;� ;D�X�C��ਭ��W��5%'�$<�Ox���K�1+���a#'L� 8�"Op�a@��:\����q�5	�v��r"O�x[U��h7А�EH��¡�V"O�Q�b�]2��S���K�2�"OP\�$�Īg�պ'�S�x��P��"O^��gd0V3�5k�oχP��x�"Ol=1��[bp���مM~R� d"O�$�Ь��(M1 #Ýy���"Oh���L�; ص��c��PX���3"O
�("��	q>�j���l6�鲣"O�sTcC�~G�q�����_6�]�V�'xў"~�K�5b�$]��G/}pHM�҃���y���b�)y�n�u#n���>�y2�_:xx�Д 	�!�du�  ��ybe��nБ���߶/�D�g�ò�yR�M�+����'R!��)�&�D��y�$J�=����Ҭ� I���yҠ���X
�B��B��ð���yB.��L6�����:��4�Wh��y_*~S
����T�e��@�X-�y��ѥ	����6���^VD�h&�ȓ��O��D�O�c>�+��C�Uw0H;�j	�
�D��)D�t�ذ�Bp��ɇ?n��E��i'D�,0�N�#�&][���p9��*D�9�.ݺW��܊D�P���,R#*D��f�U	pSh��͹`�nd��:D��ѡ�Q�@M�%�?:��l��`<D��+�+Y�-ຘ1�!��V�%��Ո���k��=fK^��Q�;~-��8f"O�y	�j��Sߤ1�͖>/�N���"O� 6�����@���2�ýs�M:�"O�D eW����b��C��@��*LO @���5>Ҿ��P��W$�s"O�P�o�j�H��� �q`"O��ak�|�>Is�&��@n@���I��D��C�'v�4�*�DÐj؀��ƺ4�v���,E�My�*ĉHy<A0g^�U�d��Fخ�s3M����)�^D�Ņ�!vt\[ΉB��U)#�W�Y��p����E�)2^*��7 =;h؆ȓ#���l��N�Dc���teZ��ȓfoD��F�q�3�Dџ�l%�tF{����K
��ؓt-�^] 5"����yc��t�P�𠕾j��D� Ǹ�yr�	bzec�E�t6e�B��y��H��2�j�E˦O�t�s,@��y�(̀=�@tI�h�(E|�{����y��ԥm`N�@,��A�|iȢ�3�y���$�q�U*�33
��Q�Hֆ�ybeS).R��P�Ç/L<��g��y�Q�	pDK��ֱ!����b���y�ؾK}`���k_�D�`��$M��y�Ñ�q��萅�7a�fpK���y�k>@<\�� VS���K��y��"r'�1:W%OHF�������ybD#�V�h�ֱ>� ċ��н�y"���@���a��f��nW�X��'�䄣��춹�")�.m��h�'�C�.Ǣ6J�U�*�&g�D�!�'.�|����

2���>Vq�	b��$;��=���%;���y4"N<���X�"O��ɂ-۞	��
GN
k� �"O4	��œDf���;a��Pz@"O����`�{ኍ!�(�0o�N���"O0�`O_Xь�
��Y1Qоi"�"O�EytF��[h�-H��
>,^P:$"O�x�[�P�Ia�ؠ��:�"O2�I�]��]�4f�ָb"O4�XA���l�ZA�ߛ�n �2"O�X�Am�J�p`˓~�<S���~�O�rh�Fa�,$}�,;�LV�e*��	�'y�)��H�A�Z�P���
�Ό{�'}���"�H�%�t�Z�x�
�'���������ag����
�'0h��TJ�r�p8vdϜ{vtA	�'�8R����� ��",���'�Yg�O.hr�; ��e��' �D��L�hL�w�E�@̈Ő�'���
cbҟ7�v̂g@�K3rd[�'E
�JGV�!�������&x�~M��'P0YPP-;�1��;w�v�Cϓ�OT��$�"e��e��o	�̛�"OP%QQ�0J˪hB�ހn�Z}[�"OhM�B�M#��o�<X�R"O5���*`o�I��i'~��c"O����g��A�6}�◿/���`�"O�P�Ԋ\=oS�xg�Ɂ��� d"ON��)�Qk2+\�C@d#�"O�uP�a����tE�uqg"ON��AǃP)���k�`Xbm��"O�lkҠԵ��� GսvDb)�T"O�Ր�[�%�a�`f\:M~U��"Ov�a ��3 �A��F����B"O�����T�#yA���9�L�p�"O� ���g吅��\b�cޞ:��Y��G{���9T�k`�'�.��U�b!�1�������M���q,T�K�!�$�|�r)��	�dPm{�@G5!�K�#�Z�P��O�W��3KĊ�ȓtLRԚ`K�h���C��vV��ȓ+�
��d
нZ�nLp���&W�J�ȓ.��E�U��"�H�QSO(X�Ň�	�<	6�ݚ|���D��%΁�p͎}�<A�;Xc�(iD�L"�<Y�#�x�<�hJ�[2�H�R"<�HQ�2fx�L�I�<9a@�+$(J�cC#_�j!P bGx�<%��c2|p�㜊�l�)�Ŕo�<Y ��6�DT���?j�N���BZT�<q��-$mp�2i�E�Ѳ�U\���̓+8�As`LR//׀yѬӏEʮ��D�Mw�'U��ڄFͣ&�t�ȓ����դ��0����X�v9d|E��S�c&|9��A5GI��g�M�S*�B�ɑ�̴��'K?�>�X-Q�:}�B��z=�0)�Y�m.H��KDnNrB�ɉq{tDx�o͵'���` }�B䉲�<0@GF�G#����O3^%2�Oʢ=�}�b��6�ժ@��zd.��kHF�<��LP'n���RBB�� �d��~���Γ=Z���3�P�^�Tӣ���pY�i�ȓ1�ђ���:ʂ�����"8��ȓ
�x讬4~���+��i|\���"Oj��N�!�j�ҁ�V*mh���"O YqԣG���X9@�������"Ob��,%S1�\#è�~L~�0 "O����
��1? �9V��R;P�j "O�|J5� {��Rn��H2��8�"O.�)�-ƾ/�)k�M�
$�!ж"O��yW$<\�p�%lR�c!4�$"O���ZEc��j��94��ZS"O�tB�#,d\���@��$�i��"O�\{�E�)3�E�A����*\X�"O����-c̘)��
�u�4P#r"O�X��p;�U*w)�/ �����"O��eD�TUl[�B�c/.���"O��I0'� Q�
��v�^ Z���"O��:���E���Q��Nr��Kf��-�	L̓}��h�6 ��[�d0�u��xE�ȓ*��\��"��S2���KT��@��Ɠq+8p�U��KG�8�cMc+>��
�'�h��g+�P��|:5O
�2j���'e�xp��M�� *�-c�R�'4f{w!�-e����G<1�1�	�'�t��bBg���I",E:-|Ѝ9���'\4�B��MS��9���#4D��'6�81EK(:¸�w���Q����'�����B�%��#'�OJX��'R�!zB�Ќf�<{�͕�3�:�	�'Eva����7a������F�1����''h� �S),R�9��%ƺ���'W4p���נ!���4-֡K	�'�97�J.�6؁p�IY����'��ӷ��q�.LrWņ�	b�3	��'�`R慼5��MP�ڥ+�H�҈b�	B~B�4C�XŒd���A���IX��yB�3�� ��4>�Q% ��y��AO�b�c��[�&�f�3���-�yLJΘ�����lbJ���y
� ����������b!8��m�U"Oj�!1�b��tJ�ËI{�(�T"O�!��Z%�^�
pi�2�.$@�|��'���< 4I����~\�h!'�2!�d�Z� <��(�;eV4�@����c�!�Õ�t�i���`�D�B0�>C�!�d0N�d@��c�cM($	6H\�F{!��V�;nQ[�!�65�4ȥ	-c�r2O�A�':ȲR��9b�h-kf"O$�����9���A�Mĩ/�8���"O�4A%��k���Fky�q"Ǒ+W�דLof�0�f3	` �5"O�L�&�B�e_ȉ ��?`�����"O�m��BV.��EB�D�L���q"O�-9� M��$�I�1/���`"O���A:M=$Y�&�L(v���"O(�S����Q�>�8�F��.�T�3�"O���Ğ�V��Eb�B�.T��b"O���$�^&D�m01�C�-�l(�"OrIk�\3^����F�6T��}:q"Ov�Z�J�7-"�M�&���Y��	F>�8�Fy���"�L**��]:Q�&D�� /¹R@J���ρ%e�Y��D$���O���>�r�n�	r�$����6埶�yrE�1>u%�Xw��ȉ"�J��y�JI(_�2��e+Q4�@�Ao���y��,}YhͰ��X�Z��4���y�kEF���X��ם���3o�4�yG�6Jwč���y��������hO���$�-f�b�q&�ڎ~�V�{'�	3�ў���65�6D���
�+�-�PF	�%zC䉣G3�D�r�24�`a��F�Q�(C�	o-l����1m�2�B�׳"LB�	�w� �HZ�_�B�*�aՐ] C�I�O�8���T�!�:�g�(4�B�ɭ��,�(�\�*��5�OUp�=�
Ó���,t2��M�J�� iU CMyr�'�(���|�հ㬚5g�8����yb��5�<
gDM�7����O7�yb��vh�����X�� ����y�DȄAѪ�V$6N�R��G���y��׃ �X�uM�'x���6�̥�y����VyX��t�͂�MF�yb�w�UF�4"B֜�T��;{�=Y�ZP�9rS.&�aS�-W80���
B4-����ôA��I^"y��ȓ�dI9�d��@ܦY�pdC��3$��ہC�S���)�#�C�IP4ܔɃo����!2�_�<o�C�	1�z�PԀT�%@���	3(8e��L](�Rj�*�,��2
��cz�ȓU��W�f�*���E 
����Sq̠ �'T�V�h��]`�Ȇȓ������\�@X9�m��bp�ȓW��0�ă�J��� ȉn�T���:�Nћ�OM	PẂ�n�,hxG"��6Va��a�!*�r��3�^�)�vB�	�������)�$��@�w��C�	G�����HX��T�6n�/�BB�	���d)�O�xH�KIiB�	-gkt�#藤Iy.�����?�B�	�C�P�mJ�=�q��.^�#�B�Ia�	�J��9��1��]�czNB�	�l��qcĝ8���1�[34NB�)� .�`FN� �ҕ���
�����"O�=k��*���*����8`��'�1Od0a�m�+:�$��w��>^�8��2"Oh��Dƚ,�R�s��+x�|@W"O|L{�^"|О]��՞[>I�"O�ևV�]��	�% ₌�G��[�O>�����H�6���P��!?�����'���Ab��x�T�K�:L��e�
ϓ�O��ӥ
4>vI��˕�:�&�
��|r�'!N�P��)Pa0�*8]�2�S�'V��C@.W����c�XH��9�'H��n���|±E��9����w"O�TN�5M�����37��D6"O���Ά�bm� 2&�lp����p��y�d��,ZLl̲��sSx�Y�����hO�c���Où�5��-��T��I棧<9��$;打LNdc�͖2|Ȭ)#�<B�/����H�3-�R��󨜝;.B� �x�hr��&6�����Z�c,C�I 1�� J�&V)%Q�!i���	e7C�I�[�H����[$	/�ȓ��+�B�+���´לn�IBP&�(�B�J��Aר\�4��M���5`B�	9>Q�����#	��"�Ŏ�z�B�b@�q��H)z�ђ" 
4B�I�z6^hA����Y�2��'Q{8B�I.��D�0]��{O�,P$���$?��Ip�â�;(�2 !d_E�<�t�G)BHr4(��m��� L:T�f����I!aP;Y:�,��@9D��(��X�g@���LM�|��R�6D�8	R�o�
��	�	D0���5D�t9��D,v��X���|8��d3D�0�E/�L1�1hvA�5`�j��1D���v�\:�(s�LR�:X174D���0M��'��["br[D5�Ç1D��F���0�6�C��7d*4%A�*D��)�i»���2��D���b�*D�ā��L�jpxXd�D	ۼ��1�&D��P�X�e��(����t�vE�l8D��Yv�\��Ҥñ#�4����"D��K��4u=�4C�*��-�'!D�ȢU+Y w.U#+A2l�^�X l�O��=E��lЩX��0 %��>�Z��t(�&�OZ��dU96�������b��F��8�!���9��ċ	+��'/��!�d�==BY2�֎E�ZQ�$��!�Ғ80H}�V�Cn���3� CE�'�ў�y҄@	va:�
�S�r&ZxZk���y�M�V%)#��	u��� %�F��O�#~�#��aXf%�EI�@=�a��@Bb�<���.c�����x$�]B��Rs�<q�-Z*v��<�b�\)���R���m�<�RN�/`�@�B��ɤL�����e�<���J?�0��e&�ؼ�$\j�<y�ٞV��!ǅ�W�bub��[fy�'�V��CFQ7& �S�̵�v����C�(#��[��M�(���,,�!��V.�(;�T+(�5X��.i!�\29#�"�$�H<FDr�(��g�!�D;"�$���	OS�� �@.pI!�D�3oW����� .���SUJE�,6!�Ā<��a-�4N1h��¦�~!�dE^-�6aI14��&O�A!�� x['Q�P��u�`����a�6"Ozuh%��1:VQh���� F�)�r"Ot,�aJ�	xy:9P��;� B�"Or�#W�KF��ȐMϔk4�2"Oz|�fҖJ�z�	;_�@J$"O�}��X0hP�)�O]5'Id�Q"OJ���:V���`��\�o)~<Pe"O4!�1_m����?�����"O���珁-��TA&h����A"OV���܍W�j��7l�9YH$�"O@|brf�]ò|C+�lA*�Z�"O�3��
qo>��i[`�X�"Oz=Q�N�I#<�1����0�lp�"O���2c����@WHI���m�f�'�1ObA(E�٤ye�s�,G�q�XP�R�8E{���ό`9�Ċ[�䍁��"h�!���6�"C�;� �v�Z�}!�DP�|5��yPO�*�F��D�� |!��A�6���!Y��5��ER�.k!�d��&6��e�
4��37DO	!���l0�ĦR,peƥ�cb��'[B�C�'TQ
C��Y�U+E%�$֨H��	Vy��ɼCu��S�N�xNjT㱁�7�C�Ih=jh�'ޖf��5��U��C�	�M�1j��LBSV\�3g�O�xC�I�HUZ�YAU�D76�±'��	�B�5dl8��F�.f�1S�B�$ٜB�ɤ����C��,i���©^��O�=�}�u�_O�JM��B\��) 0��z�<����	A"���k��KS�s�<Q0�]#\Y�-	\J�l���Kq�<�u�	�HdKw�@+O������p�<��`Z�A����c�� -Q"�k�<�&3��Y�R�J	.J���aTSx��Dx"��9F�����6Q�P�ʊ���hOq���y��ڀ
���Sg�R���5K"O٘��ک �Ls�M��b�N葀"ObAj��W$pj�9�Ӄ`�i�V"O���CAM�BCXlҀR
$�̨j�"Ol����G�Qjl ����`�Ȓ"O�]�7�ϗ/�-;�D�d*謠s"Od�� �	�b�$`D$7b����!LO���&�W+���K��9~� "O���%���U�Hcd�Dz�"O�Б6H%I ����%]���P"Oļ�a��:r����өf=�ԛ�'����R�=]]lUeI֓���'���r���gu&�$�؂��@�'�P�kEM�r���V���l���Q�T��'���O5f��,ÑPRQ�˄m����O ����+���K�H1f�"�h�"O�׉�w������"T�"O�u��'��MP�����2L�b��w"O��g��sS���r�×�\�Q�"O�P#�Ģm)�H��oX8ڴ��"O��Z��8�p��T	X�Hx�f"O\���,K Z�r�Lɸ.���c����hD��-�M��ih"B�Y�l��5@�	�y��N�W�:�9��=_�I�D���y��[�zN�[F)�X,��!(��y�G�1B(�\�֡��S�8$�d�O��y�lY��T(�	�`�����&��y�FF3'CR�s��*Zl&��Fʉ1�?I�'?�E2#X'?g�ɫ��j �p���� -��i<9%f<�b��\;�"OF�����8�Τ�'�Z�j�)e"O��zU�C$Jh�"JL"Rt��"Ov9��N-
�<P�����g/z�su"O�u�fnЯ'3�m�F�G�\=nP�2"OD8q�ހ`;�U���Y/Y���W"O����Ǐ��4i �<U��"OZ��6mC�-]%�Ӏ�J� ���"O~��A�-�v��N}z=i�"O��ڃ��Fj8�K�0 �a��"O�E�aK fhx��A/�L�*LY�"O|M��ɩq�H�`'�}�<�"O0�R�ґW���@bm]�C($��A"O�4��'��v�|�,��%�eP�"OlY@�h@/~]�y���I�f����"O<�s��	*U���  ���w�^�`�"O�dAm�;���
Qb�$3n�Y��"O��y���>�:6�S,��݇ȓCל�����G�����C#~���}G�`�6A�=;�hْ�i1yN��Y�h�vDP,rـ�z7�U)���ȓGW 1&g��� k@TD�����L�bgT-��$P7��N�ȓl�LT��ʹkT�p�Ղ M`��ʓu����L�P�x��B$N�D8bB�I=(eȘ��gI%:4�X3j��ȀC�T͸XA'�?	�H����M�Z�C�I�zQ�}��͞r�D�W.H,��B�$N7��5��J��K�H��.��B�I�t��<��M6&��S�J	l~B䉸p���j�!��
U�� a߻J�C�I�&�@��LF��֐#  �7�0C�	5"C���� �/�Ҍ� c�FC�ɱix( ���1O;��؂���"��B�I�r����F�
]&Z�c��V�{RXC䉿f��	� d��i}�mC�_�N��B�ɠL�"�y!  �E�s��	��B�;Q��t�Ѡ:.�%xg�̩�C��s� �$�Ыh�r�KBK�-��B�	�x���kP'¬�b%pq�a��B��g�uQ�͚��P�@�.�lB��8.a<�Cp$�=M�К�	V�`<:B�I1bd�-P�VYfq��`�7+�C�ɭ!�z��n�#9lz�2a�Ň<�C�	�Wv�D�힛EzP��E�s��B�I�@�i�U(M$q</sa�*T�����Їp��isƕ�H���"Ol�ٕ��Q7\t���I�Kn�X#�"Ox���ܟ}9��o�?��y��"O��-�"f�Z��T�4��(��"OB�0ī�)����1��xJ|�T"O*�0���o���cm�#"�8)F"OL�K�N�.�uf�k�n�c"Ox�(!��8̊<��Q�{n�܊�"O|`[FK��Gܬ��G��/$|d�U"O�m@���2O8\���/�4]ځ"O�4ٶ���s��<S����H{
"O�	�v��j|�q�E�NETi�0"O(b(L:g�
e�P R(7.\�qu"O���҇V(:�a�䮔r�Y6"O\��w��W��Q&DM���a�"OD�#-�+�h���f�:�"O�lH�h����J#�K�l�`�"O8���E*G4�18�j�3&5�;"O� P�	�����=��-F$��i�"O���MTgpd��(A�'��4�4"Oܩ��Hǻ
��Y
�HX��i"O �a���6�F�����..x�K�"O�y��O���
����rN�Q"ObA`�=��"K����)"OR#g��{|�pu@�&E�<dc#"Od]@��?:|��/ߠw���Hb"O0}��9�\!kD�I�b\��"OJ�9����� �	Ϡ]��T�"O�\��f\5z:h�Di_�Y�-�p"O�P/VFE���E��l2y�"O���nP�>� d�Ōh��G"Oh��5ǀ2x���J߳,�R���"Oꍙ4�����M���L?�!�"OXyZ%g\;��BQP����"O��y1Cݣ3"6��E��B�R"O^$A%a�D�@&τmf(�"O�4;�c��g�S4MQ�4�"O4��c�>-�u���#�thja"O��,u��j2hǎ%*��E@�yR�Ķ�>�p�E&��<h����y� �,�^�-� ��ʤ�y��Ƹ>2y�l)Nvf�Ҏ��y�<?ݢ�3��?A����nG�y�˖�]@����Ǭ!͢�cj��y�)��:��}i��}�(�gĝ�yB�U+I��p��0b�hD��&�6�y�c��P�j�&)�Pա�F��y�·�0IF�"t/��,��E��y���,�а�@
�8��M^�y�*	q�0�r#��)Z�n!� خ�y2BʔO�"�:�H��Kй�����yr�֪\b�beoȊm�Iх�8�yRʲm�[Ř�UsX	���
��yr_�5K�z4A�(z�> ��D!�y��p�R�z끿-�CK3�y�*�>��9"#�}x��qǉ��y�EF>,8�xU�V+e�9�Ԣ ��y��I�*�2̸��φ��ᄫA	�ybc�V�y��H�I&NTU�H��y�F�hJ�%
pbHq:��4&T��y�)���h�B=A���pS���y� M{X���팊<�� [��3�yrE��`��G� ���@�����y�8��D� o	I�����o��y�c̲Bm(8���=5'<���Ó�ybś�b���I�!-�&AA���yb�ˀ /F��a��+����+	��y"�>7*h�P�U[<|p�E�	�y��	f�D�A�iZ��zyA���yB�[�Z����QK�6^�������y�.] Nc�h"f��~U��ZU��y����!R��{�+�f��d���yB-�/E
U	M%)NْD�)�y�H�p�PcV���`gN>�yB�-rȵ#�ˊ}��(�u�L��y���8�Z�!.|z�r�%��y"&�=M����g�	�lʎ���Jߴ�y�+��+�K�D�:�,,q5@ϡ�y�(�9�Bq���X� �
,��+��y�͐,8���!����PDX��y��Z�\s)�F�̼bgF�4�yc�xA���+BXʨQ����y
� �%���D�pS1K#��@���4"O�� �"�!HӜ9`g�I6G�� �"Oz�%���q�1��D`��+W"O�|��)O	:Y>�)��ۉGIvQ��"O�u�R+�_x~��0�V<EF���"O��ZbF
F�T����S��.H!�"O<�;S�$U���nŝE��h�"O�i@Q�R�W�ⵀ�À�Z���"O�:�n&�*H��B�0�~X"OL� @���m��ڲl����A"O�}�aͳ4e�1����	A��"O�q3�D�fZ�hsf �$d�n���"ObUc�5;��-@��`�L�"�"O���4�FE��[�&�;�"OD)C���T���0�"��.��ų�"O�͈Q�ݏ R�[�X�{P�"O�y����M�c��M�a�j�"O>!�$KV��H��g��_���u"O�����GI���m�"%����"Ob�!�
%4��j^4Z5k�"O�\:���y�(�b�JdB�"O�$���,[g�d�TǊ�pԎ�!�"O�d!��?H���r#��{���1"Od����I�Vn1�u石1��#"O$���=O���P�o7��B�"O ���Z�3���iEU��%"O
��P ɢkq���'��q<:�e"O@z��[�Z:F� ��<�Fu1#"O�R�bۮjL,5��%T��E"O��ZBC �m,�XB^By� !B"O0�����Y���!�3(B\3�"O>p�Sj�e�u��H�)�uR"O$�
fG�'�r0�Ҩ��4�0yX�"O�j�KF]�Q����	0}à"O�̢UI�)L}��'�
�&"��"O��Jq�M6��p��%S�����"O����C��-~� ��˃p�ܵX�"O~�)���ir5G�/P�FR�"O���Iȟ{�`9�%2_{�=��"OF��"K�`Yud�t�,�p"O��)����z>�!� -v|�9p�"O.��t�͒%`
k�Ę4�b���"O=ѥ���(׊DrF�:2� Ԃ�"O ْ���8X��7��m{�-��"O,���7\���ʲ]�1"O E��N�!W�)B#��'"O���5p.�Ȓge �w;T��"OH�6G��MZ�2�Ğ�X�D�CG�x·iO�b?y��>$��|J��nY�yZr�6D����eH�B��۠�D,BBtc6�Ix���81��11Z�)�l�	ﾡ+�#3D�t���Q�]wL k��ۀn�J�:g�+D���V2!�����*Q�NAAt<D��q���'�  �#H�(��L;D��eD�3[��P���mcޭ�tG?D�(���N�S�����'���hUN>D����'3,GmCq�Q��	��<?�
�e���o�7r+�
���=ޠ���@y��C4N}��R:!&j�$ G��y��=��ڵJ�-�bT4@��y2�W�m��s��N�~NM��kR��y2�E�TB��X%�J<�.ؙ���9�yT�S� ���X�~�p������y���/lʼ��kQ ���B�IR��y
� ���`��au����0\Lr"O��AL8��Xv�Q.q#��p"OJҷ�6��E�T%� �"O~ي�#��P�V��c�/["&["O�HR��uڬ;IսY���q"OH ��N�l��xT�>��a"O:��vm�(`�a�dY.G�Dh�B"O�	s3�Ƿ~�F!q�j �("Ov�� ��W˄�{%J�	�T)��ቻSQ��S�D��a��| �GܲG3�X�ȓ4��Y��D��a�x��,:!���n]�T��ꆠ4�D���I&F��8�ȓ�����KՓZ�f��0G�%K�pM�ȓ�Fl:G�,E����!���Iu(����i�	�a�4����N-&�ּ�r�O$HPC�I�]S\ej��͚N�a���3S�L��*^����-�,t�h�Q���& p����L�'���/��9���h&�S�����	�'�����Aی�肄U3|��҃T��26�>E��'Y���0���yx�FJ�@Z~)�'��`�yR���a&���r0@O*'
�pEzR��,�ȟ���1��4�N<�e�"��Sc"O���g�hju���\2s�FmȰ�Ot��>���i��I�@ B8tڰL�@�7&4az���Ñ���Zu'z^�� �P��'
���^�qYY���#��ܹ�̖�n���ȓK��89�$ʛ*HaY�#�-����ȓ)�𤌁3��%�w�7D�hŅ�	v�'��$��P�uA :����f	b!*
�'\!�/�h�pv̟"�(
�'̮ #�P�Zn� :�"�:�'�L嘴��2$��a�����˗��L���<a�홿>�����b_�5���mB��HO�ʓ�y�)��	1�䚧���/���呔�!��
Z�m� �ȫHN��ѣ�c��VV�D��M[��s��9P�!ܚB��d�T��1�lU�"O&��l���r���C�T����IxX�4��n��[��Ĉ�j
/��9��/+D�`�eL#)J(QAe��<UZ���O��=E�$!�=I�.�j&m�y�j�B�L�.NC!��B	:�|s0BM�����+ʥp.!�D�a�$ɳ3��(3d8���(&�Du�d�OR����|�7�
 @Lf#"��'?�@�G؟`����EyC	b? �m V)D�O� ���I!�
=Z�{lt3�f��;a~⁹>�A-	���i�GՖt���B&	F̓��=Is��&13�d"DcْFL�A��F�'s�?��������SSg� �e��d+D��p�$�{q�pEɭ��(��)D��A�bK�N���X�F�-~h��j�2D��#e'ֻ5� �w���g���i3D������^	�]��tAɧ*O�U�D�5Q��`���̑�P�d"�Ş��8#�L�ta
�I��^)N�l��$��)C�DX�K�Q��Oƣ]�$��>��(;<O޽�G�7?\9���#4��&�'ў"}:ش<��Q�v��5e�&�� Ls\dц�[Uj�F�&��,��\�}D��/(�Ex��	&l~a2��C{�<�V��4�����C��Wg�j���F�PP���"�'Qўb?�)p�ɷG��i��n�Ή�D�:�T#���i�s:�	aehF%�~e� 
�!�D� �8�9Rm�']~��w�9�!��9mj�AF�����c0nQF�!�� 6X���(a�2�PA�� Y�x��C"O.鐐*\($?�)���ɕE�yI"O��yE�yɧ!�d�V�@��x��'�����L��:-��q�iJj����?��'�B]�f�N�8�k�I_�=�NU��'B֭��A3��Jǧ.�T�ٌ� ��?�nZ�L=�oO 	lIa��J�_��B��=���k+75 A�a��"?���5ڧ\[v|*���^��q��P%U@����j�j-�V�0�$T�P���`3�Ș�'sў�}Jd"I(W�z@qA E
l�� NJ�<�a�V�U<���$L?5h$Q1$�j�<��y'&k%�S�d6��!|����'R�	!T����5 ��[`�q���h�nC�	�sd*бW*�&q�t�A �%+}~c��̓��'F�'�h��B	�&
I�(��ɞ1Or��Y��HOj�a��޲a�}�EϧS2�,0"O�R��P��ȐE!Y)r!8t[��I^���	 (�<�D߬n����_!��&����כ.:F���L�_�C�ɧ*2���'D�^�Ѓ ΐ-A��C��!6�v���ǧ��т��,?��#=�
Ǔz	��
H�4Yۚ-Y����LчȓPޙ2��1�q �mF�J���o�{(<��枧Fj�,�V��7 ��s���O�<���R� /��#�U+��
��O�<1'&C��*�C�%0�>���Cu�<��A�*!��#ȶb*���h�<��D�a������3.����f�<Q�o�U���0�fe�g��`�<���4�j��� U�$�z���nM���x��e�p�ytQ낰�s��+�p>iH�8␡Z$i_�P��$�0! XK�<��IE���dc�B"9�CW�J�<�gHr���!�G�q��I�2�Jb�<�&��<BG��� ���b�nXy��B�0X���5�+Sm�Y0�*�Ho�B�I*�n���/�.7�fl#����t�B�ɪu��@r#�Tc�x��f�..٤B��9]�
�� ���D�L����B�	�(�ɱ
�H�p�x�L=-�B�ɪZvj�Cޥ�J!#c�7!��B�	3@x6��C
��(]��.M�~28C�	#b���b��=G��� �K-8&C��"M �ĥG�D;��J:G>B䉄T&Hբ�'.4�u�L_�C䉈S��B��g9��x�+�P��C䉲!�h*���0N-�pPu���-��C��)wt�A�o{����a��s�~C�	�;p�@� ���'��x�&C䉝E�0X+v�A�f"v�L�4UC�I����έv�j|{5�[�˨B�xr��pr���2L@�#�;�B䉆z�Z=S7��6A�> zAʋ��RC�	�S��͛�
b���6f��Q�C�ɓU��i΍E�!�wL�"Cr�B��J�͑7@��wK���E��'!
�	�nW�xjp�(g���<���'��t���:���f%¼�r�p�'?t�P��QV)J�(��T�sX���'�za���K�rwPݚ`,�=l�����'�hL���=AZ(8��٭kc���'�(��V�L�]XX���r=X���'�� �@�/C&���A��x[�h���� j0h������LY��ǳ	֬���"O��i�� �n��眒d���˷"O%:��Z�Sh�¶H�� �0v"Oz�"�O�����s��U���*#�'����"�)A�b�i!K�
{��Ư����y����*6��'~)�@�A:�nM�`遾-9���'9���s�	W[�LɆ+^�ar�'�(a���B�}5>ԪӇ�Qg�0��'�`����%]�P�T!R�E2 ��'@BQ�  V�IB�dгL]�3� ���'��ݓt��P
��*�7)U��'�J���\.~0J�
�gۍ�̬�	�']�DE홥�1��E� cN	��'�p�;���#�h�C������'�r�S"�Ez��ՇM�x;��	�'�(ܲ�љ9����cԺz����	�'f�]�;D�]��j�%��Ձ�'ג�ؓ.O�%���*F�23r��'�D��j�-Y�EXcd�t!8�
�'ch03D�^�=d,�Re�زº�	�'�ހ�'F�1 iU	���fl��'vM����:u�|�Q��"�����'��-�@c
�{n����H�r�F4��',�ѐ��*^qd!#�ĆsS����'����C�T&&�Nh2��Ȩ��
�'���k�X�'��;BCZ�[`�(�	�'����f�$e���`�V����:�'��}�%��I�A��0ۆ4��'3��S�iW�m�j	� g�z���'L�h�m^ 4�8;���v�z���'0A�Ыʲ|�Ʃ�ц�'nH����'��\���Ӌn|��{�Xj(��'KP�Cb��M�̩���ل&���R�'9���r�^�o�h;�eÌ+�D��'�0�u ��(�L�կъ
<��'�NH�"J��_2�[�

��'S����d� L��/��w����
�'�ثfɘS�L�A) &j�콡
�'�lH�&nIL��D�3bL�d��`a�'�r<�f矼�����-��u��'{���eQq2�X3�ʂ�i����']����Q�z�����m�L��'��Lh3�\B6�#GaQ>y����'�t C���Nb�;&+,=���'H&̹s�A$˄��#� ��\0�'��'��2,�v0�vXJ�@c�'����1�ޜ4��@&�S�y�	��'U�]�e�Ɍ��X��[�{ߤ��'����ӊT�z�4�Av�_OҘ�;�'��c �*dc��r��L�_�$D�e"O�X�f��C��଒+I(��x�"O0����9��ae$VM� "O �����[�悫r �@r"O戰DC2v�`�Ӱǚ�HN@� "O�,S�(�)P���kH�,2�"O����؟~�\�g��5����"O���n޿w���"��
��X$:d"O$y��/�-O�������Tp��"O $�`b�%j�V=����,{
}B"O��ЈV@����#��]�<x�!"O�И�H�8�
������0!��"O�yaI�1��I�o�l��d�""O�	,���wT1��e�b��1v#!�d\_��0��.�Z��K'kJ!�� 0����,|�P�1���b��8[%P��R�z�a{��Ⱥq��[#� $v:3��p>��$�l*�N���3��*�&ARbg�!fB䉔arp��" �:�V����"�� �+����ŀ,!�}2��z�S�a�`YģQ�[%x�OD@�B䉳�����¸���	7��z��4c!.]O*��a�O�q�t�GL�����ͻW�`�W��QH$��c�5���ȓv�Z��g-Cg�Ԅ�3��04Z�P'j�.�<x@���8� �c˺c��4�����3�L�`7�˘vX8�V� \Oڅ�r��O�uc@bCL�^��'L��T� ���"�K0,��zȀq5�
�0>Y#I�^�8B5�ju�(Hd�@ܓ;\0��C�L�b|��Q+B%�`�3���x= 擦ٚh�R��7�r�#j�
B�I�D�&�`��U�Nq�ԇ�b��}p�H����e��Hw0TP6��G�"b>i0�N|��V!� �Rx�����?_r��u&D�˃��� :LHŐĂ�3;�!I�Y3�t�C�ՍJ& 	��!���1s���?E�P�] 
�=6X��C�@:����I(�����Gm��2�)h��c�}U��Rg�I�$������;$|����-wÒ�i�o;O�僡��Ɓ��
͡]/��x��$�_*��(u�ؽ$xͨ��\�m�� �"]�Vޘ���ѱ�Ԡ�f�3G�x��� �$9�/����	<��\��D���%bW�L8b����aȈ&+@��ꑍ#t�+Ɗ�<��|�r������8`��.كdT�� ��i�����$c�!�$ζJ���ғøl�c�+v��h�4(	+9��mږ�n\P��l�-ig�":,�]��LFEy������%#�b��Q�ԉU��1�0=a�)Q���t�Y�\��ɂt^�А�#hL��5�K(�$@�'*]3�nV�$Y�HE��mℝ��H�vA�X��.�1��'X&�:W"��T@[���:F"��OĆt8��Z�cNNP��a_��}���D�k�D�e���`�MV�N"EcG�W�`�d��(�
P�|m�t �6pf�96N˦
�,�]7[�*ش���]w��êOwÏ2 @bTy��3{�ɘ��QG<�VC�3F�v �Sǆz=$;�c@4A��K�퇓?z��ǳijf$���W����~:8kS�A7��䍸�R�$��^�0�j�b�72�џ|[ŃR�`Dt9�Jɋ~�´+�.�4G�N�p�+	�
����&O�撁#�ITOyB��>�H�[�'8�)G�s��9@��M���.OʥsǤ�3cW8e���j��b�]9w@
�؜��/m��tX��0i*`��&�=XB�	%T��@+'��b��g��!Hz�J�5p'�ə�:|iIq  �i��l�j������~݂��3+�S�f}��I�h����'6,R,�o�&@�IQ$>��8�!B %Ø]��h�M���L�(U���l���vk�+=�>�?�A�
���C�cڮ�����R LH\��d��~IJ@��Ǩ}�8��#$���xb/�6i����A��X���w�<��_bnv�r�_�i�����Z�4	�E &f6�S2/x�x�I�F�u
�GѦ0��B�I�b�rب`�ݜQ�n��C� �J��	���!�+�>K4�X`�-���I6
�	��ђ���7%�"	[TBT�0�`����	��Œ�J��f�!d�O�
&�I�!S�[�����-�G���0�ڕ<0��$Ԝ
��e+V<IÛ4g��x���Q
(Xh�diވ2Eg�#z����,�o[�UXu���<j!�WO�Q��mV(���s�`N(xGE��$^F�t�Y�	��\'��"��������T�}ST9Z��;)i!��;^W8�5	��}E��eZ�hࡳ�RT��ى'�^?Q���O� bP.i��\*	�S
���"O�$��F[�\�����H�DX4�(��'l�튕ϐ�:��D��SNX��pdŕ�#��V`'&���ю=|O$yJ҉������%U�b!R��T�Sq_j5(��T|�9�'�V���/�R�ڥ��/�c�Ht���d��,�v�����j��~B��3;j,�Ǭ��k�L���`�<�%��m�L���K*Osb<�ŏ��a[����
�ʲ��'����O.�Rҡ�i�H9@��`�~@k�"O\ !��f�Q�ء~���E��,�s
0A��-��ɒ>?�az�>Cލ�0H� &�b���I�YI����L�.�6Q��
:U��E�ϗ�y��i�����J��'�Ɂ���y�ɜ~�"��"���UQ<���c�y��~��$�e)
�D����&
?�y�M�*-���A��߼�25��I��y2��(6�d�`Z$�psN�,�y
� �< ���<��JA�/6�ep!"O`k��JЩ���("�q`d"OhDj��Lʪ���3����"Ojm���~�-w���CAfi"O(	��Y���'�ޮm�j�9��DW6W7���(��%�ġ�pH�I���+P�ه��(��1;KђO��CYнpt��?1�%��8����`F_7����v,��L�>tGB#�~b�`�O�q��	nx��#_,]o2<Y�J��?�BB�I�D���S�۪p��jv���r��ʓn��Ac�اS�ӧ(�p�����FD*�� �V�m�8mc�"O�8�ɑ(N�5�W�TC��&O���(; � hu�,����(쨉��ߴ\��\S�#�^n��)������;6*�,)�!�NM9A�Z<´��ɴ5&�� �M�3n��c�`���?��� 5kԐq�/��H >�t@3����R�� �H�g�!�d 6[x�d-ЌO`}*�`�)W��	�B5N�U���{��S�O�J[<ԭ�Q��d���J�''�đ%痞vuA�u$ipl$ Rb.}"�?!���x���{��A3W� EK�J��\�L�3���xA�U��_&u�V����K��ج"c�l��ԛ0K��Hs���Ԑx�����/O Źv�ʀҘ'��@�D��\�Бë�yJ<��
�'�����cǊUAּ�S(7z����'8e�Q��;z�Hu�2��$�|�{�'{��+$H�*1u4��1�R��!=m�Ѐ��'5���l��U��*�/���ă�'4���'�ӻ����*�0Sz<��G*F76����'ɜ}������0�͚+:�(�����+58$�� O��ħ*B<���ѭP��u��'O2{��ȓq��h�g���$В.g���'Bd��3 ʸxF�]�OQ>�h���h$�L�w��i�r�!��+D���%'�(�����fso^�$���I� �ʌH&	�F�3�	�膅�`�0��[׎��X���$A➍ؐ��7���
�)Y0iv���� ��i��F$���U` %7N��C��-@dX�G�j�����Ӯ�F�ӆvS��b�G�6�h�6D��ZD�C�I�T�8+a��K+(u A�Ϣt��Y"��t��=��ӧ(����c��ppzM gӤV>�p"O�ÕN�6�����~@�P�j�p�$��`�(����5����4�j��S��>b�t����*f�!�č�6�����$��> A�1j��\&<e�W	O�-JP��D��%��D��k��l��=2�T�%�x�ׯ ��<ajP�{��X���Ҙu�����_A�<��S B�xpS���]r�Ix�<�%ș�K�0�!"��J�/{�<�D���X2��H�F�vf��KSp�<!2�D��hl �j^5X$d�Ir�<�-.x�DP��O� �,*���i�<�3�^�ufn�����q�l$p'��<���Z�N!�@L]�a�	!�Jx�<�7��H�����\� lRe	�`�<a��V�\5l�K���sH2 ��*^�<�DT�B�-)`C�!4��zw�G�<���l>@%brl|h]b��JB�<	!�-Q��[?�I����t�<�P�حd7(9[�'GkT�Z��J�<)��܋���1��b3����UK�<�EL��
��:gc�=&&�Q�[^�<A�L�?xxIݵu�\��FF�<��f�Awd���KB05�d5�D��B�<��h�)$����T�2���`KE�<����i�< q�����D�}�<1���,B��S��ʍ_��ͪ VU�<� �t�Ԧ-�ܘUlU)k��1�"O�q�C�ˇY܈QEHT�'� tZ"OTЬ�.Kڥҳ)	��Af�CW�<��+R~��Ȑ	�9����4a�o�<Q��ʖ(kx�bg�@W�A@B��d�<Iĩ�:' �� �)>fJ�arF�K�<��N+{ex��g�1�D�[E�NA�<	RGp��b·Df�+�M�C�<�#F�.-I�G�49)�&{�<q����F03uĚ(_j<@Y�L@}�<��Jصq����gS�S�t��6��\�<q���H�MF�#਄�3Gs�<q����L)���r$0�9'k�j�<��k	9Ĝ�R[Ph���b�`�<�b����җ�	䔐#	�^�<aG��,o`�ʳ�S�
���aCS[�<a� U5Js,D�b��@\�0"&�O�<	Q΍;yp9���12P�qV��E�<���@�S�4x�����ig�y��\}�<ys��$t4p0�H��<)��cT�<a� wP{�哫两�7���<�ga�#s��I�dǛ!h -	���x�<aR��1`).��3�@�s2`Yp���2s��A�{U����'�~hҤ�ȓD�t��չJ|,���4>���ȓ6_0E A��p#,�vN��+�ЅȓO��$g_�V� ��P�F�J�a�ȓbތ��a�<c�ʭ@T�J1渆�$Yz谐�۫<
��#�AɊU�H�����$��(�L$8��s�,��Xs<�u�L�?�}�T���N���z%����3^���(Կ
�4��ȓo0u��e13�����#!��ȓ7 �� B���p�A�'�0{V�؅ȓ7�Z�vĜ%:�p�ኆj�~��ȓe 6\�0ˋ �j<�ժ߇<(<�ȓ!����R$�)&C�d0@BY�u#��@�q��ж,;���!�֓1?�8�ȓ|�b��A����R�fݑ/�����)��h��N�FV ���ȓNV�{�'жL`x�&�� #�L(����31�Q��la��<D�LA��_�.lȂ\(y���ٖ�լm����Y�px�AHU!`� ���Z���9�ȓf��@�,	��)��͋{�8t��<,]:� 	44הQ11��m��M�F�8��K��fX!W��^���ȓ5�H����X��cJ3�ȓ^�f�i�Ǣd=�@o���,(�ȓu�~��'�O����HƾmT���La��	EF�<Ms���1�M�5�x �ȓ\"J4*�$�JĢFP�HH1��[Bq;d��x��Zb�ϳ�T�ȓ_؄�u@7sn�<)�M�*oz���I�,�yRA��᠔"!<�Ly��8��9Ѥn��H�An���ȓ,>%���C?U,���"J�f>1�ȓQ˰�B@Ī�*��ŏ�C�a�ȓE�0� w$O�:��iY�%]9�-�ȓG���$	�6-0Ե��iR�] ��ȓn�<nܰp�4���m�a��!�'B��x�� &@��%���5"T�A�'�^e�qǘn�A�N�~��5�	�'3�����8�|�"P�D�zV�<c	��� uZRdNT�P��`͈�����r"O�����#��)BÌ�����&"O�� ��Z� ��a�,��b"O��ȖK��@N�e@�a�B6��"O�K#��j���SE 4lՁ�"O~�R��ޣWw��J1��R���#�"O�����&� Tr,Y;JZ:��'"O��j�b�L�\>N��;#�'R*����t����,���Xa��/%Ƽ�`��J	��C䉗��X��+�6�x�KT%�d;�c��[���f>�i��2"�P�dބH~\q��F,%_�C�I'k8P� ��l�>Iq�N��8�ij�f��p˓)�T���L�$0�OC5{Q�	I>�x�����x���Ps���w�[��<q�O�?���@�^�~�}�p�'�0�;��]�Dfz�HE�X1$��<R
ϓEct�(�EY2"��(B�'�2���h�A���"ό��'%�L��'j\h���b�΄�M>�k�d�ָ����%���}�լr���@� �ĉ�3"O2e"ׄ
Jc(�ZE���:|�u�R%tA�\���TR�!��
^���0z����3�Е��͔)?��Ņ�	9o�H��3�O�l���}�0|*@�"U���q%�'Y�9�'H¥0~(r���1U ���Ш��,2�c�p���!#�7c�O|���d�A�l�I�0c�=jTG�O؄T
F�5��lڱ�^�%�}h蕁q�j	a�N&��?!��Ż�8zW���J"2) %�+AP�� ͣv�A��ӃR.���ź�*�A����4A����HҮ쳖�̵)FH�&��`�<�t��}�t���nK�0��JD�K@��'��	���F�	M�@�T@��y�\�ph��lN�$�,O����D����ȉ"4�3c�'�jex�"���L���d�x#�bF"!� �G.v�0i6 �w}2��U3l�����s�'z(Q��	�77P��GO��%;B�ȉ{f�-|Ԁ3)�H*���H�|�4�GO�p�y�(�B���;�4}��2����I:q�$��J�SƐ[vHO'�l�sgJ���zy��卻f���a�*fݡ��)X�bT9cNY!�����ЃcO�B7���e�2y��zO�أA��/�MBf��A�NH��^�HJl���Q�Ai�	4JՃQP�9�TP�Z3 �!R����_��Q��8m�ܽ�DE8�z�`�"<��JᾝK���WZ���"�sy�p�d�:����gE���Y� �%B|t�`(OF��S���*�
���F��������  �2%��6��uY�(��1z_Ѐ��#� $��0���@�t��C�:�R�ȯI�Z@aeJ^�f[�ij7��o(<�wj��T{0��D�[���!�7g�|�8T{�ӸIH�m��i��|'?]Ҁ�q~�_�n���g^�C�$��ubG��?QF@߆hV�P�O��3D?L<ux&�Ċ!�L�a.ڪ<I�͓a$��0<��� X+��j��Sjh2d��o�'j� �D�di*|�a�Q�y��1P� !�����`*�d�d�,�"hƆ#�!�X���X�E��PJ�Xh1Ɯ@�	?�RY¡v~�1yff�?:�@���R�'���"o�{:��e`��%;(t��K���3 �Q?Z́�^-&[\,�	�>��!��B`��Z�c�S�Ae���'�2��2�� m�����U�&���'�6��R�S\o2	Ӱ��Y�ĨĎ �Y2�uf2��X�e	H�$��I�s���! �<�6�FA�4��dÄ�����K(��/{�r�x���D�b|�a)�vX�AѠ'$�����-Ivl��r��&��,8�.:�ɽ;@����i�0���j*�Ӿ�v�����$�kf��O��C�	%5��ڕ/X.bѠѨE��@JfE�#�[��B��Z��~��s!$���
�`T�QxN8��*#D� �SfR#N&q���,Tj "�O"%�a$��[r�`�!���<��p�z)#nд��3�8|OEñ	>��zA�֫MT�p�%19��k�1?�$�
	�'	r9�'$N)x����Iu�8�Y�����?��2ɞV��1�~��bS%|��a
sO�7�����+�q�<a���1�Ȕ�&��>g��cE2F�8��K��n��c^�"~�I0U��j�F��L�����؛h�B�I*��$��(ߘ,�h����/�1[2�����'��<�B-G	J�F=�b��Y ��kS�v��i�͋�$D�1��]p
H@n��~*��[d"O�eW�L�0Zj8� ��X(J "O� $5�I�t��5�J*�i{g"Ol�k������R,T�|,��#�"O̠ZPF�FN8�a�k
h�a��"O�*�K�*S����t�U"O��/�'d��<�W�P� 
�h"O"���,�.�ޑBN��&t*�"O�l�Pb"n>�$N@^�0�x�"O����N� :z��R�Q�B��"O�HK�͓pE,�1p�I�H�ĈB��Τp`@�ZÓP������F����#A\�
ڱ��R��+V��\�kƅ�;WT����
`��X`�K�*�	�![I�i�7b��B�:PDbf�oR*���H�Ӝr�X��꘎EKz����]B�C�ɀ;� ��W�ut4��l�]L�˓^����J��^~pӧ(�T����])b�a��Ð^�����"O�$�EBE&<�ccS�u �@����B���'{����K'����L
5��c�:LQɓ[�Z��@@Z�h�#Hm��ճ�����@�s�j������<�C�$�/)�`ȺsD�>~>�?���M�:���q�.�IA���p�IY<���c��E�)!���4
���k=�����Y$"z�ɯC�D0Sہd��S�O� Qb%@W1���Z���"7$:�1�'R�I�p�LE+1B��4U��%>}B"�+*n�����{�Hݭ^Na�rlر|^�}2���x��,\�Z�	��q�Xݰ��k�)��Ŝa���i��~�� �d³Ir8� � �p<q B��$c������zL#"b!/'�U9Ջ D�x�v�ʹW<T���W 0��ݩ�C!D��a.�/?�����IG>�9�f?D���'��*Z,��ՋF���%ڃ�9�{��Q��'-��[ �I����D�ͱA*�|@�',��s`f���u{��P�:�6!*e��Wc|)���'}�y���<%���s��\��y�����i���o�8��'}IL!Z�'[�q,�8�C��tkء�ȓ���"��[�A��`c����';��'�n^`�OQ>i{wG��~[Ɣ�4*�w@&���9D�Ui�Qd���CQ�de@4��
���	"|�ް O�U�35U���ڐ%��(ڲ F�	ކ��$�"6�C�<b��! A@�bH@ʱl�=˾�3�����P�K�W� �:��	D�D΃�+�FUS0JHJⓥ �l��" Y��y�t��K�B�n���!�#dV���*�ؼʓ��y�Ҥ��?Dҧ(���9���'P*��Tz{�xP"O�47L��!��}��i� 6Uf��6,	S��S�j�����8���1j����e%� �(��#�ӳ9�!�ğ1h���b�(�2v�r��M)OD��a�,t� ���
���W�ĳ;ψ ��E�}��xR����8�<�'.E�:�b�)#��"i�x�<�����Y���QMn��4d�w�<yR��%w�e�)��y��%�k�p�<I1IY^ax�:�h�9/ּ`b�TW�<�S Ԃ%�ف:.j�Qs�RF�<Q�� �&}�l�RJR�T;>���`�}�<	�N#r�R��%��0S�x�#�y�<!c�V[|�D
w�C&jj�}I�D�y�<��F�x6D�K3eբz09�+�r�< g	����@Q�x �#m�<����+B�ܡ&Ù$ȴ#�g�o�<Q�:���(%�Q�/�f�b��e�<頪ˆ�ѐ޽A�1���Pe�<1Q�A3w�2��R	[2xW8��R��d�<�3.͝�m�uo�/8��}2�%SH�<a�	�"��l���_�Ӥ��s,�@�<�BN��4�>����ٹ,�
��^[�<�  �v�<f@�+DmQ���1 "O�Dف��<�rI�D�T�x��a@U"O�����d��h�����zt`�"O�]2��eJ^�0C��]!,�	�"O��À��G�����+"xtH "O00�ъݨ�~EF�=	4�LS�"O~��DѿЬ9i������"O��+�AS2�����F��'"O����ѤY3(`Yc��3z��Y�`"O�IUG=,4���#&�U�#�"OHX���d@=�$�1�P�W"O�T���Ks��hb� s����'L*����Q�e`5��E�hjp�BAB�RKr��׎��/<��)
�'��I�5�U�'�b������2m���'~:`���~`d1W�A�;�n 3�'О��V�R">��rs��, B���'�>|����){R��Y"JX�f%�' x�a�;/�`���K\�M;q��'�@���7_i��t�شE����'U�-qjr���q���S� ��� ^����CMk�H���nY�9����;��d�^�qÒ���=&�)�T}���/<������$�0 ֤F�x����J�{�B���<E�d�шa���
��_E�0ģ�U�r����O*@��˓T ���	�RR��B��6F~��8�.~Q!r$�>���!&�c>�%?M�%Ø�B���6�K,6>������]3�I6Y\`��1%ިT\a� E7[^�&�[�5'l�Ȱ,@:��@�A߈�1q�e ɧ�O����MI��J� �%@����O�Fꘘ���H��A�[@F�,ȶ�4E��h�=O���7|`��$�8z�Db�J�&�f1�ȓ�T�c�c�!`u�&H���̄�(��6aY:w㙈�.��ȓRd��.jv��2�̀G_���ȓ�<pZ�GJ��C#��4�9��VR����-�B�AV�6<z���6L�="�F�1MK�ـ�'в&P|�ȓR��t�cA�<܀I�0�JM-f��|p$�2W-Q�͡�� QT��ȓ_��Ď� �,1�E	��9�@�ȓuN �UJ��{�rA���Ŀs���ȓ=����VŦ�5�������B���fN�!M"f���I�J�X�ȓ4'����b�0*�;��*a!�ȓ6�JH ��}Vd���&�.P�ҡ��Uվ@2�`��a�XmKF��?9.<��ȓ���R��Ap�͘e I"� ŅȓT�#Wߡ%�`�8u)_�8��ȓp���H-'�b��,�-I���ȓ.@��G���:��SŃxW*��ȓX]k7�9�"��������3��"!�&h���k2n����P��}:hXHF�2ĉ�T6���ȓMT��go�+\lႵ��\��ȓ�	R�@@�\_�I�`�;sAd��ȓ6K�j��B?  ՂT�ݠd,
i�ȓ����ڡl��M[2�Cnb���ȓ+�h	�����3��]���ݴdغ��ȓME`�p���'������>[�	�ȓ"' @��],j���ڂd��A�����I�:�s�gE�*t���B�շ}+����m�\h�@�[Є�jq��U�pŅȓx�H�1IݡIE��3� B�g�"���'�D����B�[v]顦A�<�ЩW�jH �a��@A1F�@z�<A&�R1>x�QeI�*��  �FN�<� �񁖫��e�*C��A)b||P�"ON1 ���T��
���$��"O��"�C�38J� S�+M>L�4��"O��Z�
V�| �M��tD!�"O�8�R��Ty-T�i����"Oٙ2��']~I�K�82@���Q"O|��Bf|��
�(x)���"O��c�L"
�����ȓ*k �
�"OXhX�%��>:��B�E�p$"O|�b�O�bL( �`�=N`�"OB`��Ϗ
$3��ڲ-��k����"OZ4�5�
7��9*gF�:`���"O�Ȁ��E�0�B�#��,x~!b"OX����
H�ns5d_�V�X��"O���QJ�0��q0�@ "O�Ba���R�qcC� Ll�Ay�"O��[��b�D50��� `v (�&"OX�3�@�(�H�S#ܾ���@"O�Y��ܖ���[��ƽ:��� "O|�����L@$��0gj��T"O(�B��u��5FlI��u"O�qQ�䀆t*�H�J�~0\%��"O"li��É21�gݏ1���q"O�)S�&�+OP�e�G�ϛ@���"O`���"C3����2%��2V"O,��`�<o\,qe�<v4Js2"O���fҢJA@�9Ů�4q�d�K�"O�I�efa��Q�~:�iQfeΐd�!��7bu�2g˔a�B��Ę�9�!�d��l�D��� �DP����]!�E��l=��ھ/��AY� 3�!�$-��2Ϗ.�����Q"0�!�$I�(~(ת�602�"���>X�!�DQ69�j%�B�M*�fa���j!��,qL~�i�k�m�L kA�0f,!�G�S+�5���V0٬L!"ꂭW�!򤛩,M�=�f
�t�p]���!�
B��IX�˄�T�-����!�D�e<�a��� �P��߼1�!����(K�CAX蔩2�F��=�!���,��]D�d蒷�_�}�!�ď!c���D!��V�9#�v!�Ы|��y�b�3l��8�d���Cp!��	�Uir���nG�s��qzw+$QW!�Q���:t�O�w�XPq$ҁ!�!�dJ D��Y�����@#]�!�DUt TX��kZ3#2��!R
X9�!�ſ}آ�bd�ϰ@��}��ɡ)^!�$�%)s� {Ä��{{2*�h�6S!��Ԋ��` ��ޯjr���  Q!��L)
1�A=k楫��!A!�_>8Z|�	�!QH�I���a`!�K�./��� A�&�V��/�!�Ջ��Q�R�t���0b[�&u!�έn�8X�P/�4�(�H� �Pk!�$ۖJx�+.�d<����N!��b���3�x41����Sb!�d�G/�U(�lY;t&��#�O+cL!򄅕�İ�b�����_:>!�dT<u�mx�I�;:xTj�.2!�d
5d��+p�\~��X")�)�!��6k��`��fS<�uː�[�v~!�d��d�I���|(�AHH!���L�6���_��qt��<!�� �|��Z4V�� ��5b;l�Xc"O��p�#nBx�6�3k	��b�"Ov�[d��'������S�@	���c"O"��#,Z3+��CM���u �"O�u�Q�U55Ɖ�R���_���r�"O� £cU�(\!�c�	�9$l��"OM�ۆ'�@��`G�J�b���"O��������~�D`T"O
$���Z07�~܃��K�a}*��"O~�I$Ś7�p ��d=�p��"O�0�.�� �����W|x�6"O��ؠo�:��؈���^Q�]�"O@Y�'�y�v�ɐ$� R(��"O� * E��B#P2��ϛ"����t"O����'P� 4�gl�0�����"Ox�C@̈́,tu�q������ "O����-�)}����d�0r��	s"O����� [E��%O:wm���1"O�P�2A�I¨Di��ԋc\�:�"O�X��(<�\XrG��$Aʔ:"O��8�b����AD� '���"O�H�.(kjd�{���n�y+�"ObCNB�P��!�`҄�v"O4-2��(��4IY��J�"O�%���4���@OO�K�^��s"O���3�A�y�L��o��՘�"O
��'�p����_�w��!�"O}���:"���	�Q[r�Y�"O��ʚ3{�1�����B%	 "Or��U-�� �x*voZ�%�J�W"O���i�"�T��K).�|�v"O�$�îZ�����"a�IЌ���"O�E���)=�����Pђ�16"O�Q+@p�� �c�ˬ=о��"O��Sa��)Ϣ�e���=�ȵ�"Oz���I�EƲ����NE4� �"O������>@p^�����0A`%{s"OTY����i&
ݡu�)
)p�(�"O�h�`F^)��a	�^�l�""O��q&l�5K�X�8HB�I���Q6"O��R�^�4"�A�t���"OD�5̕�X�(�*��R1=p
i@�"O���o�7_��1��嚺PuAV"O<��q�Ga�}���Vr���"O��#Ӯ������L�9�)�t"O�ȳ%)�7+��1�fI�:���"O�`u��5L<0ѡ�
.���`�"O *��K" X�A��%"�,+$"OJ����#�h����2/P�(Z0"O���WA�
6�l#FHϸ1�ɗ"O��/K�#�h�1@���5SR"O�S�G�v���13�[83
  ��"O�2Q�U<+�a�8	��j�"O�eۂ[��F���N��9����"O�z-^�h���F�E�`��r"O����IuKx���G��-��;E"OV�gڷ^�zQSW��G����"O<���-�,-8q"E�Ȉx>i�2"O�q�C-�8=��m
�gJ�e����"OZ���$N�ll���'��1�*OȹbP�� DV<��B�3���9�'�����ҪMB�3"�&H xIB
�',�	D��*
?Q��C
�'Q�GO'�4`$,G8oY���� ���Ѡ~#z�q�����yxB"O����.x�9SӉƨ�RdzF"O�q�5n�<��É�%^}�$i�"O���]+?<�eF���G"O`P���KǄ���k��d��"OP�0��\J=�3吜nnY��"Oi�F�1u�r���c�&e��P�"OnͲ� �g�� y͔,H��a�"O줉r�N�X��f)��j��xK3"O�xP"�&}%�!�"�3���b"O�!���ߞLO|X�/��s�FU�S"O�-��A�
x5��O�}<d���"O�T�'+g%����*xڌ4nt�<��K�A��Sf�.�B�)�j�V�<�F�8�D��1aO �ڣK�T�<��d��ݓk*�hks$IM�<���q���]�2�P�b"��}�<9aJ)U�(s�W�0�:k��p�<���N�Dy`pi
PCH�Z0�Q�<�.[?2���Y���=�F����N�<Ic
A�S��`Q�ȯ0�xt��J�<����8H{J���³w����o�<rۧV��*2��D�2%C��Fn�<a6	��a�%+g�F��g�h�<Q�
��Kڬ��7�0_� �}�<I7 �SV�l���
�,\�m�s�|�<��J�`CbYhE��� ��;p)�{�<��	r��-�����u(��:3bc�<ѵ��|�t��V�Xm" �	c�<�6�G�FF�9��/a��(����H�<�'R�橘�@[�{��ic�{�<YSJ˔D}0�����7?PX!'�s�<	��"?����V&A3�g NI�<`AY9E_�	��Nşt�hH9F�<�ׅW�~��̳6�Փ|1�)�KAB�<I���&6�4i�F!E�e�j�z�<!3H�	! �`�fR�I��q�-L�<��$���(����j�0��w)NA�<ɱ�W���(9�.�m:z��ʆt�<A@��)���6lT:���0 l�o�<�`��:g�D�\�RYbу�(�d�<	U/�4 0  �P   G	  !  �  5  �&  [/  �5  �;  ;B  ~H  �N  U  ][  �a  �g  )n  lt  �z  h�   `� u�	����Zv)C�'ll\�0�Ez+⟈m��>���ɪ�l�D��'O�����o] �P4�ѠO����N��H'�tP�l��BY4��D��<L�;`f�K�'G�d��'TD
��a}��`��U�	Re��/LZ�ҷ��*=�p�!j%e��KǷ��a�"��Z��D�E�F"0� �ՑrǦl*��)U���,j��ɣV�:�3Q��#-z����4m���1��?���?��a� h�a��73��Y���4"�&���?i!�i��P���I3`�P�	ß��ɟVznX��ܔ +�)
7�Z��4�����OR���B�����/j3���?���=��a�5������T�!��ʲ��#�jO�+x�4��,���	s�'���Õ�Y�͟ ��k\:3b��`�j"��:T�'���'2�'��Y�d$?�j��k�d s�	��yz@yÁ�Rןh��4Td��%�|��'��7��Ѧ���4j���'�f0\M� ��B �#;.�B�'�f9"jU
�yY�a�`�J=Z}��h�	J���Q�����rT�˘�Mt�iȐ7�����-#N0�PZ(VU�"n�-d,e`'�32O��$^�и��A�a��$[-,T���5n�(,l��M��iE�\*�D�&� �pe��I��Y�W��!|��`2�͍W�6������4R�b0ْC�+R�M�j��:�� �ܷ$�>�	&��U\�0 �i�� �}K��B�@� �еi847-æɠ Oe�FÃ�������[2��*g�҉0-f�%�Kɒ��ٴr�Q:eO��S:�����2w��Y�����',��zP�%>*��iri]�W
0�9G�'��O���>���N���>m@#®��!�0G�L�+�!���]�XL�TmЦx��zW�ǂ"O��g�
-���ЀJ�K��Y�"O<-�AH�E����Pg��2p2�"O2(+'R~t(��Œ�!�Pl�"O8���C[y(����k�8!br�	�qW��~���
�,�F��GH�-p�I��
e�<q�K�&3���cE�>4�T�(_a�<���E`h���E��(�Hr�<A�G1v�V��B�b��HSl�<aug?bf���ȏ@P"���Vk�<y�*��olZ�9'ṇ�N�� a��$1I*�S�Ov�T{%o�Q&���/q��=#�"O���p��1)\M���:M��q�$"O�����0�J��D���q�F"O<Hc��H�0���P�R�t;�"O���g*H�VDÕi�f���!"O��ƬWt���g[i���Z��*��(�O|��o��.���aDۦ[�z���"O��&� �l��A��&�Ԃg"O�TY��K3spЄ��Ϊ��|�T"O�I��]v�X�ϐ)w����"O�9��j��o�8��V
�p� �'b���Mvӈ�d��YI�#B
$�2UÒ/Z� ���Qy��'���'WB<� ��/��ɇ��! �\���3����'  =�K�Ɋ6Qxax"%;}ԜpB��1tVv�� �'�����@�O�"��DKY�u�*�	Ó���ɱ�M�]����4x�3A�$@e(�QiOےE�/OJ�!�)�'��P���!3(5�-?;e�������?!VVT7�8�iC$%�D@:@����&�:4BO�:�b>����$j� ]����Ļ+��"��IJ�<��k��c� 3Bв&�l0�F_�<	'jE�|���!�/&! ����\�<� X9Q�r��k��F�N����@_�<qү̎Qt�Ub��4p��t��]�<Yg���1�c�`R7*��-��!F៴㔎/�S�O�]
`OcR��, �*&��S"O,tQ�Y���w�L�a��)"O����ɚ�C��YV��;.��!"O��p�-D� H���ǂ��.�Y�"O�h�G��c�6yF��<+����&O%�_�m�E�_ ��l�S%��\��>O�����As���^�_�.y�D<s��1�tOr<�GB_;1k�EІ�+�%�<A!�_:1m�AP���-���cAb	�5�0Չ!�'x����}�䍱T)�!oָ5Ό�y~!�$H�j�N���C���}�`!#f�X�ɰ�MKN>y��ەb��ӟpC��G% ༕k�Ă�0��ݸATҟ�I[�,���ɟ��'(�T���F��d	�� ّG���� D��PC�H(X�#���N9p%@�)���lH�q�V&̻/�P�Ո]4j�Q��g˿H	)C� �M��+0ғ_����I���'�|��H�^�Y������K>����QA�� ���N�4!��ɍ�?1B�T��yY�h�/",N�	��Y����'�Е)��'�"�'��7�!�I�0�"��)ɲ41�U�g5�T�I�@X_$҈Ct/U� ����"&1~�'��	��1.*m��9B�BP/�p��I�ETV�X�B�z�Z�Х ��-��Ŭ�:�� (A�N�KȜ���&FƬ��d���!a��O���>ڧ�y�-&��ѡ"�?�vH�g4�y��{^m���5��-���Q���O�F���V6vs�k7D�_�d�A�5�?i��?i����X�	H��?)���?	��yw�ɆyV�j�Q;T9]��"C� ��L����a*eJV �8
@�4r����|���J32�C2�ۋ*�M`S�2 �l�'�"d�m�b��0�:�{����i���'xȥFP8	�d�S���u�`������G��b�'�ў��
ۋHr�)�I����L�h�V�<��?���Їi�v(<mR_Vy¬ ��|R����ę�6s�$���ֲB����	�"*��#��P(J���O��d�O����O���c>�ZR$�� ����N31�j� a��;�Jdy�l�5$�rpmR* E�  /-��Aԋ�2]�FH���K�>�!׬O�s�X���Y�3^����i�BeDzbJC�c�T,hUCˬb4S�ME>?�E����?����>�~�d�₪)�d��C��u.��ȓ8��\[G�7�PY�����%���ڴ�?�2�ݓ���Y�W���7�
K�x� ���y�HP:|4�d!��B.e�g)�%�ybA�������ˤ4P��7��*�y��) �����19�k�"�-�ybb�v���[�1�v8iFޝ�y�B,��!��. ɡu"�!�hO�xR��S� ��$���'.�L�[�� 0C��0(��d�V�Ҩf�����B�I�+WlΧX+%��CX
�JT�V�<��bT�u@E��W�W��b��[U�<�#�P/s0LJ�� ��bG�
v�<9��(Y*Px&D�(i'�i��L���peJ=�S�OثD�M��a�Yj)<��Ŧ�v�<��펎;��+�W�7H8���g�<Q�(�%@�) K�!9:��ӰFn�<Qtkޙ��)�l��\��r�mj�<�Tg��J���.?�&t
#E�c�<�ꊥD�8 *ƥ�k� ���+�`y�G�(�p>���ΦSd���#�3GM��Kf�<�@C3A�h  -L�&���V�<�'ギQ2�=;���%���I�I�<���%^��t�d��K��IuB�A�<���؜g��)����*e��+F|x��bĹ�0T�Z�4h�Ałf�@R6�=D����?*7�eZ��AoM�d#Ŏ?D���ぎ7�� s��@��`�Pm>D�x��S�>�d��eޒ?Mn�H7D��#�셢Xp���T��˖�x#k6D�\�ʞ�;jV*ԊM$t������6�$��|E�o
	M��<P�@�-X��H�$A��y�A�/N��T�s��0[�ҕ)ٸ�y�@����L�P�A�@6P�*Ea�y�]cH�{Ĥ1H_|���[��y�6��D�ç��B�f�:�,W��y�_�E�@)��!˪'����B ���?���Km�����p��	7h�@�kM�IL�ȹ�?D�d�.��p!���>Ԏ�!��?D�T��EUP�P�V8n�8�i=D�����9�=!f��CPP���;D�ܫ2"�GNnE�e$�+V�z���<D���`R�W�v���J7\:T�j'�<!"�Ud8���A��V_H�R¬�6}�>�RB8D�� 1�G&I��(5
\-����"O�H������D0��N;~��u8"O�]0i !ܺ\A�K41p �#�"O8QK,s��q�@ ]Rpѷ�'���*�'�4���ʜP�J����F��!��'����A�'��p��-@��,�'L�a[W�ɰv��-��L�(,�
�'p�����RG�%(wh��L��ĸ	�'�D��Nd�p�RG(��x���'�R�@$�U(��5 ���h��D9{FQ?�� �>� ����m�84��F3T�LٲAZT��rV�e*�]3"O�3 ��%5�&���Ɲ
��|K1"O.�r�&<\�`���/��a�ʀK�"O��ⴊ��PY夊�6��91"O�m�gaѕ8�}Y��_�M�>�Yv�'��ҏ��;���S���VuT����#cȅ�'Rӥ�S�9�<̙�:)Z@��F�
-1�b�Y���@K>.�$��F�����e�qy8�0P��#|�����y��ԋ�L�PC�	�J ��ȓk�x1�B_� ����%n� �=�'��m��2y¦劗�~�Xs��L|�ȓk�F8�!ډ��p�W6COX��"�^A�Fܮ3���w��3D�̄ȓ
l¥�E
����e�"��K�vh��m���E� S�@�U�1��1��ɬNx8�G:P� �ʇ3f��0��%0L��B�	��x��P����*��G7HC䉇J����5�8v:e�4��8] $C�I��PֆH�&rތ	g��n�C�I�C=L�dcX�\�l
�.B�ɹ9Jtx0���]Q<�C��{;��=��Qm�O��ۖM��2O��� T'%@�+���� TJ'�єh00�ɒ׼y�!�$\�.�*������Y1��W�w�!��YHPH�OB�"���[7���!�Y;K�P԰��_�I+��$fR�zs!�dW�Q��x9`i��*u �%��7\r�U(�O?�*gmM�E� ��B�(5�����x�<a�(��;���ϟ$�4Ad�CK�<�c/�"�ɧH�+Qօ(��X{�<I��ыV�z�ys� f�>���u�<I�@�	�k�S>��ѐ�RG�<A�i���)�J�6@�҅Xg�Dy"H��p>a��@�@|�����Ը`j�����B�<�� &x�V��R���f�ja3�UB�<!�e�1	G�թ@�/PKB� ��A�<y��Iv�x%`ȧJ��p��t�<��JZ�m��,���Ԣ9r1*ƏZwx���1`����'�	s �Iӊ|��)sR�?D���	�c�F�P��˾RĞ��� D�l��D)v�hX�I�$������>D�d1£Ãv�n�����S ~�D>D��a�	����Z��� z��v�:D�4�"a�7w��u���-^��� �7ړ!2P�G�4��=���x�E��JfV�Cw��;�y"���G��X�W���ID%�f�R��y�F��z�ա�dE�4�Ձ���yB��
%�Hb�/�X��`���y�]�'^�52��PX̤qw� �y�!�#�������0V╺6�2�?�u��C�����hծI�,��h�H0lp[2�0D�lC�K�r�4���I�e�y���0D�� �<��IR
}r�@増�z�~	w"O๢��+�t��vK�9��i�"O�y��#�Mh<Lq�ʉ�m�` �0"O�����# �i��wph r\�p{W !�O8��An	N.
-��(�W]�8��"O�T���u�`���W��\�D"O��� 'D�aj9��m
7"O^��ra����eh�Y��d{$"O�v�/�����ą���˥�'Eld0�'�H�S�N�*��e���V���x�'��`���L,nd�1�f����k�'�� FE��T��2�.��yrF))������G�Q����DҬ�y�� v����GH�CJܼ�S��y (dTD]��f[�f� �22�P3�hO*�s��S#l��򡚍��Ѐ�^��C��.	1�(1C-٧\R��2)��O��C�I��C�\6���q��7i C䉾w�p��Ǘ���`��}lBB�:/6ѻn�	�~|8��=W�&B�I	�����H֓[ގ��@X�Hz��D�Cp�"~*�E��e`CE `^�l�M��yBB�b��a�0΀�Z3��34�_��y�+�l�pu��#�L$"�1#َ�yB��;@��Z.�>���8bݦ�Py��6~m0�I�`�#A�X�:��N�<���\��0�J�ƨ��Yr��HTy��֨�p>��E�pX��Ũy�4�
ǯ�R�<1"'��hR����J�!=��B���Q�<	��Yw�"�Sb��4��a�kQN�<A�ʚ�)|�=��L��hPP��~�<��k�1~�U�2��;|Ϫ%�B,Fux��"�ù���D��+����eÛ�f�4`��6D�� �W�2���Ӄ0ZDx�1D������^�",��lI6s�慺tE/D����-׌Ed��R�e�v��!"D�	�U�	��d���?+,Dr�5D�L���̍va���iøE`�P[�K1ړ:��E�t��:u��e��E�%�v�Xe�
�y2��,=�f`�3��k�|��bF�"�y"��bQ�젱�L�f�*4Q��R�yRKmɖY��<bg܅f��y�'^�N05�$/��)fɋ��yB,@0r��ҷ6V�@�H��?�� �T������q! v����0��=�m�,)D��c��~�8�@�&Q�#j�1�'�(D�d#񢄭vp1 ���"E�P��%�'D��B�o�I}x5�d�@8�1���'D�,�ť	Ԧ��Pe�#la�%CTD%D�\84�����D�]5�T����<�@��~8�x�s�՞"<eQsF�b��\Ӵ�!D�|�#��.3ژ�"
E/���W�5D�D@QOxe��1�%  �E�7�y⣂�;".���N�4��8�$��yr�^�xi,4*p�\�C�&4GS���>�è�Q?��D-�>i�F��X�N|�6k�a�<)��I�fq�͐~��騅�NV�<��#�/K�Z��v`�������X�<�5n�c��� ��w���a�JR�<���t�!bI^
����t�@M�<A��*L����Aۚi�	P�,ZB�'�.�����)<:��A�_*d��
�@իX�!��@+L��a?.���@��J)�Xɂ"Of@Qo4NH1��Z'ttq�1"O� �Ŋ�cMr���n�o�4���"O}ц�ޜm�� ���TM��"O��)�n+<�|�(�n�=5��Yh��'(L9���::W&������8J�H��Ċ]��ȓ�H	#"#�%OL�\����QE��ȓ�8���B��)5�Ms���<x� ��h
�h�� �Z�d�0���>v"�ȓ<ƹ��I:;��Ie���/��8��͆� �ٕin�aBԍ�1|�|�'�XD�J�~�JWG'p ��B�9o�dA�ȓ!N�8��Qe�� 8ӣL�92��bqx�z�.�;�\m9% ̔�v�ȓ<�f$� !�W 	���3����9D\�B�݁g;Hi�����Q��I�mLN�	*����"�:� �r����s�C�I�lX �N��P�2az��<7<C�I�~�e�0ꊝp�0��5Z:(C䉍;��`����F1�q��9��B�	!юm�QK�%��r��K�
C�=E\*�{�[x�u1i^�+�B�=��h�O؆-Y�,���ױ~�"�(	�'>����m^9J�TY� �&t�&�i�'��!Ȋ�;�r�x�"D?>:
� �'�h|��B�a
���μj�D���'E�l���Դ��3��-2^=�'�݂Wă|8ڝ)���4"���8�Gx��	޹(��۱8�ā�ႃ<��C��p��+J'J����.«I�~C�	�F��{�eIk�<���jA�t�.B䉣c]<�ȣ 
ua���A/o[B�	�1H�:#�C�LVƠ	򯄩T?�C�	�`֔)�oC��LA�_��ZP�=�O�<�bA�����O瓅vg�`�1��B@�0F�ȭ`����e"��ON�d�A^1 5��RG�Q� 	�`o���r�ƀsD�с.��%Zu�D+j�#>��ȗ�G�ȅ��+tǼ!QF��-�ug`�Nh!Ap��/��EGD�O��Ez�'�?)�ΘOϦ`UZ�N�4��'�1p�0�)Od���-� �j݃�֩:MѦ?,�}⢮<�㑕=�jjg@\#Wrt���fCByA�.`�R�'\P>��@HW͟��	�de�d�Ў��ufهȖ��I�dy�IQ��cG�1CJԥ:�����ן�b>�!�'�9�(��� C�Q0�"@z�����_�v�ɑ��kx �����؊�$�ϝb�!��텚2��a�W%E+�y�."�?�������$��p��f�
8d�)��5;��P�4D����@�U�)���95.ړG��?@�"Y�a�~�����*�N��G֟(�Iߟ�a3�P�t�!�I͟<�	ݟ�S֟��Be�s�N4A��!m�ƍ�Ч_�8�u	l
z�����n�=]j!�O��O.���Z׎�ؗK�X}v�����t��!fkߗGն܋$��".������1�x®S	��Ţ�'˪S���A��3��d��U���'�ў(ϓmҖp8f'�z����R�'9�8�ȓR#&�`C�h$�m��J�%��Sןh��4� �d�<�E��}*r�4$�!Y��P��KˈR <Y
��i�2�'0B[�b>��O"W2���تo���sU�p�hC�,	)������<�CC�gT���B��xQ���>b�ؚ��ؕ2;�%P'O���<���ܟ�Hӆ��V�P��˜3C�u�F���D{B�	'VZ\���P��ĺ1�R�y?�C��A�yynQ(yz�����.OA��:^�V�'��ɢ^�������C���y�+ʡRę�VQ'|1���L�Iោ@"+M/6 �qJ�FG��{��|J�DH�q Ԑ
��>�����F�'9Nؠ�ȉ�e���"5��S3*R��@���ױz�#>-lT8�	Ɵ��|���!0H�f!�2 ��q�q��xy�'�B��G�<BX�"�V�����)e��DpLd�t'��m�����J1ê<����?i�����|���?1"D�"% *MB5�Ʌ�tB#/ӡ�?�E߹`�B�0�M����T򧈟�����16��Cp�>.���(�=O>����'X`�p��"�|�z7؁2Ͳ0:䝊`� �^���gYV��O��S�q~
� 
Ii'��vt�&��!k�x��"O p��'/c"\�w-���퉏�ȟ��ᤫ�({�
����MS��?Y���?�o��j�D���?)��?��'�?!���v'D-�%N٩u���P�Rb���Dԏj�JM��C�"�j͟d�8�,��[  QIf�0Z֮ 2JޫW��e�E%c��e�0�.�'�M�J;�D",y  �sQ�@��c�J�	�8�����O��=��'k�}B`@�#���
��ԑs����'����RX���KT�}�$���F���S�4�'Il���#T�b��A�Q �ȶ��@LB�'K�'J�)������"D�=�â\�ᱬA�leJ}A��;I:��ϓD
��j��P�E�@-��o� �̤0��M�E��\k7������8�F����	�I0����E�rZ�z�nK���Ie�'���p�H�>��]����IpT ��:D��+���:N���ȲiN�vMX@8pi�<E�irRS�,��g����i�O8� 8qD�ق:�:a���"<Y��D�3(���OJ���� B����(G�*���<+����ǀ�>@�S�*����">���YS~>���!O�J#����F�?�R)Ɯz͐� �჎G�s�d(�P) ��I�Ms���$H��f���J*�6h��@0���O���� f���"P	���j�MF,)0�}R��<Yv�S�4`}+����+���&�Wy��'��ꓘ�Ϙ'�N���':� !�cE�UB �Ó�hO����3r*�U±,_�m���r�DB���'江n��'��%-���׊�:�D(����!�'�@�L���<aV�]9r�q��ʑv�le�%�ݫ� ��O|��O:Ł6�>�����S.�j��$P�T1V���D��F%:�Oj����h��䀁]�N<y�%� o,Hg���y���u�> �>)��]i�s���ȬZq�� 8F���&��%�?�eg�N���K��?�2Ĉ�9Xc�����ʝ]�T��_���	8\b �'��'�.1@M�<۴e\|��,�BE[Ĩ�F��vy�����ɋ�ȟ�t���ʘF�p�;QK�:��H��l?a6v�T>�-W��?݄����A >�x\�A�_�za��Km�����G�~x�$�O��C0Oxb>����Ob��(`��EE��0Z�D�O��x�'+�,��O�s��"���B�KղL�u�ed�.s\����O^s������G/�`@�i>C�r��ozRI�-��Q��!��!��R��l�'��	F�)Γ�?QuĒ�=d<�:s�(�����(�;|��I۟��'�ў�	:�S�/^�L�p��(���dy��'��0�C4o��[���?[�=�ȓh�0��c|V|<�C�v*��<N��c�C6c6X�FO�Q'~4��R7|1�t�8e�$�9�������ȓa:�,��'�D��k^�S6*	�ȓ	8��`$bӀ}�<aw�}�pC�	-zx ���Z�E7� ���X�O1�C�I>B��A�@b�h}B(yShj�RC�Y'�@�JCVy ��`UU�C�	�3,Z!��&ڬsE*|`p��'dlbC��7p��a�G�ۀ�]/66C䉽2�PuKa� >�!�ӯ^cW��ЛQl�<xbڅ�&B�*s��&�ў�c�'_-G��4P���G�4�� L�@թJ�$L�����CG�=a�)k�R�Q��̩so�	Z���<4�RV�G�4�%9�ߣ,��a�`ꄧt��*c[���M*���͖����B^�(Ҋ���DŉK>�w9Yu`�eM�{����E��v�<�&�M*w�"T��#k���$^�C�I�x<��C�K� Y�#+ʎ=ҘC�I�kd ��c��`�����oI�3�~C䉚B2���YcF\�xc�pQC�	�oװ�8Cl�1v@-�%h�Q��C�I�<�Hi�IǗq�h�P�"��I�C�ِL����$�:)�a� X|.B�I �d��ۿL�@�X��*�B�%J�&�Cu��f ���L۲e, B�	"97�s�]N� 0r���C�	�&�Ρ��k#Z3���r�ۊ'�zC������s=@$Z �)3`�C�)� �X�a/��@L��J[r��y�"O���2�R�(��������Ez,�r"OH)*q%4HX��V cb]��"OlŲ�)�8��@B��;ybz �f"OD�H4,R�H��+! ŗ%��m20"O���!�	?/�Ȱ��:
�F�T"O��k���d����g��A"O.�J#̔'�pP�ǥ/��r"OF��s,��;}nP1�&C�2���@�"O"�@`�D��[2f9�� �"Of�`��Çk�"��֨)�R��"O��T�K+!� ���<0��H+5"O�Ay���s�xY��@�e�
��@"O<C��S�o~:L��M�!��m��"O��j�Ə;~��(�aO�0H��1�"O�����Il��R�nȃp��0��"O��H���5�4Ⱥ��8?�+	Gi�<��ҏ4]P\[q�½�FB؇�!�$
�cx\C�	{�k�~s ���"On��O\q��`Q:����
�'� �2��3-���j�1B���'vŹpƐc���w�C70`�"
�'@
�����J�~�b�	 -):�E��'%&| �aI?vF�	R�HD�	X�
�'�Ȍ�G`��^�����Ĉ8n�4���'PXᐉ�-���� 'id�:�'zF�����#It��@�ޜZJ�]��'3\�ݤY)�E��&ܵK���'D Y�$�2ZH��! �$<�@5*�'r�	����,E��4�� 76��x�'��d�֫8p�֨��� +0��i�	�'(V��@�""���f�"�.!��'f}���	T�(��n݃�^X�	�'�x18���G�jE������p��'G�c&��p�:�Pi��"�%k�'�fd�`��Da�öE��	x�'J�\ �k������A\7n���[
�'J0Y��*&�<R�슫Z��	�	�'��%Q�n�)��${�n��Mx8�*	�'�f���
M�8,��I(L�
�'"f|��N�]՞l �k�o��lc
�'1��"��9G�����d��a�\��'�����P�|x��P�� W	�[�'�Ԛ�� }��=J K�� ���'ʎ�2ǭ�=������,<p�)�'$�X)Q��6��8;��V�X���'�Uj�&�[�(��c!79���

�'YL��$�>Jx|!#��*�5�	�'R��[D��C��<#�cN�$D���
�'�a��ٳ7Gv*��G"w�Z�'�)��';P��3������	�	�'ٮ����=�Z!b���
5���
�'�(UN�n�^H���>X
�Z�'ed��$A�$�&��2�ѶI�!i�'_�Q۵fǗH�*a�R��	Q��@�';��)�@θA�``��$>D@`��'�N��q�F�n�z-s��:c�h{�'I(�Z5���Id.�+�O�6h)�z�'�:{�lg^�2P�a3r��'l��s�ؚ7T��B@
Ͼ*��l�	�'=�}�A��p���喉��:�'��zv��V	J`�ƌĀ\��'q�5Q�l��Z�@&��Wh��';da0��8�T����T������ �26���fș�䓀I0�Q�u"O
���=:��p`Մ6,Z1YV"O~$+�B;.:55��&��z�"O��� �	�����U%I�M�%"O� �
�5��t׭�K|���"OE���
 �srN-�
ȹ�"O&�����m�j��@N��v��4�1"O��j԰�@%:ס/�"E�1�I�<)�A#6\�5A�ҶO���yU*}�<a)�08渀�K��P2*�aq�`�<!��@3&��A���P���3�^�<�Pn�t����3� 8�q�\�<��8�Q�n�I��x�%!T��Bc@ҟ��DI��
$,� 03J8D�Q�j��7f��a�ۇO�\�)Pk*D���mF��f+�/o�XԻ@&,D�����M	T�Z�O|dQCE.D�08E�����T��2xLF�L*D��Sw�GG�@A@��6T�ԯ<D���@�]-\�!G�X�+s��9�%9D� iQ&�a	�gV�%���S�f+D�`2�N�	NiF�T(�扸��&D�Dj�%�#\]�{��P&0���B��$D��Cq�8W��ӵ	ЕOi�lSF� D��a��*j��V-�`ec)D�������1�~��fM�R���4�,D�,�6�*-1�X1LM�__z�S�%D�<�׮R�&� ̓l[� :G�(D���D��E�X�{fl
';~6Ȉ�3D�� ���#�;&�j@r��4D���E�_��;��8,8,�ZQ	 D�����6a$��aW�A2���b�D?D�ZѠX�'p�qjR� =L�IpQ�<D���A-�:�Y�0�+|@��!ac9D��nN�A7���U%ُ�f�Ӊ)D�x
�͎�!3��3�Nn�!�w%D�4�ӊ
`P�|Y�j5D���3�r�k7̓�M4h��C�.D�zA�Q':�d5��fR�
B!q +.D��ZC��1a��D�#T]23"D���,ޣ
��R䊀mA���w�%D�8����X����w&Ho��$��l%D��� ���+3&C��t�1D��4�D^�4]s�AݱT�f�`�",D��j��3[�����""S�-@U�*D��`�m�&����O2`I�]"e�4D�(a�
��5�1*�/@�f����D�$D��(�"��(��B#j4~��W�!D�4�$�Ɇ=������(R�@rwM*D��QQ�@?��1uG�!�%Ӆo-D���`�\�'��-���K�L���d�)D��C7h��&-f������t�A��(D�\�U���S���	��C7Dn)�'D��:�C͘~(n�ڡ�L�68����(D��Bd��>�9Q��H�>>œ�+D�8���H>G��[����8њ�)D���f�܎IT�1�
R�H'D�ؘg�GF0�S2�
41����&D���D�y�jP�U�p�扉��0D���Hu��[eL��S���S2D���׆��-TS��0;^��J�+1D��yL�P��%+$D݀��u3��1D��r NAI�fx��.�whxIb �;D�X bb�!
����Q��W�2Cu@:D�� ���Ե�d��9t2��t"O 9���'J����O�BQX��"O�:�Ƅ�1�Z��Ɂ�zH~hR�"Oވ��ԅQ�����";B�r�"O�����\��U(�F�-)�ᨠ"O���b��n��s������д"OL�bmC*y��܃$X��v8�e"Ovi돎"�yҴ�4R��Ljv"OX���ݸT�|) ���,y8@a�"O�P���&9�t		0�_"1���"O�k��eo���⏌�5|�,��"O�x�NȔ[y��� �eh|%�Q"O�t#NA=%���G�~�^�q�"O�$������(�m�%����D"Ob�[��s���
2�d �C"O,�6*�3-�i�v�'m�ƭu"O�X{0�V<}ስ/�Z�r���"O���۞8�b]���%�(�"ODz��L 0b(�U۠%��s"O�1�`�$�}Cp��}�"�(�"O&��a$��q����F�U|���YF"O:ɺ�I=b}Mɕ�/��	j&"OH�����H�IL�p�X�P�"Oܤ	b��1T~܁�2oU2h�i�T"O�3���3�`�p&)�6�2!a�"O�)ңp���&Ǐ�xX�9�"OJ�K���46�-XtK��j��X�!"O��P�[!A0��dk,���"O�!�3C7E�B�C
H/�ֽ8�"O)v��PԦ������K5"O,!Z#뎯gizL0�I�L
Xɰ�"ON�
��>쁻	_�t��W"O8�cH"Q����&S�wTUiw"O�}��*U�8����ӫ �3�zYs�"O�r"oM� Gd$թ\d<n0��"O�0h�M%7�N��F�'f�4�yG"O���%!A�=d
�Qc��'G���S�"O���l[�D�Z�A��Y��"O<D� I�3�$��@��[����S"Opyq��:S��5*�/]*xpD�T"O4�s�K�3��\)7�(f�	@"O��F�[�w� ��BJ>,ZN��"OD���΍[>8�����8b���"O� S��e[r�Ca
J���aQ"O!ia�ש{�Ό�Aҋ���"O`쪳,�^�He��ΐ|wx({�"OE���6�+e��cN8��"O�嚁a�����&�./4�4J�"O �ВlIr�m[p�ǟ3$q��"O(18�
�=��U�dƞ� �"O�Q�c��Va�p��C�_���P"O�X7Ɂ�U��1f/�����"O\��B�S� $е�?Uߐ�T"O$A�$�5t+�xY���=���BP"O��Y�'F� �&�U� ��ոd"O���9ټmE��D�Yْ"O����m�\y� 3�PI[�x������3���t�T�N������	��'4ꝰ#�)�P%��'D>
E����'\��񣪃w�x�DS�l�J`��'��t��D�,?R-p ,C?Y�^,a�'�,dB���2>�!���N�z��'K�qz�&�@�0��"	-B7*u��'��Y���ӒmN#�ez��'�����ŝ;:�6d���L��vL���� �˴,Y�d���7K�K�2�23"O�jdK̲Y��-�����W�dy@�"O��9��;� �4fԲm�R���"O���dAM+@��U���q�L-��"Or��/B6j>X8GX���	{�"O�8�R��Y͘e��Vb�L�V"O:L���
^:nAzЪىLV�"O�RS�Q�H{�������"Ox�CNޕa���b�R���"O2��viٛ;E��y0 ݛ.a8��A"O�=��a�k���b$�,Pr��d"O0=2!c�(}��I�˖:9Ѝ*�"O�y�bC�=��8�"J�m��D�"O���ՃˊI-bL�S��N� H�"O��R��@|�8�#f��V}3�"O
�� �ŝ3%�h�T+�G�L@k�"Ot(�� :X�H#�ܹj�H|8�"O�M��"w���T��%D�̂�BA:�Tl�+��4 �#D�<)���r)ؙD,�;"�� �RD;D�l��eQ:<����H91l�蚣D9D�����^	bb��3��^��Sf!D�c��G>�����f޷QҪĠT#"D��s�ķ@��l�S��$�n�G�!D�\��mB$#�`q�A��m�Di
�  D���F�t�Y窀�Z�<Qs�m/D��`6�d������#_t�%P�/D����o?��f=I��сD�7D����
�V+"h��"�C�ֵ�t;D��{�&�/TD�DI���tв�Zeb&D�p�`痘{�,�9s�ˊ�z��'#D����O�wC(%��	7Kl�M���/D�����%M͖�C�)V 6b�@�g�,D����E
t��G��J�-R�'%D��v�Sfڸڤ������D!D���d��v��c��6V��p��@<D����&���q���}��S#(:D�h�DO@64
*�Ȕ�t���k�&D��bE�$ t���f�n�00D���$ ��8�� �b�X$�N=D�̹kS-1���;�'I6pA�L�`D;D�d���A��� ������N�!�L�8�
,SA�bLVL���Y
M�!򤚂o��@Ʉ.Q��L8�	�z:!�$�(*hh1�=�P�
�&!�Dݎ7�J��'(���T@ ��-el!��B;9J�d��%\�g]�����1!��W�YV�r��ȻK��R��Ө1h!�\�n��a�J�����$K 4!�d��o4�U1���Z���Je��V%!��͜g�2��E�A�tI�0R#�!�dH��� .F�*��)�ȇ �!���=��a �G�|�ʖm�y�!�TH�[��
�8�:��S	8!�	0b�HB��A���C�s#!�r�洺�Ē�0�④U�֚|!�]"l�~0ꓩN=KvLq
�nUQK!�D;�n��@�E��Qpr���I�!����B��wE͕o9�pȟ !�Ƣ%W�z����2 8j$��8!��@4.L�5��3⁳㭌!�ė�=f\ئ	ښmxn� g헥`w!�d�ڮ[�,U�}�� �A,t!�dA38<έ��㜄k>BX��!�g	!�� �(8Ō�� �5C]�m����"O�Q�mH=jsha 1Qv�d�`"O�YT$)�܁$�B(2fr��"O" ��CN��(b� q}�0""O����eE�7.΁����Yo���w"O���@���=9��Аj���6"O��cŌ�>���A kޫ��|�6"O�x��苵a�мc��� �8�"O~h�+�/g/�����ݙ:��1�'"OND�6d�_ �2��ۚ&�N��w"O�� g���&x������.:�3"O���qLA�xs8}HB��"�� �*O��0 םY�<u��
+���'�n3R@\3N�dYӻ4 �z�'%R�$�����Q#@�R�e��'��B׀�$|��-�H ,�c	�'<,yR󮄹q9�`�P�Òt��К�'"�Ss��r�a�&��eA���'W�Mb�����5Q�OP�����'��Rc��������Q.N�:�'l�=�` M8;�|��K�56�$�2�'������|�PcD�r��'��:ƪZ����Í'�vL*�'��s��ܱt�@���b�?g���	�'(��l)!�4u�皝.E"(B	�'����mY9xtP���0)�����'k����)6T�GmߊW���S�'�-�ׁ\�<J���7��]���Z�'ߨt{7�*U���c���3V��$a�'�JP�o� ZeJ��GP����'�����8D��!-LI�|��'u�xcQ	�,��l�v
�|�z���'����Җ tTI e��m�+�'+� k9Y}Z�A�O?̌0��')��@�[�u劉�đP�Z�'��� 4+�"XS�jN�<4T�@	�'��!�W�ɫ/	0��<0ZXC�'؅c��U
Ui��(�� �<�5�	�'��8��M@��y�'J	f,�J
�'���J�"�`5.	2
S��'�85�$J#;��q�[��(��'G�}�AF�3S�
��#ޥ8���[�'٨y��
=u�8y����/"2����'���S	9���#]Mɔ�C�'�p��E��boR��c��1Z�h	
�'�Q;�*A
eBL��dJ�Th@�i�'�*(x��=kI�N�Im�L��'��"v�m
�u��u JM(�'J�ڧ���8v@�td@/="�9��'M��!'�\&%4���#'5�c�'_��^�=vu�vҍ0�4%#�']�g�I�J褡�N^�/(.��
�'KT\��N��V9Ό�a�-�@�
�'J�LA�MH�L�j�hC�%JI
�'�����������CF 0rp��'�5��cذF������6`��c	�'��R���n��d�T���jl2	�'�iq5��?��P%��;c=���'�D����qZ�#��=-N!��'�¬#5 F�T?v8!5���4�����'t,3WlS�P%
��O�,�Z�P
�'��5��2��s`�4^|��'��0�ƅ'��x��W�O�I�'= �W
w���Bǋ��N`* ���� pM��c:	
r���-��n��B"Oz��F��4<zr��'���!����"O
�ф̊6sD���G�MӸ���"O<a��$1�h�rw��|WA`"O$���7��!'�!@VȰ"O�۳�V�'/F���f��j�����"O��娏v@ ڄ�Y�F� ��"O��Cb �2�Qz���<P�XX�"Ob�35�ƅG�������'"O�5�����Ru�, t�X�qy���S"Oj�s��?d�i�E��t�
�"O�ػi�Xܠ;`DF�^d�Y!5"ON��L�>s6�K0+�;Nl	�"O����L�%���b��#�0�"O�L���At��%(��K�����"Or�YU�W>&]
�2'&K�1��0�"OB������a{@���!W�jD�"O��wl��'�d`q�-_</�Nq�"O49sč�9r��h#oW�+����"O��Dgҟ0�L0��@�*2w|�	"O�Q�c��5 �)�	��z���8�"O����h��K%6��pjU�Z�1"O5@4_
���1�	[(:���	F"O\�Q/I� i�$!�$���"O�(b�%ū
�*�cDo�s���q5"O~�CD�# m�D���.,d)ʓ"Oȭ22&O�EirsFOW;85"O�li�$Y,g��qPc�#d�p�"O, �ǈ3; �j��B�u|�8�"O�@ka/P�Ie��S��p�X�G"Of4�4gVb���"�ޑ9��"O01�g�,�cB���"O� ��J�9aF+5��0C"Oέ���V�2����N8&he"OVT�c O$!���@8u|1�G"O<����Uؘ�(���A�\��#"O蜨�c��:��|)%��*����"O����D�:�p��ʀ>-p�$"OV�S��_�a�ޑ��J��F�<�z�"O|�d��Z�JdrG�� N�����"O*�𥅒�g�h�CרNU�RMh1"O܉2�@Zw�Àȇ1<)H���"On$"���7;|���L��!�w"O�0"ql$zx�#Cl��	�r��"O�4��l�s]S��5�>��"O�E��J�u�)���W�E����"OL��B RH'dI$�5o�ơ(c"O��H����x�T���H�	Cw6U��"O��I��-`2�߰U7.�I�"Op"d�W!;F�Ab2���d*�q2�"O��R!U/[��w͐�g^X�"Ot���l�h�*"��	(�"O�U���ZM�Z���ha��"O�u)���gt|�`��+f��R�"O@aՃp�H�ߎ����1"O���B�Ƕy{X���G��( �cw"O���Q)7A��˶hN&#h��"O�h�M�8��S�� ,�ܱ�"O�q#���)h����
M>;'0�"O��w'��-6,�0�	�4)�JEx"O��kb^�l�4
��
�dBr��*�!��U�0��d
�Y0U��'��v	֠I��qB�ޒq��Y�
�'�	�N��*�0!�%�4\��9
�'鲹�s W�(LD��TGτF�L��S�? p0�%.��k6�ܳ�'V/�ּZ$"O�Z!+��\��y�'ٔ+ҖD��"O�����>>�I5fۢFà} a"O��q� >Jl���e�
�����"O������B���2"V��y��	6��V�k�f$zb��n::C�	�)�H��aC�3�l��E� .ZC�I?�HDpϚ�Q��c���V��B�<0M���oU�6��K�͚I]pC�������X��e�F!6T_,B�I��`e���g�LC7C�7vLBC�I<E&Q
����xD�P�"a��g��C��� �f��<F�L5{DoD�jgB䉍8����tk,B�C�F��C�ɉe<� �F_�}I�Ր��PiJ$C�ɍX4��9g���yΘ����(>�.B䉏kD�ř�lD�`�87�c�C�I�}��\�F�ξ%(���FÇ5V�C�	��fx3Dl �>������%C�C�	��6x ���G)��.�z�hC�I�}[����ؑh��x{��XB	�B�ɨn����/��\t�ф��ҴC�	>xJ^Ac6�K����l�,	1x,�����sMU�)y��0j	+*������1� !݌$(lx�K�JX����nɮ9)�Q�8��(�M%W[���#k�	��k��0�֙��
�$�$��6Ժ�UF]*Nn��tEK�x��ȓ\4�����]�@��F�Q݅�$j��֧��khn�s���ZtL���4e���J�e!0��*]!t����ȓ�� �Ф��P)����aV�
�*��t�"x���R:��iS�d�=�����?� ��&q��� �c��фȓ9�4D+W���u2�=�uE��[3���ȓ\lY����d�T	Z0� �4P��s�W%�%��ѱ���W��%�� ��B0	�z���)ej�e�����-H�ZC��^AZ����	�c�.0�ȓF���k��?��Pi7E��`cD$�ȓu&*YXBAQ�բY�I�",y��;�.9�W��0)k�B��K����>����FJ�s�B�p0���,��Z�DaX���D<>����N�|p����6�F���"п=��٢L��<4�ԇȓk�!J�	��@��P�I��L�ȓ�F�t��7J�9(�B��䨇�c�>)���֢9�Dų1�
B0��ȓQ��9�`)H�s�Fu�"^��.l���P�yf��#X�:KoF�8��h���XX������5��]�؅ȓ ��,���IQиq�J���8��ȓ0R���g�5���ѩӢ$�6���~����E��/ΞHHd�AZ���ȓ�耦�
�����*:@��Pž��h@ S8,�)�nM�hMN-�ȓ&�������iԂ��D�!�(���i��ؓ�gղ]t�(�@��>S&ȇ�\�J��o��`���S��p-|���L㔘x�[.��J��Z�+h6��ȓKی�i`(�;yDN�"�B�?��لȓ�2�Zo�j���;#�	�N�\��]��8���7yR�BIK�P��L��1���T�+`|8�t��2>6�ԇ�S�? �s���4Tb5��V�r�!�"O��r�Rk]Zs��T��x��"O�(p*�*~t���Ih�"O����[},5�%%��2��;s"O̛��.�lL��c®�:c�"OX�a� ��=���r&b�n�N#�"O�iW�G��R���E�Nm�X�F"O����V�\�F���
�
5
���"O�b�@��%�d�Z��8Q"O>,�$�ׯx
.��A#`ج�"O2qI��*	�TD�d�ʷHp(��"OtT���C�G;*a��V�-c��[t"Oܨa5!�.^4j��u�B,-��R"O�y���S�
Xh��J�k:� ��"O^<B4��/m{lX�D��^:p�"O�eq����L�7�	�8�Y��"O�m���_%p�z�
p,6���"O8-�F���ۆ��E�܏]���W"O�������� #s)\$gQ�e"OЉ�t�ä��So�S}�q��"O���E�.��<Z�HLgL���"O$��#)�&~Ҙ;&(�`��h 2"OJy:�a�|� �9�Gϰ*崄�4"O�xW �FbԠ[�fG*;�di&"O$�⥉ē��\HW�����ˤ"O`�����#B�.AhS��25��u�4"O� ��ض-j����R�E�"OQ�wdM�[z1٦k����R"O2��tfz6�iT�
e�>ݹ�"OzmiLA�$��� t��%K�eZ�"O���@ݷ,��ŏ�)*Шx��"O��HG�Fe��s�o9�����"O�y ��	o=��H�B�6��"O|4�Q��-��'�� q�r"O���
ޅ vT|a"��㰴�&"O6a�E"PM88�dկ]����"O���r&µ�]�q��!6��aS"O05���k6*w��v�n�;�"O��yV��N�⧬W`�.�A�"Oʤ�@�L�&ox�`b��] (��&"O��rD�Ӱ, ����]�0�"O8�␌�B��u�@(@�uc�"O�1#��:Q\��hB@/%ŰQ��"O�r"(ֿC��pS�H
.��å"O�e+���$s&�%�R�Q�7�x��"O��a��"#�:݋#�֙�@�+g"O0e:sE	T!8���,�<14Z�"Ol�'L �J%�i�
�[F��7"OJ,2�:u����)�Q�dYb"O��掏&0��A��Q���"O�5bBi�hvܒ�N�@���a"OJpZ�d�,I��䭐%�Ե��"O�� #Ü�P^�Q��H�_���"OX�;�-��]����'^g�� "OmzAG�%w �5���QM����"O�s#EH�vu�)�r�>8A�]��"ON����@l)X��45����"Od��Ǎ n� 4!���4�I"O�r�φ�~�ZA�ŭĦ\pv@��"O����Z
)Ǧ$� �8]��Y���'(��D��١+�e:Ŏ�- ���D*-D��SW�@4zZ(�B'�,�t�p��,D���q[4\0-��*9������ D��QIԮ$/�\;t.[�U@�%���2D�� ,�:��ÁRn�9�˕�L�H8{�"O�Ur��	�u嚠I�
ƻ���X�"O.-0�D�D�:5c�DL���0�"O
=�`����0)K�Ã �P ۥ"O�R�#S%��T��1"�6Z�"O* ��]�Ȟ��Y�x�V"OT$���G�Jl[���J�$ə�"Oy�0R�QI\�cb� �PL.D!��4�t!)��S)%b����G�@�!��$sP���1�ݷo��}i�,�/$!�dY�w\L�KJ�$�|q5��	�!�$V�^���dP2�>1�JX�'E!�D�Z�y����bE�Bi[!���%�z�iQ�MR�K�(U#�!�dջT:ƍ��ʦW��U
�Z2:$!�Ĝ�<oV��B��iK���G!�ď+_M�H��
C�$~���e�	�!�䋈F�("T��Xh��ЄJ�
�!�D�)6�x����?l�l:��Ӕm�!�d�> 0i���E�P��5gR W_!�d�9e�JX�C	F�!Jh-a��A�!��#4p��!@"\- ��P+��=�!�$F-o�=���Q�xҎ��G ^!��3K�lY�bE=i[j�p��eN!�Ԡc:�: �_.w�lh#6gP�h�!��Y�mpPe� O�/�=�w��k�!�D��՚c��:XD�� �Ԍq`!��S3nH�dJE���iIV)��$�'*�!���4#V�0�JΆs<ZH���;�!�$F$`d4� w)ZbC>P,|�
�'�d����n��C��̯L;�x �'�!�an�|�x�tRi�|i�'���Tm�^rLa�@�H�zm:
�'�t��	Q�B�xXP�I:�v���'���#�'�9K��j����+�6%��'h����号a���k����2Lh�'
��"�ŝ�v5ȷ���S	�'��&�0ٲW�$�np���yr`�\�ZH;P�͟%�@��ʟ��yb�Z06��e���� �����yB�Z|�0"	�4Z�R�J��y��B@�d<�b��M�Z���y���S��T�D䀎�
$�1��%�y�AD�[��YQ�߶jFDA�yrBŮz�Rh�%nU�^_�ó�Q�yb��w�R��Ԫ�Yy�lRì�y���(��\[�(��>�ĳs	,�y"� �P��1ś2;Q�= cBז�y"G�5�*��A��9����F��y��V���P�gˍ2�P�B�F��yb�F.Y�x��E₣#�K�$�y�*)��; Ր ��,B�f��y"$@���P��^�A,��v�R��y(�&5�� �Bȸ0<��%ۺ�y��s� ���o�p��őƄҩ�y�-mD��qsl�<d}����+�7�y�l��3Ffh�4�ܑ&7�������y�^2�BP�5%+�8akg���y2��1�r��ā�K����˖�yr�اZ
�p�F <K��1���y�K%���0j�H�Q!�ϵ�yRD�����)jW*G��%��y��E�q��Is+�=���`f�Q��yB�Ӡ,-��)�!Y�e��1WI��y
�  ,0��ܹ~���t�8u�9��"OU���)_�`@ۭL����u"O�)H��A�(d`���f�l�;$"O��3uG�R)��٦!� �	P"O�����F|@{򏔕Q�>��"Oa��� <��M�4q�(D+��i�<q6B��FakG�)0]�a�<�I�O�6Yp��A�N�y��u�<�Ӌ���+Dנ��n$/�B�?I���@R��X.��b��5�B䉪a�h����!�VE�)edC�tְA��n� "��+�+C�.C�I5M%^�iצ �s�~��᠂<�C�	� a�Y����W�&����Ld4�B�ɺ&�9 �Tdb�L�u/���zB��"ؐ=Hql�L����ކ��B䉥��Y1L���$#�m�{��B䉨8.D�q������۲
�3ZL�C�ɣRqt|���2�������&B�ɰq�� U퐓P���bhX4Q!�ڎu$� ��	�}��h���!�d�U� W���t�����!�Ğ�AK��+��(P�'%6*�!�� �v�[�E�R�(A����!�G��ʐ�+G��U2g�[��!�d�)����o0E~`)(bc�>N�!��϶'��}����;m�Qr!���!��]�G�Jek�)S��[Ҋ�	 �!���0S��Rt�t�*uF]Nv��'~s�gC���k$�F6E%��(�'I�8��hċ �^�Q�GZ�B2�h+�'0���.�n�Ȫ��Ƕ3��h�	�'����٬n������[�@=P	�'(����%#z
��WQ�	�'�>�j��Qڀ{EI����Q�'߀��1ɑ�lHT�t�G�(�V�0�'� �T�P2y@us��.�&���'� ������	����/�>�J�'����K�\������5��!��'�بJ�OX��Ic�V�6����'�Z #���� �� y@n��.H���'q����V�)����w��Z���'=�=x��Y����z�阻)����
�'��0�aU��d1p�I��#zT�r�'m�t��T>\R`�����q�'���Dɚic@ ����	q&P�'�%�I�8�9��@��5�	�'���[��H1���j�MP܍��'�d�BN��^���ա�y�J��'�2@�@�	
^|���ʬrn4ua	�'�^@�w�]2"����:�A�	�'R.3S�Q�,Uuj	69բ���'z�eP�ބQ `��/ҳ-B�ݒ�'(v�1�G��`NJ�2E��&F�X:�'[��KG��0&ry��D�+7��A�'��!�3,2�ڨ��`	(y>�d��'�4�!�2���h#�W��4�p�'�NQ���0SF�#s�F;��ͪ�'���"H�h�Q�� '�����'��0-�\���	NMQz1j�'��dr��U�.\ 	�S&E
HP�Z�'(�YQ-�?e�	P �S�F5Ш��'�8M�Ǝ�|=<��JI�(��p��'�>��ᫍ�r�.]�vMB�p��J
��� �ĉ!(S+0���rTm�\���@R"OS�&�@gf���
�FJ�@�"OP�s$k>?�H��ugz�����"O�M#!�	>r�H�2A�N�X�*p"OFu�U�]�j)����K�>��٪�"Oh�"�(�$ {!*�h� �Ѵ"O�2��׼|H]YJ�@B<b�"Oʴ��EX!O�F=A� +x˨�8�"O���a锲{K`����=�H�Jr"OXL��΍y�ڤL�+d���83"OD�󷇈9^K�A ��&AT��"O��#hÑa耸cTj�>���"On�ӁA�O>�*0�ʅN&r'"OΑj�M�ET	�N��,k�}�"O$T�n �s����lѮP�(�w"O̹��8Dƨ]�#nѹSڌIx�"O.0k5`�h@�ӭ�x�l�$"O���VJO�=F�B�-�*&t�J�"Ov��7�ę1���!�?V��-j"O��!���6�����ys���"O���#H¦X�!`_�y�d%Y�"O�	S�ÉN8B�f+[�,��!�!"O��S�#�Vi4��#�ʫm��	�"OP�(Ԭ l�� ��H�p����$"O�{0{��|�r��e��X:�"O�d1�	�[�]"��T%y�����"O�P@���1醥"���`3p}��"O�����801��0��g�Pd9&"OnP����Ԑ��PW�:PIE"O��BMU�������x�'�ސ�R�hl���ǟ�+��Q��'4�}�G.y�F�
5X�(L [�'U�E�AL��V0y��A4�ʄ�'�>��S@�;Wl�R�EN4���p�'KN�QI�D�����DF?�d�#�'v<�X�d�<1�]�č@��R�(�'��Y�@J�.��s���tz6y��'怭@�O�=K�1r�h����'�pأ'W�Z���	�����,�'y�+��?�N�9&�C� �޽k�'f� !���7*�h���@~Bֵ�
�':�����;A���z6��a�䨲�'�2�xc��>
|���n�T�|��
�'����iʭzh���E&@�	�'�t-�G�I�I��%����,r�'��bq��/O�8��a٥p��Q	�''|!�R�Ǔf�vH@��L�y!"t��'C젉eK
�x�x�GG�w�&���'_J�Q�*� رH	�eb�J�'�ȡ���ɿ"�v\��c�91�N%c
�'~���&
"PH���! ��.��'��9C¥4w?v��PD�%*O���'dx����'����V��<O} 9�
�'wN��E�^�.���Xv�_�?UҸ�
�'W� ���	q���@6���1�t`��'�H�ђ�ם<���H�/���b�'�6����\�>Rd��F!4'�2չ�'���#��ǻQ�8%p7�y�'�ڡ�cTT&��g��$`J��	�'N)�PgW�=jD�:�`��R�x�p�'��{�A�>����q�W����'����=�htr�K_�U��C�'�h=��
De�M!�����y�'5���q���z�3s ������y
� "q��'ǣH���r�>OW�i'"O|<Å�߉�P���E�7c���Р"On�#� YM�P3�د9��`3"OrD�'�!{\Đtl�1x�Լ�1"O�I�Dg�]�B��bF��M1*O`�c���q��$Ȣȇ�*vLQ�'�8�x����ԙ�c��l���)	�'�
��S%���
�Jj%\��'ub�ۤ�N�,T�g�9t~,��'�`|k0� �q.lu��!MkkX !�'��Ygh2.8P��'
_[|iA�'�*���3}Q��ꁣ��%^���'kH��@0}�����$�L�'Ƥ�S�S�v�b����gJj�*�'nj����6�rL���d���k�'*A���C�yW~���ͅ�U��$!�'��%�fCJ�%E�pkA��N��!��'Z()Eˀu�*����^�J�C�'��ZDnQ%Qz8ba�A�I0$	��'DBl���ΪH7�-8�&�E��P�'�@m	F^���� #�/o�޵!
�'Ȱp@��3�,��֩e|$1x	�'�VIxqa�2D|�1�gNX���	�'f�9c7���Ż��
a��`r�'�tuRs��*D��ub�I&T�> �'���!� *kh��i�	��Gجuc�'�Br	��´�x3��qfщ	�'�vXcr��8L]d��5���$���'C.��҆B�T*n�+%j��<��'}"�"R$ҥ"�0���N�,��A�'�ayv�"@&�@�'@��x9��'C����A.*�.D9��P���X��'����(�)Q`T��KٍP\*`p�'؜�9R�а7���T6P�h���'�٪�L7e�������,=�����'��P#���H).�u�_�4�ua�'2� aA� !:���*���-��'L"��ׁ�-�4 @�i���D�y���*| ��#�}��:��2�y"Mϧ�P$[$cX-iZ��V�ط�y�H��1G�J�{�j�a��]�yR�	q@l�-�v"T2�k��y�H#PU�mq��Z�us(P��)���y�H�+b��*d`Ưs
ؽ��$Ћ�y2�΁��u���ä7��ԓFo�>�y2�W�N@0Zu,�73 ������y��Vo�@bl��+мDSu�ŭ�y��!]��T�2&��7���#�K��y�E�%<�k�9/���EQ��yR��fg���r/؇S���k�.Վ�y��� t���3R$�M�ꝫ&CH��yi_�6�~�D��/�ƍ�֍�yB�U�]�-#�c�#-MH5��'�y��
j^d\�wÀ��t@�1��yrkS�z��T�q�Z(e ��	��y�"J�M!2�!0cǂ
H�ʁ˚��y�.+F�jaH��-��Maŉ+�y�	�_� ���"T��������y"�ݓ��S�.Q��4 �M�y��4+.A��(�]׆%��?�yҤI�7�Ԡ"��^�Gzi��ׅ�ybc�`�|�y�%�7�@�5�@��y҃�: < S��N�/��xU䑠�y��G�"�`m��(�* k���y
� ���Հ�#������=0�2"O�5։�{�J%�CCW�]7���"O�I��9]{�<�sa��+��pf"O�B&m;z
��F|n,J"O�ES���k1�a�� �(t��Z���՟�[�EА8ߛ��I��Y3b���EW[NK�F~	qO��$�+4E*��b�ЫDI�����5n�L:�Oj��r'�W.r� ;��J7>�%���d�����I� %\��ף[I�DR����#1V0�� ������vnG���Gz�ݑ�?q��_Z�O4�FM�5/xl+��X�ʈ�P��1g�H�D'��i�Ͽ;0e9,��#�I����qS��e8�8i�4G���i��;6bXC�ɻ�0���p�'�~���O��ī<�O��'>�4c"��Ox����N2����CH�\��a�E�j�@���:JT�����Ͽk��M������2�>���צ�P��цo޸(a���6�Bٳ���6s����\c�8��!CX~n6���1%ut���44d��I��Müi���s��D� �yT`ve�F;�(��O�D%�Oz�a��҂V�x���H�������O
�m��MCH~r3�]��u�o�He(UX�!�u�8J�I˰6�Pʓ��E2`�iYay�g�%H�n;`�[�} `�uB�j�����[� �^E��ϛXĴ��G��lYz���$+s��s�i]�"kD,"f����{1gE#�8�2�F��Rt���Y?��ǩ����'Y��)�
�N�l�#�/�x$�I˕��O�����OZ�O���Y�D�	Q}r#_�7����v��7t��q�>�y�c��\\���5�
e�l��棉� ;xr\f�l}�i>q�_yb+_<�����cj.}*3��$��P�"N`�R�'a"�'B�X��'E�'�tԠq�iऍ;R�7V��{%��hW y�dg�,I������Wf����$�����ۅ9B��I�hԫT�q3��= 6��"S�2��B�,CD`HFzc��?)ߴY<�Q��M����UZ��ʸ�.�W���'��I�8�?�OB��a��,
��|���[�f�4���2�����`0�A�Ь_�Ki�H!���0�(����MCB�i��Ba�H )��O}U��n��?j��pm�?K�iS&~rqO��䚫�Y���Qz��91�V+q�~I�O}yy��	y�}
�kG�k�H�Њ�$N	�t�$���9����5��5^PD��3N�KӚ�i��Y�l�0��0�*1.�uFz����?���0���')�S�W���J[Ha��Y>N&�<p�oL��?������,L��_�&�FD3��׾SU(��R�'h7�ԦAo��6PT�q�%b�(a��|�����':%Pc�OF��|z��?����MK烝�=G�3o�
Z�Q�ܷt/~�PCà!��)�g�� }�tdb�/�"��e��r��%F�Ԉ�O�U�
I�@�{�pt��-7�� L_:)z�� )�����\c��ę�_��3���?~R�B�48R���ܟ r�4�?ы��i��9����[��1ipDU�-��!��'J��'�ў���R�K ��XE!���S��+Q�	�M�Ӵi��'��ĺ��F`��-�� �1B�~��L�I}؞+
   ����0d"̍�I���p�{1��(�O,��O����˺+���?)Eb��X�"��31���Qr?٢�4�Of�q�и1ȠH��ݝ?L�� �O@	��n
�#ڼ?�1�'Õt~�������	���$���	�t��ґb����H(��,s�vB�I�b�(�0$�,؄�@�΀kV(щ��?	�'a�`�s�xӜS����C��i�`(؜SV�䉴��Op���O��dI>3��D�O�d:^���O���,�"���p�\�ydd��'z8!�.O؈��Eb�p��S��:5�,�u�'�ܔ����?ab�A�{"}�� �^��SU�g�<�rl�%=�ac&��*�h�]|�<!�PN	2e���Y��-���<I��$�)QֽoZ�$��W�T,[DFhY���36^})v�u�C��'���'w�M8�'L1O�S4)����N�	-�l����T�j���<�DLTm�O�ڌ��b��_1��C�?O�l����$Ʃo�R�S�fpT����ƻ7�LD��P�rB�	��p��^�u��#JԓO�H���Xb�I:?��9���"*+��Mܤ6BB�b�jw	�*k�ؙ��o�>B�)� ��k���1Xk��J19���;W"O�Q�#�P)MG
%��NV
B���	C"Ob� ��UW���sd�&\��kG"O�� TH�2l��	�IfVa�R"OBEa�剩b���#Ѹ�~�	@"O�d@��D'ԠK�-�&]r�x'"O��'
�*���y��Rl2�s%"O|�Em�!
�L�@�YK�<pr�"O�\SR���{vN��S6y2�"O6L l�@QT�;CG��-�1"O�����Z#Xꐚ@g��3P�"O�%L5$6h)�b�D%a �ٳ"OZ�auf�ƙѤ'���z"Ofu#S���i:
����'?x�3P"O�:TL�/e�X��e	 5�9�1"O�Q`��	2V6�����*/(n�`�"O���(Z�!"df.s(��4"O�U(D3`���(���(�U1t"OB-� �E ���Y�F Zp��"O�x0�ڛC��1B�@��Θr�"OxD!��+v�&m�:'�ԁ�"O�m�$�@.#�%p�,���y�"O��%$��s^��d��P��d�"O4�����sV���2(����"OƩS�+E�/F�"��w�JpA�"O��j�ݾn���`W2�B�j�"Ox���]f�{�!p>e�d"O��@&G�&t�0��]��C"O�kA ��x�&Zs�T<V2���"O�4�E�@����RcS-1��R"O�f$Z�+f�����,<um�#"O��h3MLhަ�9�!H2CktU��"O4�'E�T���K@�܌%k49�"O6�2p�����
g�.U���;"Oh@�h44Ђ�o�,bc%"O�rW��C�0�[�.�4g�x {5"Oy�s��!`>�P�]9�i�!"ONR�-~GX�q�L�� 3�"O:8#�HA���'�<b�>�d"O�} 'M���R���*�>;�>�d"O� �lܷ_���B�HKO�iD"O(��d�J�lD��G�T�\б�"OB�{�O^�I��c��k��(;1"OT����� p�D�&D��0��I�"O2H�w!�l_|P��"H�0j@�"O8@H�Ő|��r2aH�2�꽱�"O0�����~�DS�D+Da�:A"O��@bm�;$vT˗�ޤo!�*R"O��!H��
���H��Đa"O�1�V<��`�w脺�!�Fyr��1H�c��|7���{�X �⌍��;5nX�<�DCPh*t�!tBw�Ra�Љ�T�	s�BA�ϓZ�Ab�)�?w����U��25�zP��	�{R�a"�(���L�e���4�k3��#��x�Ѻ	r��bu����������O6���_�'! ���!�	U�"4X�L�~K��!Q�����~ �U��f�<qb|��'D�0�m2�)ʧ��%���L+���:G��h�H��ȓ-�<C�(�Tr��J'Z�~e�H$��
�[���<���t�d�����K�
x<���$$����@a��:k|Zw���k-nHbO�	4�R�F���u�;�p`@�"O��pM�@�
Lc1$L���tq�"OyK�j��D?0��b�(�| c"O� ��XqKעUVtm9AL�P�p�"O&ř`J�%vZ�2C�H�j���"p"O�){s���x$�:@�����8�"O�]�IL�2V������
�F �"O��� B��u�ʝ�㧂�
Rr1�"O��;��L�Y8��Ɖ 	nu�4"O��� �����6� H���"O�mC�-�>)~��p3�@�Ҁ�R"OʁA$D�Z�<}���[�H�8��0"O`� ��-�9H��N�u�DT�� 
.<��ɀ8�� zVj�1rF�E G�[3m������{�O�,���A�"�(�/�(7:J�2u"O�eڀo�<-��-�.R�^ ����$Y-B�⟒��%�g�C�ބ�n�<_(Ӄ"O�"��c���]2G��n�k�Jʣ|�')�����[�d��b�^m��' ���0JמJ�]ڴ���M��U����d���"H�B!e۩[��i8��Veq!�$M�I4�R-�1P���FY�!��?8&� ��.�4�Ԁ��f݋�!�SG�������W�XP�CLٟ^�!�$Ӳ8��Ŋ6��y^��gj\�%!�$��y�I��a���)��1!�D�+(�jՂ5垈zF8�i`遧#!�L�0�l���wH��u�!�L���"~��9i'�}�!򄆓̜��3S��Y����z�!�d@�6��\��`"������!�<����5s���)�!�$L==��PG�B	}��;AO�!* !�d^��dy6c˩�����F�!�dЮFl-�����*��!�>�!򤐀~�U�ТƐNj(�ЁI�@|!�d�+c(^��4$Glr�5p2ϱWu!���, 
�I�Aˎ	�P�z᎜%	a!��Q�?�Fxv-7}�ZuI��ʶ"T!�ę�WZ�Y !L�#5����@@�O�!�ĉ�E����n?z�^�)�� �!��7XHI��,��m}hȣ�ǆ`!��\�n2j�XGl	� d:6ս7�!�˱U46�h���- N���%6�!�$\�h��|p��4m�����1&i!�d�p%�5�̀qߪ��ƀ�*y!�D;�b�ɥ�ӏ"/�`Q�l�~!�Ă�La��J���O$X�Z�՘#�!��:cȝ[0$��&���G7I��y�$��"��Sr�<q7�N�F��@�Ȃ:�4q���v�<���܈2\���ЦC�|f�"��u�I�tv�bs狷�蟊���'�q�L
���	��8K%"Of�K���#�Xp{��̠9&�q�hW�`��O\�P!0�3}��r� �4i�/Kg�)2�i���xҎ��qS��8yxX){���A(q�A)5�^��+G����tK� ki|4�&�e�y�K�"oal�&�<���	h\����J�3���k�{�<Y3@ /an�ۗD�;�Hʳkv��?�h�3k�����s�EV�b ��.,[F0�E"O<��QΙ���cs�H�Z��uʒ=�OЕ�'�5�3}¡V�L��M_�m��� �6��xB�.E�@�# �O����FmI ���$��;
b���I�|�(\k� }�����W�,"��ti7��%\��D�'d�JP��9h��R/ SU,�
�'���s��U��m�0��3Z�H:����){~L47�?�J*dOL��y�ΟW쀜G�Q�t��X�I���y
� phY�[YD9�&L<iJ�� ���(P�p������Tڢ�����>K�!� �_j�<�7	�#��(���B�G�\��!<�=`����?�	��G�DI�$�-��)�Pe*D�ě���qy��+&����*V�	�6Mn�=s�̀2�BĬ;�0�3���k|�ӈ�$lqK��̖$j6��!\�:�-��Mj�4�F�7��Yf�U�K�H��L? �D�zW���%ƛv��2��',��>}1`!�Z�vF?���!�<_�n��T�!Ky>�b�ʘ�s�ӧu���3���SB��	5M�ۅ˟ c�zp��0����p<�t��k����N\�xFDI3�C��~1�R!�k�tk�oT���`�Ʃ�T0�Ft*��'�p��$�§F�x)�ϜK�ؘRB J(<	掏�j�*�RlğD��xs
Ԭ��@�J-9���L�A�N���?et��D�R"L���!B�1�����G��|�ff�6ѫ�C��
!nm��n��X���g�G;`QT(��>�I)��	���&:ofX���ϙ0Fz��'��FM��#�k�-m�0ӎ{�Զvטhq4�X*r�}*�.���I��<��JJ\E�q�ʂ3��#�
�� ��r�MZ׬-:5+	-q"џH���/Vn���JQ�g0�w@��o|>��e�F*h(Dx����ҝt��(�� �18"���
��e �'<�v,�d�
�J�,����!��?y��N�V���n�%q�0iƈ�W�剪M�D� 32\�a�њ~�#�Y�8ט�66���ߒA�����ĨV�ƍ�	�?|@�h�ą]����d��x�£��R"4����%r6��#��<	#!J3
HX!�l�,]r�y�ƫНp��5��\�t��nԚM@0�ra�V�X�'�!�	�q<�Dg͈u�ax��*-��Dȳn4V���΅&fI�Iԧh�� ���GXPl]k�m��n[�|���l~E���d�Ie\u��	�Jx��"���}V����T���Y�VݒP�M�8�!��+Nb���'���,��t���;��@�����HH�YJ�2��;LQ��q���6c�f1��:�?�:sf�Lp�g3n�l� 2��[?1qc����'Lk��1��`gf!�&��ڼA��ZH��Ab�B4n�Y�&L�s���[e|�z���$#Ɓ�!a�>)�Gܳe��4W�X�QʟXy�@�(ly�	�P=�����(Ol�@���'�|�C�H�-hWR��W>:��A�� �+-�p)M �z�ף*k �&D��0<1E� 0H\�S��(��)3��C�݀� ��'&��i�����/<�%��._��l`���k�<���P�f푰��9/3n��s�Mp?�3c�����h�*�kD��YZ=�sGDj���Yd"O�ڣ`�w?<Q����!6��|�q"O����ɸX�H��T�M��A�"Oji�bI0�BmZ�	�V���B"OVT���U!P��i�(��$�d��"Od)�H�j�����I2�xt� "O6���dK�k�L���-����U�7"Ov40��9m��eClIt�l�Õ"O�X� �̆}�P��@E�Y�hQ �"O^4��%��XURЂ&F��D 8�"O���B��?pX�H�C#Ӱ;�a��"O� ���-(�Ƹ$3B�RA��"O�A�A�)3YR��C���L�"On�	�mD,Db"eg��*����b"O�`��,�� ��z!nJ�U+t��W"O@a�e�E����[#/E�H[V"O�p fNܒb�q*��O2*X�"O@`���G�vY����;>�`�h�"O*t�r�)u���s�Ĝ|��|S�"O��g �7	ty���LxP�xw"O�Dj�L��2/��7bY���d�D"O��éޮWG��C'��2`�~L�"O�h��J$X�Xeڑ-�(�B|�g"O� 㐊R�\EBtK�)E�4u7"O��$�(n�h�3,��S����1"OrP�B,)CN`@�7�L�)A"O�a�2 �fiJ2N��tȂ�"O���G�d���'��B�n7D�P�)
'DSHA�"�"kj$K�E8D��z�ѵ �*Q�����*4�5D���A��Q��5��ψp�Q�3D�� �ܱ�)сJ����e��T�b"OT�3U��/T�~��1�Ϧ|G��E"O�q�P�.߸I��Y%}��}��"OT�8@-8^|H9�i[q, �3"O���dj�))�0�q"@�gx�q�"O�z�L�&n��M�q�K2��4�v"O�D��%�J�I���S�]	�c@"Ob5����5g���&���5K"Ov�`P� �_M<4��A�T��``"OR���Y=m���BR�; ���@d"O"��,�4i����튮$y���#"O�THG��l�dS���(+Z��"O�zP�]�o��Fm�qF���"OfY2	��1^��,�/+Fj�"O����U�/��,KSZ�"Ol�)L�5(�M�ĀP6g���P"ONX� !f�bH�v�ť"��I@"O����'בU�ީ��m��~Ո]�"Op�1 �#18����C�;�� �"O"�(Q�(;*��1�&v���"O�������:%$��_�٫"O��5HJ�B���r�GբA"O�t�T�$��x��2�2��"O����A;[p�;fR���TÂ"O���ѧ޴b�G��T��"O�GI�]4P�%�ȚP.�"OƱ�! y�Ȉ%��ln�p8�"Oh�1�� t�ra !��)ZWl��c"OZ���n�Q�
���)�;k72p��"O�1��	߅���7#G�K���yr��z��]qK�: ��\���
�y�IGj5U��;'Ԏ�ٗl��yR���!�b���l6,�����y"�,3\|T#�X�G*)@!�S��y(�(jxy1%�x��0:Ʀ��y)��f�ap����<R��z��yb  ��̝#��A6<˖���e��yR$��oZR���agNڊtr�ͅ�IC}rd�B�~DQՊ���٠q�I��y�JUb�	Q�i��l�D��HH�y����\�Ҕ�3OL�8����4���y Ԡamf��OR�4���CT���y�b��e����Ɓ�	D�>�	�'̬T��#��k��|hFɋ�	�'��LY�%�:X���� �J�'$�3�18z�����Ӭ��	��'���e� �X�'O�E���'���{�CM.��yӠ�ݎ��L��'6p���E@�R>���k�<76�lJ
�'ϮZ4BN���5��\45l�As
�'y����<	��c"F��6i0�Y	�'�T-�b�����ҡZcd���'c��HV-#�޸�#dQ$�Z�"O��r��B���1��Q:AL@�"O>E���ɢ>��D"6h��W)`�g"O�,	�%D�J:�f߆1'�M��"O(jQ*��?c�4�F�g�d��"O�S0����xY�ӆ��.�x`��"O`���<��� ( �H� �"O
�Ge��&�\Kæ�u}��""OU����.)���[�A;��y�R"O�$��i�g��"vH��Hq�"O�m���&4�NKM��<�g"O���-sf )�#f�,��A�"O� �ö
��YR�l���Qܜ��"O�Ma��ηr��5Xgǉy�*%)R"O�<˳�\��T�� ��=�n!�g"O��w(ci,ɋ7bQ?�|���"O��)P��P�P�O�3Q�����"OJ 8dfV �b�S@������"O�ay�Aӫs;�y��6:�DH�"OTUP�FF'n�6�sF�Vլɻ"O��5"Н��$0��<�X��"O| �Uƙc� ��+�X���Q"O\�02MV�6)� :�`޶O��}��"O�����хP�4�CCnFW3(Y�"O"ɛ��U.ܮ��G��oB�@C"O�]�e�V�n5&}���%4�@k6"O�|�'�'��`hE��fZ 	*G"O�L+�ӢO�x��Î(!�(�"Oq�f�̊iu~M0�H��;�����"O�mcr�?S!���AǕ;��Q"O���"O�7�&� '���\�P�"OT����؄,�����e��2��%"O�M�"�X�'QJTړoX=H��	�"O����#nFJ��UEGф�;W"O\��A���1�e�<��PY�"O�hB����L>RQ�̞�M���t"OP�a�NثZ��|�G��tv��"O0X	"�W.�tL���N
-tb�"O8:) ���yyS�G�V]���E"O ��T�Q. w��r��$?�A�E"O�U:���� ,U�7#Z|W"O���,]�U���1'mT�"O`M� �_˒��1G;]Ա	f"OԤ`Q �6�l=��=V{�Ę"O"��rJ�	B�����R	fo�}�"O:	i�o��u�LLj��H0m�B���"O���R�u� ��t � �d��"O���#��^�pM�	�M�4Ғ�|B�'�bB�r�H	�6���y4��+�'�|t�5k��~���t
�_�<�A,�rL��R@ѩ,K^ ��N�<a˜S>�)� � #T~�+C�G�<�ϔ��Z�C��8}�ƽ �g}�<�eJ	�VP�gG�4���a�_P�<1DJ�"����<.�|)c�BN�<9sE�{�4D���L�IXШ��AGI�<�!�*I�*�C�[�d�Y�)HM�<�bU$o���2��g}Pui6dt�<a0��/�@��+D�d|z9�G�Z�<���B�[9	�fD�t�MXD���+�(X87���g��ɝ
0�dh�ȓ/7nF��w��m1�J�h���e�'�D��E̩Gc����ۮ^z���'KV����+k�4�6!ΎE��'���`�/�4BT�hJ�-O�%V<�i	�'u�+���42�.Cq�Q6m� ���'X�r
�:D������]:~�
�'�T�F�v\�k��O�O6���'�yz�ě)C�՚�M����� �'���昢We)G��)�Fz�'��M9��V�)k�3��7��}��':nqd�����Xsܨu�j}��'92�7-ͩd~ ���e�p��'��z����ڙ��+ζY�����'D���A��}�va���VN�	�'�����/#$VbB@�E��P���� ��@6m�&�2]�BDԟ2rZ,ڥ"O�i	B��uS�81� ²;U2��"Oh���>Z%�5�o�9
@d�{#"O0�A.G40LP�N��U=� E"Obh:D���T��a��_�:���"Oz��fIL4kr]˔7Bٚ�i"O�Q����!h&��#�O�`��a��"Op= �G�1z�89�IQN2�#�"O���[�-�蹛v	0�R��"OB�2¨�	T��&���Y"�"O.�*b����?�ܘZ��!4��P�Ν	P@)91J�Gb�5�b3<O�7�:��##Uvz�""2��`XBh^ed^B�	~L8��O�?����D�� C��=��S3�&���,��g[x�/�'L�\B�	�3^)(Rk�Hx�%��Ba*O6q���ՓW)l({�c��?�d���"O,80���=q�9�!��V��@p�"O6}j!��\U�q�C�Q�!����"O�	֌ưz�ZQC@�6��u�A"O��(�&
$&�J,j�AT*I�
͉�"O����p���j�^�^� �"O���qH������˂�`*4�G^������/_�1q��6@ExD Y8�C�	�HB@[����89{�,�y�dC�#zB`a�Q��}�+�Qm_�B䉞)�J�A��o���"�C�)"�B��R8�pC�=:IbMpᎍ�&����%�$O_����	6{���
&���cd!��p�6�P��X�X���p�J3X�!򤑟Z�peЦ`�T��T �7L!���Ns�T���%S��j��ؐ/�!��@
���y�
M?Ch�W�AU�!�d�hJ�M��a�����,��!��+F�LaIaL� �%j�!���Z��` �'��U�g��#�!�D�����1�Õ4}��M(���K!�	O�x T��aC�Di�۶-!��
��l�X�B"$d�mT!i-!򤆄�0œ%J�-�ȉ��)]�c!��)I��y$,�?{��mRU	C'i!�S�4��
b�S
�2�G�Q!�$R2�T����R"A�Ap�M�rY!�S�>�$a�/��y� ��R"K!��J=}�t4��D�J�Qx�E5rI!򤖜I����O_E t���$I/!�D�8`�Щ;�!�-�(�'m�Oy!�D�gY���b�C���=0�N�>5W!��^`��J  �m{���$�ŏ�!���8*���:v��nv S���~t!�ą3x�a{�l�l��A�A7i!���L�`�&"U�0=��'���P�!��ſi�E�
�T�8-�r�W?�!�[��j�O٪Zr�1윭*!���*\	ラH
/e�eR�h��5#!�U�J:��r���,hma%�#b!򄛱 DyJ�J^����DڪC!�d�3.N���D����S��B>%!�d}>|4�cq�����g�08!�DI�c�ŰT��+*�%bE��7,!�1Jj�D��nC�R�J��O1#!���f� �ie� �����^>e!��б$*ʡ���D�d�i���!�ݭ�<�aoɠ,G��g��{�!�� P���S�&e�l
�I�2&W�y�"O|���V n}�Qk�h�=)TA!F"O،i�F�;3�����g��w2��"OR������$h�H� $^�)�1�"O�U���P|�%Z�\�D���"O����M�{h��pPa��L=�"O����(#�@I�5A9��Aa�"O�|��iܬ 
J5�@@D"�*8H�"O��`�A o�����@�.F0�S�"O�#U"R;:]ۇ����E ""O=r����l4�PNڶ~R�ѓ"O� ��B�`�h)iDK�O�D�#"Oj8��F�,2�U�Eg�o�U��"O�U����(~����fR$m�(5b"Or!3��l��!���?vNP�"O°"&�נS�l�H�
�)8VU�V"O��#��t@���WK�W<�R�"O����Lf�=���U�4��s"O���g�&^[2�9F��a�}��"O�1 ��X�k�`KB���4�N8s�"O&Ixg�8�0p�Q/�.>r�[D"O��I���vp��2NA�3ؐQ�"O 	C���2�`I���@g��a�B"O�M:'E�i���ؕ�� ��"O�0!� mΌ($ �о�`�"O�k�"�9j�j�u	� K�P���"O���=eQ���&���h���"Od�C����ys�͗`�N��f"O����*�BO��9�3"O��K%�p\��K��\���"O�M�&愊? < QK[�#��i�"O�HR��pfv��J�<9s$Ha�"O0�3�ʐ��4̠�(D$]��"O8���o�:+u���#��BP�C�"O<�ɧ�
0��䐲e�� ��p�"OhT�c*:!о��#^% �쓃"O�@��\1)I�ȪvbZj�y�F"O�I GdN#MJ�8+g��}R���"O4u��ce���#G��|ȷ"OT��	B7x�����n�6̨݅4�!�d֩*_����/L�80� �.�!�d��"�.�)�!�"-�┲�1!򄅶T��%�C�ƄҚ���(&!�$�>5j�D��K�F�8�q��C��!��~���z�غ3��1'��"L!�$��]���7I[6W��p���RD!�X�"lz�qD���������8!�$ҋQخ�˴cB�B48�P��YZ!��߆O�&��c�M2}�5yկE;Z�!�dF�F�`�w�ҤrdD�1�E8tJ!�D��I؄�����;ZX�Pv���qG!�Ę�z��rE��;W�1��I��|-!��F�����ΗM:�0���S�!� �GؖmYcN� |=��� ƀ�!��d�&�i@���Q&�4{�瓕d�!�$ۄ^���Da!�.�n���"Op�ʖ�ݭ~��+f�A-P��<�w"O����N-�9J�d�g�93w"O��"�菙 �(P��"�ݘ"O�� 4�H���P��C�eex��"O�%bAO��	 � �n42\�E"O���'k�� q�^�>��`�"O�mc����� ��ȸ'w��"Op@�Ũ�/jր�1'�A ��Ě@"O� [W�*>u�"Ύ���*"O9�5��N|P}�u*E�
h����"OR���]�ol%�7�L.UCv"O�JuG�@����CHJ�#���"O98�!�$�^� H��g�}sG"O*tZ�m�&��[GɃ����a"O�)!�hR1?��8FC΀Aր�j�"O���Ŝ.'ZI�-W�J�J��"O
���A
�H�v �Ԇ��g&5�#"O�\��^�)׊�q�z��4Z"O���@Z�➠��CŤ0�6u��"O�` �@�%%;^�[��M�>D��sv"O�aP��)#;�i�a��(%0h#Q"O��Q@G�s��24eC;`7<-Jw"O�{�iV�/����X�W2�`�"O�X�E�ՍC��)���U"a'"Oص�@�E�B�v�A�ϛ�Q���"O��(��Q�t�3�G&.\�"O~jq;3,I��LR�'2��e"O.谳Oɢ*�T2��Sj��r�"O�u��"	uR��ʢ1���XA"O�`S�ͤ��Z��˨,�L�d"O�1���u�@�%M�+.3�r"Oơ�U(�77xc,Q�x�'"O��(���j�QL�X���"O�d(�`��^B.��a�3`ȴ�d"Oph�#ș	�58��7���V"O"���@�p*䰒���ڔ�%"O�Ԙ1��	o�
䩟�K�@<�3"O4�� R&f���B��L�ֱC�"O��@��@:�&���!�`�ib"O��9Q�̲f�x{�)D^�X9��"O ���B�1=8m��a�j߆�#7"O���$ۥ@#�;�Đk78��"O��!��b�16/϶k)`)xC"O �C���@� ����n1#"O���p	81:�[@�d��9��"ORM	A.@���P�V�1�n �"O(A��5 *���Ĉ)B�J���"O��x��
�v���8W���H�ZA"O��C�i�h�M�H0$"�"O:u�@��%�4qD.;��C�"Ov$b2,	���$2�*.�Ba�e"O��c"תyr�8���'�V��&"O��1� }z��&%]�"O�Ha�_��D�:bo��MK���&"OҼ24�\�O��\�!���m���"A"O��R%(Tw�e�S��w���"O�@��@�9^��T�����ő�"O�k��Ś>c��&]�k���J�"O��e�e��	�+W�C�2�SS"O���TO�xcZI��)B�����"O�5��'�/n��J�9>��=W"O���f�Fp#�T9����l}p���"O��å
R�s�¥�B]�2��$"OV]���@4�(��g��L��ْ�"Ol�C�(:Z:黳o>|����"O:-��
�n��}Г�
C��%9�"O�x�%N�
x��̚� Q).z��p"O�Ir
�dt20*w��6}Ѡ!"O�����3�h�з��1Z��"O@I ��vAfLs�T!�y�"O��[�茱��B��9[�ԡ�"OԀ ���l��(��_Ixxh�"O� �,'�^�=��MC'�:h�a"O���B�=!%T�P%�3s͔	"O4r�$qk����D�8�,8P�"O< ��8��X�'a��m��\z2"O�H�d��[�<I �@W�n�\�i "O$	�6&�"�\���o�h��Q"O��PR! "|�ɻ�-���"O��2
G�R�LT;�+Ȩl��E��"O��h��K�N�n��K�m�.a�"O���TK,]
�ʊN�>m��"O.� �"B2�e";� M{g"O�2%�+�e��Z�b��Q"O�ܺ%��0�ތ)%DҊnCLR�"Op����&ȼ��ă5l�4���	i�O\*�K��6��d�Q��0��MH�')��j�c�3��as�	��PL�9��'��p���� �֙��V* �����j�+R)�r��m�$-��JzY�ȓ5�Y��l�8&� V��n섇�d�\S�H�z_Ν��j�qu�u��c�4��! ��NT��Wf�"ar0'�����;E���qeOD/$L�4`W�
9D�vC�	e�Џ��\x ׶y0N���r����Xݜ(��0@���}7F��$ePd�'���Sj�l(�
r˸H�`�J8o�FC�I37z�1��^I���AΣ]�8C�I>P�Nк"���}�vc�o�C�I�jA�E�bN�f��D#U�˓�?Y	�����3��P�����.9�(Y�ȓl���3�.�@���mK�8N���,O���ĄV�Vp��n� zM6�E{�O"Qѯ�:]���qOё>�|��
�'�%����$/)�x�����	�)�	�'e�a�@GX0+�H��o��Yp$�
�'_�p�� �YPzDB� ʤz�=�
�'�;FL\�Z��p(�>y�
m)
�'��p�!����h4Hp
F`�&Ű	�'��Rsτ��T�8�)Z��и�'���ۤ�٭G����"-X,a�,��'m6�;�o�$gV�{�j�.t,����'�VuH7��e���b@��m��)�'����疗{0��ɾaj�x�
�'O�x��N^��4Z�(-�X�	�'��<���Ⱥ1͞X�i�B�9�'Uh`�&Yp�E��������'e�A���O@@����?ql�)�'�V�h7yST�g� �^a��'��̚�"2�U�f�E�'�����'�	���2��)���4-��Q�'����>S楩��S*4��'���xa�ƝR�ș	�ރ(T��a�'����� �XȐd�������'�ʤ2e퐣z�t��g�##N0 ��"O�U��D^n)�S��PM�\r�"O�8Â��;p��E�Fjk�"O�����^>�ZX	�E�h8����'%��'֕i�h�*�����G��ʌ��)����/LH���/L.e����)���y��R�0� �eΝ-L�H�F��'�y�L�ph�R�M&#�0Iم�M �y���'c�����6Ns�-��BJ�y"��u�pZ�F��C��0�B��y�+"���C0c�>Co��9$H���?���hOQ>I"�o�qنo�[��h�7�!��0|� V=��>F�0�����&R�L���D.�S��0X}��݄)��r����!��7�h͚���1�$��1�!�;�-��)�}����f����!�dق$b�*�˚?�����T$+�!�Ik��%��"Yv���X >��|��(���Ag%�,��[���/j��-�$��R�O4�`�N�&k�� �L��PZ�jN>������f`NȢ7@O0X���i��!�d��k
jyA�a�<!�Ԑ����7Y�!�؎D���u��j�z ꓈UW!�ě�G��e��I��-+��(�[/A�!�D�('�j�r�@S�5b}�!�ټb����5�g?�uz�K��=����G�^���hO�o�\]�cεf�F�B�+շ����/v����/Մz1ah��ԍ��e��h��3�U��Y98#�L��4 ���m+�!C"��:�x���^n(����(A����"LAa'ִ���P~򋙴c���C����
�� ������&��O���ac�&5�6(:�+�!~��R�|B�)�S��l*�FаȈ!��7}��B�I��٘�� +TɚX�""K,��C�	 $�n���rR�xI5e�)U3�H�
�'���񔄂�4��p��FQ��(x
�'�0Ч�^�6,�XP�o������'Z�����޷"��$36j��"�
�B�'��9PE�
Ō,ƍ�'"b ��'�dEI7��U����	�W��x�'W ړf��,�Ҡ"U�3:��Tx
�'�h*C ��/������0�LU
�'�-�Teϲ)�}s�`�8?�LA	�'����,�0.��Q���[� ��L;���+�p�h� �+�8 5���HE�6"O��ҧ�<S"@
A�;aH:���"O��p�� ��yd��C���`"O5�6��yh4��!�.b]+"O�|���M1c�	A �=K4U{�"Oz��׀ʛT�<��E10���"O>Ei,�/M4Naaf_)0"��j��'M�	Vy��Ӿxs�
��H��Q�0ˍ6�!�$ך�.!d���]�:L���� q!򄊯�$�*4N޳y��͢'茭$�'�ў�>�b�$H�3(��zh6D�����U�M$LP�N��d�@G4D���.Z��\ɉ���D�(#-'D�<S�.^?
�hq4� 4� i#|O�b�Xc�N+I^@�Q��M~��ɐ�3D���T@U�ʵA�ܻ#"����0D���U*��kp��0"�O��H+.D�T��)�+ÀM1DaM�ZD�Ф8D��A2'D~��*C��]W*��$`:D��j�Oӆ�<aඏ	*sb<�0,%D�@'��I��|��c՛Ng
@�#D������ ��;Db�"V����"&D��RU�\ւ���T�e<�R(.D�p� F0%6nU{��љK>��b��O�=E�cB?�4�''��6��([F�!�;%`,�!���'
j��Ǘ�r�!�$}HH��������t��a!�d.&����8�����Ы�!��Y�C<ؑ&�p��T��&G�i@�O:���#uG�=X@��<q�x�����3
��՚��� !��Aqx��Q���d+�S�π �ItlI�.�0h9��80*��Y"O����I�h*�A�"��%r)���7"O�M���1)xּ�f /z�0P"�"O�Ed��U�b���
+w��e�"O���fDn���3��M�B�{$"O@}��,�9	��Q0�G ^��|s�ONA��nT�	_fJ0$���	�0m4D�0��He`08�D�X�I(�)	6c2D���!�K��<J1jU5�P��/D�`pի��Q�(�aԸn�Ȣ�-D�̘�(X$U�Q3�%/&���I*D��ђ��;'�VU�E�8#4�ۃM"D�`��k���p %�k<���'i!�O��䃁D��*�p0�j�◵HB��5pr�M;eN
�G2�|��C� '2B�	7f�����b��*�>^S�C�ɦP��ӨܶsV�iU�O�w��C䉾4R�X��Ү ��iT�6Y�B�ɥa*K�[b�U�#DЬB^JeyV"O�42��� ��0Zcʄ#����"O��H"L\�"	��B�$��q�"O��9�
��m���QD���; d�!�"O�$�7��S���b�ذ��"Oݛ�!�b/��2v!��x�Z"O��S�*ܙ?R4��^����P"O�a��CT7��EM$�8i�V"O�4 �śq�F��W.�$V��h"O����^8`&�A���)－�W"O@�+�˄���٣�ʍ�8��'��9P���8(�f}�I2Xj����'�)3�_�Wؐ9�S�@cRq�')v�B0���IQ����!�(UʴJ�'�!ڱ��>jܐ��Y�!74�0
�'�n�f�B<x[��1�X�
�'�"�+�ȅ*A�� ��Ĵ@�X`�' N��@nS�Z���A$ŬJ�5!�'P(�1�C�a��d8�$P�P�T���'֪�� 1e�ՀU��-Ml�`�
�'�Qq̀eI��ۑ׻O�n�
�'s5Hՠ��@�M�PG��|:H�X�'��!���܀M<
	Y@K8t�����'����B�ec,�!�@�Yf�4��'����n��u�d�h��$#���'̮�u/Z�]��݉�fډ+n��{�'z1``��]Y�y���-�����'␽A�^-D�$�рI�L�襁�'?&X��GM�\KTt�ԁ�{����
�'��� A
4���#�V�l� `
�'��y*d�ƽ��S�n�yts	�'@���N����h�%��o�L���'�0Yx� �gs��qp
��7����'�H���dO$�.�2Aǈ�2D�J�'pv�S�F� 1����>���'���1��n�^z�O��7�T��'��y��\�VH*�1`.½x����'t�	�nS�G��U�$�r����'�&��G/8�mb�.R^Z`[�'�jgi� Q6*0#�
A��UB�'<$����նe��� D1)Ɯ �'������I� �"M�4-d��'jV�a�!�H��p����1*(�
�'����`���|}�s��2\8@j
�'H��5-F:%E���3Ōz�L��	�'Wn���j�x�5����zY�Q���� ��7�C�_�� ��,+�TMk"O,)j�.�$0jZm�VnBm�� �t"O�u�c��17`BA��i�eP6�'�1Ocd��	*�(�,D6O���"On��5��u�n�S�E��U[�"O~���-\;\���6%��ym�E§�|��)� ����uj '�<!s��o[|B��'0f�H�'�M�g�:9�AgβXZ8B�	S�j́ �ƞn���B���**B�	?9�(̘Cꇨ+��� 2��4b��C�`�l�A��� G=��]�Q4�C�I'�n� ��.N���yg�[�D�XB�%E��Х��I���J� Z�V,T�O��=�}�1'�ltH�1�=OJ��D�C�<1�᝙%V�ţ�ȁ�q�*e���G�<I��K�]Y��s0bƅ)�01��O�n�<9��G(EW&�����A~�qK��_�<)�Ꙟ\7 ��gET�N�(�«�t�<1� �{�|��!�#o)Pd�%%s�<Q�BH�%
�3�,�h����fyb�)ʧ+����eK٠zH�hY�Jˠ+ap|�ȓB�(����� ���~� m�ȓG�p��F�:> [�n�2U��(�ȓ����&`ťlm�@: e@�6�M�ȓ���1�I� {�ZK&������(�rΟ9w�^���hQ��܆�\�~ԠUJQ�^Gz�Վ�.'"P��{���{�b��iC4��'���@U��Y(�ԃ�Ӽz��,�S�ǊA���ȓ=�$)�ȿ��T㴀O��h܄ȓD��蔋�JV��2�@O���x��e+X���n��k��)"�%HD��g������%e�|@hƂU�#z����}<���N8�A�
� ���	��t�<)!���Zl��jS��j=2�o	j�<Y����&�ع8���/��H�b�f�<����~��d{V���?�~��0��}�<)�V22�5��o 62�x��M�R�<)ǓY���,�_"���K�<iͅ�X���L����e�fFğE{����2|������D6e�X�0��BB�	!h����I%n��
��ͅ%8B�	."<���H��Jl�a���k|�C�ɾ|r����%�� �T��&D��K\�C�	�T
�00��g�PL�� �w�B�	�:�l�
�.ķ�K���;�����,�x�R����ԞL�t[׍�'t+���y����X�x�� �3�H�@0����t��*(D��	�&^�> 8���
&�|8V<D��IM�E`Phڃ��ɥ�9D����IV�D���$�׀�v��& *D���S�֠
B)y&EX9%�&$��'D��
W�ˢ'ɚ5�W�U5U`�6'#D���\
�Jݡ�H�,e1�䰧�=D���� ��<��	Q�4��I�GG(D�8�w�[�$"HT�bA�-�V�Ȥ�%D�$��O��� K��W3l����6D����*��2sq��Рmi23�&D��F��-��<���� ��-87�$D�PH��¹�F����FX����#$D�\X��V�>�ɰ�3�M���-D�8�l�)7Ā�XG�
�;v��BD'(D�Xa���
�T�Ul�q�`�I�&D�x���fJ:��e�C�0,x�:Pf#D�� ��u��+t5� ���%���8�"O�U�C�U 4�|�A4��:yDT�w"OD��̌�SU�{᧞)/c��b��'(1OJdA3E��z>j�# �!pJ̤JP�|��'\�����@���
���"���'��M��h�(p���&�+�����'�<l� *C5e� ��.�2T�����'��x�A�NȾ�ʄd��di�
�'ޕb��=Lc����� $wR�	
�'880��W�� �9?/H�$"O��B��G<H�����BŕBUXT�p��!��џ��'�R��qE���}��Ȝ.r����'=��[�/[+R��y���xJZ)X�'`�1� �V�$	����l�R9�'#�Rb��2��Aу�F��'7�}�G�L1����#bCN�fY�'�� 25)�(5o�]rS�F�wX���';ĵ�'�C~(���I��n��)�(O��OV�?��'{�8�v�X$�ޅp��� 1�ֈK	��O�}���P:�`8�ZZX��`"O���sǗ:kr�])bb�0dy��"O
�@��Վ=��졡O��]G�|��"O��А. �7،�醏�\,L��"O���#�H�8'�Z5���wL�@E"O4Qؗ�J�j�
����n�H4���'�ў"|r�'���S�g�W��1����>IF����O�}�E`�
%;�$��	Z�l}�(*c"O(���_BŌ
�iЉr P�"O\8�dR�F��Xq`	�(9.<q"O�������5��-%KC|�"O� ;3E
�5�@��ˣh�����|��)�S�'��D8 �X�}�	� �P ���I'�T5 I�%�����eG-�\���	^̓n8��!���W"�!7��=m��l�ȓH�	�3�Z9�9�C��\��݅ȓ	�6	sh��*�LP*�V�0��d��q���S�|Bd:���9:��ȓ=:���G�ɍD�>$�t�J�0R�F���8�j�&a�e.�����Q�g��㟈�Ig�'���_3 �R��P)D�|X�B��&f������I`���'�p����w�lT�S�-<�D��'b9Q�� �g�j���K.t�	�'�tap�=$x�򭈒q@*��'�B����N�H��!�M	�@0�Z
�'�x�Q�L (����F���x����
�'l"�TgI�f]���eo�8^���C�b�'�:��@�O�譱�IφWqdp)O�O��}�A�����L�4����'[)�"Յȓ	�X����~�\�x��-`�"�� �q׆����(p7$'Tf�ȓ(�6��e����ĳ"���ۓ@ D�t"Ĥ�������D�R��d�� D��:\�12���Y>��g�?L\!�dȓ`�2E*d�c%�|��	ay"�'��O��?��{�
Y���7�:$X(��(\~9�B�i�� 7!�<U/Pa��3����B�N�N:�����N�H\�e�ȓi�N�#�
@�s�N>~Q0��ȓt"��Q���)������O��2���`N�c�#�T�{�@�9�v���y����IH�)>��#�JlJ�'���>\JB�S��|�`�BuI�/H�C�Ʌ$�)����T��Jv��{��y��v�z�"T�g4�"��V�Y]�y��S�? "�#��9j��(�a���]:06�'����D*��;�Z�Q�L�!oDp�e2D��a3��!S$�p7S(.|؉��0D��s��4�D��b�7/�F8�-D��p�j��D��BCJ�)�
@#��'��hO�	�a6����Dgs��J���4r��5�|��I�v���h�81hܼHj1D�t�t�ן�и��a 2f�Yw�/D�,03���c~�yZ2"K�z��P(��)��0<%��9ykN��ҍ-���@{�<��@P'�`�TKO�Bm�!��Py��'�O�#<�D[.A
��'��J=pLx��R�<Y�8X�p)W�ïm��#M�<�$�݈@���M��m���� Cn�<i%F��\���+_+>9[f�V^���hO�Wf�dP�J+l0 �Q�A�6۰M�ȓd(q�0�٥$�-�u�B�P��!�ȓ b@Q�#8ߖp2�
�HJf���ٟ��?E�D`�9y}`hs��j%��1R&K�|�Ig��x#Q�*-��˦�p��h��7D�,�fK�Z5��!��	ʆ��І9D��K�
�	�ԋ�����y��4D�(�2�B�?/�����NF׆0i�'3D��9Gh�����KZE,�Y7I6D�����.�x$����W�2k.D��8@�9xY���T)�`��Mh���O���S��}� ӊ\\*�K�:mr�B�T�<!�։;Tlp��7��R�R�<��D�A�V�����;G<e�a%Vf�<)Oۉ,�T1��1F�\"�_�<�� ?����"[*a�����q�<!��P�q�|uP$C�(Y�`�w��x�?!���Oݑ��kNC�ӒP=r��t"Oh���Z$%��@#�P�bV!F$!�Y�4�Ƚ�pܔ$��r�C�Q!�D�2@r@����N%쮥2��G!��"�4���Z�
M��L�pb!�W�=g<8���S�#��1KY;LN!�TsWk	�<<���۞/K�}r�'��� J.ҹ��G����a����&��)�'��H  @�i�� ��iS/l���p�'�VՁS��!LW|��7�EZl4��
�'���*!S�ց�D�?��%��'X>�kw��4G�b8:��̤DAf���'����@$�l%���$G4�ѻ�'麔���"
�Ͳ3�A}Zl�I�'����@a	��C��',0������d-�O����!o��)&
�\i�"Od=�UnL�E~��r��FU���"O���׃	 �M�ӆB�m����"O*�3f�Y+�zИ�ԗ2�pA	u"OD;ec:��u�
A�CXd�A"O(��%oѭ���Q "U^j�!�$˥,�*hi�'n�9��ҪOD!�D0܀A���S���Bf✝g4!�$��p���`b�@�y��`p�aA�|!�$I��h<#�$��8��D#A?4�!�D۽u/�U��H��]:�L&�2u�!�dʍ-Lqe�U�pw��2uϐ���'+a|b&�%��1� G����cf���y��P����큠.� ���O5�y"��4�h��b�����0.�yr��a�$�J .�{� ������y�Y4����G۷?��U`r�ȴ�y
� Rs`�:��ڀ��?{�T� t"O�Y ��-�(�QǧV�T�fW�X%���ቮj� t���@��M27�XDrB�	0*2��#CFB�pf�-CgD;lt�C�-���Ċe�z�r��C�I�%��c��\Q:f�k��B�,ל���b�#g]ty�T�U�"��B��%7Pd)��Y -�l�6BB�B�4 _���7fM�9V���T�m4~��!��=���y�l	m���J�
,�Ĺ֧��y�M�&p|0��!�N��`�6bT��y���o�F�铠I�%�X��sB���yb#H�%a0��!�Z����s�i��y��N-*�#LWZ�3F�.&�vE��'�.�C���.^�m�Sa�% ����'�e��H��e!Ҽx�M\�S0����?y�'�ҍ0��!
jd��Ɵ�I%����'⌅�v�X�I��,�u�RA�<*�'�.�Z	T�K]'<�d��z�<i���}ݮ@�*�0)d����Ys�<��$E)3���ITÚ+�\lF�c�<I��h?d��7	�q���&O`��C���Iw�J���Cc��zi
cc0�t�)�O��	8B���G�I�~�PS�й}��B�I t�b�`O�t�`��d���tB��;'�!)��M�U{B	G)֘C�	�-
� ���#���yB!�1��B䉢 ��uAQ�ĳG�hC4L��}��C�;m*<����0d�$������C�	�EI0D��Q�M>�C���:�C�I�M�x�=�$����p��B�Ƀx�������$ש�:p��C�Ʉ0����ѪM�`�� �&��r��C�	�v�Zȡ$a��1���7!�3Q�pB�I��=���&of11��� LҤB䉨%U��� �k��r��fZ�B䉣p�t���o�8yt)yu��O�\C�I�9p��Т���Acg��C�	�`Q�!���\.Uc�D�Z��B��.78P{a$p�ܪw�ФO�C�I�_���YB�' ��kƀ�TR�B�	UO���0�CY�.ț���H.�C�	4f�
����͂N*t�����_BC�I3~��Hcu
Cd6�9���64 @C䉑|Eȣ�˻X{�� �Λ@|B�		��@�"߲k��P�
L�vH�B�	p�����N(G��\��B�	�` .��DM��T�c��7hVB�ɛN�Y��U�(gJ�)C� �B�Ʉv��\1F�?g�tk��m��C�	�ej1�#��1;�Q�5�^�[q�C�+�>�s���
�Ԍ�$�'YcfC�I��X8�uA��܄�q�C (8C�� � ��$QT�m��D�z��B�I�ʀГP��JM�� 6iO;|2B䉡v����'�X�J�Q�̓�B�ɦ���ҡo�0(�iU
��B�	@�p��d�D	 �Q�4�bl�B���:��"�_�,l�q���8^��B��%��t��A�9y1�-*5m��i�^B�I�f����!���'��4B�I�M���SbP�B0��SVl� B^C䉺Av���XH�^H�C���B�	:S�Z�ŮA�,�7��=�|B�)� �L�7!��z��{�#/j���"ODX�o�7N@�H�#NE}���O��r �J]4��� R��BЁ�];!�\�&���S"�H/tZ��q� ��z1!��$1����
U<@X�jj�55.!�^#t d"3�)��o�~!�d��Q��ň�Ε��^!� k]�?�!�$���:�����L��8���y�!򤉛�4��!ٱ0��R���qsa~�-
�?aU�ݏu��0�$�f~����=�y"�L�r�C��!8I��s�K��yB�T�S����G��/�R\&�y�D� J��Y�6�G�)�x�i��F&�y�/A%P���#�B��h[s��'�y2Iͳ&��\(��־-��/
&�y���*�ڭ�X<��x�@h̐�0<y"�
ҟP$�|��#��w�E����=[�t P##V�<��^�|E����N 	�8i˷��N�<�nR6:�j�؆�	�9��(��C�<u+�?�|8��a�1D�p@H�}�<��HTkZ���E����\}�<	��n޽)�n)b����Vz�<��Y1^z�0P!�[&9��[1��x�<��K(f��x!��8+�ec���_�<y��V!��� ��	���rRl�]�<�V�U|~� /@�:,�j�A�A�<����'��y���e�1:�a�z�<A�G�2c������4BC0h@!�AR�<i�
����Ө�B�<���Di�<YÍD�
in-�	J�<Q��ƪf�<tbC&�d5�U G����M�}�<�P��O_b�C↜�Q���Q[S�<�� �"78d(�ڙP��H"`��R�<�A��2�\�'�À"2�ŀG�Q�<0����u�2����
�����N�<���/MAVQ@���@e��a/I�<�D6hd�I��{�2U�o�N�<yag��(Kz ��nY+䙴��A�<u�Ӡk,~��� 0k89C��z�<1.�d3�	:D
P�il�����p�<Tf ]�Q�rk�X��x�<Q�%C�*����3*�/���) Mu�<�@��T�s��W�tp�2�Yh�<q�B ��x�s�fЯ:ʎ,��o�o�<�2�]-@��u���@�H�~��k�e�<!D���ʅĂ/�� ;q�R�aD p�ȓ�X�)2�x�B���G���D��?��	j�ǔ���R���qN �ȓ� �:����\H� ��>��ȓ,�����&k���%�̭[P��� ��l�Va�qA�<;�	ȟD8,�ȓgb�h�$)�<[�S�F�T!��n0���`!	�e��5;���
Rj�Y��"dHԻB�!��`ju'L�++���6"~�9u�n�ʢ��y����D�9�wL�mxV��"�z�%��_��Y��%~����C�[ %�80��{��y�gR�,.���Ȓ4F�b���kЕ�⌘x,����(����y� ��5ij\i����-:�=�ȓ|���[t��̼\��������,>�8suC´x��4�C�R4Hrp���:ġ'GCWl�bbh�$	�8��T�4��"E�1�`N+r�����S�? *���O��Tm �&�0���
�"Of�[� %A�T�X���W~�]�"O^xPw���U��e!ƃM;;�d��"O�s�(�pXuB�oў9܄=�"O���I	D|i�u�d� X��"O����/ujȣm��T���04"O�x�%^-N(�4S��<� �p"O�,JP.Y�1��h���\$j�(&"O�0��薍i��IS)�&M�Ըg"O0���BEHk���A�k�<e"O|� ���.U�ؒ&)E(HD}x!"O2QX�5]��|P ]�3�V]��"O.A�	�
|;!fK
Œ��g"OV����Hk��wE�/Q��"O���k˃Bɨ��q�Xcp��"O:H�dI��艺N[#<R���"O,�@Ѯ�L/��MTJB^	�"O��8�IE V>�K��U�Z@���1"O���qJnB"e�P+P,H��"O�!�y���)�� �}��$Xp�!D�x"3���7I�]J�چB��D�%2D�D�&@	;h�p��ʙ ����E0D�������a��G6xC��S@�-D� �.
p8"0E�@ߌ��m*D��FB�50��|A�	sؒq9�`=D�·�ų[�`�gkQ�?�^a�B >D��Qb
�9#g
ѧ�.�-B�=D��5 �!͖�p�*K�E .� �:D��A�G�<� �v�ތJ�d4`��:D�B�h�(��u)�7Njd�Re�9D��gC�� �|�XFK���R��sB,D��)d-�	(��3O�;5E��T/5D�P"��ɺ�	�A�-V�ģs�.D�[���N��L#jۦ �
P��7D�kq	\>(�B'JY50����K2D�|{��ν�&��/�]�I¥�.D�<��"�D�R|s��,EB�Ƈ*D� �p\�*�z�GW6PI
���%D� �@�T.y�E�'��7պ��#D��S����O��C@����N�q�H"D�l��F��>��E��42RD+�?D��y��%f	B���؄3,8�!<D��5�e 혔�S�*_�P��/D�|���K0.2X�Q�o��@�V�*D�$Y�n�2��� �<TRG)#D��A�HV$�Z��v
hx���!J!D����,��]9�-�����!,D�`�@mJ;d�b䉗��	D��E���)D��:��\���x#�9���i�%D��k�Ã8L��W�&]����@O"D��!DF����2FO������;D��"G�J<���q4�))O��c7D�`����� Kɂ�K���(�E�5D���P��i��� ���-a��`kw'2D�<2�#��b$�R�-�v��	,D� *��7�����i�V��g�(D��xDd�6�f�
1Iݲu�T�P��$D�L�d��N�q{���a�~-9Aa!D��RхA7A�Mq�Æ9�h�B�=D���!�Ĝ`�b��Ʉ�8�R�=D�a4����25 ԱN�\��l%D�f�\�b� ��TW'b!��>D�˳b�'g9��W�Q�rx�bN?D���N�3��<��@�F�4�'(>D�� *�K�>*(��k���E�6�&"O��c3�҆aKR�{�\	(��`"O�dq�oʴ\�
���1uu���!"Oޜ�0���
x>�;��tb�m��"O���qgA� K��o�\4��"O�=��-�lJܢf��&Z�)H�"O,}Ƈ �X �ɐ�02�"O�]��dS�A���*E��-y��ԋ�"OZ�B�A�9 |2��e�VK�
�PV"O��{�&�)tw��$C� �@��`"O��P����Px0D˥�!����g"OL��W�H�!�@(�AL�s�tq�"O�!��K�`L�@ݹ_�h� "O�L���~m��x�l�dcN��P"O��щ�o���@�	�M��H��"O��B���.BŚ���J��
h�a"O؄�$��2*�.i(�	Lj\��ц"O~�{cȃ3z�,"w��'G�`#�"OT
�O��e��3��y/��bR"Ot؈�Q��E: �[�Q1pQ+�"On���/�
8KX�@�4@ؽɤ"O��@T�*D��(d�\�B0�`(�"O~�D8]�l��ԩ�R	�u�"O��ZqnT4t�Fi�ǩ�j��d
%"O��p�%I��^̚'��#v�8 T"O&� ��vw�0�� T� �`�"OyP0��T``@ɯ,�v 0�"O�qS�"�^�4��s.D�m��P"Oy���k�<���L)�0��f"Ob�"���C�z���MV�k�Ɖ1�"O	*�]~u`ɣ%M�;ͦ���"O�\2�)d�P��[��Bu!�"O0�S���#Y����j��Vb쳶"O�	07�^�R0Hp�7��. (Vr�"On �VnH.���;�OT�3#�-9�"O.h �A &�mїn�|��""ON���a�:i<;f�RP B�"O��SV�$2��D�Ŧ�#����"O�8�K�DP��Qr��d�5"O�9�"�Y l6��@��R|�kR"O����T�Q���3bO1"=K6"O��k�IJ'�x��':�(��"O��AҤRǤ��`�.I�2��"O��ҕ�Q,�:�,���"Ol�
@ᐼ�Wh�v�B�"O���W�GY���鋥p|Ը�"Old��� �@�b�Y���#R؈���"O@}9��P�B,�K&���X�9��"O��y ��6�(m�@���|�ࡳ�"OB��A�(,��d��[��Šb"O��h@(*vbpuY��:pv��9g"O��yя߷Qv��J�5D�X1"O�=xuo�
i� ��-qjq�"OT	��cx0��=9�Ġ�7"OtU��IQg6@낁��m}�Ӆ"O2i"4)݋��J͸����.D���sᑳO��,kQ�Ƒn�b`��)+D�|��f�d��r ���`p|	�qi&D�X2���q0��*e��.x��i(D�L0�k�&ZeA'%}�$�2D��Ig�$s{
���\ ch�	x�0D��1r���=%.h��V���+F�/D�X��+7v�TcB�ҝ)䍳��,D�k��� u$)��ϔv�A���-D�� �ѡ�і�x��2G�)`�tDy�"O\첵��N�x8������r�"O�I��bAZ8�P��'(t1��"O.y�%,��7���
���,��i!u"O�2�G�6t�ɪ-���k�"Oҽ�Bۈ7��M5C=Q��q�Q"O�҃/N!Ocv���X
/��s"O�5!5C�M�<X�a(�v�ے"O0-j��M���*�C�Rpa��"O���a�)�j Jϗ�Q
�r"OV-b%�V�E�$m�1�X��"O�5B���H���a�l��y����"O�``��ϬtTlJL�7� ��"O>h��E��7�A�:����2"Oƴ����-*��RB!}�%)�"OT�PErě��R#z@lh�"O�e��
5�>���eM�:O��x#"O�D�%���5��5� A���b�"O�r`*�����:u��p��"O`Q6lF�Y�f�I%�I�/�I("O�t
a�#;�6�<��r�a���yraN-���Tf]��lJ����y"�ٳ9�"��#/����R� ���y���G��Ƥ @dm*�����yRJ�3�,�x�"Xy�}	��yB+��u\$ȶ�����5�й�y����^=�LP�-E�����B���yr�7#�b|3PNV�N� �*���y"�i��hJ��9P��"'��y���0��HC�-٠K�Lܚ��H��y(��;xBuRp�>p������H��y��4�����J��*�y��
�ydQ�&����KD=�.��h���y"
B�"�Y�1	U�1m"�)�j��y5��7K���ٺ�%��y2&ɔ~��-�U�N W�ē�eL��ybm�������q�4�H��yb��9��)9��
��J$����yB�̻G?>FE�Ld�b��ɢ�y"�ˍx��ˢ��E����jN#�yB�O�݄X�/8U���4`��y��\�Z�	�fN�?���ȧ-��y�+�X�NШs�R(2x(DS0!��yB(6�,uxī��,l�B�e��y"�ǭjZ�|��a�8Q��������y�a!PL��	�I<�9c&L&�y"��[���q�[!,��JW.)�y��/����㌈;R��I4a��y$�5c���Y7bٹF�A�'��yrh�5�f�����;!h�*�g�y"�ǘM�J8��œ4/�)4`��yr��&I���ibDɷ&�4��Ƚ�yb ބ{1re�̎$�.�B�-��y4�L]¥O�(FP+ �3�y�aQ�Hl�\#�k�5��r�!��yrmW"#'pEb�H׸31L��#�y�-�30�4�jf%P�u/�=H��)�y�mܝ~�Z���
l��h��W��0?�-O�I�v"W�	�`)"���[�H<ST�`��������D,6&.�`2��~lB��`�pyWfER��D��i�
�Jb�\��ɣhY�aB�	�X��8;D�Ph">Y��i�>?栁�#��IJ�����T)!��H,��� ��L�����KO<��7�S�π � ��f��2� �*%�lZpO��v�V�G�
h�bZ�:j�}Z�GnyB�)�',���a�c��=�!�2��|Ɇ�II~B»$���3�F�n�|b���yR(�~�Ĵ��InU�P��+���y��=<��EAǡ�+m�؀ C?�y�^�z�$����a)��1�	�,�?ً��S�Y�ژ@�m�\%$Wp�����f/)ck�$RX�@���C�504`&�O�㞼D~���%-4ЅA�lɒ?�0�W��D��䓎��|%a��I� |z��[B<��*OJ�.T��!A��V=����j����D �S�Of���7�9~�8))�h�$����'U8ٲD��(Uށ�f�:~}X�������9�)�'K�*8���[qD�lV7H86��'+�x�U�S�=�f�z%��2B<Tq/O(��䉵b��@��%�$Y�*l#B�C�1O��=�O�rj]�Ns�t1�[',v)0a��y�˥v�2�zF��9NbL�+�8�0<9��d��D�@�3�c?�i6`��2V!���6S�d� F��46'��`�<�r�)�'k�~�pP��	��ܪ�ā3qL
�s	�'LJ�c�`��AC��bd�^>|�P���'E�\���8Um&8k3���+ X �'�^xa��N�TK��R�6��%��'΍���Քv���µ�K�j*� �'_���F-3||�c�F�(<��'������-&��Q(ǁU%;�>����'�!ۆ�9'X%�6
�:C
���'F������R	���6%<N�l�	�'�@���KQ��{̔�9�x��';n����?Q��UN>�z1��'ʦ,�&�>fO �a�gI�j���K�'�E��dU�[�5x0A��b�U	�'���1�&9A��Ф�9V�[Z�'�|Q��T�U�'���^�6y2	�'�g�Zd�v|���ݬF<@a�	�'*�!��*
��8t�Ա8+n��
�'$���[0`����*3<��p
�'�:=ʤ�)n�d��Q"wL�aK<9�]��Z�lݢq�<��5��4�� �ȓP |�8�B�-<8�%c�8]�T��'0a~��%�n���<qef��g��>��>Q���y�Z�z��bKчk{�0[��O�����O$$
דm^A�S�Z�p��D+����h�tD��I?H�6���'B18�Έ4�~X��'�Yפ��h��I���-��Ī�'��rg�b��E��癮'W��a�'����l�2t���0e��b8h+'o D�L�#Ҡ �L�B��S�xV.���+�O��O���I�-{��P�v�҅P�,8F�x��'L|8y�D�XӘ���iƀ[>����~��U�,�DS�i˜`p^�!�B�;�y�F� �bM@��*U$�� H���O�v� ���;@�]�������V~�'F2�� UdD�1E�>} Bdc���ybm�XD�����vľ0R����0<	���'�~5��J��sR��qMܬ5e�82	Ǔ�HO�t����'��A1�Q�?gb`I��	y.�>��d��'��ai���%����b#J@��y��L� "'�=�{�H9,�.�R��$}B�xb��	�E�q�J�/1�L�w�|8dm�n���m�3j{`eW��#c�~��r�VR
B��19`���רZ���X�S�;{����b��� lA��H6"��P�7�Q�k�|�c+<4���`NE�v����c��A�����3<Ov��}R琟BJ������O�̼Br�Ϳ�y�.ɒ1'~A�_4�8*"��èO,	qB&ҧh�j��s�!;x�p�Z�9Ҽ��q�$$lO��0f�E�\ �BP�2~H�>����	�)qZ��E�ғ��q�m�\!�$Z��8� �mX*�����M�qX!�DČ������O�:I~P:"
�J!��8j��y�|��)�A�P�Ie���fx06�
�6��
[�S��:�"O����~��傪k����#���{B�'(��%��Sgd��&�
����	��?ar�iFt�*����%{'�-D�R�'��:�"	���1�T�� 	Ǔ�HO���p��!��e��ϭK%T��"O�yꡎ���eӐ��O\�rW�>IT�)�S�~���w�,"��y�圊*d���d/ғu�>	���ˠ ��ۦ �B���ȓQRi�����1L���t��[�J!�'_�F�)��)t�Uj�7 ����f��N�JB�Ir�6�s�&A��\$��Gn��"<Q	�*XM�a� �ȁ]<~�5�ȓ5� x���d�\`WIN8��i��-�,��g��m2�KE%#�F�E}�;Ox�|d�.`��2�@�h������@�<I�fZ�H��y���v6c�@~�<�E�/UG��S�|�0�D�P�<��p�T@'n	q�HL3���N�<��@�u������X+  DH�<!g��	�2D�@MP�Ǥ�j�C�<!�'%|4�GƏ8��UJ��H�<��iA���j���'�0B�JDF�<I�Ɣ�_�ź���KW��3�Vw��hO�O����I�j�!��Ӓ*���0�'� ��5��&�d}Cf�!��u�-OO���@?վ�j� �^Ap���$�!��;� ���_bPa0�"L�t����>y�(2E��A᝝xxjpp�eqX��O�1�$e�w�2�0gW�a���"O�Q{ӌE�LR|�&ؒ
 ���"O�����O�yP%�]:��L�e"O~\��1�]���/氰jcR�8��	;�ѱ"��<�D��͚/@B䉤�����쌟n-����"�6=����M��h��P�l�#g:�9D N`�j�����V�'�󉉈b��Tr��Ҡ���M�|�!�d�<��uɄ�29�p��Sl�8ǆU�ӫZZ�S��?��b�.��T˅�^�ln(! ���l�<A�C�`Ā�(�w�R	��c}E�,��D,�S�d[*��cg��Ia�(X��>�#�� P3@<�.��׬A7*��;D��:#�R�LF����c�*>6�p(�D;D��R+آK�)�'�!߮<ST�8D��#���v;J�Ν�!�	p�	,D�<RN����2�H\b-����n=D��V�[�pZ�
%"�0z �Y�&.D��V�N�e�\���3m4a�.D���f�Ճ9��� ƿb�I �"*D��:���,���!D�	��ȋ��:D���M��c�ni�5.�#Zy�l�r�,D��y�kQ'|y����#!��;�*,D���ϭ}z��k�^��#$C(D��ƣ�|2�
#�P'?8�-���;D�� j����ճ)��%BE��41�A�"OH��A@\D�j0��<J�Τ�"O-#��ڞdVT�ˤ�ŕ��5��"O�]:F�\Bs���ԋ:sشh{�"O����*N5<���	��,�kD"O�(��]�i P\���Ԑ�2�"O��b4	���x���
I�6�"O@�D�E^�n��
C��"�+�"O�I�D��[y`���ǖ���1a�"O�`�WyQ�x� J��Qb�"OX���)7R�I#���/z��P"O��X�gC�	��E{1 ƈ ���ZW"OQ{@NʠWN�s�P�"{�LY�"O�����S�-T��p5-�ӈ5��"O����#�e끪:5�Xe�3"O����N�(~��&��[��(R�"Oz�bA7���ť["6��1r�"O�)�,Ӌsn̻&d���b�"Ovi*7%��{;�tI�o
�����r"O�% PF�(4Y��iۤh;��"O�D���B�:iI��(ڻ7�9��"O,��$�D��1I��
���t��"Od8J����2��2���!KZ4I�"O�Q V��4q�
���I	:XLQ�"O�\��b��p�
Lv+p���"O4���бN���d�U*�4�A�"O���%Os\$(䈍,d
h��0O\,��'�E���:V`׃=�����	M�I�jV�fi�qEɁ*�<B�	�`����P e�A���!&B�	<d��(H��߃�A�P �9Ee>C�Ɋ%�̥���4E��	���ޥ��B�g��嘶B
��ux!^��B�	�JO���!��iR��E�_pC��::w�<:�F[(A�Ċ�{,C�	�-�`5����Aft�F"
,;��C�	�;T8Z%��<P�*u@�
�bC�	גg��sv��`�V�?z$X�"OpPBt���q��5r2@��I2 �@�"O��b5o�$|��Q�@Ϫw�:P��"O�0�ፅ���aYЉ�p�"�q�"O"��*��{�@=�-�<@��4�D"O�lYT�E�e��EەW�h(�a�"O�M�c�0?�RH��� :ĭH""OFig#�R��@O�M��:�"Ob9#8B��`�/S�t��UJ�"O���ʟ�zp,%������y"�=
�X��1�I$=<�P(�'
Z@k�b�9f��s�8\e��'�*�Mt
�K��+0|��'�����ή{���5��j�j�'�x�1�мYs�8�'�K_�-��'�p�3r���B��N�A�mP�'�n�8V��.j:|��R�O-�]�'b���e�S8���h� ��K����	�'$��g��:�ph	���VѨ	�'� y�ϊ |^�X����2ZzB�'��Pq��%��B���@4T:�'��؀�\�s�\D�"���xۄ��'�`�ȶ!SRU`����$X� ��'(0��`�-,����4JˊQǂ���'���9B@
j~L#
�qR\x�
�'e�Q��%���&Ui������
�'�F,���K	p�р���t�HC	�'!0h�t���2\E�W��;c�H	���� �D�� ݞD"<8��J�dzB"O��`	J20�XI(A"�q[8���"OҌR�ȝ��A� ��0ۦ"Ont�3cX/^�Δڑ�E�a��X�"O�l ��9��-�&��-_tmJ�����#�ʚB�'���8�h
_J<�Jw�?9JR��ȓ����V�9�L�c ,��͓8dѰ�耥m3ҧ�����O�3:IX��hMR��yP1"OR)����vn�Y��������W���6���	X�B�.S_��)�
B�l��P�V&��$�7�O�4 !K��G�4p�tn�c�I!�GVm����4��N�C��^<��C�Ɨ&N]��U$R*��=a�a�|��X�QE	�ҘO
|�����D��f��YG
�
�'@H 8�KPad��%[2/�%���2�
���Ɨ�P�1�*O?��2/�N����,B��4���bg�<9��'y;r D&Ȓlv�$��by2�И%G�顳,Q@�ax"�v����/��0�8������>ѕ#�$��91���w�NpC'E���`1����8���a�'H���p��'C�D�3�#Gz�����+�4 ��)P�&�b>Ia)C.��|2��~W���$c!D���0]"0���V�P�T�1z�$�e�C��f���>E����,_=@�J�R2z,
��@,�y�H�%mK(�y�C�Oz��������ɰ"�����_MX��(p�PV����` 0�(R`%4D�h�B
�
P����}��-�0M3D�#�H#b�闢/# ���,D� *5�(e��"!�DR��j�l+D���p��$5���5#_9명�ei+D���g��1bb�p�뛭d0��v�7D�8�H\(k{`Ƞ!�V���F9D�L"�d�88�@������-�rO3D�<�R ��U��1�U�5��j�A3D�,���\->�E���hd��r�-"D��R(����B�-}{��A#D������K.���D%V��\���-D��!�C1hܨ:p.!M'�|JK*D���j�7:������̐m�Fh��@<D��PPGIl�2l1!M(]����:D���� c@��A��
��bޞ;��"&$ިvzӧ��BΘrZ~�Jp�J�S\���f���yrˍ�VZ6(�0�^K*�D������y�%���䅙��Km�y��*IMR!Sn�J1���R�R��=�4I�/�&m��IT�K�<�#�͎�N��IzA�Lupx�C��3$�h0�*7��큥��,!��v*)��4B�^���#d
��#�	�$:Ժt[����b�M�7!򤁴"*Up�J�*2Ꜥڤe�(T��"Sr�̙r�n�j?1���O0p�DOY(rZN`i� ?b@���-D����PYנ8y�ʎ�0B2�R3��OѨՍK����h���+��<�k �5�\�S񍛖v��J�$]��`A����BF��a+��h�Z�Ԧ"4�B�[mM�=_T4���Ao�$�=����'�B��2�,X�T>�v����P0�K$(T`,��~JS)}��S/T/���Q���<��G��<�J�jߓVv�a1�{ݞ�zRJSe7�4J1���&���-�&���1�	WP��4�&Q��Måύ!>!��B&��/d5j���cFB�<A�C��9�<K�H��7�q�#H���9�CN�A���R�!��>��6C��=�2��S����є)��0��/�$<����dN2X��|���R�����GR�@��K-p0�H`�Xފ�6F�=U��'��>�	><��Q�feE�b�$#qJ�
h�>��qq-߄{tXA��IO�i}���g�;k����0+��y�]���C�_����D�4ҚY��&��{+>���ELo��Q#�-�6Yiر�OT�ӳi�Ҹ[!�=?���B�շ�M�
�6g�&] ^�\0�0�b�<I� �<�N�x�׃'�����8����#-z	�ILhv�E �<ϛVDŭK6���3�D�e�2A��
K~�q�'���pdVR��oZ6��T"�.2C|�R�eL���Y��ύ�a�x�-O>`���F�j�1�1O� HT�t�$T��a�!h��6#Yr��$��H$���	F���O'$u�QhI6?!Fr0m�7y(M��bJ=��H��"���<�i��'��m^�8�r�͝{f]��i)f�~�ٵ.}2?��ٸc�"Z���S���J�������aҷ{k(8�@�(�!�[���z"I=A[ I�*QR�bܡ#���{�%A'�A0M<񧨋��'Y���y�o���@��uW���}b��1X���oء<`E2��Y�A� 1t"��^��c�()4BY����ē&�h9����d�rX�#��2�t`FxBf��NH6�b0�	B���0�ٴ86	
G�ˎh]DC�	^�B-q�&(c��᫕�P1�hT���"~�ɡ]P�s���X���k��R�`�XC�I�:?�<���P���CB�uK>C�I^;�TāW?v����g��lVB䉡p]n�{P聪i��U�Q��0��C�I�=$|��ѩ"���B�K�U-�C䉀{L8�y`B?rFD����>Z��#;g�����s�B)ӆJ����4�B�-'�)�S�p1�(4�/A�.�!�˳D��C�ɱr#��Ⲏ�6��!aRe��#$�'�$q��! �c>c��QdJ)Wܦ���Ł<H����6�Ob�31��]ZeZUMU�.8ءY�OH� v|Qx��&հ?q I cT�y����F�n�(�H�j�'I	��%JL?Z�JL�\Ĩ	��A�`,��P�H+%�Ơ�U�'^ZM����g���
��F��&�'��)#DEW�#:Ƹ��>i�,!Hh�Aɟ�m�E&��,���S�EF�-+�A��"O�إ �(�RT+�]��h@L?aP!�̘��'Ddʧ=Wf�#ꄿ��ݑ�V`c��׍QQ�h�S�	�
��$B=AM^�:�%�I��"ej�H	�tE�'PVE��ΐ��԰��!IR�m*5�Q�J�Fy�%�<�nUI�Y�ڵx�bĄ�O�ٻAm��b$�5�}�H���=�H�i�)��Q*�e���=�<�
6n�u�.L8Qł{8�Hs	�	��u �H%Z��؆� h5��nK>�� %�����4A�W�*0����On`��;����f��/���C�5�䪡"O�}��N��������J�� �5h���IH?��$��]��m�%ٟV\��ǧup��
�w���G�@zq)�F�d3&a�	@R���_��&!řk��0�W�$����ќcV�Y����0ij]"��̃}��Y��N�Y#
��j.���6"�b�V�E~b͛S�&Dc��O��{�0`���K�V�=����G�Xx�M�n��,R�E�"�J��DW.*����т��OJH��aGX9Rp�Bˈ,L���DX?��K�YC��0�jE�#(���S(��-
D>�ʶ����k�E��y2	�6P`�""�I(��!bb1�M�&�L ZD����<=JT@rf�Ro����J��O�H�íT5*V=h����"JL���UPxI�� ��;�ڽ	G%��	�=�e��+��p�rP4����2[�n<�P� �"�Z6�(�3$!i���1����'�� ã�MӺ��|�3�Jݠ� ��$#8��[�3�\��S
A�WB�|j"H�6�<��er%�e� =7����Xц�v�VXQ اO�)�,�.&��4�G&Y#S��]	b�Z�s�G,T&e� M��e�<W�Е{bǘ��y� ִ^}rͳ��ߡH�ȃ��yfY�u��?oR��4) >p�A���V5\wj��v%��ɘOC����/I1{@�A�!ʮEf�ѫ�#@^L�r��b���	�?�B�YPO]��0��*�"Aʱ�㍔����kC?c�\ґ�=���fW5(��<�VeY)Id��@(N�ٸ'0BA`��Q�0��I�~"��/hV���pM4c&`�镥ѥc�"pK[�	��ls��p>�2�ɗOZ��!�iC�%�]�zfy!�K�/���'�8خ;&]8e1'T�A��{����?�1-�P\ &��''��i�dj�4j�D��ȓK���C S�~; � �²
��o��uet��o��E�h8�������	�|9"�>��@U�8����,ef�Xf*6|O2��r&���$�{�8��ՠH�U��ya��/�Z,�(�\y��Y.��}&�8Ӧ�O1t�,�:�&�`�f"4��R���1�*�h�,"�0�@���j4��l�0�a}�B�Z�2Q4�]�S�B�i���"��<Y�'P�L�A�͢>�w�m�ލ��ޥ�e���DN�<��eR�N���B�$r-1g	B̓&z9#a牂������U� U�0�Hی�҉��"OR�U�50��j�(�p�2ā1jU YtqO����Y���5DO<�q�CMڡ�����1D��  �Q�:��,)A΍"��iZ@"OvxÐ�&K���DK�9%J��"OHd#$��"y�x��vй�"Of�k�E��+�h�ЪٳE���"ODq���Ch��F�@�8���"O����gT^	j'��j��"O2P��>�Ȉˑ,Q�1�&�"O�qb�oX/_0`e��썑b�vR�"O~h�O�?`g����-�`�"O������q���I�V y��m�$"O
,���4^|f��g��g��t�"O�Ѳ�d}�x�VE�;pT�"O��kf.E�N3�l�D,ԉo$�u��"Oȵb�K�(�*U�ݍQ��Bc"OAC!�NI���JأhW�f"O��CWa�`��Q���	TC�`�U"Oą���$�j9��) ,Un �c "O����M�y��Y���a^�=('"O&�� *L<"M�*�Gގ{�hM�*O� �a���.�KDL����$��'&���I&c:R1��N��!4٢�'�P��D@�%E��ls��ЙX�x��'�="��ݠ7b@���ͺi��`�'�p!��a��a�x��˝1-��'��|��eQ5_d�q� O l^.��
�'�Љ�U�SQ�J�`�	gv\��'��L�G�9�Bh�E-غB�����'�b��q��v�n�
�E�68�d��'�P<[�)�-g:�çn[,
���	�'G��0C�ϤQ_��#r&Y<yN����'7@�Ra�

`$����rSΠ��'U��U�oF�!��G�����'����e��6� ���af�Wv�<I�(ރTb�M�c��:��	'��T�<!�TA-�*�a�?BX�=B��H�<����3�t*q�^OR�H��@�<)d��^*AJ�Aվ2H�@��e�<q�n��}Â��!ǹ�b�@�N�t�<I����*���c��?tp�����}�<��L�/�|L���;BoXy���{�<i�.�?u<���kN�<������q�<AA�*s�i�tN^�V�>���$�Z�<!�C�F~z��C;6��R�[l�<	����s���b�ˏ�0�B��C�<�0A�'wNl0P1��^��\��Kd�<A�
C�d}R����TQS��}�<���3���k#^�i��xSKt�<�QǄ<@�
ɦ��d�1�TN�<���I��@t�L�t b�T��v�<�%ξ9bb�����S�f���_{�<���]�A$�d&΍nh|�@F
�t�<yw��LK�&�2D@��6������b�X5�(]�2x��R�"�F�ȓ!1�Q����1�
�6�>yN�܅ȓA�4�ᖃ?d�K�#�O���ȓd����\ke i�����`��� 8�ȶe��=��9��;y�P�ȓH��9���*R��%y���5}���ȓY��L���K8`޵����2%�q��X��X3�V��@��o�5P|,��!EI���<Vu0�g'7�l��ȓ~^*��G��3�NH����dS
�ȓO��=*v]�g�L9��T�=��r�j��eꀸ^I��p"��r�Й��S�?  �˲��5�4x�ыE�WZt �"O���"�ܼ�pפ�9/$<�#"O�`p��PQ�\@�"E�#c���"OBm�2e�ut X�V���a��,h�"OB�S�F.:���Q�D����|�"O�}�􊅝6 a0���y?.̩B"O^��E�^:�8�!H�P�r�"Oh�0��9�0xZ1ᑙ�����"O���,�3	&�@���x�c���.N��4�� R�L�x����L?B�*hj$�6E�����iB�Px�Nޏs��8���2&vZ�7������"CLҧ��2x u���[|�Җ�iZ�h�"O�h�)NE�����M�,E�icU�l�vbV�5�Y���U���(�%h89��5��]2vF5�O�M�3o��Tp��ąq,�Q�K�e�����Rd�HB��ZL��'L J��Lc��M�z�=�qa�sp�9s�dҢ��O]�|q�]?��Ec�.Ș!�d�J�'f]8�e�!"p��"���3�$���bYX4B�g[+$>�++O?3���>��ip��X�8t�g��n�<�ס�%G��P@��,T@�L����~y���0N�H1I���a�ax⭅�:>��#�I�KZ��x��Z���>i� Z�<�N���\u��1���!O_�8I"Nw�q��'��e��%N*+j.�r_�I,hͳ��䒥i_n}��*
I:�b>q���?[�V9��"G�Z�$|0��3D�զM�z4�5c��6Lqڙ#�r�����t�:|��>E���X7#L��mH-����F�S2�y"#�iXa�GT%�@�Х���ɨH��؁�oX���qF���|rӦWj"Y��1D�@k�ò`k�xҤ�F��I[W�2D�4�V�]�z	�5ڰ�޳q����#D7D�@����
╙�G�=�h��uC;D�$�����R�T�QQ+ܹh�t��<D���n��6��Lڶ[�w�,J�:D��QC�ϚN�41��׸!9:��1'9D�Li���;6������:c��*�A D��(���)y"�X"� Y�L����>D�xs��Z�C�,�p�a�#C�n�I=D�l��"�A8Ιhw
�\,��
$D�x��4Z� YkNF�Y�
.D�(��X�2� MY�^�&k���d(,D����
+��赍S�Y���1D��s#ٺ=E(h��]7���V�(D�8#�]0}��L� �Wl�����Rk��
H��~ӧ����ˌ����H�y��᠂��y���N�<�z��u b&V��y"��)Nt�8 �ҡ g�y�	D$)��=Z�*Ѯ`��q�ˇ��=f��`�d`��ĥ+��� �H/oƀ����	���Iӭ,$����#��l�Ǖ7U"���)��tqpI���0?�5����x�����O�2�(J�CБ]�!�d�g������J�,abS�[&%�,� v阨LŶ4��A�f?����O��q����-B�J��s�̡�"O�|�Va���l�񳅇�
v��?�`)ҍE��й2�\&g2��$��]]��j�a�)>G(AJa��yk�{R$ҥ�xh�w���XZ4%R#�%.� cC���G�ܑB��"4p
Y���d1��(�#�/,��G��%��AYgf!�	3*�� �G�7=*N@B��i��"*
 #T�
?�(��ի���2@����"|O�#��3M2č���)��y���0!J �T�M��8���'orP�T-��jv�7�K5Wd���G1
.R�Qv�T�!�DF�Zi��@S�^��7垏W��f�>$��u`P�~S��8u
ǚ^m��O�ؗOh�qQ�ޜ{�r���*U�@ߓ��1%��Gm�yYr�� ��Ik�	ȫwQ��D��O���aRn6e���'��>�I�V��P�T��$m��s�,�°�lZ� 5S�����:1�v�jR�
�*�`���0���2F*�('������"o������c����K�j�V=�2�L�2�R��FͿ+Y��O��{Z�l �+T~����Z*�M� 橁�#��wl����]*.�U"O\��W"G!A�h��Z�0*� cv�''z"���.㼑2B�0b-H��"G��`���'b�����!�Ɖ�+fԨ��2|m�8آL�`ܛ��@7E��[�B�4�-�ճ
�hk$�=*f7M�: T�*����#e���:\�t���,�O���@��A�8J���0tp#d8=����VJ�+����!ƵUJҜ�s�N?m��{)�L��Ay��8>e�b!R���h�4�t��'�_�+� �Iw�M�YA(Lz�0O�Xz�;1�6QH$F@D?��0`"OJ�x�/Q]WB�����O���*��'�-��eՊyx5�����ē��RH|z�fҸNn`zf�|��4�ť�t��T���_[v]k��i�dl�Q�Y�Z����Rf������&�	>�����L<1tm��miz���)\a�0�0b�u�'Bܚ6H�v��>����+��x#C�G6�؉�#�;D�PCFc�>a�ZPI&K�?5�hM��(�d6B���%�)����T$.T���"��&-�^E��A7D�D�����1�<���ϑ� }c�6D�t;���,?aB%�b%ʔc�*5D�h�ӈ�
m�"��V,L��j0�<D�py%M۾>B=1AW�^��V�4D�D��mW(Y<�=���`�j��u2D�����y����F��q�nA�0}(z����=��Ǎ[��x�JԮU���r'�j�<�!��3p�6�E
�*??��
�$���q �c>c�X0U����@Hqs4�9��,�O�P5 �{�q ���V�2�#�
[�q�G�����?a4.Ѵ$��A�Ù9p0�1r�]x�'���� L�ܑK|
4���$]�%�̗l.R	��O�<�D�I9pX���d�j����-Q?��D�$��e+4�F�����'����6A�Lu�EH���bäB��
h�����L�G�`iBA��e����.Oq�%%�W��Q�J?��w�K4�]��(3l<9kV�)�O�A[B��(�HX�!I�]\�`�!I?:�Z�������DSMv�\�"�ÇS�gG4h-Q���'ϖ.^.Tx��p��f�~5�f���$9�L���C��7?�Y+uH�7a�5I��
2zkv��)A�L�i�Q�՗�h���P
�4Y�!�	-}~�z�"O8ݠ5�8#�J�)�.�;`E�{4�3?�D] rʞ �(0��b'֦9�;���"43��S!��p?�c�[���Q1�?i[:�s�D��pi�RG͝�B��*j�R�(�'���1ʃ�q�R"?Y���F44� ����� �H���΁".�H1P���y"��Z>4�hcB�2��9C�J�R�>`��c6$��1c����F��'�p���TbM��@�6@X���'�"�x�g�z�µ�����)fe�ڴ�x�/�8�p>iљEg������4��8�/M���aW�Ō="B��V3O��Ag��|s܂�W�Uw�qC"O�]�шC�!��Ѳ�bllL˥�DK05>�͂s,Z�ǈ�qJ���

����P}K�Y�d"Ox��ՎF9,V2<��*�&N�lŠ1��]�|��B�>��(��l׫�<��'z5���%]c&�q�E����Y	�'��l��)Y���� �ƭj\@J0���hvh���͌�h���f��ɧ�O5|
`�C(B� ��'�@�~�	"���!S ��G����{��l�E
ȶ�����㙌W2�nM���3�x��O�|s�4�p��FL���rd���_\Zb$&���h���b�#M&8�|���X�nB*6�Lғ��6�>���ش�.%"��<���jބQ{a�r�����i��2�]�E �!���Ǿ&��D@E�J�t�l8R%�t�!��F�O�0e��G�|Y�lأ�W�G����'.w�鸆oq���R蒌��)[v��Wʕ���PJ$ʅB���$��uC�T �Ot���ePpL�@�&f*�h��F�y[إOP p�,�3}"k�ג�S��C5$|V���ϗ��xR�˾U}�c�BQ�[�@��P���A4��uǁ:r(݆�I`��X��E2[_��`�,O�k����ŲYY�Xм���'2����e���0a�OB��.��	��� L���,R�8�8�˛`�:���b�0�&�$��1kDD.�:Y�L�b��<=�ڨ��Na!Deۄ9�zHI�D89���4�Qr�\�|�'��@q�U	��+� v��Y��'IDex�Á��2�X�2̒�'߶|�0�� �24��dG [��z�'J6ʒ*K�i�����iΩQKԡ��'Q\|z��
]xjh+v ��S��=0�'P,�R�%�?w�t8��Ԣ����'����		�AŊ�de��<�q��'�r)���sw
U��a��ȇ��'Ć�3&���qD�5 M߀H��'�"� �!t2�*Gʔ+zah�'��`�#�G�H��j�ʬ/�,��'VXiK���=�X�nm^��'8���k�c8B��j��M�Z��'�@2�+�B���1t�^;)�E�'#J�
�H?'�,��0K<,.h��'�^��ƪZ�	� �*�/�XlUh�'�ZM� Ádqdb��!|���'|6����� k�Ⱥ���':���'��i��AlE%�aR��'D�l���-6�p�Də�J�կ:D����-�.��j�M���6D�TS3��Ϣ�� ꍌ)��e��8D���@�R6{;�����<8���J�)8D���ʝ'(8l����5�iK�h%D�$��L�t9��:�jڐ2y�����/D�(f�U,K�Tɋ�$�"�8k��!D� `��� ���GOԡd��8�a?D��3C��#>#����EYv��F?�y�A�X�� ɂ�Ҽ=��j���y� L	I�Y�S▋��8�3�
��y�C%lhL�YA)A��M�rH��yR��;y�){e�ͮ5XRu�n�*�yb'Z1P)��"sŔ�)�h�
����Ohe��f�<����ѥH�9O��E"O�PP�Еz+�q�S#B14J�"O�P�
ʪr�:����89-0� G"O"��*݂�H9*fb��h"� 9�"O|��T�X�&ؒ�o��%0"O��r�o܍e�uCP�H�$��4"O��cD�,!�p9���)zX��"O.Q:7d��j�eNYQJ�\ۆ"O�4ja���Y�4pCʡrQ��J�<�2� D��c���2ZB��(E`E�<�4 +)�^�q�2'�2 �D��}�<����5������^{�ux �D^�<�`+Y0G���C��L���f�c�<��%�\�,��rir�xp6��b�<a�%]	p�їN�"V�ؼ�R�g�<�Sd�2y�d��5��� �VCa�j�<����ڊ��c�� m嶸J�Ś@�<ibbƤM�L��̎�<�^8:��X�8�"S�@���M�'��7^f�ː"ԈF�A�'�F4�?�u��1(@�`��Y|�l@��#}�A��eKvf�1o�������� 6df���&/?E�.L�n�Z�˃0KԠ��6M��p Q��)u/�8�'��O`���ځh��#2���0�^�\��Њ]�<5*���>Y�j��0|�p)@?_i����9�)AgZ�� ���&J�O|��ْtW���~BN?E(ֆA�SЬ�*�eŨq���۵MblP3=OT�W�:�)�S�{֊�b�
�F$`P �><D�B�I�y�(J�Fٌ7�Le����0��B�	'I��b��M*^����0��(a��B�ɕv�"ȹ %�+P�<�U�d/�B�0o��D�Q#�.@4�Ġ�LrB�)� �d��ĴS��(�� 7/�I""O����
d�p�R�o�"�m�f"O�|��@.��|SE��"�����"O��E� (��:��oDR�:"O�h9���[�pd�ʙ��x��"O�� _�a�������)^.(x�"O^��Bͦ	R|s�b��*[(8K�"O�q+��Ϛ>��G�ΎUL>�!"O�	��D'R$�C�OkS>uȳ"O0���$s]JF�$x�!ӳ"O�{�b�8��-_?�a�R"Oeq�L�LVh�6��`�"O�t04��r��,��E�p���3�"O�l��`-�~����$sE��`"O�|�N�{�4���N58�5"Oa� ��;.���iCE�쭰�"O��a�i�@��]�eJ�T�� �"O��S�X�,����4k�:���X"O<aCdFO$
^ƱG���,0E�""OبqS�V p��P�Ń&D��!hf"O��W$ܩX�,P��0&5�"OZ�zg��:���5��`*�"O~�za�~�̸J��$S���"O��:7���5)��B��-!�$ǚ�h9�a\�^Ub0{�@��K�!�$A6=�smP8>Q���#@�:&�!��X�jtX���{<��f/�81�!�7Nt��f�-�u�o��!���i�]�5g "�[�Ȃ�n�!��G�p�fN2W���S�&�!�آgfڐё�4���\!�ĉ�nK��ţ �D�a`  D"!�� �^]\�m��JHġ�3IM�<!����L��''\�:B�A��
�?�!��L	g]B��SC��d-2�
>�!�
!�Z�§
,j�@�` ק8�!�)�pQ��I�3
y��dI�3p!���yg� �цV9{W�؊T��)e!�D	*2�楪��DML�	w�N�b�!�Մ澽��D��>��Q�n��g@!�D��<!��F�&9�#'(� #!򤅕�2��o���"(�?!�dڬ+=�\"B�'�D�s�V8!�W�v0L�q��݆:А5�Uk!��3GdF0�u���!p�C?X!�DȊOK���f�ؠ/�t@딾8B!��
D0��t� ��]��J�&)�!�d^:c�P���)��~�l��')Z�Y!��ˍf�@M8AE�/)����IA�#
!�O=b�&9�X;b�6�y��1\�!�$� 2a��ȥc3ڨa���G�!�DE��V����A�_A^�"��D��!��!��9�#C�K_�H+2���s�!�$Y}�0�4GD40R�I�Fې2�!�D�68�x�3�ŉ�o_Ve�G��l�!�#]�Ӆ��-/^����^=;�!�D���h`���i�X@F̛�Zߡ���.k+tJ$%��L�VI���yR$�U�$R"�+[Z{"Yb�'�����,R
>6�i��C�3U�V���'�f
'�!CpT�4�J,Br����'����T M0F����Ά�4xft0�'u6��۰9�x�&ؔ��e��'�H(�U��&�����JM"�t���� Ly��JV?Ő�8��K��4�1"Oڼ��J��j�~�#,�R��a�"O�8C�N�G Vh�� VC~ @�"O����!5NF�|���N1ffQkV"OB��Ο���� 1���"O�lA�vCPг� �c��6D��ia�&0v��I�(�8���5D��"&�I4l�� ��EIl'fș��8D���"Lf��X�2C�6.{�`y5�)D�l�VI�x�\(:�G%A��@s��(D�Y �˒ �x��.a��i{a@*D����L�-7��)R�7I�U�@,D������-�Zp�QϿ{��z�b<D������D
2��^JJE.D� ��`ՀUK��p���v�v�hDL,D�ܒf0�0�?	a4L���4D���E�ؕ'�Y��FX1 ,x�e�0D�Hz�Ie�&�k�DD9��,!D�t�Ы���T4���y��1�a D�(z@`�S���V.P�r��kF�<D���%_*P���������� �>D�܋Ԇ3+���	�
�H��Rv(/D�,��l��C{JT��M���"/D���-ŞH:V� @���I҆-,D���0�D�I�t��$�(Wy0��(D��	a,Q=u��50P�d�&/�*v�!�$�&-)���E�\e����Mۏi�!��� N "9je��>"�	�"�%%�!�d�4Rɴr�C�9nذ�[ ��,n�!� �"�0	�"���ۗ@O�a/!��̊i��q����3��\�So.�!�L�h��I���
�T��ar6�@�/!�O) ���,Y�]�Ƽ��.�$�!�$E�8^ɡ��9St�e���}�!�D�u��M�Am_|V���A�z�!��f5� DJ^?<]�z�'��Ux!��G�l�~p��O�pL p�DL�pr!�D�?s�:L;�I�i�w	c�!�dP�(EV�JF���^��т�@��!�d�X�0�(��A��fd�7��@|!��8/J���X5�dq��$�VB!��
	<�[tcM�Hu�{		(!�䟾F1x�ҠUh���D6,!�ڦ='� ����
������W'!�$�[�6�1�a-. x�hV퐾7A!� X���I�,ݦv��1�➙)6!�䂳$���"V06��=׏�"!�$OY�L���>d�|�1nҘt!���n�"8�'͘Y�@i�#��P`!�$M�=��2ajM+�j�X�	��|[!�D9al0�R�^N�]��&ư�!�$�4G�{�d�&[�|��d$�;{B!�)A��y2 I KȈ���LL4e@!�ė0(\���k��P�05x�œE�!��A�̠9��i��q�Z�F�!��ѓ=��H�!�Q�d��FiU�)�!��,HȔ;f��[r�-�U�ѽg�!�DT�@�&��eN�Wд�&��.!��W9{Y8��cUp�y�O��r�!�c�ԈhM&:��t���!�D�� ��*$'2��01D�ɟ�!�Df ��r��^@�"��`���e�!�d��#�3V
J2��-J�J+!�$ ҍ�Hw��!��Q�{!�� \���M�.� `�Ңr�&� "O��CA�F6�hy��!@ M肤�"OPq��.
��1��N]`�"O��j&N�L��t BnΥQ��zF"OU�r��Z�B�)1MH4bo� S�"O�xi�ȝN�uU�ϱsi���"O���h0F�+�ʗ	1[����"O��`7�ǃ��8H�iJ�}Fp�ђ"Ov{d�P)R�n1��.֋q@�$j�"O�(�G�B�+�rIr����~)���"O��d��'VLJ.@ٹ�"O�PۧDü/pNX�QP�[�"OrD�F�{M:m2gH�/BBlq�"O� b��#$����P��1<'��r5"O�`�"��eB��� �X*T�"O�Ы�j�&P�Q�`I�@Y(r"O\��5���p�er��53F��"O@-�߳G�5���7��#"O���Կ2��@ �O�0� ��u"O���僙�&��<���ʸ�I�"O�����$vd��pU���F��"O����<vbث����Ͱ�"O��%@Ыn��|��J�ˤl�"O��M��EX�eڐNb��)��"OX��gMġ\҉R��$��<�v"O*��bn0<:�C�����-�G"O*��` ��,ԐPM['mZ�]A�"O��r��rу��I��	�"OPX5iӃp� �S ���
prw"O��C�$�A=�1���!,k�"O"(r�'ĸ5a�x@�c�� �r-@G"Oh݃��U8��2Y�9=,��"O��[@M�	J��)�&ݏ>�x "OX���IU�3l��4T?F���"OȀ�3�F��B1���Ѣ���A"OD�K��V��)P�,E�~�	"On P2j4U�-��
�UE�!�yReZ�
DM�I��CN��y�M!�Q�G�7u�U�F��y"��5G��k�
K�F�p�h7�[<�y��b=
���7E��Xf`���y���(G����a$�<<�a�Pj�#�y2/�,�N�k������͉�y2�H�uV6��a�F������dL��yD�6e
�lxP��gf���uM��y�	����E�����Y/�y"����f�@v�	�Y�\�cO���y���xڠ���<�r*�yr!�SLx�KU����~���+��y���O�e�*�:5�a��J�y�e4�$��-��0��9 ��@�y�jJ�Kl�P����=�H�$����y�ǓJ�ݪ�dX78z����\�y"8}t ��d��8/q^uz3�Y��y� �sc*�Z��)�\�ђ)�%�yR@��1:�t:��%*E�& ��y�Q�S 0 �l��;A\Y�9�y��M/xq�OG�8x|�pE��y�"�<6E�boQ5v,1�X��y�G�K�p��̍='I��0U��y��;r��1��U�Q�d�Q��y�<9��1%F�TC��Sb���y�(�l�<sg�!�����C��yRaϚq�!�4��>$��W ~�Dȇ�S�?+�ş   �   �  <  |  s  �)  5  <@  K  �V  �a  ,m  'v  z}  `�  ��  �  4�  v�  ��  ��  B�  ��  �  L�  ��  "�  ��  �  R�  ��  ��  ��  K�  � �  H �% - �3 %: g@ uD  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�Y�G{���˾R5$�Qb+�jBƅ�7��Oi!���l8��Ӄ]*W>�\����]O!�ė��ތ F�8#"J��7Lb!���P~��#���(%l�(.ԜoI!�d�0c>��=`�r$,�
�!��LP!���6HٮsX~��!ݺ�!�Ĕ�m��G꟯i�̥sQ �W�!򤃛]Q���D�o��Z`A03�!��R�6j�l��B�^ ū@��;Ol!�P9��$`b��e&Ī���c@!򄊡jX�QTυ#i��A(PhˢF"!�D/2��`pB�]�6�`�6��9!�dEE����BݙB~�tK�`I�W�!�DV�=�i�H�!(^n8�䏔$g�!�$��mMX���9OT���n��O�!���-
l��WoР>J���NE�ni!��K�4�VYP�ɑ����+L�xT!�$�4<{��J��! �PhX6*ʨI�!�Ff^��PR*C�lʹ����F!�ͪ&�����'�4j�\���(�8\!��/�:��������bN	i!�$�<PⱫ��53���{J!��@�S�vL���?ʀ4sW��*t!�DT��`Iȧf yƬ`�c�]�#�!�D�p�,l G�.x��ᲆ�T<@Q!�@7_�����=�"|p0��-N!�"F^�cbI��i��,�g�:'�!�0�@1g�żm]�,�Ҭ�
3�!�d����(�qKrأR+�<q�!�ںO`�i�눏`�p�5mܒ<�!�d?B�>�1f��~�>�#���0b)!�$C6h���@焐K�и��)4!�� 4IAI�R@`�g� @K�C'"O�ِ��3|�V9Y%hS?<v��"O�y���<9�t��'��X=�"O�a��Q�/k ����$�Lu��"O08DF��D��6.M02㼠���5D��")U+e$l�ȶcX�6���Hu*8D�T�N�,N�n��4h>~��ǈ+D��@� Aƒ���eT�VD4��%D���q'�
1��Z&�Q�9h� 6D� ��a��1k��T% ���J)D��(�f�4��US L��1�z]���4D�p�3ϐ�ѡ��R/BI���&2D��I��.��s���p�� -Y����@�Ta��ցE��1 �oÓ�y��SZh&/\�SIRݲ2��y���(@��Sʀ�9̸3�j#�yB�ZM�z��?~�t�>�y�NÙ[8,�kWG!hQ�\�C��+�y��/����C�úkl�Y�-�yҎE G���롃�f�P}��eɱ�yBbӣ6OI��G�s�@�a�NI�y���(�=�"#�1lu�l�7' �y���8l<v1C�G͌eI^yD犠�yHг w�Ժ�=S]��������y�c�'�8*QE�K߾ț ���y�]*�������9,�ٸ o�#�y��M�j��D�2|¤{�G��y"#̽���h�A�a�Z��1Ů�y�)�s�0	���\Z�����yr�	z�H���+1��	Pj�3�y��XZXt�-�%`��ʤ`%�yR�IJ�P�����XWI /�y2���U?E���Ԍ|�j�!���y�c'�V��p�P��Bh7�J�y�:v% �𥑮r?l�i��y���T[�)Qg��}�`P1���%�yR���.���8�C["#�v��AOV��yBn�b=�A�X<� ����M�y�eD�_"J���t2a�5�̂�y�*��X`Ht���:�xED���y���1�J�Bc�"��,zu"OH5�5����\�B�ʄA��=��"O| [A�Ȯg��c/,�,��"OBy�hP3&>(��AI*�H�s"O��Ru���d�B�@(�&���"O�j�"�	�S �W�0�P"O������n[�}���>K�Ь�G"O���#��q�)ڒ@#Gt���"O��S��CT'��kR�Q�11��)@"O60�«�j_���hٶ4#�"O|P�d�I�j@@�2���4�,"O�@S��W���@�����TwB�(C"O��C�C׫Ix�Qi2���H�X�6"O�ɱ�dZ�{��ͫ�/��	l����"OY�!/\  ZR��BHW)+pD�ٗ"O�q�@C�lx�#cgިk���P�"O�lK�&T<T�����o�t�2�� "O|iA�,���٧��#&�YzU"O\ȲX*��9[V�C��|@r"O�-�Q�j ��	���`V�lA"Ox�ۡ,�:m�d��qJ�i��h"OD8bC ��\��c'/0f���)V"O� �/<]���z���F:z!�E"O^���'�����+�"ԋ$(�S"O� �x{U�jHXAY�̓v�x2�"Oࡓ�O�B"؈ �Z�6�1�"O�Y$�ِ$���RS���>-vd��"O�����?Kr�HA���X�=��"O4A$!8<���M��L�`��'z��'��'7��'��'��'tj�1���<w���G�B���'\��'cr�'?��'a��'"�'R.@q��y�|$�QՁx�ځ g�'��'~��'��'�2�'���'6�0�M��
���U��1�� p�'�r�'n��'R�'2�'���'�Dq���+K>��`�3������ş�������џp��ݟ�����4qlڌ^Q�<��W P�t�ǂ������ԟ(�	���Iʟd����\�I������Ԫ�^�h�c�I���3��P�	�����ޟ<�I�,�I̟����h�7ɘ�!���4&��W�����JΟ$�	ڟ������	��	�$��̟{�f\�`��<h�c�� �x|��iP�������$��ƟX��ٟ��	џT�����I�Ε�!�����P��
V����D��ޟ����@�	���Iʟ��I��|�&��D�d�r���>�D�$������ ���0����d�Iß��I��$��6&��,H��[�e�6!W/_���ş��	џ��	�t��ȟ,���,۲�%M	����[�ТZ��Y�������h������	����7�M;��?Y�R��"��8a �i`��0k�	۟8�����d�hG�N:`pLC¤׵����&K����_3�v�4���O>�&��O+
ͫV�� Wɐ�����O �$ڛl�07-+?a�O���5�$�<iZ�]z�)�=U)5/�)��'T"_�lE�DƷ�h �a��8P��u 6m�0�1O��?5�����@���b�h5��k �;gᕅ�?1��y"R�b>iѦ�S��Γ6!���֌��u&֝�$c�"~b���yrB�O$,��4����-Rg���J^�fL����]�)D�$�<AO>�i�Z�j�y����ة��V�U����b	��]�O���'���'��T>�05Ù���fѐ\��b#1?���bj ���FF̧bk��F�?I���gb2e"��F6�E�� ��<��S��y�,T��Sv�n^0P@�H��yB�|�!qӝ�@Rݴ�������y����\;]��Eh�D�,�y��'���'N��1��ic�	�|�#�O��)4n�!
6�%���w�=å�X��]y�O�r�'%��'3�i�3J^�<�W�Ւx��dC�B]�R��	!�M��V��?����?�M~��}�n���G��rS�4`�ǻ�Nu�$[�������$�b>yr�O��0f�X���
R`�3x���mZ|~�*Ȋ]����������;�
�j�#1�0��$�.;qf���O����O��4�|�
C��Ǖ8��-jN��	����!�3fc��t�*� 8�O��D�O��$��I_��ఫШ1뤔�'b�1\�Ĩ(%x�V�!�,�3s2ʧ��KT�S�U� �h- �c��0��<Q��?A���?1���?���o^�Jn�9�F�U�_c�hh@��8a���'���l��8)6�<a��iR�'�aI�� 3�@�x�ט~u\��P�|��'�O���h��i?�ɠDҨ�L�6]���"uIР��~]"��+~�O|��|����?	�N�
��S�l����"�C�Hb�����?�,O@�l�e�j�'R�Y>9���%�X��b�H��6�cw� ?y�U� ��۟�%��'6����'��ec�t1�O�p��k��Uq��,�޴��4��i��'g�'5�a(�F���|�cv��]�v�rv�'T��'o����OS�	�M��L,���b6�O�s�T���(1z�����?!��i�Oة�'t�d��8��H}�Z��V���'��Ġ��i;�	�f�:�����&�P�Ju&U�Ev4��b��fu�D�<i���?���?����?�*�2��GLؘh_̱�!�*q,�C� ��I;u��� ��Ɵl&?牟�M�;L�I�l���BǄ0u4��Ο`��z�)�(p40�m��<93Hڟ-����HE$P����<�"A�8"�^�DT��䓢�4����"X
�h�(�dZ]K0��/�O���O~���<���i��)��' "�'��|rp��:D֐yR��[��9ѥ�Du}r�'���|�\c�]�� 
���1ሂ��$U)vy{�`�^c>����O��d��G`���
�y�:��d��!���$�O���O��D!�'�?��!�~DŒ�O(:����?i�i*Z���'�c�X��]�h�=��J�ce$ٲpĚ5�x�����	�� ��Gצ!�'�,�&��eʀ)SF�iAL��lJ� C����$�O���Or�$�O��	�b��婒h̎$��PE��B��)�f*��R�r�'�R��d�'�`��gfG?IAn�#��[�~�Q�O�>	���?	M>�|B����L�jq�q�Ũqb C�_�CҌ��4��$]kM+�'1�'��	�$@hq[��ᐝ�g����D�	�$��ݟ��i>9�'G�7m�{����2F����� իmP�re�������?yZ�@���|��4ik�4��@S�(��(��#B���tB�����)�'�20��m��?�}��{�? ���2I\�*9l`���:rP"6O����O���O��D�O"�?u�� �-$1��@U*`e�!w�W֟��I�l�ߴ;q���*OPunf�	�2��	�@D2iM�[ �	%���	ʟ�/ƘmZB~Zw��Q[d��\��ϼSUXy��nٰD��L�g�	py��'�R�'���K�jz��׫A�9�@�@�pr�'��I�M��	��?1���?!(��� ��ׁl�|���_'-9�������O��$:�)rf���t#�&Y��N�X	�g�챂��_?|j�eX+O��C��?I�A$���(+t>2���(�Й��O.N���d�O����O���i�<93�i��E�b���Z���J��	�t4��N*��	2�M��J�>y��j�ё%��|���gR�R���?�3����M+�O���v��)S���B�8���2���8��U���ςrH��<Q���?����?a��?�)��pԬA�:Vn�b(ܚa��9�b�ͦUі�
myb�'s�O�R&m��n �k�l��ǂB�����47����O��O1�|�j&,u�6�ɨ;�*)� ��2n�RE[pH���c�,��۰n��d*���<ͧ�?�v �-��P���^O1R�I4��?	���?!����N���E��������,J'����p�ZԫƟqh���b�Mc��h[����l��]�'_� y�e�0lD8cG㍓���`����W�(��|���O���OD��3�֥BlR�i���/0�%���O
���O����O$�}"�MDd��5L|�Y�-=��I��G����/<���'�61�i޵C��ìZf��+t؛4,!�w��æ���ٟ4��mU�9�'fҨ�t ��?����5L��(�)����pJ� [��'��i>��I��<����4��"f�`);���5��v���)���'K�6�Ӕ~t��D�O���/���O��k�+�	�j�r��a.qKG��x}R�'�R�|��T���K?�4+�4P�`�`@�l�ݘ�i
�˓����n���&���'� 1��`QRq�䊶��
]lc�'_��'�r��dQ��;ݴ;4�Y�:�&� i�B��k��&Z٨��:��v���d}��'���'mژj"iF�Yd���e�^8� �*ڃ:��6�����ǆ6��t�	��Hɚ��5#;��jP����5O��D�Oh�d�O&���Ot�?E�-�;C��j5��ؾA���՟��I�P�4�n�ͧ�?���i�'h\��C.�!�%��$��\�uI!���?���|�#M���M�OҸ ��g�И��D�7FrF��al
 	x�Q�'��'���`���	.Q�*��H�D�ԣ� �UR���ϟ�'47�[t��?�)�z���)�0�VT v��%� �R����O����O6�O��;GM,��a
F�-H�q+&�V`�d�st�B�>LvD�"�ey�O��,�	�"��'�ҁ�`Ӝ�88�a���O Ɓ��' "�'��O��ɷ�M���O�T��s��X�(ڕb�,�0X-O��o�o��^��	��0`�ȷ{iJ4j�� *U<}9�oßl�ɹ�$�l�C~��^������W���\����a$x�a�i�)��$�<���?���?���?�+�5��ّP��5;���9��y!�	W��a��"��������8��ŵ�y�.4&�}H�7)�H3��6J��'Bɧ�OO|��űi�d�<"���*�c`���!	�zi�䎭b?��q�' �'��I��@���*T%��#����ƌ (N���ܟl�Iן��'C�7mVG����O���,��"OfaWc+�p��e=�	�����O��d3�d��s�>a��M�\�N��]��ɐ8D;F�P��|�f켟��I)#f8d�~2�t��@ʇ@�&�I̟\��ȟ���G�O'��O�*����	,�r�#��6U�Al�1�E�Of�$�ߦm�?ͻ�5B���)̳�nuɶXA�4Oz�D�OV����*6�$?Q�[2*WX�	-��zQ#��2ڜ�js+­e}`�xI>a+O��ON���O���O�=������P%���˓�R%QT�<ɔ�iӸD���'�b�'��O�"�?4�ai�h��zb( �f�2 J(듆?����S�'|F1�%��JCkT6d�N1r ��MC�O�JĈD��~��|R��	�n��zh"7A�Aj ��Dܟ�	���	ߟ�Suyblv�(I�v��O<8�v�Y�]i̝
��\�Y�3C�OV�n�y��a��Iោ�	Ɵ�j��@�" Y2
KH@�D�O E�J�mZ`~Bh�>���'��ֿC����L�+p�	Z�I(��<!��?���?����?щ��
ܟM�f��Կ�E�N� L3� �럌�I��iݴ��ͧ�?��i@�'Z%���*��T�'�Ŕa#�ͰՑ|"�'c�O�@�/�MK�O<�J���6a�*�	���-3|~0� ��2s�h3�'��'s���h�	ߟX�I���j�ƴI���PӯO6.% ��I��'��6M^.j�"��Ov�D�|��a��_l��V���V�6���ECR~2�>����?�M>�O����a��>��MQ(7�� C�N)�\	�#A #s��i>McU�'��y'�����X�!ؕXC�*.��d��K�ğ���ş����b>y�'V7�r�RT;Պ�<n$u)�#X�?���
G��<���i��O>u�'<bK�."�T���'N�M�d�P�:v�'���13�i�i�=ʦ���?e��^�� ���ʃ��u��MC�b���zC5O6ʓ�?)���?���?�����]�@������'�Щ���W2>e�m��Ti���'������'Ԗ7=�������K��A@��N(�Z�A��O���8��iT�z�7�j��s��A?"��K�SM|J ��-z� �#L:Dt�$0��<���?1Cb$�8��H(B��8H"K��?���?����d�Ԧ�kf��4��ڟز5M�.X����FP�{)�u�m��zy��Ο��Id�n�VY��D�m̺��W�ѡn��4��u9"��9TȀ�|j2)�O܀��_�N9���s��,ї��3(W�A3���?���?A��h�r�$�e� x�-�66܅yU��,���Φ��r������I��M���w R�cBFJ<
:<��ϿS@-8�'��'B��	�E�Ɲ�����P�iF�D�j��r���a6��$ �1{���O�ʓ�?9��?Q��?I�l��D8(�*9����҂�%V4�2/O��n�3\��=�	��(�	\���D�q���P%�Z#O�4O�aCu-H����O��D;���M�|l���7�y���Z	O� ���Ҁz+�M8,O8�S��X��?�7�9���<i�$�����l�9��y�b�>�?y���?���?�'���yQ�@_ʟ�P��͆A�������Q��l���{��	ܴ��'��?�-O>��Q�Z�X|��9t*H�y3<�ȗ�!'�7�=?���Y�
�h����'���c�KF*i+��:���H��Y�<i���?A���?Q���?�����(�\���%s�B� ��^�P�2�'��(b��+:�����!&�HY�hռ<�|ѳu-߷p�8d�2h�V���d�i>-��i���'S�Z�#[ x�2��c�{��-
 �E72�	���䓙�4�x��O��dμ,
.Q悈9�$������b�$�O ʓ~����\��r�'�\>Ȇ,��@�fyY$b$kH���??��X���	��%��' >mQ�E�<��,�!Wu8�[ "�$�D�k�4��4����'"�'o�� �M(��<�2,Ƌ;��E�F�'�r�'����O�剗�M���*1��D�3R���`��>u4�+O��l�]�3�I��ĸ�.Ϝ=�mۃ�se�cU���ɒK��m�d~Rg�5A��4��[�	�.�L0�/E�X����n+��<A��?���?����?�,�h�I���> ��
��3f�V(��@Ӧ�@������	ȟ�$?����M�;B�v�Q��=(�H����*gG#��?�J>�|�A�+�M��'�����)���;�N6R�R�'_�9���y?�O>q,O�	�O�e0���j��^���S!�O|���O��D�<y��iX��'�B�'��Ї%X�>;>��VD]�Q�����D�]}��'�r�|"�v���z�i�y�3#�Y����Ә2�(�C�Գ[�4��, ���^���$#,Dɐ!.��AGKN �d�O����O��&ڧ�?�EEݼ[�p�	���?E � ��ô�?94�i�\X{"�'ج6�0�i޵!�ʈ&h� �
�d�4r�xR`y�h��Zy"�X�TU�f��HsA�Њ& ����6�v�F��4��T	v5&�$�'���':��'k��'����_c�,�D�-�B�r�\�H��4*��i�,O���,���O���6!X�p�d����.{Z�tjդ�_}"�'�r�|��ԥ�4 Pr'+ѥuB呅14+P���'?��6l���P%�'���&���'z3F)6~,\��!�'/ ����'�r�'R����]��	۴5�hq[�N
Zd���9��h���G8�$���K��V��`}��'���@;��+ n�;Sΐ��Pc�/�R�ZV���'��J�E��?��r��4�w"@�DE,uo6��� _$A"��'L�'>��'"�'Z���xV�����S��#3U 	����O���O8�nK�6����|�P�~�b�n�"a����"��)��'�"������'ԛ&����Pd�2�c�<��a�̥(��Z�����|W�<�	ߟ��I۟�zd �Cj�R��X2Mh����4��iy"�c�vm���OB�d�O$ʧ/�`�Ӥx��Ya`E�;-v���'����?����S�4f�\������W���1f���vbF��� '��擟�����6�D� !��Y��-ήF�������l���O��d�Ot��<�4�i㼔��#Z;�
5Q�f��'&����9;剂�M+�"f�>y��P��:Aɖ j~�B��8$�|
*O �y�b���� 	Q�F��$�(O���2l��b�j��6�U���#2O�ʓ�?Q��?A��?)�����J�HZn0S�
�������Tn��~@�	���	U�s�p�����s�ې;��@����;yg������5�?����TOO�YK�v4O(�9��� ����9c�x���=O��/���?��>���<���?���F�?�X���&h�5���1�?y��?�����CȦ���LƟd�IƟ�8GF�1w��I!���,[��N��Q	�	ǟ`��E�=r��m�\3�bC�-��6X��	[PE�M~�3'�ODE���K�X}��������!�B�?��'�'���S�x:��>/�|	�#�q\đ��� #ش�bp���?�W�i��O�.C7�i�A&	�����c@O/.m�$�O�D�Onaʑ#k���qyzp��?� �����-��SLߵI��T	��$�d�<)��?���?!��?�0@�;80(���Y�EB�i�ɟ���Qʦ�1Є�˟���ޟ����Ży �X���@���a-_��I���L�)擉\I��ˠ#&�*�b�L� 4�Ȱ�Lꦥ�'�J8�dB?�L>9)O�i�A��8�pS^���D�Ь�?q���?!��?ͧ�����N���`�7Z�>�Z�&��1se�`�'�S��X��4��'>�ꓣ?����?�A�X�9�H�+)C��E�ఖ���M3�OB��cF��(�t��Ԁ�0;�$��^p���m\��OR�D�O��d�OH��4�S1C�-���N�J'��dK�@R� �	ӟ�����M��|B��N����|2l�#Nu�T�SHŅ���sa�-��'�b���tB�<*ƛV�����:D>������fq�!�g�œb&6�K��O��O�˓�?���?a��~g<�AC�ȲU�z"@�Zw�$���?/Om�Q8��������o���ȗ:��ōA&3�`��������C}��'Hr�|ʟ�H��Ř.�z���i�j�9�d��H*��h�(_�LI�i>1���'��&���(ð!�E�3�*
�����T�d��ɟ�	��b>a�'�\����6�RJ5��jU��J��A�Q�'�b�h��8(�O
��3O2��I�V9��Pw��h�&2��?I�Å��M��O�mSO�O�t�&�,T�\�ё��tMH�H�'��	⟼�I���I����IV��'�
L� �鐣ɴC��Q1NB�,N�6-�0*v���O��d.�9OAlz޽�׈Պ^� �-S:46�9���러�I@�)�847p!l��<y7�%�h9����y.AQ�<1���"[����1�䓢�4�����*3����ɝ�.���	X���O���O�˓p����̓���'W�w�$�p�A�hx��I���O�<�'�r�'��'�){�(B�pԊ0D�ˉ@�.��O��I�)��7�!�nP���O`a ��!J�5�FQ�Jx�w��O���O(�d�<E�t�'ᦘ����6��l(��5;o�ar��'f~7MB�D2˓DQ���4�0Š����1�$�!����~YV�QC=O��D�O�ZB�7�5?�U�_z�@?,ڑ,#j�Q��A�f:�X��K �$�<ͧ�?����?����?�����\�Nyc��_������������E�c��vy"�'m�O��i��Um��PP!�!D�0ohj꓊?������Q/o� ��6���}�:p���/�M#�	�!��I�w�Xt�g�'��'�`�'��t���]/j�* ³ ���P8r�'[r�'7����dP��شV�<���lo���VJ�>���`ac�Y0�����Y����d[i}��'���'�f��w%M�Y�(D�A�5ղ�`��&_�6��Pˢ��#Yi��?�	��p��^B�ur��Q%gOp�(0<O����O���O���Of�?1�s*�zo�Y�2�82���{���,�IןX�ڴ-.v1�'�?���i��'b���ڴTCV � e*3� 	�y"�'P�	v,��lb~2&�'AҺ9a��S�8�``�T+�`iP���ҟ40��|�]��������I���0Pcլɢ ��#]� u�u����۟(�Ity��dӎHȢ*�O��D�O,�'qxL}:��;����R�:(�8��'���?����S�d���O��(A��KWo�mr��?����t�7N֛擟�ӦK���-�ԮR3"S�ϒ��b��EQ�'���'����OV�I��M���$/z|�����tA�֍�l% �y#I�<Q4�i��O��'�Rb��h5�����5=V:-�E�V��剠$�llZJ~B�̓.d�H���\L�I�"8�����4���"�T"
����jy��'�B�'�R�'�B\>�H@�e�&X�̺-c*e�⛒�M��ŋ��?A���?�K~R��X���w��f�uT:�r�(k���'&b�|��dc�t�?O�J��)l�ȁ�ՅP��PP6Ol�L^�~��|_�$�	�������N�~<x���j�.���k@ٟl��՟ ��\y��uӌ�jPB�O��$�Of�;e��+ ����Ǜ�gcxJq�&������O��D;��Q�n��|S��!0lz��$�/Ft�	?B0ؼ#�Ŋ�_��c>�+��'��5�I;Vv�Aj �e��t`�I�<��������������Q��y����z���a���0��h���*A#"�y�2�Q��O�������?ͻH���Ŧ�9^�8)9�BR6K%^e͓�?����?��OF��MC�OȨ��M��������U��D�U��.�xb�'E��؟���(���ɯI�����m-T��Y���0�^zy�`}�6�`�<a����'�?��iR�$=�t B�*y�(Q&�9(��������`�)���H)ϐ$"{n(**�@#����@���Y�'? 5@bˋC?�L>�-O�hIq�R�N@u�$��`���M�O��D�Ox���O�)�<i@�i��i�&�'^F��GFE�*��D�q�I�w�Fl؟' P6-5�	����O��D�O��y���_��j�	��e��"��Z��7�9?���V"-���!������do�"ھd�AI�4�ޡq�fa�(�	��IΟ�������"�!mNT�`��vW���@a��?���?�v�i���O��hӸ�O"���2����EDY/5u�y��.#�D�O��4��qEoeӨ��|D� D��c�C+$˾q��Mע.V�A�b.�.�~�|�R���(��Οs�䈖W�y�%��%8زٱ� X��0�Ilyr�h�J�bb�Oh�D�O��'U|v=!��ʒ^�X�t�C�2*Z�'�4꓂?Q���S�DɎc���'�U�.��H# ����0��A)p�X]j�\�據�ҩYa�	/R���f��\Jb!p��>^������	ǟ��)�SQy҈r�Ƭy�/�8&�y�!UYxPsg�*G���d�O�n�B�����Ɵ䙇̔�;F���p+F8�T��S,Xny��?�������
���M�Hyr�T�t�=���O e��J�I���y�X���I�T�I����֟$�O����U,
Z�p��/C"�jU�nӊ�pP�O����OB���D	���CK��`���u$��K�cP�2����ԟ�&�b>s§�ئY��Z$��3��9�%U>(͓D�,��si�O�PZM>�+O��O�����;}�0<�q��^�8D�O��d�OX�$�<��i��0��'Z��'-�݋@"x�}S ^1:^T([���J}B�'b�Oʱ���Y�P�)*���G��Й�$R4	��i9�i)�Ak�h<�����ॡ�;'��#7��X��`�b�ڟ��I�0��ڟ�E���'n�4��ѝ0^�Z���7�%�'Kx7C�ʖ�d�O�mP�ӼC O� �*x������q�͇�<���?���j�n��4���F�t`Bm��'p2��a�,��~�<0ۣ)Q���Ó'?���<�'�?����?Q���?����/ZY�
�	nfJtd����D䦩����p�	Ο�'?y�	�c�ܭ���#@c����.�ʀ(�O��d�Op�O1� ��éOJp�i;�Ȕ>��]RԨ�A�i�Z�t���K�Ƶ��'���'�d\AN�.z��!%�sbvXC6�'�b�'����Z��H�4w��$C��oM���t ��]JL�t�Z�� ���&���A}"�'o��'Ά�G��h����8N��!��yN����rV��6ai�)*�	��Z����Ֆ ,T���~}L)CP9O^���O����O"���OT�?�"2��1!���P/C�'����L����۟t��4>�lϧ�?YP�i�'��9�˫��i(@(��sWj�pV�|B�'��O�M�¸i��	'e�����^ƀ	��)<hp�:(þq���`�	~y�O���'�2���)�ҍ&�̗�t]Jd텅x��'��ɹ�M��o���?���?�.��d��HeY慛��Nd`�r��l�OT��=�)�A��y��!6�8�h#� �L�&nݗJQ )O�8�?1D�-��E�L�T5C�HBm�  [�5(��d�O����O2��<��iL�аu#W�'�	���b4�H�Ci��[5�	��M����>��i����gB(�cOE0:�
Q����?�ӂ�(�M��O��3Bې�I?�Y���L�d0f&R?^
��yD}�8�'���',��'L��'5��_�صrB��F���C�B׺a�E{ܴ
��Y��?9����<��y��G%b�I��ׇ=|���U,ӈ#�R�'ɧ�O�j]���i��bQ,�B������t�r��3/��-<*h���*��Ob�S�jC.in\P�7(��a�&�r����0<��iS���'[��'79�'�#AW�	1��l�25�� V}"�'��|�z'iɃ,�18����2L.��$Y�:�B��	�MS4��d��R?���m��3��:��m�Rh�]�\��w�ma��;e����썅\̸L��8_�f-���!�M��w�pA( ͞9L*�r,@ 	��9!�'P��'����&J�V����	��%���F^�
��h8�B@�s2]��|\�8Dr&�g�!��J+6���nA��dU٦�;��������ڟx�*�/:]�� �G�+8�5���&��	ٟ\�	e�)�ӈZq����
�`�j�R�HP��5�����.O�0`E�K�~�|�U�ĳ��ݏ}.ĸ"�$��,�h)��%�O~�m��p�R��	!8��Y�LkE�x�R�לVǄ�ɂ�M�2f�>����?1��:ʭQ�Z�<o��P���>j~<ە���M+�O��)�l��V+&�I��<�qOL9��C�&C��0�;O�����d�D��7�D>?�%E��6�d�OV��]ަI!�5z��i��'�Q�s%��mOb%zᇎ
����|��'��Ou\��Ʋi��	�`�d��OϸP�l�ڒ�I+�A�r�A�Z���<���<1�B�
�Uu����O�t9DphG�J��OJ�m�a�Tŕ'4�Q>�ñ��9`�Jq�2�)k�	�N1?��U���ޟ�'�������N�<F�^�F�Y�I���PL�8&lUC��:��4�.����ꢓO^�2CJ�����$�+;)<���O<=n�%D��+�׎b�l@ڕBA�v�R��$�����	��M��i�>9����;Ԁ�6��`�>������?1��^�MS�O5 ����U����i;/Z.-�kɾ\��Ӈ+k���'��{�C��c R��f�w���Q��)|�6^�4�����Or��'�S7�Mϻ@Бa'"�% ���ZPbN;������?J>�|J����M뛧� H�@��L�BCV����W�w(�(&>O��*6D(�~ҝ|�[�p����0��.
�r�҅�`��/?�S�#���������	qyb�z�v<��'�<Q��:��$�shW1H�4Ja�6<<=����>���?YM>	u'̗�p����@�� ��Y~"l
;� <�p�i�ғ��EX�'�g$"v�1zN�7uЉ`@�n6��'w��'���Sݟ�P����w��e ���]�"LV̟��޴��0���?���i#�O������[�(�:_�V%����d�O��$�O6�Bd�x�~�T	��Qi�?��JĢ_�,�ĥM�] YyS��B�	Cy��'��'J��'M�Bʱ}��vhͷ<qΈ�b�]�j剭�M�aM��?��?qL~��e�yʲ(ٺH<���b�ܼ�rV�D����$�b>u��$�j���h �E��D��zP�o����dF "����'0�'r�I�m��p��bC!Z�@<J�n�8�9��ɟ��	�L�i>Q�'��6�Ъy����8
/r�Q�Z�7�P�/ �B�B��ݦi�?�eW���I蟌��b�f%H��S�D��� ���*v��ئ��'�NT:t��?����t�w�4�=WFR��p�V�t"ސ8�'B��'���'%��'h�2�97�J��*|[1n��i+6� ��O���OԸl�9���ן0��4��l�X�{łG!#4��X�L�b��=�N>Y���?�'e[�dk�4�����٣�Fݧ?�"E�jЖ�@'�"m���������O6���O��>��83+�2�����~\�d�O�ʓl6��@b�'^>����FC�Z}`2%]��n�`�u�8������O��)��?]����&���+�zV�����SJ�Z4ī��O��ᗧ��E���J�|b!I�Ga>�9��Y��b0[1d�F��')��'m��^��,�h�!!Ꮔ4�&��"�PT�@D��;W��$�Oȸm�j���`�O�G�k��S�daL���	�q����O��R�ai��w��U��?�'�ƙ�RŞ'a��q�`\�L�P8�'Q�IX�I�|�����M�t�[�h؆�S�w�Ms�u֮7�
��x���O���=���O(�oz޵������E�Qa ��LP��"[��l��D�)��&|â�mZ�<��P$mXi�w�W"�\����<����u�t��������O��d�$�i"%�ў_����Q;%��d�Ox�d�O~�U����ݮ���'R���!0�&�R2W�|�GC�)]�'\�M�>	��?�J>��	8N�6�S��W0�&TJ��t~�ٹ`���g"��!�O����	�!Z��F�qA�x��a�.V7�J��	�
��'Wr�'P��s�}�r�{�e`Qa4f��A�f�ԟ�8޴\�"H"��?1 �i!�'}�w��b˟�|}>���.ۘS�e��'��'���%��&���]�S�y��*!&~����ׁk2�,[0�לz*ԩ��|bX���Iߟ����h��ϟ0��O�\�4��&qT��
&�y��dӔ�����O��D�Ov����$·c.��0J�.�lׁ�1�T�C�Q������%�b>��%���D6�a���{�ɉ�="�nڢ��dN�l��1�'z�'v�IjC�]*�kϳ@�U"�	̣Y�����ݦ�8!�OϟD�U&R%���e��XJ��$�j��A�4��'���?����?��,� ;^<���&��8���P;xD�؛ٴ���n�!���`������J5���bL�f5�a���ޚ<��?�O����E'@����!�8�,� 	�<�> �fC������ަ�%�Ȣ� �B��}HgJ��$�� �Gl�ޟ��i>��a`ۦ��u����@ A&�A��IN���B��,��|�R���?�џr��ih�����4�x�'��6
~����Oj��|�֡E�(��}��J����;S��}~2ǵ>9���?�J>�OR-Cp��(c@<�L=}
Z���!�"nR��p�i���|��J��('��)T��u�T3���/��xRT
O��nڢl�d{է��a-�M t�#0}8mI�&��l���MS���>���
�T�d�۰=�n��Ɗ_�ح����?ٴǒ"�M��O<��4�M���d_�<��&��"�2a4�P��e�	rk�Idy��'��'�R�'�V>�J�]0?	����vE�1"pg���M+�A5�?����?M~��r��w��� ��U���kD�E���'@�O1��H��ff�T��5g�V$XC�>�Vl��N`���	�%v0<��
� }8�E�)^���)���
����&�Q�@ �D�'b��(y�%vPR�䐇<A2	�+���������=/8�)�#Z1O�t�B)�1''�1#`Y���y<�(F��'3�(p���/,��	�f��,.�n�5�9�X�`D�Dq.50�jT�PGґ�C�
����h�5IT��&W�yM�IP�����T�KT�%{C_�>�xX�Bo�+C1�d�� Z�M%�����:s�@5��c-%5ʬh�+��L�����Vf�e#����o��y7�#@����b�ݔ�,6�O��D�z���!w��o^��ͽ��<n���P&�������Pg����O ܸ��)y��9�F����ıi���'��	��l|X������OH�� "R��4�]6�L�)�eT�a�T0$�����`J"'�K����h��g���pD]�1G�Lk��3�M�(O��i&��æ	��Ɵ��I�?k�OkL�)O ��t��0�f$�S��J���'�B-��ub�|2�� 6�0��H�Jʠ� �ߍH�LEa�i&�1�%y�P���O@���&)�'���-tV�,"i�cZu{��V�r�J%Zشr��������O�"/�	6�@��_h(���X�J�7��O��$�O�PA�[x}W���	?Y,	91�N���F�s����#d�q$�ȳ�J�<��'�?���?AB�NX�F<��h�(�����$F����'8%�	�>�(O�d7��ƺ|�p��7$�Jȑ$��,/`�	�[���Ծ8�O\���OX��<qd@#W�l MFAt��J�12�\�l�'�R�|��'�r�J�Ph���T�RJ�@��G�@�%�G�'
��ӟ��Iɟ,�'�6�
T p>�Q�L� �Qs�*\��H[��qӖ˓�?IO>I��?	BPt}"�

ɴH!E�Z�@څ������D�O��d�O��a��Tk�S?9��

'8�hp��w�V0�@�ڹ|̖�Z۴�?O>���?�����'-R�*��IsF�PP#_�y��=rߴ�?������ſS����O!�'?�4���Q�X5�D�S:�]ʠ�2BOv�d�Oly���:�IPr6��>�0��6�Q�<ڶ�#����'-����j�@�d�O2�����ק5���#A*��b�`��&�i�F��Ms��?�®<��'q���c"b�7Q9� d�	f�Ř��i���	&Lj�r���O����TD%���(t��m i�&��E8��y������M�)��?�W�Q&�ӡ���W�A�����';��'�����4�4�\�������ƩZ� ��MM%9��,���rӈ�d+��e��Od������Gf+�xx�����. ��ye�q����ޚY6�~���m��2�! ����}�"ɱ@㍧EK�����x�n���$�Of��O�8#4ș�E��w����
56�U�5�Ϝ=^�'k"�'x�'j�i�U��԰3�
{�^ x�>l��{�F�$3�D�O"��?Q�D����t�(�V �T��)vb�X
 H���Ms��?1���'��Ix�7M޹P�����'�a�YY2�
J?��ܟ4�IޟT�'�DpҢ�/�iT�_}��j��S" @0��7p�Z�l�p&�����t�'�'=°��e�ԣ��P�`E�.�Pl��D�'*"`Ȉa��Sߟ����?�X�G�%8E�K�M���`�R']�.O@��<��V��u7���	(sL�e��������d�O�p�u��O����O��,�ӺK��o����KG+=O�T���ݦ��	Sy�I���O�OA̜	A.�F��颴��-���:شvz�8��?����?9�'��?�	�LC1`^L��A�-Hp�4�w�ϛ���J�w��b>��� `Ή�rG�&'��s���F�1��4�?���?�w��#׉��$�''���,.f2t֝6�rxb�l��~���'B�'�\�g~B�'��$�!I��[�,S�qvm+AlE�<��F�'#4c$R�������L��I��~u"��#�z�إ�A��ēL���<	�����O �S��iZ�AZ�j�(>��=�2�	?T�ʓ�?����'���O�(���7"��;�Ęm�*b�i�I��O��d�O���<Y�!R���ӊ,��:�iٔJ��Y��G	W��IٟT��u�	Yy�O�B�ݱ0�d�	M�0P|d� HN0[���?���?�*O�� WOⓌ"5j�Sc��N͚�a�=.�����4�?YM>+O�i�O��O�Z@�$g�&�� !���2>�Z�4�?�.OV�De,"�'�?�����N0�b��j�Z�1���=l�̐%���I_yҀˬ�O��9f������D����;hG��\�LSuDԵ�M�tT?���?�P�O��ʢ�U18ǌ��.ŵfJ-�M�*Ot�d�O@$>�&?7m�i� �'ة��<bR�R�k+�6b�� X�6��O����O&�	V\�i>MoڣT�F���#Y��X1���h���'���'1ɧ���h���цE�$`�L˺W3����
^.�M��?!��D���-O�Z���An�����t�z�C�>�f�Gx��(���O>���OE@%�ڞi�(ٱ��(�1:�
Ц]�	ߖ���O�ʓ�?q)O�����h�fN5I�B�z�ύ�Iv��+�i�B��y��'D2�'$��'�剔kG�U���mxx�Q�)Q�	�5��Y����<a����OH���O�͑�,$k�EC�/�<Y��#g��,e�	���	ޟ8�	y�d��k޾�S�p�@�SPmʵXGHP�Gϗ�|8�6��<1�����O����O(T(�>O���5F�q����@ʻ#���� � զ���П|�	Ο�'��H���~r����h��!ʍ0�(p�"��	��K��M�����O`��O�ԣ2O��D�O�(I_����
>�r( �)ǖ��7-�ON�D�<���Ԥ[Y����d�	�?=�Ł>|C��]7g�M���8����O��D�O�)�6O��O��S�B`�A:%��}>4 cf��47-�<ar�P�a����'j2�'d��c�>�;*Ϧ;b�Q&4�\�]�@�4,n���8���Y��	F�	]ܧ%�L�M�:= ��SOL���4}�zD���i���'"�O.����d�4-P�x��iC4\�ܰ���:�l��l���Yy��'e���k��3�@ ��tsU�N@���o�<��Пp�#����<����~b�=5�x�h&F5YB�-c1.��M�O>�g��<�O���'*Z� b�h5�U aT�8HwQM�aQ��i��������d�Oʓ�?�� @܁RFB��S�� ��#���*P�'�ᣞ'j����L��۟��'f"���
� �BI�f�2��X(�]
qG������O�ʓ�?���?	�#����}����"m����C�4�N���?���?A��?�(O:���(P�|b���+NP��a�9j @�IUƦ��'�2P���I�0���6���CL�))�g������
L3m��@�O���O��$�<�u�S7&��S֟,)G呲f��2�'�S�2�"�c߱�M[�����O��D�O"��4On�'2 ra�I"q}��Rg!�(SG�,)޴�?����D�д�O�2�'��E�Yﮁ����4� ��W'���?����?Ajc~�]���'H&��������=+�!ݚ5��Xlby��(�6��O ���O�	�Z}Zw�&b<��B�)̦e�l���B֊�M;���?�f
�<I����3��=�R`D�Ȼ`�r�Є凥@�H6 o�(m��@��ퟠ�;���<I�"BM0�
�dƻ:��H��Vw���h�����<���t�'�4�`�M0�� {`/3;�����sӒ�$�O��D	�|�0}�'���ʟ,�c��'AI<'�N!
Fj]�r�o�۟ �'��K�����O��$�O��Kv`��[����pc%��P������	lL[�O8˓�?.O:��Ƥy�E%��z�hY�����z�A�A\����Ee����Ο(������y���"0���BҢ(�|�sf��4VC�0
��>9,OD��<1���?�i��e ���RP���S!+�J��a���<���?a���?�����1�ͧLYP%�=3�L����<�>�l�hy��'���d�Iϟ��Ʊ~F��"L�h���C�'r@"�s��@æ��Iß��I��'��e�!��~j���7*ɜ)X����ۼY�A�W�릡��Oyr�'|��'>>��O��I�3���1'�-h���*Ǩ�"@7M�O��$�<)�͜��O���O��in�0=ѸA#t&�9t�.l�E�0���O���ٝ
����:���?���k�-7hp��9(�ݚ��l�~�=� ���i���'�?����I=P�68C��
*�94��yY5�i���'��r�'��'�q�$I���I�R X��"I6b�v�Bb�iN� �aӊ���O����-$�$�ɅM<P�����XP�d�#R�7��"ڴw��9������Ox2
ݝY�<XRhV�L��r��ئ���ǟ��ɮ+L� K<���?��'7��ЁP�/�f#�K�UT-�ڴ��g��|�S�$�'���'y� �Ǣ�DiٳCO ?j�� G|��Dӷz���>�����S7�,��lڷ!Α��L���v}be�y�V����Пx%?��ӭC;v.J��6�$3f�ԉ9�8���}b�'��'�r�':Zt�.ц ��!����Y������?��]�|�	ҟT��wy�(T�`��S�d��f��X���ø�,��P���	�t&���I��z-r��S��H�>��X� *�m�px�����Oj�$�O��Cj�A������O�={ڨx�$_D@ఊ��1?I�7M�O��O��d�Or��T?O�'�ШB����#�����'ܮl�ڴ�?Y���Q	bi�,'>e�I�?�B6Ӆ\b�|!���cΔ�����ē�?!��j�< �������K��dbe�
�]ZBiP���Mk+O&Ż �Y򦝡��0�d��l(�'r:�+�eѨu׎��R�nC��x�4�?���	,�?�I>��t��8�j��r.ԋr��iF�
��M��-}X�F�'h��'[�$`+���8Dt�2��ф41�5ka��3I,%`�4zg�Dϓ����O b�\�"�:庲�S�+o\	��dR���7-�Oʓj(���/O��?	�'r�����0[���蝫7�U��(��OF��'���n��hPS�+[$IQ@��:`�"7M�O�1�eeRd}"/�~���?�K�X V@Ǝ��	�jQ��X�1�d4���Ov�D�O���O�%��X�xU��F��1�Qg�4�>��?A��?yH>I���~�J�?V�F�ps�C��u�t�M0%	W~��'C�R���I1�"9��Z|ڨ0�m�o�p��ӆA��P�n�ٟ��I֟p$���	Vyr���M[��4Rt�q���z� A8� �|}b�'\��'�剢'ґ�H|
BB#d� pA�2!��C�!B�s�'>�'���Iof�<I#O�~��KO�z��7-�O���<�a��7Gm�O�2�Ovܔ��цg�![%��=�,Q���9�d�O��Ƅr����K�(٦�\�K. ���R�V8��m�SyR��WZ�6��O����O��ITZ}Zw���:�&˂E�2��!k�u��@ڴ�?Q�R�h�͓KB�s���}��C<j�F����S)�6���
Ӧ�aV\��M���?�����[�l�'#�����x�Zͳ�!.)��l�G�e����O��?y�I1p��y+B�H7j`h9��	i�r�!ܴ�?����?q���B��Iwy��'��՝*�.8�d�X�tt|i��ǣ>t�6�'���(x���)����?��*�Fm�Q�� ,��Sv�S���c�i0���7~2����$�OBʓ�?�10��xiFFQpӼey�b��;�Ɖl���Ky���'U�'�2R��#E��t�:p'ˊ8Pi8B흩�	S�O�˓�?�.O��d�O���A�d��|C$�8bU4�Z�m *8�8OF�d�O�d�O�D�<�գ[�>�� 
$*sb��s����c˫M�.�pS�im�	ܟ �'lb�'q"��*�y��ěs&8�PTm6	��Y����,��7��O����O�d�<�"�K�p����֘)B?����[�S0�����.��7��O^��?A���?�se��<�-Or�P�D\�xI�X0e�H�C�d���9�	ş�'I�Q"h�~z���?	�'<�>,��c�CX�Cpx��[���Iߟ��I-���	ȟ��	՟���A��b@h�uc�(@EJ"
ynZ^y�n��Rm6M�O��D�O��C}Zw������N��(i�R�h�Pܴ�?������?��?I���(ܭr�z!�^
tI�p�@�?ٔ���0g��
A����cH O1D��0�0D���r)?79�!@��)\��,Q���/�j��Sb�@d̢�,�^�)R�+5#�����'@ښ�!��%�:�V B�9��Z��#�@|
@@;b
�x#H�o��i����0|a��"G�-�Lp����-�0�J�B1v9Z@ �	�U����I.%ư0�2DT2_��e�D&�ܟ��ϟd�I��u'�'��5��K�EU���q{��	1͘M+R���83���1��S^�X0jմ<�AG~R�A��]�p+ڀI�`�˖FЍN���� ��=?��-�G�[�[IG�ę9� #=I7�޵1-j�z"ӵR���3(T*�b���⟘G{R���BA�����]�)\	(!�M���6�&"W���z�1OI�'��! G ��O@�$���.�蕞x%^%����%}
���O~�JP��OX��m>Mh�Ϛ�3���s�Y��~��?��� v�A�w���p �p<)��+1^`0�(�sy��L�]}��z�M�	����
�H.�x�Q��?I����	��t�JY�I�x�BQ���k�1Ot����6�V�ؒBݪ'R��J�Ka�!�D�I�s`P�g@&h��+	;f����|�@�'ӈ�� ί>����iH�f�����!�b@��%#�]P�b�6�j�$�O��r�B�%a"ʥ�~���|�-�D!.�LI���D>����>'�Kv*I( ���|���ɖ0:,δH�Ο*��tI&YP�<V �	ܟF�T�'}������zQtq��&� L`P@�	�'�Z`W�1iD��rV���	�ґ��;ҍ٧z��Y�G��f� 8���A.�M���?����Xe�3�?���?a�Ӽ;4�]!sAq� (T/H�r����Tm�%+�MF�p��/�1y4˲cҋbS��:��ϯ>����'�t�BvB�g�ɣ|�R虵 �3Iy��y�o��E�D��|~� ߌ�?�}�Iϟ �ɐ����fG�!M�L@$�8."M%� ��I�}/�uԂE�@�hٰ�fq3 �~���'ɧ�i�<�f
� GH�'�Z�޴�&L�"�J��Q�[��?����?���|
���?	�O���eg�0M�r g��%t�1���cv�7�'Q���䣐�0 �b�%<,�Pf�	rJJ1���'HH1	�_+Z�\EY��؊ D��5����?����?���D�O��X҃o�Gj�IP�c�f�)4g%D�LkF +�"�Y`/W�JJ	�!.�5�M;���������a�q�� �>�{���\!��?y-b�!g�:p��k6'A�!�$�@lHC���!0��I��S�T�!�$����� ㊰i�H��U	!�8-��@qN�-`j�:�M]�^�!��2H�fH��m ���&L4?!��Y�:�3��.U�,z�"��mT!��և��D�U;
qP"t��M�!�d�a"�r 2=�4ѫD1�!�D3Z�ȇ�N����7D��%�!���&$C��9&�P�tNP�CD
NG!��RO���p*��Ts�pW�A�`4!��9f갥�a!�)w�N 	�!ʏ+(!�䎂Xh��hp��P�/3y!�D�SK^��uƞ*&�2s��	,x!��a�L�t�P�l��ゟ��!��é6���4S�4���ǝ�$�!�Ę�[�8�R�A�L�\�� �A��!򤎷`n*T�& �Yk2!R�aԁ|�!�F+|M�d��:w^ P����%�!�$�;�d[b#N#2L*��*9l�!��D�uBr�q�	�#ScD�L�!򄅠M����G�U�N��	��M�!�ZnFT� &�hQ��!R�!�� �M2�K�Pk��i�o�c�^��C"O�t���ޢ�f0�g[�V���I�"O��: MZ�
�q�C�Bu�IB�"OR�6����Z�R�F$,V��d"O�d!��*ME
�J�7eENX�""O�+�ڧ'�]�%	�):l���"O�����0$���(7�̿�t�"O�ّ��ܰ�Y�" �P��چ"O.��4���ѭ�'A�  ��v�<a�CV?U��ZS+�Z��6�g�<�d[$p�tA�
��G$���	c�<��C���@}����3��93$Mu�<)3f�S���"� 	$r���%[r�<b���(�
A�ƀ�b3b!�tnk�<Q���:,�M��慔;Ŏ�Y��i�<�Ɋ.��kq��|&c��Wz�<��	-s��s�ÊR���q�s�<y���}�vf�1#�^�jbH�c�<��d1B�x��$ޫVQ���'�i�<i%�ۑ �걨d�N'���c�MZK�<A1��2W��h�U)L<]�����K�Q�<A�ܑW%��f��F	0�FS��yR��+=M�A�W�_8�|�ħ��y�HY�v�H���اb�j5yt�ٍ�y��)"��yw-NR�NL�ҥ�y�ƞ'1	�I�9*���+�y�KʅH��̑�%'B�"��O��yM�{�Ptkt!ЩHN@�5@+�y�e\��Mڵ�F��3�'P�y
T; �p�� �ǳrW�q��2�y"H� 330u�D�S;d����E��y�A2FҺ	rK�%WRЌ�e���y"��#j��l��IKo�`bi���y�I�4a����Ɯ��-�&EӢ�y�6,� ��f�`d	ֆ_��y"R�q�@f���尕(�	�y�-�%��1J���s�`��ȓh�xe�N�g�j�ضk];rЅ���$��N��ղ#f͑x����R-�F�B%�䙓t��<�� ��h�E�1
�b���:��5�ȓU4L��bƝJg*��@Ɋ-�P���0���i���F�����M�9F�Їȓ{ ����I�j֐����V�`��nD,)#hF51((�2��ʁ"^Q��h�p<�c`ʲp���14jT�kZ���c��Qg�҃)�r}1�׼5��ȓ����Ҍ`|�D)�e0���ȓ\lX�s�m�Y�P�д���t��?a�㓬��?M��i�N���q,�2�Z�
�#D���So�J�n��S!ٻ@�$=)"��8�ư�ܴVr:;�O��g�'K�ܙ��$�t50䮛�Aɢ ��`Y ��V#fD��E��=�$��PD�6����I�KW�����'tJ�q���S���A;3}�=�M�<0��
�z�x�WUF � uB�Cv0�"禮|�BA�'�e!�%�6])D� #.Pj�<��J
̠ !��_�y��JSI\�h�"�(V�����m���B�t	p���'0����Owk�0X@�;���^ۨi��MΨ�xrg� <tQ�Tf"P\@��s��9�V `��	�.��A�	,Y���d`}�	J�p�z���|�$��g@uc 㐔g_N�9�B'�0<9�1|O4�t��t���(�E�)N��P�RgMGRhEC���4Ӓ � g�>��+0?��9O��'Q�[r��BO�MT��C���z5�<u��	E�_t���+A��r�������h֚9'0;Q���j�h�WA:(,��3�B��xb��9X��8�ذm�����	�T�����º���2��T�c��;P��xgٲiC(�ԧ�[Wř�'<9qIR�_a����U<YQɁw�? �<:�-�f�adf�;5�6��Ց)���Fe�/"�V��`!���6.�n115�:��$=��`��MԬ*�>�	B.��(�ax��b�T��W 9�Er������P@f�ԥ1jrk �hz"�x�ey���<9Ó.�t��F��}�x�t�Y�|���'�z���R9�MHщ��a�	�R��8O��T����p��s����G��#�"O��7�M�O�|�1B�ǳD�m2�G֛�Z����G;c��<J6��6��O�=H2��V}R��m\�ٹ��Q0;F�)���?�$���G�e����jA
��MA�>��I"CTi�����0XuY��_�d�DdG~r�)Ҹ"Pc�xx�u�	�Q���&�Y*7�ꍲ��bn��U�뛴`��\���T'p�aY1�uN��
���%|�a�U�В�.�0!DE�3�G���Dފmք~5bD�`�W�a4d��"Da�o���M�{Y2�)vЄ&�C�	�`̀�)�$�r#���E�/*~l��ؾr�2"3�i����Gɗ]��:Z}���+OBA�d��~:8�1U�6vs>�2
O��	��@�5��#%U>�B���(���T���<PV�z��Ó3�����Y�{ڦ$��v���I�;Z�,��6��9�:�AXFoP/���`*R<�'g!�43c��|z�1:0&؎eL8	w'-�	3���K�Ĝ�SL��c���xܧH[Ε:ġ�(>�,5A�	V�t���ȓi��);V)�M�����Q�>Fd��2���#¡�d,>��D4�g?qQeB�Dq�4H2��O٢	)��N�<)��0���k�W[�U�Q��<�e��0ax�I���<9�A)=c�߿�rXQaK�gX�䲦ʆ<�:i�a���Ip��Kq*@�-Q��y��ހ��%y@g]9EP��aR&�"O���J$�'���;��H��� �PhC�v�p��
����K8p�YrFn̶V%��ȓaF�Xc��U0 �$<���/O���ȓ'�L����;C"���
ѵ�(Q��!�Np#r�D�\Aޜ�6MV�=��ȓ~8�pa4�ʺ+�&X�E�ŉlhL��H��y�Z�(�D�Ӡ�P�Z��E�~����?e `����b��]�ȓ/��1�´M���b�%�
D���|�M���'��ݐQ�V[
�ʤlW%�fu����y`�8�y�%�,H���lÉE�(�6�م�y�
ϤI%^���h_�7a̪�"��(O�P�A
Φ͈�$dX��Ɠ[�98t%Q�J���"O��$fߟ'mp���nY�N컇nX(Dj��9R���O��
b+�(rN����'Q2'�>x��"O(H{tiN<1���%`��@lZdR��᭏,�0>Ѡf�%�,)�em�= �`��$�G�<� �f��x3� �5�ّ��@�<���̟N��8�%�zi�Ap)�B�<����:;Knh��A�4G|�P�$�B�<��a��3��H2e*J� �#4b�@�<�@� ~8���2l��UR`�o	W�<���
%�d�t�� ���NT�<Y���;9&�|+Ď% i� ����M�<�`I�j)�I2qH�*�Z�Q) H�<�t(��!Ą�,b��L��G�<�I[�n��Pr� u5^��VC�~�<��!� �j��t��I/����b�<	���).�8��$Yp�Bԛ���[�<�v.N)cT�u#X]�FT;���S�<q��%�p�*O4.U�IӁ��f�<�����FM�% �~�� C5([^�<���Y����d5:� ���S�<yҩ�3��q��ذ,�`bg�Z�<�ƃ&|��&IvF�`�O�V�<aƭ��.�&XXt��S�H}J��X�<y�-�9c4��!"��=TV.�8#J�<���]�d$Yq�OO�g��M���DC�<u�0%�֡���zR��I����<� N���I,��z�E��b �2�"O��4eHs��`��%C�	y�"OT���(��ɱ�/׈ā9k�"O� ˀ'x� ��͕*�˵"OhȈ&�͑ \��P��9"OXMz�NX5
���Y�� )�b�x�"O}�&�/C-�I@k�%�|y�4"OvZ���lH�́S�C@���+�"O6�x �E&Xl�0�4H�<��]k�"O&ESF���Ib��g	�qFh�{!"On�1�F�$�\�Ȑ�ú:=���v"OԤCH
�Jv�T#%�9q"O�T	��(��	��'O�i��iqf"OB�ԽL�N�:���"�"B"Ol�%,��Nd���jA%}��"O��]2��1�A:���#�σ�y"-�3�*�I�ɕ1/�(Đd���y�ġ��JW/�qB�M�cA?�y���"Fx-kF�X� ,�g�4�y"bZ�T��#e���C`l�J��ǒ�y��ϴC�nwA�6S����G�
�yrO��8.2�C.KL���v���y�,N6,t�y�2i5o����'��'�y���-�0Z,��g	�˓��y�k�a�Q�&�N�w&�UV��]�ȓe7,��SQE�;��'s��?�*�Q�/�& +&�Z`K�H���ȓL�x�q��Ăx�!�2N�<]�ȓ�����B�H�ł4�ٮ��L��D�I���XA:�r�2^8a��-�Z����6jj�Z�) ,x��\�ȓ/�u�b��CI��l��[7��2t�eJw��f�~I[� �1�n]��Z�4]؆�ʓl/�Bv$_�#ŀ4�ȓ���"P4�آ��̗E���ȓTz$�1�"�"v(�Z��:=&ĄȓI�����ڧe�}:T�T$��I��V- A�˔;hI����F��\Q�M�ȓL����Zu�\R�!Ĵ)�d��ȓ.����1f�'0�j�h�&_��2`�ȓ^b��0���,��jѬK����/ �(���H�
�b���)Ѭt�Їȓr��	D匳i�h�h��\�V�X��HT�0��
m�Af \|�E��'�(����[9(MX�h�$0�
�ȓ  ��¢��6�|���Z�T��Ɇ�=0�Xe0T�z�*��ŔwHNԆ�,��3)V���	�$�Z
%d��� �p������nivp�,�%¤��	�t�0�jN��9�tC۠��H��A�	1"�,�@L3@I�e�d�ȓ:��[РH8v� �֯��	����k񎭻á kb��!@�D�Td1�ȓL�R͘D��1
�i�`��W����M�~(�	��BD�
EoV�)*���2�&,�l\V���n��4��dq��� Ied8�7�G�-2X)��i�D�r�bX�F]���`ߜE���Bc�E������>%�C��3��`��!�6љ��2R��8 �X�p�؍��=�$,BEȆ�[1�4�'*^�9�ʥ�ȓ%+&<��Ş3Ԑ�H1'�*n8<̇ȓ4	@A�UA�%^*tA`�n�* b�|��n�.�I013��3�!$-�\��S�? ��Z��_-�Ұ��ΐ#R��ݣ�"Od�{�CT�/d��2���'r�8��"O~)i���>-mE���%W�!�""O��k��L��!ȧ'�`=��pq"O�`�%�G��"̲T��%{��!�"O�0�pM0�2Y� mz�p�%"Of%@a�A�r+�ÑnrF1#�"OԍW��-|�� (��&n|ꩣ�"Ov|R�V�?�5�ś6Fn��q�"Of (w�٤m��C��<iF�W"Oj��`�q�ѡ"�T �@"Of�+SoF j��T!���<%[�"O��
��0z	�k��+32	��"O���4M��d�	�4u��t"O��
7M̿��He�'�@�"O,ň dU��XU��q��%��"O�����*{It��)����B7"O��We҉!�||[�H\	f��p�"O��p�#ߛ:���I曇�Rex�"O�d� UǊ=�&��p�Q`"O� ҧ�n�$TZ�W,,�]��"OL}��琉!���`*F8ڢ$3�"O�́��أo�E�p	X�N*��Ct"O��P�,�|��'D�>�`!"Ol!j��T�I%(��M�X��P�"O�`�ǆ*���B�T�u�kF"Oƽ�R��\i�QX��Ai�}�P"O�a�Ꮭ�bF�kh��aM��s�"OvDaG���2��Я�++����
`�<9���/��|#�/N1M� I �F�<7%'R�Z"E2[�h�Gc
F�<�§LA ���e�`~(B�@�<��-M�@DT0R��F,mH	
�f�x�<��E�1B0�e��Ą�v ���Z�<��`�46�,��U��1����7�N@�<i�*G=iNv=���U-H� ���f�<��%Y;=��!u���~ ##f^�<Y�jԒ.�@(�R��]��u[���\�<�G�ƃIy��� �� ORm�Ҥ�X�<92a\�%����r㞞�M��B���yR�P:���gF�.����HH��y�I��]�ՋY6"�$�Q���y����nT!�B����8� �fG��y"lY�eJ��c�����eHA��y�]���m�z�D�s�� �y2��68WJ�gOӀt�t������y�'�e`��� �W�d�FAY� Ӟ�y��
4mǲH� �۠����y"@Ň_���Tkβ�LiZ�C!�ybB�-�E��b�n��,�=�y��	�F�ZP���	�il��z����y�C�ii�Dx�OZv|�����y��ݍ}�|ZR���Q�D�yb��	)��`R
J[Q�-SC���y-�*<V�+�-�OՖ���L��y�b�4]{$,Y;s��,�ĪQ(�y"
 *����0dz�\�%I���y��,��(��j�(@,����ܛ�yM�3����F̾C(�f���y��T�c<Pr6k��eJշ�y""��u@L Ȅ��#���҃l���y2�R�.#F�Y���,6p9#����yRe�2<P��-��:84X8nT��y�oc���0�ݱ*5&R`�	���p>�  ��Ơ�(����Fݵ�m�"O����ݶ>!`��c�K
~
<��T"O�ahP�_I�� +�
�Z%��"OBE�t'��U�ء�OM�
�<H3�"O��B�ٌw�,в���	10h��i)���Z�9q>��@�}c�ူBV! �!��nW"�Ԯ��4U���䡊��!��R�Y��mz�Z@T�]���a!�D�)ô�@�f�18I,d�с�+p!��+�إ��a9�Pp��7DT!�D;P�0�A�_�^t�`��5:!�$��~���ZU�܄��A�یY!���*�
��E	�9�tt�%��o|!��Śc>�I�4��h��S2�=a_!�dO%�daE�)����c�7[!����Xe��&C�vt�a�\�1�!�dW�<UD\����EYʸБLW�]o!��:>m0�a�*�aM�1EL �f!�H�G.�+Ѝ,X~�QFŒ�:_!�$�2�m!� �".��QJ7!�!��'J�h�c0����XB��RA�!��oTę����&Vhͪ�Ə4e�!�d��0!�w �^��˷��!� �������L�V�%hϽk�!�O�xA�ݛU�^t~رs7��*�!�d�R��q��S=my�c�(�5E!��Âkb���g9N
�� �g}!��E8��	�ib ���u�!�d�TH!����)Abĝ+"�Ă�!�d_�5Y(�Y���DxT�x�݀,w!��S�@#��x��܉f�iP�-92�!�$��_����@eN�%���S�!򤚈�8M�W�=5Yr�#�0�!�䕧z��-���I {10}�#B��!�d	*`�*�ڱ�ȑ��*��ۧ^m!�$��2v%2�V,�l�QP�C8V�!�O>I�t|I.\�h¶NƼ�!�d���]:��D��6.F�:0m�[�<aנ�3^ؑ��m��^sX8iB�O�<����,���������I�T��I�<ߡ5<�����4S�����E�<�t�Ǽ#8D3��U�d��8�L�}�<)�L��:��1/�z�|��WI�x�<��S7	6�K1-FV����v�<�#�6Ux�"���9���Yg��B�	2(�Y 0l��EL����* �g�LB�I��[r)�^��zV%�w%B��)I�x�kA"�s��W�<0B䉇8հ|0w��9y���s�ȬB8�B�� u��qЯ�(z/� �'� {�B�I�{���ʔc���Q�A|9�C�I9fҀdBV���b(���
RB�v\�d��L�-1�!��/�)$]&B�I3R*�j�n�-(����sD�,V"<iϓ:�P�+�N������^�C��i��g�㤉V�Qt�P��gZ� 2>��ȓpU@@o�9�(���ړl?6܇ȓma���	�M��IZ;Ygt��C���	UӾ�b�0�A��kXX�ȓZr�)��kN�oRp���e�/ �*e��	k�'���a���:|��]���k�d��"Ol�����H��0�ʵi��Xxr"Odݚ�a�g�)r5dR<P�d�"O4 )��X{v���E�|с2"O� �M֋�?0@�9��Ц=�|�jC"Oh-ٶ�B�aFa�ᅼP�����"OH�ɕB��y/���f!�szP\�"O
���N�S3N�9AϯA!1"Oxa�f�y�ܔIt ��O�=��"O�{��� H��A��:%vej"O�Q�r���
���9Gϑ.r����"O�1S�	�+��;��XK���J�"O�p��G�]z,)���l�R���"O���Z >�ب�D C;M;=��"OBQ�S�߃~e� <*���"Ot�*�%I0:V<)�QČ(l��t"O<�; ]*E�AQCc�b�d� �"O�����^�~|b�@����`�4"Ob����7��m�'�v��Y �"O.yE��S�8��w��K��9C'"O�@"��ַ�ң"�-Y��4 �"OF8��-G�x�0M�p���1�ʍ`�"ON�Y2�ӿ:7�LzFb�n�6L{�"OR%����&v�xDcLQ#tJ���"O0<J��8Z��=Y���@h����"O�ɋ���.~����*��#nڬ�"O�M:�Q&yt��"'��Q 8 �"O�kSk�z�Z2-VcZ��#"O��2.H5.t��E�8I���q"OD�D%�e�D�aR���b<K4"Ot�"�� Vh9k$䅡v�ٚQ"O��c�T"M�4hu�����l3"ODj��S�*�X1�⓾5���V"O8��D�B�h���`}�.���"O8h�F�Ʃ5��AM��5@({'"Ol��G/�0N�T���N�E �40w"O��Q��w.��酨
�٨�"O�q��mR;J�8����4o�Ls"O D��QE��i�kP�[�m��"O��#�!����)I�O0X�ش"O�6#^���ޚ<NEҤÍ�3!�ĕ�@^��)G#�,,�	����'���aD'B�����	?aZH��'/*�@�l�l3�h��ٱ2g<t��'*�a3�,P$?"T�Ud�?10����'� �K�`Pþ<�QK�t���J�'�Ta30g��^3:���a���i�'������8�-��L:1%@�I	�'�|�c���0~��S�&S.Y0���'*��M��y.��auG�0�A��'�\�ł{ӒĚ5L�=}�c�'�*�I��B�5H&�z�� 4O}��
�'����*�?h&Y�s�Z�@*X�!
�' ։zQ��{�\�zC�ɇ0-���	�'�ᒻ�!��Ĥ(�p,k���yRàf�(|�3��N�SO���y2&�2��5&D�?�K�.���yҢS5v�j�K`n:Rra6 A��y��2��آ#�F��u'̎�yၣ5B{wM�1Q�B�n�6�y"#�s)��r#�D)���TƋ��yrFM�	��M����eɊ�y��"��� �`����yւ	�y�o��a�ð�L8�Τ{D�Q��y���Iup�+�	��6��9�F 	��y�K��	r�y�`(�(r 9�f���y�g��Mm���)תl�"���.�y,Xm!d؀NR$r/������y
� J�8I��Z�xE������k�"O
m"FL$[�L�B�ΉO|�\�!"O�:PDP%��� Ͽ�
���"O�$�%B�A@UC$"y��4"Oգ��E�x�z�{���=Vb,8("Oxt�i��D��Q�k�:|Qv�*�"O��G�e
��Zk��!Jn�Rp"O@��'�\�vyr9����04���"O���QM�$4�Y�&U�1��"O ����Y%BB���� �.$�P�"O���"���
�]" ��y�Zݳ�"O�]+��*��`��W�i����s"O*�k��ۋB�X���甛W�� �"O����Çz^
���E�u�^��"O2� �A�ȒH���8��!��"O<��⋘�a!n,��m�)�l�C"O��ĭB�:��$��b��4i�"O�U�T[]�-�o�-�m��"O���R!K<[x��sg.Q	�<
�"O�$XR�3tvx� 7+�8F�"�0'"O��NgU�����1&�܍h�"O*T{ ✀F-@�d�64@�1�"Ov�k��X��0���8Kf���"O�bjEsBm�%K���p�U"O��V��^�6��%���O�<LZ"O�u C�˞oa��/�,-ovсw"O*)0d"!2~z�#��"Qe�@��"Ob�2��L��D
>Y���E"O^D�Wk_�Z`P�;R%WRVf�H�"O��3c�P㖁��D(|1���"O��0��@�V���bX	:��C&"OVI����u�����!�Aװ�d"O���b�?8��E���Tʹ<��"O�hJ5��5. e�7 E�U���d"O�Dr�K+���-P3i���ӱ"O>	�uĞ(5a�K��s�z%��"O��1\&9�,p9���=o���e"O�4��$.]��U��DP�{���+�"O
q��l��P�ԀK��$OV�M�<i�'צ=t� YF`�X����L�<Ab��30t���-\�+��kp��m�<����J�N� �h�3j�؈��Fh�<)�-�<E-BH����Ch�ɻ��a�<��)�#��u�IZ�3� K#�E�<1D�A�,���4�p��\����<�1�Ӻ9��C�N��h�^��R�x�<Q���r̶Ɋc��vB����Lu�<1�I�u��"ʔ�� �Ik�<�2M�m>�l����,�XgO�<�p'�F�� P�3��Ñ,�K�<�'L�JZ��p�NS�!}B��1GIl�<Y��Y�L}>��a��",�j��!+V�<��_�>&�0�
�%S��kF�[~�<�2���*r�b���mh����I f�<w`�(o��9Rp��'� %��Lv�<I�cȶC��
�&M ���b�ğZ�<��h�92Nu�ፉ6<9�s��V�<q�ǈ�^�!'#D*?����3 �S�<y�b.s\f��`�ӻ#���Hd��L�<Y&H�E��s��9����FJ�<�3d�
%��I.�_���$ I�<��nW���a��T�EB�ı� G�<����0��	��@(c�Kn�}�<��M��Ar�Y�2mM�
|b0:��q�<� �<�1�E�20(p'�@�G[¬��"O����b^n��s��=K��3�"O���aK Q�v�J�b�i%f]�U"O��0���5 �F���Sw�pX�"O@+��Ќ?�$�0���ke��v"O���qm\�C�����/�[a��C�"O�d��Kηf<�bvn�;u<kt"O ����#ea�m	���b��8�S"OȄ��MZ,&X [a�U��A�"O ��� M�s`���	�?�ڍ��"O����
ё;��
�+׋�Z�bC"O��C����B��[�5��ڥ"O���񆘺a$��'�ǘ4�`%�"OЭR�M;�
�ң ��I���"OF@���J3�$�I���(s"O��c��RG ~��R胢� �v"O�X���<u����7��ʜ�� "O���Gە����GVS�H�+%"OB�x׏�5i���D�Q�@��E�$"OL,9�m0$5�a��]rG�)D��S��B1M���F�D)��.%D��H0bX$`i��c�T
��E->D����d��~���F:p��P)�7D����#�/��9��$ܣ��8#�8D���C��k|��	Y�,�X,1 8D���d&U9:�н�Ə��YD$pe�2D��@�(��/����(W�3x6X(&�=D�$k"�@�����)Ѽ�j�K�B<D��k��"fO�<�r�B�Vq�y��E:D�(�ŀ�6,����R��,R���2D�X�F* 9c���E�^�R�h1D� ��ʽ!X�%_�V_�=��)-D�К�h�:%ΚP�ٯ��Rb,D��s�!I�a:<ͳS�X	R� ��'D�X��BXX&�HC�W����� D� *�d�.�NY1�� �����-0D� А�7]��@	�n�I��m-D�H1��Τ{5�e��l��A�x}�q�,D�XJr �?b~Fx�� �-��-؀/8D�x/=+��#u�سv�
`5l�)|�!�ۛm���\�Y���:�^�2�!�$��}^,*l
)�Q�dX��!�"�D���+$�*�LV�W�!��%+,h-��N�+|"���� �!�d�%l=̱�F���d�!��&�!�$�-6���#���#H�h�F�e!�$B2K>@G�Y�d<Y���?�!���qx�TH�+ģ������I7݄��&�ї��Ⰵ�Ҡ�(]���b!��ZS�R,x�8���D�x4T���v��qs��5}P������ȓ�N1{
܂E�xyILu���ȓE��[�� "5�� 无���6%J�f-X�%�h| !,\���y�̱��J�Ml����&E3�x��W��=i��S�5NTh�"P�g�4�ȓ
jq�wFBku�E� %�*h�ȓ$�8�*$͞�wtΡ�R+�'��X��r�a*t�ʈry\ݨ%�T3����B�(sE[�[u\Y�.N���ȓr%��3OĄ>�ٸf�Ũ-�|�ȓ"z��a�5/Q�r&�*yT�@����<�#e��N�PN���(�EI ~�<�AX�?�MP��ͷ�`�Z�@Lx�<�  	��^�dr�x�/يL́�@"O4�C�!G�����@�
��"O)!�JtB:�y.2ޒ�D"O��"�
6XXd,`@.��$� �z"O��"�<h�dQ�퉶���w"O���8l�bI6�\!R�"Ĳw"O�"�mX!]ָYp�V:� �Hd"O�a� Ȼ3�ldnڻ�8�+r�9D���4-iBTZ4�S*̕��8D�Ӷ��q�H[pB1�� �5D��C$�·(����D�DԌ|J��?D���ˈh�4s5A5L�N�{��"D�Hi���vmN�2�G*"D�!�K�%w��z�"M:)Z����3D��K3+WU;h��A �UB��p$3D��cR��3(�LY��M�',���C%`0D��qo�/b0���.����j8D��Ќ��]�*���)ǫ4Z}�3c8D��7��5k^0�����(mJ�{s�5D�Li� �+`~^:E��K~�PT�4D�����/: �"e��H���y2�	�1@9  �:A��aW����y�	R6hW�!����i�hq�����y�H�jP�P�.��d�25"#ݴ�yҩA� ��a[�)�Z �$�%5�y��B:w�ƙ�`l �]� � 4F��y2`�W��M�Hζ'�.�	S���y�'��-���*6�%jZ�C�gT��y������!U�X$�NŹ�O��y�Q'i���q������y+ �y�C+`+��z�B9ιk@�J-�y�!h�f���Im��O��y���!�u�6�_�)�
���y"��v���'��/Ң�Rڻ�y�O�J,��ID�|��8�K�.�yBm�5�H���������9�ybO3,ܞ��"�V�ݲ������yB�֎G��s4�7}cNa���4�y��8-�\�1�N�q�j�sN7�y�΁/Uܴ�P�G��U�`z���y/֊2 ��DA
K+≻n�!�y���i���M�m�]@k���y�`C6-��ܯr_8<I���yү
({�lH�E2p[8�����yRE��o�V�R�g=v�D�d"ڝ�y�ś�v`��v!�*�t}DZ��yd�-y/����33����
��y«�;J̮,�t��+�޽ �A� �y��&�,rg��m��`ccCɸ�yr��,>�ƨáN�Y��[�L���y���,
OB|AGC�P��a`�
���y�)�=1NM�e�Ñ3�H�B��_��yr�Z}����f��&����A@���Pyb�X �Vd�w�r[��G�<��hV�L=��R
 �V�H!g�J�<i��K�� � 
�uZ���I��O֮:T$�� �K0,*��݇�9v����C�&e���7��,,X�����#�ڼD\� X��lB�ԇ�S%�A�K�3"�-{�D��J����I[~ҭ܋{R�'��2^��P[s���yb�~#0�̸j@Y�'���y�#B6����E��4�qAB
ѿ�y�@
/��k���pA;�I�!�y
� D�p$�=+D�ʀD_�O:M҆"Ob�Xdf�;"���'Ɣ_R|�"Oj�Цh���p�A�Z����D"O���SE�z�:aF��(
��d�IZ�O{l�X�
��N� ؚv]�v���'��@��o�.5�B5��N�Z`�<��'4����*EX0�v��Yf(Ⱥ�'2�ċC\ߚ��TC��S����'��p*Dvl�<�Ƒ�9�����'`���JI�dB�.F]i�H�'���2/D.��9P�F3�h�p�'���s�.��L��"E턽E��(	�'\�$�ɕ��ܲSI��<��)��'�� X�-��y�Q��ٝ<��u�
�'�l��*ښn��D;��?-����'EX�`ٻ+wvɻ��ѭ,= ���'Lҥ�#�/Fo����G'*����° -z��EBU6. J��d�c�!�D��	�i�@ӠY��eJ���7�!�däP�쬚��Df��Aےd�'�!�סJ.(t �ԏ���YT�\5�!��ɫQ"�u▉<n���䀔x!��U�f��l���6}�liפ�r!�&4����*�8T��{��bp�}��'{�\�$���.��^;������2i�!�ğ�\:<�hn��3��bS�X�J�!���3T����$�~0:|:��\�!�Č$)[�mJÛ�t����
Pl!���_jB�nÂ.r`�Bd���|6!��Fy���HTm��pL*�PF.��8!�ď:3�����D	��iR ��?�!��(��ᘰ�?/͌0c�.r�!�Ą�P,��U���A�
�!�d	pi���u���0�����@,�!�dӔ<�h��&�	�zt
���!�DY�>�yCT�";�*�۷jJ �!�	q�`�qƣQf��R��Y7!���9O�:���d}}n���(��!��[���ȀnZ
e�s0*�2!�(L�t�/��>L�q����!q�!���p�M�P�ǽDe:�"K�Y�!�
R^D�T+P�H]�� P�!�$��I?��Y�L�,),P�Fږ9�!��W�Ҥ�'�)t�<`����HG!򤂛H��9Ӄ��xbdD[��;B!��Пp��8wl���ɦ���9O�*WIC�6d����k��a`"O:X�� ��C��� c�?⸙��"O��T��8��g��d�F�/�y"���	�`4�a:�N�ԋ�/�yR�T`��h'��!7h �
��y2ϓ�Βxb�P�^`��m��y���	��ģ��=\J��1�A���y"DS���=����CHDC�	��y�F��C"�ZAf�??S�-� /�
�yo2`_��¥AI�v�� oҟ�y"�վ=�:�x2���>v�ZcnM6�y�k��@�ly`�# :����2A���y�ܝ1���P*N�/��S��*�y�L�
�(����'ҮeJ"� D�$���̦oJ� "Ç�Dm���uC<D�Ȅ)M�X�j�E���}�Ȓ�4D����A��e
�C!e��qBy��/D����`F?`�H ���!���$l!D�� X�CR��C�pX�1O���lhR"OfQ �N��80�MS�;��,�F"O(x�!�!X�ᙑ�^�<�V�9b"O�H���Z(~���,�]4�P"OL��VL�SԚ�:Dk�xްP�"O*��#V5_���au逤/j�2�"OrP��"�'��@��5v�j�"OZer�ëB�d�9�lĘE��(��"O��	C�M*N�Fd�kT�
��"O©�E�J��9��L�r7�D8LO�e9S.��^L��"o2rJ�%��"O�svi���j��v���:4T:�"O��	D�����Ù�G0Ҹ�"O�� �D�E�|�bA�jث�"O~��r%�:j#l�4��?>!Ne�Q"O�ث��_*N�bl�����"OPy�� ���*v��i%
iY@"O�[ �*��c�>+��I�"O�ux��ɐ*�8��f��A�6Iq�"O���)B8���r���Тq"O���E��`��9�pG�"��	�"O I�q/��O&�11����\bD�t"O2@k�Jվ4���Z'�<{M���"OZI�p'_�ywLy���L�:Q�HS��|r�'-�9�%���k�,`�EAߖ��Q[�'dZ�'��<>#�i �((�.=Q�'�JÒg��0����- �h;U($�|��'�ND����"G��^�H��'i(�)�8y�}�&g]+ ��hr�'Mv�r#OF�l�qG��Di$��'��t��I�
�90���C&����'�D
t���лc���7��]:�'@�U��,���1�I�)4�t��'���Jbl��<熡�d�4_Y�ExK>1�8X��coÏS��	�"�A�|u�ȓYk8e�0�����ȋ�C�5�ȓ4� �q�斬\��
�D�P��ȓF�|���-ÞV���2QOS�
���%��3�eԜ���@�+] ��ȓ(��eB/-�L�"@Ƞ �f݅ȓu"���K�>20rP��q�|���V)�4��-��$����-|� ��ȓ=]:��iT=R�*A���&d�V��ȓ+)�)��٤?�$���a *�����c�@�Z���2|h͂%卞J��1�	����bu��뗵H�H'.Ѩ �t�k�'.D���VŖ��'�= p�IA�&D���'��8ޢt�&��!)810m%D�̉��ĬqF��'n��z�%D��3��P:���S�F�
 �)��("D���
�	_�� ��$0ش(��>D���1$�<%N��B�8Yt8
�n<D��6�@�#��|8��j
dD�W�;D�����L<5����4'����4D��sb��|�� q�b�tc��6��?)���O֢�!� ����� ��PB�'��		�!��Q'�y�p�@�x!Y�'��ⵡJ�":��b�˰P@��P�'�X��J!����I�T,1�'�	0!$��\�ve��EG�>|v�p�'->Q����ep4�����BfT���'��yJ��o�j��oF�6�����d5�B��xCc��~�ĉ��N8�(��ȓh�� f��8i��QIW�B6E$���S�? z��adۛo��@�#�&��y"O�xGE�6:��Є��\���9LO&�����USBd��ճS����1"O�R���%�����=\���"O�䑁/��'����-	��Z�A�����o�')�H��D�۵qI�l�D��0E��ńȓ4��!PC��
	��#����X�m��er��'Z�}��p�p/S�B,��lz�x�#W�M)�b'��$P*�܇�O`���eL�30�CƩ�!CF�Ї�ybU0���$:���#bI l�}��@�4��T2�`Sc��C�ҭ$�F{��*�Р�pu_+^q��*��yr��>O�qPa�ٞRy\�`U�X
�yə	�:���
]�AV����E��y2��Zx
��p�(p=�(Q���y���F�ё�;MT���b	��y�$Э!=�������3�2�*j��y�lH�fH�R���=��5���y҉�.�0(jQF�2�vݪ@����y�Ɂ��D�3�^7.*�� ���y��PaEX4�� %�6l�b�܉�yB�� :r�S2�2�8!C�H��ybFX���B�c��flD�-�y2��8Du*a�F�ij���w��y�D_ND$8��I�S�j�kֈ@��y"�׵[�Eq���I~�-��̤�yl�%<�̄kB,�B��0(����'���t(N�����i�:#O���ȓ'�����Kfp04�@H̝A�0�E{��OcJ��$�6��0���F����	�'dB�3�O�/@�h�$��<����'�8��F�5Y�������~��a�'׶]S�@݇�nYa�ٯ�,���'3�@�3���lw(��F* 0Z��'Hi�޴G�U���$`>�8�'��ABBl��g4���r��g�� p
�'��pӮ�"m%�ib��d�J$��'�t�%OŊ�T!b�G.K�H���'\ ѩ�a�{�x-��Kβ=��ي�D3�[����˝>��2�(5�h���'�����N�L�=�t���p��ȓ�lUs�d��U��`����+i��ȓh,�����L!�X�`)��.��ȓBΝjg��D�l��e )�x��@��Bv�نs�U�D�D� �2m��<m����γ]�<����z &U��o�P�k�`������i_v �H��6�L���� v�S��ٙa+�0��1[а0�FS�]�c�oH�5��ԅȓV�
ؒ��ҥ1��9��ە-���	`�'���R#(�^zzuB�߹�x]B
�'�]�H���ZٙÑ�A�u�	�'�L�i�n@!T�&ea����Ի	�'3N];PE�P���QLB����	�'��
� (3�<Q豪V5{��l+	�'�x�H3لI^�A�ԇxNN���'Ѣ1�g+��{�мc�wH^<�	�'6���aT
H�a�(�{�&1I
�'8 %B��R�L82���q���	�'�|�+񢕂C�ay��_9V�y�	�'��A�*Y2g���C��O)S	�'(B��D� kdP��-�+�pR	�'~D�"�C��W1� P
0Ǯ�B	��� 4̓�G� ��!I���#%\�PE{��+'͢%�wH�� �"��t��z�!�T:N�"���#a늕1gʍ�3�!�Dطm��9p3éQn�	�v���\!�S{^@�fK\+0�i�c�\;9
!��Y�H�C�d��htC�6!���k�̀)t��4�h�c�D!��&qpvtjQ��N��#3��
9.�r2O���p�T�a���R����,u	`"O���7�גK�	�I���W"O�h���$Q��Qe�,�v�	�'�R5O�"�$C.��}�wƑA�0�s�"O=cC/�&i����OE�n���"OH��e^}�z|[�m�!�\9�5"O���2h�1Μ��%��Hƨ�Qc�'���|�X �Y�Z �;���{2!��
S����#�/>|х�V�!�d}2�$�2LM�  � �G倦y}џpD����2E� A� +Y�Lr#���yR@�4r�T�sf�8%�0�!DcV��y*PHmz��2(I+MPU3遡�ybgո_\<\2�
�f��1��O��yrˡrјr-S�	�Fi�Jʹ���hOq��y��	�/ḁ���F�j1n8{�"O 2��	"��P�fτ�F���'��8WE.�I���|�(�CkR�k�!�$��3� �↸^|l�F�Oe�!���2BΑʰ�V�j���	�^!�$��T4�W�Y�����hX�R!��(;R(�!Fz�.�Y���=!�d�&~����Ryм�z&]�!�
�z�0yhfȎ-�Q�9�!�L>J��a� ��NР�G��+,�!��X����Ŭ�.I:��4�!��8�4ݱ2E��OՌ S�$+x!�ݫfx��nOI�Δ�q)�	cr!򄆖T��Hʷυw0��rThFW!�DJJ%�$��Ïh&�R���TX!�L��I�`*$�p�"��Pyb�D�y���g+�,?x�]@�aD��y�ӷ'X`F��ڔ�`Ϥ�y⍖b��р�mQx�B�����y"�5�V��,�`��0�-
>��'�O�c�2��I�5�L ���f"�(77D�ʒ��hr��8$�H1�S�44��p�HG'z�R���W���Ԁ�p�<�0�/5aRC
O�D<����l�<�%�OH�����J[m�HY�I�N�<����1
ʘ`Y�Ɂ#��!���H�<���յw�z�i�R&8԰Xq#AI����<y�j<fH���ԐE��ŜY�<)U �t"�!���(N���HLX�<y��^4����@dHS���_�<1DD�^� 43�
�}ـ1K�ȟZ�<����C�2	6�0a�0[��+D�,���$J��R��[�4�Z�.D���Da�j>�3�M�7?�N�K� D��Z�H��8@���eԆ-<B"<D�TR��y��%�3)�$��Q�c9|O�b��&ȿ5��)Jb�ſ�x�+5��V�'U�ɥ�� ��j�cЀ�+�����DC�I���:7��"\a����!*\>C��2i��@�� RL��5�P�\��C�	z#��ҳ�_�[:Y��J���C�)� �r��G�Tu�VH{G��"O�p�v	G�v6,I�����q�θ�C"O�\��M+�: �
�~��sb�|��'��G{�\�Ҍ��f*�$i���6F�!��^9u�|�a�39�T� EM!��ݭ)��X�,O��<!#w䛈H^!�䂚p� ��e�]�x��UxF��!�$�Uf�d����'�ra #h��2O)��O�$�}hR(ӿ/H��!B"O�)�G�
|&�H
��
-�,�"O��v,��6hȔ�LG���k�"OB�R,�.�.a���8��}�s"On���G�"	u�5����3B@��t"O"�v��@�,US�f�q.�TKB"O�U�nݲ`q�q���� �"O~h�ħpfZ���. )��"O��$�W�j�Fui�Mǂ�f}��"O~@��
2Ak��Y3��"��Y�u"O�<�� &�2���̢y�H�"O"�h#�4�01�Aݛfmn���"Oj�C2#�8l�f�c�
T�g����IX>�cd���`�LX��A	���$D�`P�@&Nhji�iH�q,��rV!�D�O���>)�q�J3��ɵ�K51��? !�ĜP��X�o�Z�P���	Z$s�!�$��E1Z�
��'Ѳ�3�h�:5�!�(Cn��bB�� �L�%h̕9�!��ʖ&A�G�I�%� aȲ�Y��!��6d=�˔�>dG�ЉG��72ў��ቕYZ\b���p�`�����	"��=!
�',��Y�N�,(f/��p���}m
��!ϊ`���Dn��K����ȓ� U�w$�Ty��+�[�R��]��;2zX�K]���O!s���ȓE��A��X{�≺V�9O�Ňȓk߫�4{n�j!@��z��x�a�IC�s0Ă�A��0�o��S�Z����<Q�
g�����C�Phk@�;ݬm����<���)����b'U�DF���dC�I/ؒT�%�.&L`5��/A!bC�ɑ�؀��G�9+u2��/whB�ɋ�Ҡ@�z�\��f�P�7FB䉚t���w���V2��c�'v~B�4���cA�My� �C��|K��=��K]u3$T�6��&��|U�ȓk�V����(W.uA!(�(+$y�ȓ���Y'�;خq����OM셄ȓ�\�Q�-��p����$]�䕅ȓ<޴��N2L0����!1�<���*S��C�m�y�D!Yn��
�'�p�Zf���2�LD��Ė"mܚ	�'�	�1%8h���R�Z�hD���'pVl�FA�:r�d�q��J]��c�'�t}8s�½]���Iڀ0%��'��-G�\	��
<׎�'uN�2F��2M�a`r��"/�Db��:�'O�*�@��x��`�ͅ(0@8ͅ�?`�/�*p�2)+P�6���1Xv�����6I�L9*!�-QJ9�ȓ��̂�F���s��a>}��"O�x��G%舕����aL(��T"O  ���
�P�a��� eT��"O"0B�� ��m�o��Z�"O��p@�M�l�$@���M�Q{U"O� ��Q)��gL��pG�lE�`"O�<�"*F!1�]s�lH0QE�Y02�'�1O�li׮�<a�����˃�o*��ʰ"Oh9�eD�,F%ޑ��͘�(�=1"O�)��&��W^�a{��S*�s�"O��3� ��$E��ɒkΝN$����	G�Ob ��6H���TV0 �6�;
�'Nh��i�DTPɰ⨊3"��Y�	ϓ�O�4IF�C�"��i3��ר=�^-���|�'#``	�3Q�@|��.����'3$H��Ș�D�Ҥj� ��!�'��<�q��_(L�2�]Ya��'B�;���"13�D����%�N� 	�'��S1�K �^�� �="'�9x��!�$*j��n�!8��\|xt�#D{�ID�'=1Od|��i�2�~�I�oW8-J\EpT�FB��#�`��]2�B�!ƌ??$!�d���� ��j���D%�y!�dB�or��Q	�vL0[u��3!�dn�����&<o��a��ܵF!�$�E��y)�Y~mP��D��l�!��թg<��D��'^ UICn��N�!�$>O4�A�sOє�Ľ*�mT�8͡� 1E���$-���m	����y�����Hy�_u����`\�y�o�-$J�����ɵ�\��y2�5k"��4b��|#�U��F�.��>��O�aPm��&�����
�~�lY�"O��z��=[��=����h��b"OlLI�݅v���q#։OkN��"O�x����2@HT�5bU����"Od!͋�I>�Y"F�6���P�"O�E���rh�p��#T�2 Z�"OX(�炣==E��@B�yt��Ye"ODt:WO�y=�� �!	�@Xԉi@"O��Q7)����aΐ�d)�"O6t�t#φH6�p�՛6��X1�"O�p�ς�K�޽��D�a� l�3"Oj��1�I�iWZ�r!AI=`˺DaD"OI+�D,$��o�b�^=2�"Of욧o�)-��"�S,'�����"O`�Å�M%;
�}�wd�" �d�`"O\��f��pD�K��J�F���'�ў"~2�`_0yڜ��d*r(́� ���'�azrf��%�8��B�Ĕ~+���u�O��yRo��tx��3��o40��ӇO�y�'�8~��D-ŵd�.�j��j�	�'�X�Ȗ&JOE�aр�D82%jM>!���?��7v$��7���9�a�)oXI�ȓXY�Ԑ��x,j�Y�
R��F��_搅S'�Rz���pI��)�C䉆)���A�aܹCw-��$�B䉖s[��0�Z:O#�5(��	n0`C�I�U�
�3�Ԁ;�8�b�l�0��B�I�}��A��ȕ�JS4��odh��'e���H�D��z��P��N@�)OR����=���h�˗e���6bA�}��� q�	�@!qA@��]~nhI��6D����j�'G pHQJ�$7Zx�k/D��h�CI�O>��x4�H(��j�-D���뒌Yy��#�C3X5Н��J+D�d��k�(�R$� : �T����(D��9�Z3T�P�c!J�3�8I�"D�`�Ђ�Z�|�F�^�F��s�� D�� ,ѩddÄF3lQ*ao�y���d"O	�)Z6�9�v-SV��1�"O١�GjՒ�.8'����"O�<�3J	�$q�dB�G��p5J�"O��3%�Y�?���b�6�A�"O,���� >g���`��*y�Xkw"Oj���K��.�<�㄀�/U�`bb"OH��EN�f�L͙C�/-���"O�}��m�IK�+{��:����yr��.3!����X�x�}Q�+7�y��@�UԐ![b��� ��������y҂>Ċ<I��xi��K�%D��y".Ϯx�mcT�k���C$�р�yҀ׳O�<A��#p���o<��=��y �k�ɡ֢N(��-1�����?�S�Oa2�C�^�<��Q�G`ʃ�f�
�'X�葂K�
Xl�RתQ%�@
�'�@ $?�j�Ag!��v�ހH	�'�Fd�1�
p�9�6�o�J`
�'n��0Nۣk8�xx���s��܇ʓp�����I���"�؅���CC�'�ў�G{��3FE�@)WÇ�.A`�%��|�ў��'p�|���\�u�,�Y�íaA��3��6D����䛙9�0dS�KB�qfb���4D��r��˜���!f��v�p	�E2D�`H/ɤV����j!Jv��!$D��I&�ŨR�\�6�n~���n"D��C���H��	"���4#�Tq��/"��8�Sܧ��Iª��x�S��%U*^X��]�92�ʊ�"��S�@�}DX�ȓ�Z�9��2)I$0�`��L}�l�ȓ�N���ަ"�M	��֣9HƬ�ȓ��eǀ�@`	�"��9I�z��ȓ4���!#��H��� 'd�UP�-��u�'B��éߨvۊ�6��ZؒO�=�}J��6ux�y6����<�d��Z�<�P�.�&dȩ*�����Rn�<�r�϶A�X��գ<!0�ı��Ej�<YDo� ��14�V:�X�!ŀ~�<y��<;�5��15ܴ�zrMz�<��jI>�&Ah�Uhv�ʡ�MA�<�A�ՙ(�MKB�ͻ�#�w��0=���E3Z����
�@�A���p�<i�(�+I�!��F�	:�ĬQ�<�4��� m^8o~�ȑ�w�<�`HĹ|f|,��F��U��a$��I�<�r�0P�OD;�H�B�G�W�J�ȓ@�^��B=�V\�bE�gY�`��F�Y� �]U���`1��-8�P	/O.��?��'�rV΂?;F Pd�-L�Շ��m�'x̀هK�.+"*�j���TM��'i�!��b�~@�*��x�����'�>�I`��Ft�!'�Z! �b5��'���w�1#�~qŢU�wِ���'�=��	�8Q[Ĩ�$G>j���)�'W*�Z3��5OR��0�A�<<U�	�'�l8#Re
9�B� ��v�����D�O�"|�O�	�n11Bj	6�
@�q�<�u��7��m�Dڳ���� ��p�<Q�͖jт��*Y\rTbIj�<�҅ۃr�����@�*i"�m"�BNe�<�`��G�.=���B�.�Ѵ��a�<���C���4��6x��)�%蟨���Ywv��" !P�n!c�'�-�X%��S�? t�IȂ�2Z��V��<��q"O�u0��t8q���;XR��#"O�!���b�~1y��[����b"O<�3�oP]�<���+�̑$"O���R��u2Y1㊅@���C"O��U	F�~0�(p/�/�����"O��JX����3*�!f<��A"@��y�E�<e�D�?�-k�f�C��(M������ڷx>��)�ds�C�I�G�`�M��@S&9����7��C��]��Gh���d��R�� P�C䉀O"�9X��A�1:�3ER4ɜC�I=:�<i�Z�<H���A�6|.�B��O�p�5�Ƨ<mh��U?�B�	>h@��j�,�cP���@З�B�ɏEP�!��T�O�0c�g͇G��B�ɳi���A&���Q%T���	=[�dB�	�g�P�a��?�&��Q�4k�\B�	�:��䲖��Y�|���lA^B���0�@0Q�	��5��b��C�9_�4�@��Z�|���E����C�	�K��Ś�LN�1�p��	��C�	lL�R��N�+gDwF�1I�C�&hUx�;$O�[���gd���\C��G��f�Q�X�#7f�(V�<C�I>q*
�Rv��xQ4`K��S=	8C�ɂ&C�y�C�e��v�8'��B�I�h��x{
�n&�%
Q��B�ɷZ܌8�O�������^(C�I�P�<Aj0f�+%0e�+��B�I)U���X�c��0 ��Q�fU�C�ɱc[*q�WM)p�Xyr�̒M/dC�ɥ)x`i���$	Q��	G1�PC䉨)XT$�G�E�07<ە�P�C�I�k,`��N\�{ ��Rą�P��C�ɰ)�f)8�"��y]���%�^$0�C�ɚ6`j����$Tw�Q臣Жr�C�1&�8]�S파r4�[��P�sB�	g�Nq` "��+��#	���B�	8o.l}C*FZH���4�-�DB�#x:Ԩ���]	Z.nT���I��C�I�}��r��=��(C/@<$�B䉷K�\9SM,�d�X3�.l�C�	9O���:�h���dؠ��t0lC�ɼ2�b��gh��k��{b�B�a�jC�	>1EY����|r1�g�8�4C�I�R�H�����\90t'�u�C�I�S��ZTe�?2Hl�p'ȥp�B�	�'Z0���*ܔ�(w�G�Y�B䉧2h�4�@�O-^t0�4�"R��B�� 9r"�����Q�ت�hޠo��B䉲9/���ҍ�),��="DAݵh-|B�ɉS�� �]K�2�s&�۶A�~B�I� Ş|ˆ#�1=��r����+&B�ɵ@&�4(@�O�
��ܘW�xc\����D8���\�\���&6���3:!���=H�̺�T%l]T��lXu��ǔ�2�X�j�A�A�a���X�k�荒5$�3@�G��M�ȓ{hiۑ�P�mE�(h'̌5q> ��ȓw}��y��,�]�/~<����:E��N��w2�����o�H��ȓ!/L�[�̓E1�)C��!�݄���d
�O?:@r(sGn'Y��d��S�? Z �6 R����1Gˉ�0���I"O^�����gȊU�%�ۤ �Ա"OR���}4B5@�D����B"O�]�H؏a��䅼Z}��"O.iʤ'F"_���� (�3w<|{�"O�@8d!W�N��ɑ<\l81"O0m��� B�(MōZ�q����"O|�"s� r�(������"OR1(�"�+z|�e�F�z�:�+6"O`fkʟM���c`$�:d]��"O�����O0�����	H"Ox�*�
б5Uq��>pQ�1"OX�i�
W
��j#g�54"O���ǧz!��!Щeݐ�"O���LՕsQ�Q��(��PQ"OF��
V3q}�9	㢈&|���"O��ʅ�?�M(ӡI3s�&Tp�"O2|��N	�� ȵj3HJ��B"Oj�S`�!rVE{�LZ8+�9(�"O��@��Q�v��sU�Y�^),��T"O��c�"׭y�����!5��d"O��q�	
d��I�%W1�E�"O^TtǞj�0$�B�şsŐ� "OHM2�K��'v�$dг�N4b"O�S�L�� ��I{E� a�"Op�᳄P���H@+.���"O�A��hR�Aw�ݙ(G�!�A �"O
�ek�9X��-KeFI�-q�ԑ�"ONK���L�4$��#ҡ
�r!s�"O)��+A��L�b�QraHd"Ob\��I]	*�4MR� �vU��%"Oq2�-Z�0�؋Ձ��=N���R"O�ED��8hA[3.�1'"O�)! ��+}(��Fo���xX�"Of��S@K�$"np��J< �`E��"O0�7�$YׂyCMѫ#���s�"O8@�7}���s��S�����"O�̋�@��:���ť�A�"O=�F��h<@8Qc �`̲�Z�"O|�2��K<8ed
P��)oP��b�"O^�sqB�f�t���}Np�s�"O���Cַl����!��+����0"O�D@��=�`��R�
� �D`�C"O\�J/�,�
U{�.�2��,hq"O�,k�hU���#���:�
T "O��3�R��r��ìQl���"O���1�I1m�䤈�oɰ)Y��"OH�9N�LK��0vF�LZ�0"O��5(xP�P�5��Gh
m��"O�����Y{�|7�ҳS�j9�"O���O�s��Y�,T�U�L�G"O�Q#〉v&��aC�T�|�<E�"O�����s��� �I4�Q�T"O4���bɜ.�����ΚON@9	w"O��g���H�!�p�?c2`� �"Ov��nPyL���N�:`�B$"O�Eh�yY��I3�&1���2"O�L�$ɑ +�X@�X�N�HV"O�I�#��F���q+ֹ����"O� �Jʾn��`�R��4i�4W�V�<��� {Rj=A&�D�,��S�I�<�$@�hIF�6ȍ�xfA��G�|�<A�.2 `+� �Lz���-@�<a��8F����I�22B�:%��}�<� ����H�
�bA� %�4ŤlC2"O���Cђ?v�]�E h\ زS"O.�����l��Ł�d�Q0$�)"O��8��}�,��Bޝt���P"O��#4nˏz=�Q�k62��%��"O\Dؗ�Z��1y �V��<Ó"Ox��JS� 0!��T@l��"O��!6�
s�ޤK#�?%H���&"OZA�'�\�}��� Q��YU"O ��Pd�J5>�R�/SA$MBr"O8���8x�|
�-C:Q-�(
%"O�%b*��G葪&�[�q@d �"O4���!Ay|%"�KEo^B9�"O ��ǧ��Bn���/kR��aA"O�	�2囇^�$�8-�=E�6y�P"OR��u�6�ֹ�g�G�J�^X��"OZ��𮏠P��,�9�����"O.�[qT�)f��: ��b�ny�"O�8۰��9�.]���Sg��ԛ6"Oބ:�C��c�l�H&�@�6�)�"O`�*R)$lV�B
��R��0 "OVA�m�,^>H���I��Q�2	*D"O�T��l�'α��-Y�:A�r"OJ��W$)@Q\�鱌�-�a"�"O
��r�8dt���G!�j�z��"O����a��;���{�%��+t�ur�"O2K�m���E��D�2f<|ae"Oh<���@%RU�T�vP�5"O|<8�,�4Q���r �Hjj��"O��i©8qU:��p�C09i^��"O�)v��A�D��D#]7y���"Or̺3���1,쬓�,fX����"ON��2!�5�"fǇ\P���"O廦g�3X�B��՛
7�*1"O@z��P�QM@�A@��F8d�!�DʏR4T�&,��B��I1G��!�DΖy�9�A;R̸�I5�!����	�B��/�P���ͳ�!�� �:��4��X6��@`ۮ!�!����P�2�U����t�]�n�!��$n�E�a(B� �U���!�{������*� �U�!�!�ٯ{|���-�Nl��[�eO��!�E�X,�8�m�GV4������!�T�!f��:cIt�F��?
!�C+	�8Ma2��1B2�#a�p!�ə7u4�3�h�'ya|1�R��69T!����,�c����hc�tF�'|�V�)�:]jdY���.�8�vo�C�,C�$B�H�BԣL5�Xg,+�<㟨��I�(��$zw U¤�CSB8:C�I�*Z�Y��$�̙  T�4C�	�R�pa@��ՙ20����	�;YV C�Iy���*����>,�w(�4C�.5({�iݪ.�����NB䉶��l��Ji�f���lEG�DB�	�+~���`�M�C��&�����>�4%Z"52�}С�@$�ʓ�U{�� �'��`�1@�g�|袠J�Z�Q�'θx���6�E#��:�1��'A��C��s5z5B���?��3�'�
���E�B��s�\�9��ջ�'�~E��'N�4�<��!Đd)|Ez�'ʸٳ&�Y�z�B�	�*5^�x�r��� �=�ʍ/.$H�ҡ�>K��U�"O,A�"[�(�6����#V�ށ1�"O!�W��-�%ɟw��"O~4�I�#��Y9��B�MC$@�"OD��Dع��̋ ��%[&�ӣ"O�,;!���I�R���Oٍ&�Y��"O����������q��j�q[6"O��r��D�+����ѭ�A�*���"O���㎊�<'r�)q�![����	.~�Q��VA@�ȁ� �i0�pi�EA,?��9��i5��P��I?g6liF��݇�jcHtr��	���[�ꑮx�����mj�[�G�ͮqc`�N)3^<��K9 1:�bV
m�9s���%J�� ��I{�$g]��X#' ^Ӽꆎ�8, ZC�	�SOXXƤ+���6�2^�b��D<�V��e���K�@#�\�`k˒a+@ ��Iu�'d�e+L�-	�Ŗ��1Z
�'K�512C*<� Q�DK:E�>��P��$�>E��'��! jJ�[{�q�0��5�,���'���y��ڇ\��X����6� ��dڡ�HO���r���b��w�K#�̡3����B�Ҷ��(Q�1p�[�a�ц��	���'��?��e?�z� �3~X� �	*LO����ͬ@vH���]�1;a�;��`��"<��y"� Ô� 	�g�̕b�i���yR�Q��=c$��I\�9玀!�y�kC>C���q��ˑGs2�+Y��0<َ�d*&�U#�$p��8��e!��	�9;��\WI���W�%h!�D'*t|���:2J05�&�R7{g!��,O̊�P¯�-YB��B�G�Y`��c�'�̉��>��\C���	{��i����<�'�1��x&FC�&e�-+7�K	�PS�"O@�R�p,�h��c
N�!��i����<�۴��?7-^:��Eh׋Z�]���re�&88!�D��p�j�"@	�咴�@e�&0�Q�T��	,���{��Z8%����p�	 �C�	w��h��M,b8��3��z���$�S�OK(���B(I�� 1�Ԝ[ Ԝ�"O�`:uB���^$1��ӣf���"O�`SOڄ+��ʄL�~gY��O��	D��<�L<ͧ@F��2M�l���C�ئ���	i?Q�"�5RK.!:�å8�RT#N�P�d�hOq�,�ǧ�z&��\�\�����'�`�)�N��B�:T�xC�Ol���<Iߓ0����3?��᪀c�r�F}���E���A�e[��t	���${�C�ɴ�^� ��W/\�;3�Ɔ*��B䉅���J9j�B�S�@8o�B�%~ �Qg�T#$����b�OSBB�IRdTq���&-�YJDcD�K��C�I��i8�NM>sI�ģĬL�(z�c�HF{���ǅBN�!7 m�H�p�gI�yRѻT�
��m�(e��A����'!h���Ib���xp�O9)�q��ŕp���$&�S�O��V� xU1�l�T4Z�� ���y����l	�p�\H��9����~b����O,#=��F��{R��C*�Ds���-U}8�$J�4i2�+i�ġ���M�$�D���1��:�S�'oA�H#a�;�ģp.�/�ƸGy�
v>m��k�S�ʬ�E�)�@��?D�hsC��}�ڹ����8���d;D��K��U+Q��+�C�)��3�:D�� ~Xi�;R���z֡R=g���"OH�j�eK-�T��^�R�����"O�)a�H�m����� <�4R��xR�'�9�b�ͺ0�����
.=)�(���?��O�,�R/[�S��I��k�
��'@ܱ9�!��3y*p����+1^\@��$-��?�n3C@�p��!��P�B;3�DC�	'{wXi0Q�Ԑ]K*��5I
'V#?Y��(ڧ+w��IA@ȟ{���f@C�,���L����w G6���:�n�'[�`��'aў�}:s&�8fHe5(��p��M���XK�<ai��Y�t�㋜�P���21�WH�<��ő���u`VnʉJ�Z�!ԫVH��$�'��	.�9���=��e����=+,B��
N�����/ݒ���Jb��c�ϓ��'��'�J]!,^+_K�����04�L�Ǔ�HO<8(��!9����+Y�uf@��"O�x؁$Vf�~i��	�.X,�}��Io�����E������#w� )�׀G+y�!�$�
�)�-��1���A'�!�R��|!ˀ`�ot��C"�/@�!���MM��oμZFHM8E�L=l����I�\��(�N����s�&øB�	�n�аk�F�{~�3��C?F�v6�:�d��ݖ|i��p" �F���m!D���*\�,���$S��<Ѧ�*D� ɇ�ʔn��P�T��T���&*D����)��-�A����d��F&D�xh��)�����(�"4�׭.D�l#`�]�1����fQD��#d�!D��Qt�I�9�r��V��I�f��M�Dh<1a�ӻV(��/ȸ-^*�x#�p8�H�OT���.�7[�$�:����<<�"D�t*fB�$wh�!P�+\�zk�$D�Pɷ�{� ��j4��)��!D�Ăq!�4H7�|B�̓g�8�f*-D� �jͧjI�h���^G[z���I(D�T�r�O�W&���dK+YD�1�Q�#D����K.B�	[�kC<PLV��2+#D��[E�ށuN`�Vi�n.�i5D���$/��䐸��ߘp�^��w'4D��{���37���q��L�VY� �0D����a׬W����A�?��#��/D�,K�F��U�L�@r엽D0Hu�#8D��)��]M�����?�x![1K5D��!l4!���*#J�	u4!���.D�D��$�)#��m�L��,-+qO2D�XpV��6G�2���&W>�vm/D���p.����0@�F!j�h��d,D�T��Ǜ*� �C�y���*D��@���zfv�8�,@�3�H��*D���� �?s�X�����-Q�q��#D�4�B]�	��x�V ���5D��z)�/X��$��%�F�x��6D���gEz�#�ɖ6��I`J*D����0i�lX;Q�8>8s�I(D�P�@g�-����"���7�P���:D�<�@��1(S���t�3:��:��8D� �B��e�����:W���a�+D�+�b�:X���e��f����Ѧ(D� K�ÃU��Y��"��%����	�'��<STd�3ʜP��E0*Dp��'�!̗�6���f�%xD	�'���e�	H�J����ݖ�4���� 
q�0�[�q����iQ8�dR�"O�XC�F�3�4m��J�"��"O�����T�tB��`ߦn���"O�q��`Y�R5j<��i�:���h��':��ĩ\�Q�f� bl% VT$[p�:[���u�I�Rx�%q	�'Tf��5�� � 0A0oU�Uz�dH�'4�Qb@�oZ��G@3|���c�'�\-
��'��l�_|ذ���'Q:��6��S'ĩ�f���-���	�'r�A�R�Ak��B��U�
���'S 4�0cX�'�&1�L��E��'V��է�����V,�\�'0�q�S�D�l���@�Ў]��'{���6d jL� �_H,�l��'~0�� �<�\Q���Z�2��A�'F �)Ѐ�<ꖔz��R07_ĳ�'�R�Qgc�%E�ġ A��%�.� �'�*�� �!q���լ6�:�`�'�ށPM�;�|��������
�'��kek�XT����r���!
�'��]=-6�$y��I�y*���'�X��k &o�1G��5%@1��'��9�d�= ���P�Ϩ\�B�r�'���Ġ޿-�����l۸B1�Y�
�'+� *�N�}˨�z&�L�;�FmJ
�'~�)��,�%x �yq 
�*�nt��'uh�H��u�v�iP���Āqz�'P�I��h���w (c%��q�'��l��U�X����M�"�|P�
�'D�T����;��)�e݌�-X�'�dA��h�쑰��[:fHY�'�����Z�P�\� !�(UH�'������V6��z�#Qr44A�'HHt�Mۜ� !��l��C
�'�=���V��i�J^?[���'m4 ��� C0�����Fp����'��@�B�<4�^h�c�7
h�x��'; ��ǈ�5^��5�s!6 ��a��'�P�;�'�^���V9|[*���'��$0fJ��/>J,��mz�(9B�'���MO�x���V��/�f���'OȽ �&Inf�� �M2��*�'w��'M�#��Q�' �;��A��'�ʵ����<z���i͝4:���'�l���(ܵ|:��)6&�<7:���'w��P�G�pa�i�%�
��U�'g )�d��as���0g�xa��'<<p�[E���ؕjX\p$i��'b ,�	��ٔ�Hz���'=�IS3��<������#A�����'�F��!�хC����*�A*�T��'��� ��)"��Pࣦ��1ˠ�[
�'��E�b���Rt����<7e,	`�'��AR�DM�a�����A�u� H
�'�.��c���ҍ	�(H�]�� �	�'H2��M��Z������4��
�'(������_*m��B�K�4�
�'��A���ޙn" �\91R)�W�)D��{��Fg�*aD�85�TY�P�)D��!�`ί2�]i�c�5�"�9d'D�,�K%o"����.�JBj11'0D���#`�$.�84m�Y�$Z��5D�Tf�	�,���Ώ8��p�F	?D���dɀl?����/��B�8D�� |]�)�D��2ė�b���v"O��J�d@�r���2O$}=���"O�]Bfd�`�
 �&C�')���B"O���A�H�Rf� l+$,���'���H[
���?i��$����B��00']�B��Dz���F~�����GQ��b����g�S��,Q��S�M��]��GԻE
�8��X8xB��>f7�h%��z��B�jW9n�TH��\�U�2h�/O�Y{A)��pX�&>�'�t�z���!vz�Qq
_9?,|+�����M�R���JAhR�h/���S�՛[�Ơ�GaĲ�2��v�X)�0>y֎R ?�� r@0=ހ٠�ˉS}r�و��FLƥ\L�8�O3� ��̎4f:<�Z�4�v����5>�P=�
�$Z^ʥr�"O���"�/zO&�I���4����ъ^.6��I��t<3m�;;g���ҟ���26��˳6�Bq�үS%=��+��r��{��'��!*�m�>x�@�B��5��	g+*���Gh(Y�)�a��q�R���h�{�N�r��4��>��5}���]^���Ǌ����ؘ�ڿ����'�J�2�P� &0���IP�N=��@���>j֐�q�N@�]�܁�&n*z�6�l�s7�'��ijp�;G$n���)c6�M;�'�6�[$V%��z��X5��aΧG&d� �ب`0�E+��Y'{���d%Lt��`b�،P��\��ݟL'��#&x�Z�Ѣ��!��{��K�5r}���ަy�W�|��@9  �,M���E%B&|-�W�H��Ɓtf8uq%m�r�����c��}���a�|8�fͶ_���8 �ؽK\"�*�� �T�����$%C.}���̵Y��h��Y�I^*��ת�<ѱ���EX%�׌47t�! E�'r|���$}L1��C�[l���7P?�y�6��0@V�0���F�-#�ߖh��ɮ��
�-�0�џ�{-�R�������Y����5OP �k2]d�0��^-x^�7�ڋ�n�Cfk�W�4圻b�J�`֯�F��S��PC��z��0�Z��kvXP�
x�VB�}�xYZ0捲`;�m8�n�%i,B�gI֦n��]bP�spɚ�Tr�M��Ok�o������&�4KM	J@�}"+M�HF�5�Fi�!yF�t)��T���k��7�(��d�7�V����X�Cs���QS����j�F��	��V��1�k^�]7�y�F��2]���w#"�p
�gc��|U�}�$L�4��ɰ�GA��t�ڗ�W�N��/\����ʱ�W���$��rL��'O�l��KA>D�P�4�ʐ~<��2O�c��4Ii�$�G�/�`��K�<N�H��?u�b�)f)��@���:H�� ޴V�^�r�
O���/�3?fȤX�EEc���;�!���~-���	rQJ�HvͼV�S�躼���:?�4E��1�H��$Ǝ8޸��1��A���s'�Ll\*�(�%i4}i�g��v�x�!$%Ǧ�q�F@R${r���֟@Pax� �	T���`d�9W�,d�9��O�Ȁ�
:J^��ӥ�gJ���2���hRJ=}��3�n$%S堚��x�c�Mb����:ƺ�3qk���D���|�av]�^/>��p��5�2;�N�]�'M-p! �^+�b`�R$M(s��t�ȓ0N����O(*:|(��A�R��[#�\�Dm����BC���5�	}����'�b��#ϐ�?�$XU	�&qD����'�f��s�m�r���Y%l�����l:	�&iƞ*���`raVxk\$���+�,����O�G�h�2n�`�p��D�?�ъQ+ԺW�q�����	@��pq���@�&I�ӣG�+L��!�?$����- ޒ�6�=M@(�� 1�IK��)(t�ߵX{r;�ӱT���34/O~<0�é��VC䉠mY�9I��?*t{� �=���6ř�G�\ٛ�@��~�\��ϑ^�$b�΀-�ƈY��-D��[Ƨ�|l5���)	��O�<�G�בj���pៈ��<��C���M�f�E=HMH�a�ϐ{��Г�DD�E���@_�
X2���N�>��CkW
~B ��Oܝ�# NК$DB�>+V��Qቪ3@����-�%Y�����V��c�h �1G\��y�k�'�`V_H�ɖ`L�~P�-Z�K&�j�ˀeTn��S��?A'Ȉu3��!c�%V�Q��x�<y��|�~���׮o�N���w~2a._�&���'�P�� T��y!�$�N���d�~QRE�;��S�j�Qy,m�Ї�5z�VC�ɱW'�}�Z�z��$f��B�ɌT1x+��[:�f	R̛�Z�B�	����Y�E�Bd���[�JVB�I�en !��?%/���j���B�II�����' ~��S�O�<��C�)� ��)w�Q�>��mV��("Oڀ� �ӨW��&�6@�"O�Y�e��@����ao�*V���"O>h;c�	I�}*�%�(bQ����"Ox���^=yb��Ό�[��@��B�,b
H(Ó_�N���FE�-���)!'�+�����_�F�z��Q�6�:����Y��R���E��`� �����Y������#5�6hE2��y�h����gⓠh��FR� L��!��77&B�.@Y�q�!��h�a�K �+2�ʓW T�1��,|�ҧ(��-h$!��Gwlܨ �B�+�H:@"O�hqU�����Wh[��xЁV�䐹=���� �-���X����C�h�;iE��1C��l������IA%�0�n�p���_\,}#D���S虇�It�(�`fѦ6�����K�E�̢?�`cB��T�C�#�i�u��W+�͞����35^!򤗌 �6�1pg�7�B(���<e9�I�[��=Z�ڕi��S�Oz��󆤏G�jҢ!73G�y��'�`+�@��%x4��ٿ\G��:�*&}"i��|����%���{2ኜ;�~	�M<Bl�����=�x"��94��,R9^ZDhJ���#KRū��0���k(.`�K!b�>��Bo׽�p<�!o�@>�b�h�W'^�!QD�r��	;g�����9D��1cmE�*&\xfC	��U���4D��0�C�_��,A�Ǩng�S�3D�@U.�ʰ�h���;uX��.;��xw�'���Vf��,ގ����	;E�I�'�����]54X��@�%34�[��C�+N�U@��'��e+�ϥ
Vnq E�E�M�>�j���\�>�$D��!���ħ�}v�9%���� gc8���\34Yj�K�2J���f���S�f,�'� �+P�xF�OQ>�cϔ19�x!�ֆ�L^v	r�H$D�hm'J7�P��ى!U�Em�����3Vʢ�K�3�ɘv�B��1(�9.�CQe۸$u@��D�u�Z��KUlV$��)G6���D�;�Zq���sT\Ѓb�.R�����ޥ�.4GR�ϋH�PK䣋z�S# �a���:k_HP{q
Ѷ/�C䉀i��P�UcՉ0`la����FH�˓T#Π�%mG#jӧ(��Y��	r@�� �膐)w"O �8�gL�/��hK�O�(qߎ]h0H�H�$�S����0��� (ښc��6U��l�r�٨px!��� *�^!���J�,;~�B/�q.���FU*���d��P���Um놴�G��<R�x�k�eV���<A�O:t�F����)g�0�Qu�GU�<�T)I�M0���RJ!;ڤH�⧆R�<i�	�YP!�#ef0�7�LS�<1G�<\B���RKP~84	�NPN�<��Q6�x�qd�r��� !F�<�1��R�dQ�1�H�=h4ᘱ�B�<�VO�w�V�@�B@=SÐ���a�<IE+��m�	���F�9��s��P�<�2h��	/���#;w(�3)Sp�<���]<!
�B�0U���+��s�<��O_�7'J}���.[�B]�K`�<A∅q�t���nҢA�Ċ��e�<����7iz�r4��4(�
��i�<�i��uI�p�e�m���j�<a��&b�� Kg.HVF\RA��N�<��#�q!���D�2f^�y�/E�<c`	);SNLxg&E�Mb:}�1i�|�<iU�S9"ijL�eǇE�Ĉh�O�<�Qd��(A! #B-`F���˜`�<��#����k��Q�a���v�<���-���͙bN^���IHn�<� �9�FøE�$��E�S�(<�""Oڭ�N��Pe��b��pR����"O�=a���X`)R���h�p�"O*Y�P�,�n���gI�i���;a"OZ��d@�7�H�{�%U�`��P"O�����٥NQ)�%S�9Z���"O<T�Ю3Z�t�Zq�ηA8K&�y�f �'�2'D�	��Rq䑋�yRj<v��Ud (
�����y&��I��y��8/�!��G��y���D9nx�`�(f�Uau���ygS����+4����q���y�	�}>��{�cK� ,�0���X��y�$�)�1��k���A����yBj<	Ș�8 �N�zo#�yr䇇Zބ��I��~��X��Տ�y�M�E���x��-]D����ė��y��y�F��#����H�	��Y��yb-ʘ�\��֙kA��	�3�y��`G� cĈ�8cF�C6)_�y�H���)��_�g��U9CD*�yBC�
`�2}��Qi�8KgE �y�D��"�����O�D�~��D��y�C�J.iP4�O9���0U��)�y���!����hͧI6����A���yBk�cSj|q�jK�7�} b��y��l��9%F7a��D��y���pT���E�t�c���y��'\�s��2ւA0��Ң�y�kƬn,�<ĪUf�tU�D��y�ĄFƮ�%�@�m�� �F�yc�	K���ׯN�V��l�&!ԡ�yR�LY��l��6W�z���mF��y� ZU��IU��M"� �e��ybOD�#z�<8�H�=?�V�xċ��yҏ���<
��ȗ\��(PC���yRK��\��Ћ�ƳW�ܰâ�U��y�`��*�X�!wf�X�3b����yZ�z�Z��$P<���+�e��\g��I�*M R�l�Ң.�[<���.W���F<\��a: 
g�8�ȓr�t�Av��y��+:�ه�~'hY�VIDu��AA��;/\��ȓL�.�;%J ?�q��|��]�ȓR�vtK���^��b� MW2��ȓ�AEDY�Ft)!U*͝#/�Մȓ,ƒ�r�H�Z�p��R 
�̆�3��;%��$ƀ���ĥ+iD���$n��;BB.�v��BJ�=�1���:+��uh�0��Ʈ>����ȓ&T	sF-���g�J(2�u��
{4<h�C����fQ�!��фȓo��PH7a��KHV�@��/)��!�ȓD��x!�Ďo~�x+W���4wZ����W=M~�5"OD�v�ۊ*o����W����G"O<�[� � ��ulϊ<���7"O�����5?/�+�99�1C!"O�t1�ů�=����$��q��"OX!W/ݙ;~��"��pZ"O�,X���v������-�TA�a"O�1�잪8�����
渹B"ODP�	O�*L�8��L�=�ұ�"Oժ�٬dӒ��j��.����c"O� Z!�R��n>5���UE�(�c�"O
<��ōP����􇙿0U��qf"O,�#��ԫ
B���I�6E%�w"OE��J%�vI���Аp<p�t"O�)�7Ć2�Qa2��/,��X;�"O6��q%�]���C�^�+����t"OPbr�J
t��8âT���� �"OH\�']-�0�!\7M�9!��'?x��͓uO�I�Y"({V�
)L�W�F:A�B�ɪ,�8a�Q�r< ���3hYlb���aE�j\f����S�j'^]�eeM����j̛n�rB�I&I+�� ��j����*���u�:�(H�.O�Ӗ
"�3}�M��K�H�����0^���sڠ��xRIĴ�R���ڸK�`P�䇂�>]LT�h��KF���d�'�,�㖎�5i�,�AL�?i�L�	�4l����M�9c�X��'�%iT)I="��BL�x��3	�'���*�A�a�S�#ܒu�B�(H>A��\�s�Z�HpoʭÈ�L�	H6	�T(*5�O82i.`X�"O0�b'J0,���5!�M�Z,hP��-pδ�r,��[���t�)��j� �nE����M޾ 	�Y��I�����O^�`���+?�A�o��J�����U�ȹ�R�7�Ҁ�di��B2J��$�Ϯ4�ą�.O�
q�L���O��#����z�p�I_�0�`$	:3r�g�2mD|q�$�Q ؕ"F۲g��Q[��D���?�1*�*,@:��dĐ_��H�a���|��R��ND��ȅr1�j�+/H.������t�W�[�N��55Ҹu,��z�s'�n�<ᦋ�>,0
�`��?�T�T��$o�D����шq`���a�@%H�.@�?(:� ��]?�@�,OZ��"�C�(�4�.+f�Iq�'`
��FK�m�L�Z��^�#�taV�z{ɐ���Ԙ�"��WF}�$ �؜�d�UP�'�F8;�]�c�vPs"�6�Vq��{Bb��W��LREbY8S��4C�S��Eө��sm�<6���w"цlV�5��4М�����7!���
��*֬D?"�ܐ���/�>X1��P�a�J�3b)mݍ0�&J)	VDPz�س�����VF�F}l����
�
vT��O�8&_�]����F� +l��2��NO������٩n\�R��+F�h�_�p��@U�5jT%��W��`���%xG�렣
�d
lҰ� �f��IdN(Jt���+8@Pf��5��8��! ��spCm�"	A+O���o�f����E�F:�H�
��W+���Eo�7��	*.@N���#��?aԤZ���
/F��dUJ��b�"B*�Z��$"D�n�0s|d�J�o(<�6��4�8��(߈<㦌k��eq�KA�6����mI0h�\�%?9����p~��{�rXhE�܋��%.���?�B��}�<P:ȁ�FЬ�c�7U�T9�cI�'0�0�č:;�D35�բ�0<i�޷\�J �blW @ZX�*U�'�x�{A䋲Xa�	+S΄:4-Z 6/\U���$]�� ���c_�J�O��y3u�ZxRw��.T �3R�0K�I\?5�L	�΋/t�a�����|
���<��|�tc�:��uVœN�<ӈڭ4���G�.@6A�![�4���sJz�~�䓵c��$?�R��u~�@���-*��̛CU�hc���x��@	I�(`��.>8�& M�Z����Č��aA���l�`���_y8�10�y@�G�f����6�H�y��xB��1K��zj�3$��M/l�Ԉ�ǼP�H��V��.7� ��v$�)_!�0^~�S��Ԟm��=�3��w±O�Ă����1F�P�O��Qy��d`{K"_;B��E�
�ތ3�"OARO ��㷩�<Z��SG�L!��qQ2��9{�0���h��W�q8lq7 ��G���yGd�a�!�$�^�� @W9k�9��C�#���
`��f���:>8��ɤ4[�b��W
>��c爠O	����:p��4@ѧ2Q�d[r�ɛ����$I��7�B$�fn���x�K��&�4�z��ׯY��Z�G��O ���g'GRA:��	o�g�H"'��wq�`u�� C�.l���Jq��A��Єˁ��x�C��PhH�q��)�)�矘�#ŇU:8]X�#]�����l;D�<��+q�n��ADH��423O6?����	0��a�@;�5P� 6 *d�F�Vx����_���� �GC�lh�ł8T��H�KBV�!�?_�j�@�	�?B62��;!�� >h����
y�(⮀�#�8�P�"O�Y�d��ҵ���L�l����1"O���p�.Sw�c�Jō Bj\+e"O��J�O����`7�H>l�\���"O8�`ՠ�l�ΙAI98�y"O�T��#Ǔ=��4#AIC������"O�%�Dd�3B*j���@(&�:���"O⡨�Dąo�}: �ϛݾ�{5"O��C0�E�HW����A�P�B���ƨa����	Ó^�<PELƽl���Hr`�.S����^�4 '�ӱY��9�a�V	Lu�@,ܸr�4����x�����@�F8he"Ѐe�J�D���d�U+���I�S�L	z�P��Q�:�@�fĭq�\B�,��a�cD�={�< (���.*!��ॣ ���e��ҧ(��YV
2x>�y
�2�U0�"O(�˶�ڧkT�#����8�d���-}�d�t{8��U�;��$\� �*� �@��7��C���⋜�%����B�e�D	9qiؤz�+T�Y�-s:8��ɾG�Z1�  4A%a�S�̢?y�@>4��$D5��ʹa � 3�U�f-����+X!�E;�T��.Z4bʌ����+,]剻jטyx���t��S�Oxh�1H�q�̩
�C�	;����'K����	e�:�2�N6:䀖d)}rj �bh�Q���{�d�c�~P)ǉ�p�ґ�P����x�$'a��9e��B��<S��&=̬1q��N�RG��G.l$�t&d�o�^�E��=�p<)��p��c�D�B�0jQ��X�֠IqRi���$D�0S	�n~L3ţ[$M_2Ms�,D�D ��$ j�B���
=�TH�A-D��J'K�3J�}��Ҩ;ܤtI�*=�oP��B��'���^�ʽܴ#����O�1 ���#��J��S��0��)������?�thO�&NZex�F I,��1+�i�'�,Y��� �$>U��V/z�MX�cA��� �Q
2D�|A��"��%��M�?
3j��TB�<��̊4 �<옵�2}��I˸d���sA^_�*�C��&Z�!�	,E�Y����Uݠ1e���p�b��O�U�JI���qOf����L[XIK"�I�_T� �f�'dl��hюlA�=ئ!��*���ełZTݘf$ZC؟\ c ^:j�D)�v �>8��Yx�&�y�Yreh[���]�4�^�\�,���R��Ic�"O�M�w*ѯ`T����t�N�;7_�X�"�8
����>E�DC�gۢ���I#k�)��Q��y'��av�8�O����`j�`ֿnr��' ���&�|��ϸ'�~�S�X�(�(���I�nj��	�'�z�3���PR���OW�ڪY#1��%o*x5�'��d�7	��g�����C�T$y	Ǔt�R���:��9�00����#�Y�Q�؅s�2B�I$W��E�u�)��Xe�)L�ZB��L|�%�3h�h���U�7�&B��͸ i�@.p3�@�۔P��Շ�n@�E���U�\N�0�KK�m��h�ȓ��d�b�V�
AHڗ��,)\�ԅȓBxdP���G�������z��ȓ� ���O�"���#0�[�J'<d�ȓII��r�À��q��/Rw�̄�dڌa���^t�2%�2;b���ȓ*`8�¢I̧um����<��(�ȓy�D�b �s��䒡iB�Z2q��+�zѩ&�!of� �V?air���[��L�$EC.p�� �!�>h
�$��Qhr5��E�(�d�c�#�\\�,�ȓ��V�E�������Ea���[]�e��J4/+�$�tj�U|:\��S�? �%�ӂ3(1�ىSGP�M��A"O,����]$2>=;�>\��+""O�1�뇴3(�P Sf��6<����"O���b��0:=����ft�{0"OH8��7ؚ�Y��g��@i�"O�d�m0���5��<��XC"O��mU	6Bq�Cd߲�"O�J����y�f�2�IW?`�\��&"O\�h#��$$�T�$J�*��D�"OD���nà���j�
PX�1�"Op=q��S��DU+�)��H#���"Ols��[�Q��l�Ub�V/�4�W�'u��R���(I��SU�Z Sߔ�s��Y�.~\d����53�`���'V��B���&̍�`��0No�Xd"Ox2�G�;7b���g�0H�Ti��"OD����	#��yxƄ]��,ɫ�"O�$�1��9�+Q��o��	�"Ò��&��eNX�T/�!`��J"O�0�QaD&~����^�#�0"O�mK%m�zd.R�4�����	=�HO��$�jJ�)]@��J��3��	�P�L�
m*1r�S�'���#7(��	�>RR&�Y�@�v�5z��`^��+5E]y��II�uMVI���ǴNc�`1R�٬Nn� S�Dդ^~H�'�8��� ��� QiX�6���+DD�1o�D	�윏��	�"�v�q��?�i�&i�-0qȒ@��|8�FL�1T4Tb�O� ��ƃ	6cx��
�'LM�"�U� ���3�Q�y�5�'�@ �P1��ȻN>������g��\ 
�1p�=�&o�I}�B�Pь��=E�$�ٔI��[᧓W�����%V;�y��Qz�����k +En5��'��:��S��6D�@Q�MB��p��l�9���'D���b`?M�$[E��7���3�$D��z�Η�Ń�ć����5F.D��C���$K:��6Ʉ*Q�,㑃-D�,��B
u��C� D�E<Ը!�+D��{�Wz.���m��9�s)D� ��]Y�N@{��[<��ܢЌ:D��8t��;����v�X�hk|�@	4D���V��)��1$�X�
G.�c��3D���2 &4N��4�,�$�&&D�4�ܮPHv�;i��v2���, D�@ㅚ�!����b�/� 5��<D��)�O/ ���G�}+J>D�@���'ܰ(�t$� g��3!/D� �"�Cy��:����j1iG�8D����+�d����)F�_�n(�B8D����{"�sD*C�Wn���B6D��	� S5S�*QZuk�x�zMh�4D�@q����S,�{�A�DR��0�H7D���f1�`1yӦ��wnt�9�*D��p'�4dҢ�IF��C#V��4�"D�ل��=L�֤��D;OW$1�1B;D�xzCb�6?�[�CiP�H��]�v�+D��h&�1��,a6�A$��2�*D��J֬�.q*���B�(7�`;�k<D�����{D%CvmT�,	�pc�'D��+�oCC1�mb��M0@���r�/D��A�ϖiEyӧ��	�hi���"D�dZ�`��zs(�j����N�;ь?D�\�C�4;E�1{n�IlިIRa>D��c�/E8�T����@�1�$R�� D��x�%O��y�Q J8�j@�d�<D��˥&�P�Y{@G�%��q"	?D�x���$<�L��7j�
���"D�ԲSDʡKR8�C�' =]1�@9�D?D�� �,�cIR'@ܸ'�_�;h0]�"O pD�87L)b&��)h�`��"O(@�f��Q�.9��� �cHfA��"O��t��h��xsm]�F��"OP�ڴ��+����,B��P#"O��hR���J)�İ#)!CR"On}�A��	\B`|(CH��T �$B�"Ol�cCa�c�6�.�R�"O�m+5`Ҙr2v�S��)t��2B"O<�+�L�"ר�*S-�� 邭��"O(��@@�.Ka0a!�,��E�nx�`"O�Id�A�!���d��,ժE�D"OV�ť�)4AN`���]��@t�""O�QukA�+�.��0���{�$]A2"O��%&�\��y� $�lI�"O� @�D �
0�շF�n��"O̚�Ojb�pѠ�9&t�h�v"Op����84��ҷ�*B[�9�"O�͠#�%~��)z�OK�Kq�{�"O���dW�^t��0�G�ϊ��b"O�h�@%-i�n����BQ���S"O��1�ܔF1�a�&�Ƣ43��!E"O�\�gC
NRh�
 �7#^�"O�t�G�7g�$b��<�"O-��]|	v Qf9<
\z7"Oze�aE-Z�DD�.R���%QK�<��f�1N^��8alѷl�2�PN�O�<AEO�+ʠTˠ`�FLn2Ӂd�<��j�,��iQ�ķO��Hy���\�<�4 U�JMQ���כ�]Z!�D�<#;T��I�H�l��J�T !�Ɋ=s�`P¢�#:$�yb���~!�d��G:H� Q	��G|�%XCaM$i�!���m�DbpU N$]���P�����A6o.J$�ǉ$�"�⬈�y����4�Х��	Q�E{e�)�yr(ĉx_�d�T��-O���o�y�a�4�!3 ��!�HZ�m�$�yB!�O��hA�.u�����X:�yB��7D���I�S�y�,��6��+�y���c��Y$�wt�!
�Py�ˋ>]hѸv�Y��X\`��Rp�<��ᅀ.��X���'|X�HVi�<�B��1H?�Qi$D�X���[tIJq�<�b��-~l՚���9z�Y��̑b�<Bn�J�C-�?�T��!�G�<a�j��رW�U�f����a�E�<�N�-X����b�Ab0��1-C�<Q�낂r�
A�a�^�(�J���c�<��V�%��q`%ǞsD�P0I�c�<��L�[]HsQ�"A�4���Le�<q�^�k���ɵ[7Z\ѫT��k�<a�P,/���2ȚwZ�-2��p�<�̢2 ��С�\ z�|9ƨ�h�<��@ߞi��km��=|�BG��d�<�d"��S�<[#b
��2��%d�a�<��'Q����Pj��ug����e[�<�E�<E���@�OO�>�m�T�<Y�-�'���z���u�R�[��YZ�<��T�����!n��\�X�R�V�<Q�I�7%�>@����'�|9�QR�<�ʒ�9�H�C��B$bh;Cv�<�&,��z���#��yZ���*�o�<���]1x��A!�Z�m�@c�[i�<� H��î�?f*.b���C�I�"O�q�T��5@ZVa v-D�+;�=R@"O`���W"?>�Q���݇L*��R"O����$x� !�ϖI"(�g"O�@sp)C !x�1!�7:v�|P�"O��#��DF�|Y�J�9AA>��'"O@x�G�W,�X��U(	�M+&T�R"O�:�/�K�6�Y�)�,���y�"O��dʹz0��H��o�� 0%"Ox��Q[x�|z1���h�z���"Ol�XO']��#�j�2���"O���Vg7t`����ڎN�
HA�"Ol݃�f<H���ZD�ɖ3����"O�|K�!,���61?�԰Y�"O��ã��y�h��&ުb�����"Op�r�Č12Eh��_�4�X{�"O~�B�k�w��p"�
��U��"O��͕1e���G��|�n��"O^�R�)�2a�0���1[D��"O!��kÞU��l	ƥ�|��v"O¤�SD؄/�:��7d�d�cG"O��Q�@O�q��!%y`�B�"OD�qr�٢]���H FXj	½��"O,�u���V@�S�M� ����"O��[�@A ]r�@�'�T�E"O �#�$0������,�PA��"O^�˒⃅"ul����]GF|yC"O��S�/ٙ]S���D�hV4!S�"OtD�6���jF�+zh"O�!䦙�yil���*��<���[Q"O�W�� =�(�F���`��5O�\�<q�J�Ȝ��
��7`H�"U�<�RoQ�^?�E��?x-�C�F�<iș�*햅�� ѕX�:�	%OP^�<Q����wy�k_�HCL���\p�<х�?aΕ�َ8���a�![n�<�ؕf��ya�E�|���$i�j�<�G� Exp����$3���_�<�"T1"_
	i�ȅ-2��n�Z�<�p/�v�#���9� ��J_n�<iV�^>=\H��K${ܚ0VO@l�<aը GvbY�V�ψ[b����R�<��D�F��`�_/��r��N�<�⌗l�R�����;��)�!B�<6a��4�< 'E��.�uk B�<!� �2Ԝ����6I�Q��"]@�<���:a�\HV��V�~�0���p�<g�Jhd�C�F�s��l��#Ul�<ɅH�)�R@���nխg�Yr�"O�V���0���MS�P�8(�"O��hc	�	fBB`'k�#p��j�"OB��'@�
{'����7����"Oi��D� _fda"`��#�\5ڤ"Ov�zf��H��	/�tt2�"OFT"�n�>?�8�2σ%w�p��v"OeA/�4����P��/�.�8%"OH��.U
�4htC��W�rmX"O�M�b^!Y�4�QC�	��a"Oh,@�f*y��M�S�ʩH��h"OX�������H�!��9��١"OH�3�ڧ�(�!k>3TDD��"O�!aG�X2,U<�0�I;IT�\
4"O�e�.A�!G"|;6�Т=~a�"O�t���:@c4��ף�m#N���"O� ڰ��Ȫ�,��֠8"�e��"OF�6�4W Z��d
C���"O���되=��Iʱb#x<��"OT��mEsI����k^!й@�"OJ�� h���� ��#=f	:�"Oly���O����1��7��p"O4�Ra�̩	�@��G��`�Y`�"O��R5d��>z�$�֮�6��d�G"O��AI�0`���s䋡S�B	��"ǑK%�@�A�ܜ����@�P�i "O��S�-H�n܀UO��6�����"O������LI�9���E}xx| 7"O���6D��DEd�΁�^���"O��%̉z�� ���^�\ &"O�-P@f�9.5ryȵ1QT$���"OT�P���,ܪ�`��a�rU"O�D�&�#�J�(����q�8�"O�� M��]��͢��G��~d:D"O�Q��TY(�Uӵ��_�"�Bc"O6,K+ې$��<���̭:���xw"Oj�h�

�Q׌X
��
;�����"O`=��S!��D�3���r&"O�9��*֭~��o� @c�`�q"O�a�UL�0�o�\q< :�"O�hsq(D�9;Xh�U��uYH��"O"���O\<-����D�Ԧ7=�]�r"O������#;�貁`�'hD�1K�"O���H\Lߎ����\"];!�"O��x��B�^���Q5���J.؍��"O����/D�IC��&$^�V"OL�	%	S	H�r	7���T�f-{�"OSWJ�~p9K׍	�d�֬JQ"O�  G���{�8�9�+A��` �"O5��LĞ�
0a�Kʝ^�p��3"O��͖�8��agJ��N��0"Of�!WG�Z�>}�hײ����"Od ).!W#�S!B��k�LmP0"Oj��ǊJ�K����@��O��Q�"O�����T5YN�`� #��y3�"O��dO�'䙐7��eH2]آ"Ov#��2{z��R�ͷ 88i��"O�L�`   ��   �  O  �  �  `*  �5  >A  �L  �X  �c  $o  �w  p~  &�  Ǝ  �  W�  ��  ܧ  /�  ��  �  k�  ��  y�  ��  &�  h�  ��  ��  }�  ]�  � � � � �!  * �1 "9 d? �E QI  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(��I|�O���#�H�R!��њ]��p��'_��uʆ�vӲ�R�c�*m�'�*L��܉�` ��ڭ\�����$֮w4I�1O�,��g�W�b-h4��Ӽ9�HMB�tX���;%�2���IЦ�Fx��2R^zmC`� �p��#�ȵ�yRO����!�L�q�tR� K��$"% �"|���6U3��B0)зez��%�~�<)0��.)�#U��4��뵥�T�<��۞@J9������
�ĥ�F�<���R�}��%�	2a ��`j�<�d��W��aP��ۆ&Z<�j�g���'o(�TA0g�]j�ȺS�����'���G U*=�~@�g��J��p`�'X���	B�z��X3'�R�m�4u�	�':��D�K���@ W/�S<������ �\q�C1������h=�A�#"O8��N� Gv����^�g �<#��>���tl@aM�/Dc��2X���ȓp_�B�"'���BQ �萄��N5[�œ�J�lU���V ��-D}�����Q��*�	��ȴ�� �C�I�qv�d��+̅Z�����슃'�B䉌�����"� TU��gɭ 6#>��C?�'w�6��![�.v���a(3�i��j�X��`	O̙K�aX���YΓ�hO?!F��*e�@y�FP�@�XɫA0D��:4��(N���q�S�/�����,D��z�K��U�TǄ�'TI�9�+$��g0��9�� �:�����o ����9P�M���4t\�\����ayR�O֒O�0���xb�Ӷ���V�{�"OQ4�B�|;z��&T���S�pG{��	�d�\@A �K���)��/�!��>P� L"��"GBi��&K/}�ttFz��9O�I��rL,y`��hX�xp��'��+K�Q�����T��������1��]m��<)�]~��ʆ�&O`�3�X'>��1��	k}�K>!B�;q@ηn��l����yRaA�90�����Zcz����Y���OL�~:��N�8aޜ�A($}�q��a�c�<��R;/xВ��E-�:ѡf�c�<Y�Y0�����j��u�C��i�<��#=uL-R��	�+($Q�E�]�<񳋟�%D��O�g��,P�I[�<��g�&�:�r&l��G�.a��&A@�<6��_N^�R��:���� �y�<�w�ґH�yz �3�`��� �j�<i7�}�2٣QO�p����2��q�<�5�̏�xq��T,�s�F�<�#��![����UN�t˞�b!W�<��k���≨��Q &Р��|�<�ƤS��ڑ�UF�JIj3�Mq�<���ߣ��� �M�1vN�Y©v�<�q#����g�)��!��v�<ag��R�F�� �>���Вd�V�<�����Ttހ	�[\��,3aL�i�<�a�C�2��-�I��T��x���F�<q3 �jT�㶦ւa�j0I�~�<a��WB�<�S�	?sC����j�o�<�"��P�:���=bJ��&��n�<�/�"��ړş6K2zD��c m�<�6�P�*���^�B�ވ��ŋ}�<I���1�0��#�3c�R͒��LS�<�$o�^ľQ�ԀR;1�:�Ns�<�d�)0��f�g�����/DG�<i���B���UB_�&���SFG�<i���b��C�Hܭc�����<�k��FWL�#�M�%j(X�FE�<�ä���8�d��&J ��DoV�<s�T�\���9�2M���Q�<��/	�P�RfD�<��l�F��e�<���G�#�H�1�K(v�d�4By�<qB�"J14Y��͏%�B���t�<�PHZ�:0v�a�U�E��!Y��p�<A&	�W�� ���~tb|��o�j�<Y@��.k�:��m�9pt
Q�5%f�<Q�4F�(�3�����k�'�F�<����r��t��v�J�{F�{�<!ݚa��	���.����d.�z�<� v�B_�0�q�� �f�2���"O�}p�4�V%Y7b��i�!("O(h�`�lB���5�B�	��""OJ5�f炖l��1��Åw ��Ҵ"O�IȒ��&$.i�Vo>)#�ı�'M2�'�B�']b�'V��'P��':L�Ye	�#?�T�*�j����ͻF�'���'���'N��'���'���'��q��(�.mZ���x��1r��'�R�'���'SR�'.��'���'�:�`I޽f��PmK;�8h�t�'�b�'�"�'?��'b�'���'���# ��4a�R�QB�Ɣ�f�'}��'���'q��'�r�'���'s.�[ukF<7aq����`%6���'���'2�'��'w��'/B�'��p�D܊o6~Z3�E$#d����'���'b�'-B�'��'�"�'�8}�#ެN:�J�MI�?	����'Q�'��'��'b��'7��'B���
I�s�t���ع5sx����'�B�'"�';��'/R�'�b�' ��J]�<�K��ӧc%tQq��'��'0�'�"�'*��'/�'�b,!a� YH�,ܲ4��>�?����?���?)��?����?���?���� #�d���B ;�
1�A��?���?i���?1��?y��?A���?�r+�
�\��,O=4���+� W�?Q��?���?����?9��k��V�'���Y�i�"qR�)�	�~��5ET�3����?�)O1��I��M#�O�(���h⦇Vvb�S�"��'��6�.�i>�	ݟ�P��f�~�d��Vp~�S�M�ڟ�	�a�zym�[~�<�:��S\�IDL��i��.�� Ƴ"��<�����/ڧ��sU�8!�0�밯��J][S�i���y������]
)����t��r5���Z22��������i�4Ҳ6-y����]�[�Rsd�(��v��̓5Fr�Rp�����'�N���W>hӚ����� SΤ�R�'��	g�,�M�K�N̓n��.-k�̺ �QI~��{�Mw��t�������	�<ѮO�x���[�"�Y�#�V,1,dhǒ���I=F� ���/�S�GҎOݟ��	¸� �J�/V8�SmxyT�<�)��<)�C�*����c��O���3�+�<��i-��1�O�Yl�G��|2�ꙷhHQ���N^���Q&��<���?Y��Sܞ ��4���`>���'煏�\�}�"�L�m[l0Bt���b]"�Of��|"��?y��?a�t
�2T/�D]�)�Ĝ;]���p-O�5lZ/u�����4��b�����$d�*PR�*"i�͹�*X9����ڦ�*����S�'U*��P�h%��N�B������x[���<)��*1���6���򤆱Z��rF5�����	FL�$�O����O^�4�0�Sg��*�7�
#�Fɑ���v~��-W<-Ab�v�����O��l��M+B�i�F���� ��h�An͸7��!�#�H?����L�F#,l�����$9!��ɭ+ ��$��YoN`8t5O����O��D�OP�d�Ot�?a����h�3�K&3���v/���@��d�ٴFk��.O2�m�t�Ie���H#��Ք����Ncs��YN<ᴽi=�7=�TP�u�4�3ʒ���	=2��x���N4E0pe���DR?��d�'����4�:���On���{�ƥ(�	QZ̈���兦y�@���O^��2�4R�7�'���'&��5d)̱d���WF�qY1C�)\d�$����M���i(O�3@(\X�-��&�����,&8!Ԋ��pn����l(?�':���dې��a�l��ӡ�.�r�P�&#�j����?���?��S�'��Q����ANW��p0�kb��ӣB9y�v���˟T��4��'J�2�b�Zܼ}Q���<;P��+�O�~��7���EqpN����'ܾ�Su���?駟��k�(QKnD�&&�}��Q��>O��?���?����?�����	A�Q�F8c2�P?Vu�b���$ �oھj��������B�������Ӳ	I�@���$�d4{�:m����a�4�&�b>%�t��Ʀ�Γ^)��	g���㉌./�(�l�Q a��O���J>1)O���O`����,	�ʜ�׉H�W���X���O�D�O���<&�i������'t��'���@Ř	
��)S�`�#R���'��_Y}�'M��|�j�jz�/hP�YRGQC.��#�OJ�.�ƌ	*�8��O�Ę�	:z��+\#Y�1p읊/��(���_��'�"�'}���	�V�%0�U*�ʅS-$d�U�؟��ش��]���?�c�i3�O��8"b�%�3S�%�F��W�+1��d�¦�ٴS�V�DQ`�&���Jפ��Vj�E�
9��1�F5	E��D.G4BP.�$������'�2�'���'��;QG)S�����+p0�R'^����4M6�Y����?I����<1chٯ>Y��p�CE�M�6h��<�����X�I7��S�']Ԃ��o	�<�(*A%��w=j@q���h����'�z���G�П,���|�W��ا)�2f\�H�G�5b@�*� _����I͟��I��zy��r�r䊓O�OB�⩌�H!�U�����a�O�TnZy��4���ß��	
�M�S-��W��)+��K0���Y4y�%3�4����J��\3����Op� ��QHV�(�8ĉ�'8R����9O`���O���O���O��?ɘ��ي�@���@��}d�5Ӣ#U̟���ٟ@Zݴj掠�)O�og�=�����ߊ��@(�"rm��eO/���5���|�d
���MC�O��!Fm��{4Ht�IR��#��52������v� ���<y.O�	�Oz���O~���gW@c��q
���t��O`�d�<q��i�"4�'G"�'�������1��.���yd�^���8K�I� �	���S����n�ja�rF ��:���E.V�P ��C\�L�:�O�	8�?�u��O��Ӓf��HЌ�����,}i�{�ͅ���������b>=�'��6݁xFr���,5Zɢ�s�`B�#��btD�O��D���]�?�^�����~蘉ȇ��>u�^%��`�
o����
�M�B�߲�M[�OR�V�:�*H?�0dFԽ^i2i�qӈBt��{�ؗ'"��'2�'br�'��S{�j���
��$:��bo��[���0�4
@�+���?	����Ou@7=��E��=WE�<:�G�&�4�� m�O���Nc�)��&'���l�<QÅ-x�|�AG�H!|���d��<��nʷ~�dG/����4�^���%����˼>���YG�����O��D�O��ac�6	\�L���'^��
K��j�,�qQ&�JQ� C��O���'E��'Y"OHIǎ��`e�X�@L��P�咟�����h!~p���/�i$��Oɟ�Y4��9�HTbA�ֻ���ȟ0����T�	џpE�D�'n�0@ʂ�b���E�%uL �P�'M6��C�����O�hn�R�Ӽk o��z�r3ρ2V'
�##�h?���M#U�i��{$�iC�ɩU�A�A�O~&h0b'� �$��e��g���A�G�F�	Wy�O,��'r��'4k׭s�l�9cc�9j�ve�F��%��	��M����?Q��?�I~�Fe�p@$õj�$����1X��$W�T�Iޟ��H<�|��V� o(E�&�8=֪-:���4�̜H�fS@~B�1-|���	� ��'}�?;Jh����/C.A
B�~���ԟp�I�d�i>Օ'�"6-�	u����3	���P�y05!�W�j���Ŧ	�?IP���	֟�j�4 <��g�n�B���k��/ �������M;�O��Ф�����$�w��=���C�j�����nǴ�rQy�'	��'��'��'��ء�.~|
ђ�b�.;�X+c��O��$�O�0nZ�E2N8�'�F7-.��H�?�d��F��(7V�o��N��&��#ڴa5��OL�}��i^�I�X��C�e�b�Yy#�K�x��Y�T�?fTb��U�Iy�O�2�'��gU[lr�H�կ|9I7 9ri�'�I�MKdOǭ�?)���?(�z���G�M�f`�3�Öj��Ý��x�OmZ��M#�xʟ��¤�\��uBB+�~���+5�Z/�>L��.W'.��i>���'H�a%��R`Q�]^X8Cb"Z9h�4��Z�p�I����Iԟb>�'�t6Mȿa��`j�"�\#�	�,Q�+���?���
����D�u}�t�J�[v�P�`�0�j�ı0��!Ū���1�ڴ7����4��$ѕ:��:����S�[8��Do��{J]H"kN�h/D��zyb�'I�'���'
T>UHWk�m��2a�ΦV����C�̗�M�vHT�?����?�H~��Xj��w�b8� ̌U�
����`Sj=�#af�։mZ���Ş��|2�t�;���m@qQM������P���hC�j��,TF��Ly�O��c��m_�qG���h���4�F�[ ��'��'�剉�M�4���?I��?�S�0"3\��q�ŤA{����	I!��'���?���Ez�'�I@��ەM�������>o�� �O"�1�!�F�KA�Ʉ�?1A��OLD:�ǌ�>f(��c!-$�^����O����O`���O~�}*��uV���Ūՙ��H�Ɉ%^)�t8�����M�	��	��M���wr��R��1���8A!_�f��R�'��'�7MC"j�6M7?���K9at����,�"a�C k-j��n�
PЩ�J>�.O�	�O����Ov���OB���+P��pˑ܀WFy�Dj�<A��i�pI� Z���IX�Ο �pHR5,Bp�C����e�h���B�����O��\�)�S�	=�e����<j�� �߄�T��V��j���$��O�ՒO>�,O�����ٮ\:�x��
2���K�
�O���O����O�)�<���i,n `��'dؗ�*Sx���GL�ܸ�YvF��?1B�i��O�L�'M��'a�@.|�B$�����0�H�&w�:8T�i���"q��u���O�q���+2�4����VV�X�����d�O��D�O����O��d5�ӵ0A�LI�c��K>�d���ےF�nQ��՟��	��M�-����$�M%��1�@�JsP�Cw ɡ75�)�Z�ēm�F�h����hϛ����1�KE�n��s�ڎm��D(�f'i�2��@�'٠�$�З��4�'�b�'�|�e��g��R�	��5>@1�'�"^�y�4,Q��:��?��������$"��H�L�v��FѹqD�����O�6��b�|���&.	�I8�#�6d(!�A�EL�8m��n�<�)��dD]؟S��|�璾C"p�2�
6*@ 1e �(M��'�R�'>���Q��8޴	��$���'��$A��W�9������?y�.ϛ��dvy�i�\��J.By��U�S��S��e�J�m�z8l�}~b
:Bm�z�� 0���"S��"�.��K�X�:�>OP��?����?����?�����	Ї,���� ��p���b��$̔=m��=x�,�	��x�	b�s�({������-v�5�a�A1�!h����?a��5���Ok�����i���G�/���4c�B2�X$@�D>�,i3ؒ�G6�O��|2�X���"��O�[,I�Ei�<a�� P���?i��?�/O� mZ&1�	���I�G���PC�=�B�!�%Z�Z��U�?q Z�hH�4j!b�x���5A���HWf].�pB�AB���$̺�=��%��@���)�������M�̚T�C��_�F�c�Z(5����O��D�O���*�'�?�IӀ91�m���#��0�*3�?��i�VUsD�'���p�r��]�b�\��IH�(�R�gڢ-X���	�M� �'����S�[b�柟�BTo�$/W���&%��t'���
"�֕m��$��'4�'���'l��'�`�:$��a��MC�N˅NMvy�0]��ݴ5HqJ��?����O<�6�'a���&��JƲ�BE �<y���?�N>%?��P��:sAL9��OO2���r��'yu��2�ĞQybOȻv����I{�'��	 }.��ʦ�N
/Ҽ���+.E�T�'�'��O����M��*�?y�gN�7y@Ձ��2`�|�� �?��iY�O���'`�7�������4D���:�	��W\��A/�K�Ę�#X8�M�O$qX�������w���3�\*i,`�yVi��&@���'b�'���'�RQ�b>Z��B w��SCM�0���:dE� �	��`�ٴE<V��O��6M:��*&�*!����\�.m �t}����xr�'e�O���i��	%UH�!ae�0�Xq����߆���Q���P�IXy�O���'z"�*N2��0�H��a��Ȳ��U�T���'��I�M۵�Z'���Oʧ[��E1�/
�kMdX"MgQ^��'ȴ��?�4G�ɧ�)�z 8-x㨝,q��J� Tcfdq H��\�jǕ��ӕ"��v�	�D^�q1�Z{��!�?Np��Iџ�������)�Sgy""{��X����&:,��_�{V)@�����vқ��d^q}�'�� ��"�M-��'��J9�'$�6��1T��7m.?9Fئax��-���V-'����S&yP9PǭӅ�y�X�4�	����I�\�Iȟ��O{6<jW@�N�;R�Dq�@Xci�zի�#�O����O�������ͦ�ݺC��(�&Ѩy�AT�7,��ៜ&�b>9j�.�զy͓bL@�ToT�Nb��.\�H��̓@��ux$��O�u�L>I,O�	�O��#����1�2Щ|xV����OP�D�OZ�$�<ǳi6y���'�B�'���葭
�}�d��aU1'!��;t��GQ}��'i��|r�ޖWT԰��W�"�ʕ��4��D���XqA�ïlj1�8\Y��ij��Dٞo3,H����pXT��;����Ob���OP�$>ڧ�?q#d�($�|c�g�'	�¡&B0�?�@�iTt���'9�j�4���h�� ���m( ���J��9�M��ii�7�@*Ү6!?i�9��I�D̂��E#�6�*`1��T+d�Y���<ͧ�?����?���?�F�)&�]��߶ol��
���ʦ{��L���	П�$?��I�M�"�@��/������3D2�`�O��$�O\�%�b>u���(K�A�b뇻.������:[&�B�5?���}�>�d	�����E*	qDt`ta�;>��4�Eʗ7]v�$�O,���O&�4�l�]�6��./��Y�D�$R���(mBb���i)=l�p�6����OD�lھ�MC�i�\)0�P5�Z�㧌*G��=�3.��Z�敟��7#�W������x��tE�
�t 2�� l��
�4OV���On�$�O����O��?�#��<���9�i��>r`���������ڟ<j�4^Ũy@/O��la�	#`�b=R!�)F�|0teԸH�N<����?�'_�,�rߴ���0}����'J*A�a+w��x�jAx�.��?��8��<ͧ�?i���?�D�K�_lF�oڣ!~|�CuQ6�?����D�������dy��'��ӥL6�P��5T$�}˃��!()��d�����\�	@�)�W�� WZPXQ�Y.R�(�	���z�r�C0�����ġGǟ4KW�|2C]N����5� #Y�I`s#����'�"�'���\����4`�ҥZ�#��Fw^Pb�]��5����?a������z}��'!��F�F*Ϧ=XK��%<V�q�'@���Ŀi���Y�l���Od�_�|��C�5Ґ%DM�#;�<̓��d�O����O��d�Of�ĩ|:��ev�TWiNV$�Ҥ{��-T5
�����%?u�I?�M�;F�舚�L*?.���#[�tБ`���?�J>�|z���&�M��'����+�=u�, ��Jױ_n���'��R��Bß4�U�|�[��S��|#�O�ZZE��,8�n�j l���8�Iܟ��	ayB�|�"4pd�O�d�OH�*���n ɺ5�Y�r�v���%�	)����O�d9��ͅY+����	H`���©X��2C����@�S�b>����'���	�'pzlj0&A-:���v���;�D�������ߟ��	T�OM=x_z���4[��ɹ�H�4}*�m���u��O��GܦU�?ͻF,�Z��
]
p�q���)-����?�ڴ��vc�p枟Ш��đG�4�7� �p�5FڷJ�n}1ǅ��H@��Z�)�$�<�'�?���?i���?y �L&C�D����F��t$U+��$����``O���I��'?���*9UrMy�L�x�NK1@�%�`�*+O��d�O��O�O�VB�Y�G�@����ØzJ\cs��6�y��_��)��(��[m�gy��3�t�B���; d��"�Z�*�r�'���'�O��I�?A����,�Vl�;D�6Ha·c7�8+-����ܴ��'�˓�?1�4AЛ�ŧh��{�l�*��`��fޭ"q:U ��i�I�y��cQ�O�q���.�>��ш��_]=��c��,��O��D�O*���O��;�S�vNtx��ʔ�tp���D ʡ�i�'2��yӾ5���?���4��5;t�ɦLޓu�f�Bsd�x{�1��|R�'y��O7�(Y�i��ɛ��\�b%�$�H��EgT1O�x���/\�D~�Sy�O�R�'W����c��!��?F�J�A	;R�'2�7�M�%臱�?����?�,�$3p��{�BJA1"05�4��@b�O��D�OT�O�142��Tֿ7�p�H��A:H�C#&ȿ~-8�z�-?ͧw�P�����Y�*91�-�mĮX�v��8>|�����?����?1�S�'���Q:�&f�ƌ�P��M(ر�e��!Vnh��؟<aܴ��'P6�A����V�[Aˋ2bN�Ԋf����6-����ƝƦ�'TY���?���F1�!����5�ƌ ,�����0O@ʓ�?q���?����?����	�Ȱ���!V�aU��:v�Po�?�����˟���Q�s������{FFך%�����ƅ?5���S ޡwg����O�O1�ZY1'�eӮ�	�
V(\���Ʒ!¡0ĉ�
����ul C��'��'��'���'nD��rK0{'�M��B��@ZS�'��'�2Y��@�4($�����?I�����#����i1 ���R�$J��k�>����?H>1�
�E��B��#Q����jK~B�F�5ٶ��7�U��Oδ���
>����[��H��(�Z���C��E�B�'���'�S��ST�ќC? X����>F6q� ���̸�4# h1�+O�unZN�ӼÅǟ"$�)��q����A��<!���?Q��i6����in�I�t�5�P�O�|lDoէ+�8$ �E��|�4̊f�Fy�O���'["�'�2'ʆYBTP�!D��h����)��^�	�MC������$�O��?)R��J��ʎ
(�|��@����Ц�a���Şg�H���� E���(���!���  ��t�rM.O��K��A��?�5e1�D�<Q�b�'NX�Kդ!Ф	h])J�d�O��D�O�4���$��v ��%N�.��t���ʌv�2ŋpGñol�l�6� ��O�ln�=�?��4x�}�G-�Ƥ����<�@���J�M+�OL�B#���Q�)����Dq�E�M�t�T8�Q߀�Z��3O��D�O����O���O
�?�B*��b��,	u��+��!�$IE���	П���4P���'�?�b�i��'�Ơ�A�.��<punݐb:�)�5(,��X���޴�z4Bˌ�M�'rh��p[Ƀ,/gj!�4��蜵�%	������|BY������,�	��P��lQi䞈۶^nV�I�!������py��m��J�h�O��$�O �'8h}��Z�S� ���N-`.���'����?����S���	I��]d��%��%o'y���A�x�|�8�O�)���?�q�$��c�3���*���BӺ_�n�D�O��d�Ot��<F�i΢�Ղȁv+��� 	�����Ð1_/��'�6-?�������O|űC`�ަUc�@���E@ ��O���E"�6??��@��c���)$�/J%t}tq�
��)�:�{3G��y�W�H�	۟��	ٟ��I㟼�O.T�� L��;� ���ղ�!�:2����;��'"����'6=�52���J����a�#~7�B6��O��D0���	vA�7mv����n�z�0�� ���5���f�t���W�#��Ic��Oy�OgRʁ�W�Db5bI3}|Q��E�@���'8"�'B�	=�M�É�>�?	��?�!��A���J����b��b"����'S���?I����+p.X��Β4��q��k�Ф�'jH�#ΰ!�0�ɏ�T%���g�'��h�l�6"��{ ����;R�'���'���'��>��	��-��(����āS��|�����M�iL��?���;��4�&�3GT�H=�%����]��b�3O����O�Uo�n�*0oZH~B�Z�{�F��S�8I���7���;�z9!&B�u�Za��|V�������֟���ܟ웅"ϪT�`9��H��6���rqH�pyB�h�DkD.�O����O����B�/��8�bH߂,�� ���?8h�':R�'��O1���M�?�B�&�Ӯ���rK� n�D@�#��D9��: ��GH�{yB�
�WC��9�Bĝ6�A$\(uR�'2�'��Oe�I�M�q�:�?!qF��Z���� )u|�����?aдi��O&h�'J�'!�㞧
��#�%�I_�d�	@���x�i��I' m����O�q�x��H�Q�=sBK�d��a�GfĘ���OZ���O8���O��$*�3c�|h	W�	�L��Y*���&Ae�=�	֟0����?�&#z>e���M�N>��$�{�pI�7���0/��AX3jL�'AZ6��Ʀ�S~�qn�z~��I� �(�"m
-~�lbUK,ά�BV��#�?q��(��<�'�?����?�F)ɒ-+ #r0VtvMٲ�*�?)����$���C�A�Yy�'Y�ӣ	C�`U��5�N���DN� |�	/�M{�i\O��F���dF��K�]�!ŏ1o�Jei�f���$�4a6?ͧ����,��K�*�Y��[:MA�'�8�
�����?���?��Ş����eI*�+X~�e�_hh���=Π��g	ky��y���XҮO�oډ�zqI�	.o�H!A�"ez��4*K��cK%6�֒�DYB�],e��~�pk !-���UJK�Y
�0�Œ�<*Od���O����O����OR˧_-pX��M�,���U�6���׷i����'��'��O�2�a��W,I���Ǿ���B�M�mOx�m��M���x��I�R	��1O�	 �Þr�p���o�S�`�1�3O6�2
�.�?��)6�$�<�'�?�$�E,u����t��x�`�a����?)��?�������ћ��]��|�I�IU#�j�t�dhP
R�(:�`VR��r�O���OB�&�ĺ�G�.m���r�'���9S�>?���E&!|Hq�i̧#v���)�?�FE�YnL��N P�� ��Ï��?	���?����?�����O��z��#�f�Eƙ�*�|��C�O.�mڛ��4��ϟݴ���yG*J�/��xr���+�l�f@��yB�'��fӨMˀex��|4�a��h���}A�L9qH �%�
X��zc������4�����O6���OD���9�\9HCiVsY❻��5,&
˓|)�V�ޞT�B�'�R���'�r	#q@Z�.�>�ҬӌUIpٙ�˵>)���?	��x��d����XȺv錢���̎P�]�́#�����3 J�Od�L>(O������>�n%�tDO�o��L����OZ�d�O����O�i�<y�i��rp�'@�-��1(���{��yw8�1�'8�7m3��	�����������M�4o�}����B`�HȈ93���
VR��4��D��r*�c��c�.��$�����$i��'ƫ8���"�&F��d�O����O*�$�O���$�S�$���Ss��:-kP@sc��:;�L��	����	'�M�"k��|���zM���|"/�)BXՈg��tæ%�1IW�S��O�Hoڌ�M�'D�L�cٴ���^0�ZT
b!�!� ����]\�R���?��( �d�<ͧ�?���?�ÌR�vT���/� �0����?����ঝC ��$��ԟ<�OG��jS!6�Ȍ�­�(3l�O��'��6�⦩�L<�O?���e��"�
(C�F�T�鰵�\u`�sb��7��4��Ģ�e�ԒObA�S�%3�T���"X������K�O��$�O���O1� ˓} �V$A*Z��qq%� ���;�@Ni�=�%�'sb.}����O�,o�,Yb0IV�#mNjM���� #�d���4$ț��\�f?�V��0A�
Q�mF���~r�IP9���!R,åz���A���<�+O����O*���O��$�Of˧��R0���]Ere�ǔq9J"�i����'���'�O��Ob��׃;��P�C���TC�Mw�� ���D�O�'�b>U�
ϦE�|y�1@s�ؙuR����74 ��͓5w8����O"pKK>�/O�)�O���tϘI��3�AˮX��lB�)�O����O��Ġ<ie�i�Zʐ�'��'D .�>c�8闤�2C�"x����A}�'�Ҕ|�㉵�\����|e�U:�.ۿ��d^3}� -�GP�z1�)���p��,F`
h����s�(4S���G�Ot���OV���O �}R����a)S�!#?�T��֑z�٩����fC�j���'&.7�%�i��맏��ti	�L��Q|z ������4#��-t�f��F�r�h�o������ܑ�p�ߐ��ԠA�0u]2�p�HѰ����4�4���O����Oz����B��rf�o��I��  3�ʓ<c���Q�B�'-r��T�'���r���5%�p�`}i��<���Mc'�|J~*����Goj�Q�̐�/��eJ�
B&�j�&O~�;�*d�I-+�'��	$�!B(T�%P�y���%?A8Y�	柼��џ��i>��'��d��Ns�덥m�ِ�F��F�����N���yr-r��⟖ay2�'��&�m���qb��#j1�8�'�OqXUhdl��
y�6-,?IU!��<{��	8�S�ߝH�����2`S�C�TY�es�,��ޟ���џ��I֟���Fރr)�D�U�z�~�2FLP��?���?�ջiC!S��pܴ��j*�� ��O�zG,�.���醒x��'^�ON��־i���5����	)��
�ύ;?>��'$P� ��i��|y�O�2�'�"�O#a�����M��2�`@Q�	�)b�'��I4�M;���0�?���?�,��0�
�<$B�*Q�1���O0�d�O��O��'�rm��͈�<�LA���_�l���q�)W�f-~$���>?ͧw�P������,��գD$FI���;;i�hq��?���?Q�Ş���JЦU�5K��b���`��vϠ!i��I�02v���ߟ���4��'<���?��˩�x�y"��(Hc���v�HH��ȟd������'!�a�e\�?��:�"�c/q8�PZ�)>5���G1O:��?���?���?)���򉀼l�`5�.��X�6Q�T,F&vf��n>m��-�	����A�S柸p����%�%1�H�`�;:F���E�?Q���S�'	i$
�4�y
� JT����\V}ԭ_>lW�4"�3O��AgE���?�vE(��<�'�?���QԒ �F�+[����iS�?I���?�����d��ғ�U�x����g�M%ǖMRE��/oX,$8���s�p�I��M���'܉'E��P�).3��QI$��<Њ���OP��T�(L酠!��8�?����OL=��I�*y�h�a�N�0WLdY�N�O*��O��D�O£}
��!��IP�ڱ_�̵doR=��LC��"�6�Wv���'l6m(�iށ��SQ�舋��<��#��w���4���i0t�i���=�ʩt�O&0�"�I�Q��`��I��Ѹ��Ty��KyB�'��'��'��ӳ
��PSH[�;��M�S�HI���2�M;P��?����?1L~��N�ڭ�S�ۺ�9'���L ��TY�\�޴�"�x���*�lm �J��Q1�A���>1�̘P��J��	3ds���'(�&��'sz%�.ݗ.�2X�pǛ[;����'�R�'Ib���]�p�4W$؁��SQu�C�^�٢�v�Ǭl�͓5Û���uyR�'��jj��F2�0r��Ȃ|���#�B�f5�6+?&B�M >��'���0AO���8��I�4�{t�c�$�	̟ �I����ݟ��R5(O *�\#hJ�\��hZa���?���?�7�i��;�Z�l�ܴ��b��A�Jրr�Tx��]�'ЈbF�|��'%��O_4��i�I0K~ � �NL
pVI�D+L�($�_ �"��D��Oy�Od��'"�� 'V2H#q���$u����3g��'N�ɀ�M����?i���?)*���a�<��H�Bf�,1JFY[���D)�OFPoڿ�M3'�xʟ�X�5�*6x���T;R@�ip����Qb�X�GN�i>�Y�'���&��� Iêqad��r��1;��4�'AV蟨�Iɟ�	�b>�'��6�X�����.]6 =,�0E\&(����`)�O����䦭�?�TX�|�4Q}�8J�ȝ_J����Z�_�Č��im7-_�^ 7�'?I�H�PZ�	8�$!B<tC�!a��2���	A��yrT�H���L�	ޟL�I�p�O+�l�u!I-,)ꍡ5D�6�l�g�n)��e�O��$�OD����D�Ԧ�]?C�	�BC�Q�r�`Af*$s�u9�4QW�I4��q��7Ms����U�f���W���� w�@P�f�#"ɏM�	my�O,�GI8�x��D�(?<a�Ff?��'���'��	8�M+6n���d�OBm91�V/j4ܩx�&.�|�� B5�I����惡Y�4l��'9v��ק�'|�a�W�x����O�#���c�j�����?�O�uؠ�Ö`h8���!u=�"T��OB���O����O��}���E����_A��!&��acl�������.-pR �s��OP��R���?�;w;����QN�@\Y�Y|ʌΓ*o��/u��m�k@En�O~���  ����'7�ZAv � �8�0���5S��|rZ��џ,��������0�T�C�W��VO_0sP���Q"�\y2rӢ���-�O��$�OJ����S�0'�M��c��-�:e�c-�.���'{7�֦5I<�|��eΐ2��=a�f߯g�D�N]�_��9)��G~"-��\��m�	���'���$U��� �b �5�\	ز��|��L�IП��Пp�i>�'6�TY\"���' ��ȩ���:7���«��R����L٦��?�#W���	����ܴ}z��[&�_0n���I�%O`T�%�?�M+�O�<aT���B����@*B������"w�y��o�,`u�5/L8r��qҗÝ|�n�a��W�BǪT�v�,k-��agm�8HVՋ�*G.^��h��˖<c�4%�5�ɲKd!�5K�8#� �G�D����%Yx�	ɣHR��u�6�֧llJ]�@	��2�Ř1�S��6�j�%Ҋ�hL�"JW��d�Y��ѭxD���Ŀά��"�K ![ٸ��Z]n�ڃ���&��T��d��m�m �f�#$2ˣ�N.=c~9xf�Nu>a���*
��$��a68�(K�1d��@b����)�	֟��^���'\�S͟���xƴ�r��Әe;0`ߜS@�p�󄊨J.�'>m�	Ɵ��ɖXj�(6��Щ��>�l��6!�{y������<I����cy69��ȴZ���K�g&x�@��c]�`դ��@����?a��?���?gJ�'w2<D $���x��3�fS�vy����?(O���=���O��d��m�³��5�8�C�B�@��� R�C������������џ`�m�H����_`��.�	+��H�q�'|��'̓0N��(�4_V��`����-h�c�-RW6��'}��'|�Q�TȲ&����O��u'(�Lg\�uh��:�b�ꦁ��]����D��=���[�2`����F��,
C�˦%�	D�'b���Wå~���?���~-D�A��;]y���U �:~�EB7�x"�'t�J���O���5F�x� )u��3dEe9�7�<�)ԡPa���'C��'���F�>��(���摆F,^�sg/;hV m��8�ɧ8�&��	�[���ָOwT}�(
�b�U���ͽN�PL�ٴ��A9A�i�2�'���O�.����M�_"�!��R�! ��EQU]J@nZ9wZ"<��T�'7��g��:he���S;2�.� �K{���d�O��dH=7E�d�'��X�DҸV�m��*�[8%��5�*z�D��F����wh�t�Op��'�Zc�V��*۳6X!��<��A޴�?���J+ =�Ieyb�'#ɧ5�h�>�`hXa�TBR�Jv������'w�l�O����OP���<��� �Y�d��?
�69��bϘm��	B���*���Ty��'w�'���'��iV���f�*m�᭞2=$�a�0x��F9�y��'\��'k�	x�z8��O�f�zE%�9`)B]چ�1F���ش����OʓO����OҨZg뵟�k��ۣE�@�cόIc��h%��>���?����򤃈 {��O��ۨ6�\-�Ƣ��0V �P�G.�6��O�O^���OA����O5��]�L��X�d�֘�B��;v�`S��gӨ�D�O
ʓ3]�uI`\?�I���S�bDɘ�bl��J�O�R�&� J<����?���U;��'2����:��2L�p��X ��%j+�VR�$"��Z��MC���?����j P��X7f�d%9�`�8.:!�7a�i 7�O��3�"�<�}��$��d�4̲5jG�H�ڸ����ߦE���0�Ms���?����B0[���'H�Ђˑ�2��)w�o�����<(���O0�������W��|J2�[!y���b�F�W��iub�'_2��
q]:���D�O��ɼkܰ�{��A	od��N1_c�|R�KV��ן��Iޟt��"%��� /�3H����j���MK��7zFa:0Y�|�'�BR�x�i�-��%Z&Y&����E�м�F-�>�dK��䓭?����?�-O�$1�m]oT�,�AN�0���W�����%���	ӟ $����u'A��oB�|ʷϝ#5�d](�L���M����O���Of˓���b1�԰a�S������~� c�Z�h�����$�l���$�'A Y.m~�(Q�M����j4E����	ɟ���@�'=Z�`��?�I?��qSvg�3�t3����K��m��@$�D�����'��%��%��S`5�a��iY�oZݟp�	`y"��c�����D�k�]�8�u�V�I��2 ���mƉ'�I��t�I~�s�֝�)�@ݒ�mQ6:pk��ĭsJ��?B
�?��?����(O�.ӥp�Ib�� 3n\�p�?!��'M�I4w? "<%>Q�����r�0K ���`�~b��O�D�O������S���^���$�@lU�P;�ۍ_� �^���Dx��	��H6�eXF�<�DYG��eIڽo����럜Iw		{yʟL�'-��� � `�Z���XpV*x� �1Pᱟ:�䲟@h��X6!��P���۪0i�E!��xӦ��3$ِ˓���o��$İ�&� ?,�P����E�xR�ƍҘ'��T���I�%��X��Q>3�F(��d��wXhxG��ey�'���D�O��I�l�J��4h��$���;>O7M��
m�I��	ǟ�'�Z��sJp>K�>���X�5�ܬ�'mȓqs��֟��I|��Vy�O���#!�n�7��<�H��LD}���?���?/O6QʕC�i�S�[	t�i�5���{�A�?�F��4�?������ON�'�?�J?!(�+�Y�v`j����L �\��j��d�<	�M��-���$�O���(Z�!WC��� ���m� t���x�'�B� �H���y��(��$M@�\pk�A8Sz�K�i���%$F��ڴA�ʟ<�S���Jt�1H��!���C��N��VY��b������O|�I~n�=M�P�ǏH<j,����0zH�6M�,d���$�Ol���OT�I�<�O�$P�ǜ�f0�ӁCV��L# d�5ɂa�9�1O?A1珖&+��2�A�\
�������Ms���D��h/j�S�4�>!פT�L���d��t��Uz��ɩ�1O��{)V�Sʟ������*!�i D��%��X�����H�+�Ms��d
"`� �x�O�R�|�fe���b!*�1,(�
ĥ� |9��V�a�����?�*Op���\\}.
�Ճ��\j	�e��.������e��?����@)`�c�$`/p��E&��6z�A�4-�	���'W��'+�?�i�|� ��?u��0� ʔ%htu�@l��]�'1�Z�X������	��u�|�V��.ꀀp��Q�#�R�*2����M�s�n���?Y*O���%�Q�4��5I��;t�Yc���z�CPʟ��M�����d�O>�D�O*�:';O�����@p3�6\��`!d�7 �H�"�j�l�D�O�ʓXe,���W?-���$�Ӡ?jn��tHH	M/~�+��4�ڑ�OH�d�O��%M0�<a�͈�������Oq0�i'?�|�ـ����M�.Oz8��Ʀ����t�I�?a٨O���H�*�R��o�p�`�5���'B򪞘�y��'��	wܧY��8�$C+i�R�5D�?M	P4nګ��Hs�4�?���?��'���Zyb�.x�$�0sc�-�ڥ�Э/��6�8z\�1��8�����d��o���"�ʳ`�䡂d��M���?q��h��5_�ܖ'x�O�A�!�N�`�n�����w�4��\� �'Ŕ���O���O����Ot���-!�Щ�Ɗ�+�H��Q�릑��."�޸*�O���?�-O���Ɛ��f�H�5�VU#����#f>�R T� ��x�����I˟���Py�M[/}R�y{��_16��YS/�C�J�اj�>�-O��$�<���?���q}@40qFg^��!�_"SG��Y "�<1���?�됡�?9����$�@�ƍ�'k�99���RڰM�w�U( �"$lsy��'��I��	�L�mp�8sB�)�F\�%��R`��h���0�M3��?Y��?.O���ςi���'�� N,3�KH�2"��Ȱo�6a��أ�i'bW��I����	�k���Iq�dJ�8��ըT��r׀ !���0q��F�'�B^��T�O&����O��d����z�m�_m qkf˵~��EO�i}�'Y��'��58�'��	�>G��':���굀Y� 0Z�
u̟2e�inXy� �)cB�7��O����O��I�r}ZwF�1�G�i�j�n�i d�hߴ�?)��>@͓�?y.On�>u8
�	S��!��ڢ>(�@��|�`Q������ǟ8�I�?Y��O,�L�@�v)�Dq*$jH�KUp�0��i ���O,���O?r���Q��N�|�,	��N@��l7-�O���:�FA�ej����O���f��+WF�A�Δ�b� L07�#����^o�?��	ԟ$�''IV�XƁJ854<�'�Ήn\�Ln�ʟ��N�8��$�<������Ok��).�j��J\57��CM�:���<&|������I֟���˟��'v���	5,p�0��,D*�#��	zt�O���OʒO���O��un����@��	���!U���<	���?������ Eb<�'bX^�a���@����8m��\�'��'?�'��'���%�'�x�)���Z�Jl���#32��6�>����?9���DH�l&>5A�F�Mt����(��K�����
�MK�����?A��_��͓��:Rj���Wu��؂u�P�oy�6��O`�ĺ<!�]6�OS��OBj�c3G����LA4K�Z�!��(�D�O��d)%p�$8��?�w�=,f
��cJ/�f!�׉fӬʓ6.�|��i�h꧳?���c��I�bY�㵀͕|����� &�B6�O�$�'\����8��=�Se=��K7E/Kx)"��$�.6L,Y�*�lџ�I�`�S;�ē�?��̙a���� )�O�r�!�&���lݎn|����O.�Q�O=Y�(�#! (�I�!���	�I� �I�i6d��}��'H�Ė�I`Jl�q��F��=����(�|Rb��y"Y� �� �i�5���[�xS\�@�é_`�`*�yӼ�d�43idm�>Q�����+�&�(C�D�s���qIF�n�g}��I�yZ���Iܟ��	hy�ۦ<Z`����^�.;��f	/Q��@�#j6��O��d6���O��d]2}��E閼7�|�Ӈg�BL���s
=���O��d�Ol˓]?�5y�:�zA�EN�~Y�[���"z1"��x��'T�'���'ՔQW�'m�HjĪ�5jT<5`�ЬI.��&�>���?q���к,�L&>�jE�
Fc�0C*я9�8P���S��M[�����?Q�?�ؼ�����IH��)	���q�Ұ��lާHF6-�O����<�d%K$8��O���O��顁	�6m��9�/;m�	�!I0��O���δJ��5�d�?�{�jD�J[����/�:j�>|3 "s�Z�|~U���i2맯?��'e�	8F:Y�Wϗ��L�i�$�/4 7��O��L*=�D&��0�S�u���4mA{e�h��6�ʤw�(�oZȟ@��⟐����'��i�0 \0p�a��I�J>�3UIk�Y3�1O:�O�?I�I�pj$����C��c�5YT�)rڴ�?���y��<9M�On�d����
�� `��r�	X���t�h�Z�O\�!1�Q�矼��韼&a�{P��C熣fE:�IK.�M[�'�ذ�x��'r�|Zc�xԻP�S.\\&�I�4�x�OP,qV5O���?�����Jڸ� ��ߢ-[pz��ʨ~q�10��TڱO��$!���O�����aX�2�!0}�\��R�� *T2�դ�O�˓�?)���?�.O(9{Q%��|b�/�c���02�E!,]0�jBi}"�'L��|2�'M2�&�y>\2��Po@(����!��%3L��?���?�)O���� �]� ]�5���y�TP���A�E���4�hO��dV:fv��+}�o�D�a��HN"6ġ)܊[�'`�X�x�\e|D������k��Q�8 �ά1�Z=��E�e*�O���!A���'�T?AC��b6�c�#�>d6�y�3�f��˓
WD%��i�l�'�?i�'���Kdp�d��p=�4���KO2��?�l$�?AH>�~���ޚd^1�$EB��T�Qł��y:	B����ߟL��?��	͟�O�֤B��E��p��D_�_�	��{ӂ тmJ�11O>��Iil��c&�:}4��I��-��ز�4�?����?a�?���z���']rC�+np���ݽf%��s��7y�c�0�bd=�	˟h����T�1iB�Yz��d$�,�ʜ��,\����4*b�'��Iȟ�$�Л�e��$��qj�a�:C����-58� ��\��Ο,�Iqyb+��J�ܜ�V�z�Tp�D̠P�񠤤�>/O�$�<���?�~E�83D郪S�Nxr�wG��{Ć7������I����'v���w�m>m{� 	b0������:`h�.l�ʓ�?i(O�$�O����� ,�Ĩ���Z�hW�0�7LH?e��l؟���ԟT��SyB�+���'�?	�n�6
�B�!�T$2]�l &\�V�'/�I��	ݟ��0�y��O� ��Tҵ��;B������M����?1(O�`��D���'�b�O�"  # �-(M1��OA���ŧ>!��?�\J(<�����?����^	�2���J�8n-��hiӘ˓0g^��F�i�B�'���O#n�Ӻ� hT�VGK�4	��AH(X�\0� �i�r�'�� ڞ'�]���}��E �0�3�J�(�bp���Ϧ�"a@��M���?����_�Ĕ'*(� ���cy�@	]6���baj�6HK�;O.���<�����'�`Qq♡#}�̋5�%Z�%��/g�����O��D9dv
��'}��֟X�(U� 0!��j^�t�G�rDn�ӟ��'ڈ*�����Or��?ib�$W(���)�F�� ��iuӔ��
�= ��'��I͟L�'�Zc=���K�; Pv���`ųqj�8�Oph��=O����O���O��d�<Y�B���\��U�u��d�C �-xFP���'W�]���	ϟX�I>r,��t#ؕ7�@������}�D��۟� ���Y*�NH��)�	!r�@��SJ#f���b'� oh!���#�%�#)K�C݊M���]0^IqO^d���X�'Y�H���NV�Xzf�H�����R�������To�hZWd�
�$`*!��3�r%V���Q>!���(FR(�p�Y[�����c�8���k��z�� ������ل_�9	���#t��)��7R�Œ���h�<�@E�/���G�irh��������p���#|�%�2�S�*�3��˟\�I&
��~�S��O�x��9��� ����֪4}��w���O ���,I�F~�,C�l� �q�I��I�J�O��d"�I9�	�p����S��+_��2���M�1O��(<O �	"�I����BF�&c�sR�'�"=á�-z�f_�\Z�j�%�0�����F�>�y��Dş<�I����iޅ�� y��f�çW#�A��ٓ#�{�Q��c�*��@b>�OF�k�)ޞm�2�����1J�T����� �C}r)��:0��}&��HrDJ�Mq��ٔ�ʘGgeC�Hß��'��0���|����H�b��c��h;~mz%� S0!�$� ��L{!l�7�4�����	��HO�Scyb�G�I3:0����)#6P�c�T��I+�	-zH�'���'1:�]֟ �I�|j�+Z���0�Z(S�*
�*^���@+���᱋�(r̢��	��J�x7fٳXЄy0�L�)Аa��@ց���t�Te�	ϓC֙�&G����� ��@�ֹ�e�JП��IA�'�O�����$7H`qc��1 :̜[C"OT3�0[z��jB++��(��T}2Q�h,���M���?�� ���-�D	��ːLHD�̭�?I��X*��?i�O�l�Ғ'	�5��'E��X��^� O$\�d�@��8�8�S���0s�Z�ē��h��,Qq�|ՙ0���l�XI��3Dy(���Oz��O$-`Ũ�}e�X���ɓhyj(XRƲ<����������M���9G���W\v��3Odn��C�9�ʟ�C���fBʜ(��	a�����1�Qh�l���34�%K� �"O�,{CM�:�4AB�Q�A�Й�"O|��FI_�^�X)K�J-9
�DA�"O)�'O�bX<	��K*$� P"Oz�s�F�.|�Mk��%���"O\����R+ؕR���L�|-�0"O��E�O��<�(F��$#a&�S�"O
1�VA�D����U�5"�"Ox�R�/2)�NqCS"��e5�@�C"O���,�t&2��ӊE�9�PH2t"O:)�$E�Egz���J�B�$���"Ov9T���h[��xc)�!���"Op% ��$Y� a)���m�r�"O`� �F�8� ��g,�%F�����"O��*���z�H1�)҄��%�"O�$�I�2�A���� ]~�D��"OP0���?��X
���i�-��"O�P��dŴw��9��_14���"O`M�G�X};��m� L��"OΜ�3�ċBn�(gI�G�^XJt"O�y�뎳K��SW�hx��"O�H��$T� ˂p4���`Y#"O^��0�I�'ttS��O�R6~ld"OTpҔ.�{�!
l؟%�Đ��"O^�s�,�i$���\�����"O���%H3��p'�ёj��p9�"OH�r�'d0p�&HB7i�R�X�"O�-Be��
tS&����R"O� �x�
�6
Q�}�1�\�Y�`��s"O$x*��!l��]Rd�l�`���"Oƙ+���(�|����1�P���"O�#%$�`d&�@�OJ�l�ptk�"O�m �["D4�ű���)R¾��"O�`#ҖA��ũ%�o�h��"O���!�Z�f����@���C"O�jB�H�!�HiS�h(��ˀ"OA�&�۱8��1ۺ�R�rE"O\\��/-�������^1pF"ON������&� x�`Q[���Aw"O�eB�Kx�6I�w_�T|�p"Oh��N�&�����K=�I��"O���0+N*����`k� β�Bf"OD���KVt�4H�'�ĆH�a�"OH�YH���]yԬ_	Zƹ#�"O�آŔ2;L;u\�2����Q"O��jL	�.qTmb�������"O�]��|5�1�wM��|Ɗ�)�"OP��&䖯T�@�[�n�$9��s�"O�u!E���K�F�>�� ��"O�a�!�]7�a���,�0�"O�a2�hا8WF}s��)j�X!��DL/�� G�tmM	�$:%�/W<�a��ʎ�yR�]8�|zJϘM��48���i���A�d;�g?	�ܛd��;��ϥ2�ZZEF�M�<A��/k�$��ᛜk��9`�(���vj@��0?�s�A`�U�S&�?��"��3|O�Y�c-�iy��$�:���5e>�����y2�۫lDy��4M�I�	��'� a��a3��9Q���8��Y$��	7`Y��#{����9)
}!�Ɂ&O�Hs2�ٚ��'��>�ɕNJ��`��
"��:&��f֮C�ɧ;^\�y��9�l��oD��牜S2L�����%�d�^��t����P�J�ȓ\�� H�c����Bӗa�,�ȓLx��*���1���1��������z���`y����Y�6��q�ȓP1��A�MX�h,J��r{DA`�<�Q��U$���p�*�qPt�Tg�<��c
� +�C!�L'4	��0jN�<1BK�hl��2��K�I+B�QD�<!ザzR�B�
�E1���5NA�<qD&��.��̳s�_�6X���"O�eRP�E$v��`�	ހ`b��""On�Q�+�G�F(�0 f,��"O�2���7o�%#UA׎k���X��>	ƪ����=R��@L�#g̗"ȑJb�H��� �bI�����~X�%�	�+шx!d�/D�*�n�z�,0!�P�|��#+,������I��=�[�dT�A�R3\�`�
�'�)Q#V�Wi�陑K�1v��u��'��
S��S<nz�mH%ɖ�R�,��K�B��C�IRI^�z�!A"%&��ۇ�</Vh�'B\�7�'n���2Ʌ�a�����V��yr���Ey��ʃ�7iX�,�Pb�y��԰qN,�$�]F��B�'�&�y�KTFD��)�ãPN���O?�y2L�r厌H�&�N��\S/Q2�y��� >���H��@Ƭ����y�˛�jgV�)���.�,����y���U�����D,+S�]��BT�y���7�����ܤ*b��y2hO���C���X���eV����� z���%!f��Y�2�K�Dц0�"O�ea
_�_.��R�U�"�"�Ѱ"O��{7@J�mF0��ҥR�zBM��"Of�*�lT�s�8��E@�4�6@ a"O��(	�!_�s��$@�L<+�"O�-0�+�$���j���>#(���"O<u1%�4U(�aC`>8k��s#�'xୃrV���q�\�L��v��J��H�&7D��%n�7-n`%����è�Hg6�^i��p'B,�D�^eq�G��9�Nd��a��A��i�ȓ^�����*XlH� +(zD�!gM<i0�"~Γo&�����	�([��T\��~�z��	� ��J��_�)͓hpb��>�O��*#E;�)`�i�#uG�q���'&9Ps�
����^�L�F��JZ)/���"O�	��~�]�%(��\v�� �$��]�:�0#�
��h���;��;0�,]��G�%��P"O�lr�M�9߲M9t.X����'���ߴi��A��@˧/Y�O��kt�D�L[)��R,B[�Ј��'�i㕇��7�(��͓�>e�y���Y,NT踱�͔�9\<�W.�j��Ą�,��IѤm��V�b��dG��OQ*#=����:w�I���N ��a���h|�I�x&�c�iͻv"�+d+�!�dZcꙩ�ӮUR����Z�4Ǜf�Rw}�A�1�RZ<P]i��ȔFF<�E�\cK.���e^�n�Z8@�Ԕ�����'Dl��A�P3��i�fT�B��`A��]$4��oQ�r�V�i���������'������LL(�%�5)\P�	�*ڨ�x�K&~L�:W��
N@Y36@B�@0���3��Ph���u� ����TW���WA�f��i�3Mء$��4b��C�o�����v�ћ"�@#R ��c@!x|��A)�㐃�4�y�İ<��@�r�`�h��=�M�"6��b�&�V��x����!�>�|�1C�8(�d��\�t@c�J|�t��ȓKи=�ALπL6���ࣈ�W��Y� ��]D�-���I*O���;N�e���	�ggb��ʕ�8���\�~�(���X=F�8{�>G���`�%�!"~l��Ql�;�0�oZ�Z춅:@�'��Hå#�a�^U S�F;H����z��@p�h��T����-E�!
�a�.^�0����2D�(���7�-�Xxa����=UJ"<��Z)eY �~ڷ䎩��r�S!�e���Z8��ȇ�)�I�T��	�eW�o��-[������I�A� !�qO?�ɄN��S�a�/�Ai���G6��H����>�r`тI�4k�����(fQ��	6�����p>vh�X��g�³C������ ��4�>�*<mږ�V�9L|�̟�Ė�M��I��Ɨp�ذ���C�Zv�~ң�=>6L�4l��~4k'��1vnfl���CF����W�6�za�n�֟��3�ɐ%�������K���8�e�$?qQ����"����X�'�AY�r�Q��OXY8���5{��L�h4>��CdU�ؑg��Dk�	K'�b��gc����_���,��+S�An��	=8~��Bbn��2p�e��q��O2EZd��?�P�@n�`�GO�RC���Mz���(&��|�fֳW�f�:�-�2d�>y�1b�q�f<y�d�SX�'�v8�4��Pp�ʠG�hX�	�
g�f�iG�'�ڐGMЩi�he8Ma1��bg	��F6�̓��`Q�}̓3QtA�6�ij�i�)rhd2We�;j� )́�p�^����d�'�&��P�2A�
��
n,A0�$v�d�N�#Dt&�c^V���BP��s��6J����&B��Q���'@�O��S/�-y��jw�ؐnfҍS1X���3�E�F�u1�f��Vrͫ�&?�`*�uC,�U���:�ܢ��L�BUUG�::ti�բ�*h`ː#$|O�����-r��/\��8q˸l�������Byb��1�21��jKܨ���%�*E���R��?[�m1"�P���?)�-�
\�ȡ̤u�X�K�kذ������<�@L[����T����n4�Ԥ�1dH�H�x�� V. V*p��H�W�h!�� ,��E�i��cm^Lp���{ �58���J��I#����7�ڠ���T�Fhg�i���ZTxZ�؅��8b-T�B(M����?a7��s�L�PB�=�\щ��RV����r&�����]�R���Q�L, �Eo؜/�0j� O��ԊC�@/4���vh�f�(��'�&�d�;���)�� E/�=�I>)�����e
� �� ��ƚ|?9䈯�2�oW�}&Y�%n2���)f�p(<�7+ � j���놺��܊� ߵl_8�" ���/w��W�՝x��\��]�|�q����!i��|�m=h܈���G�xsp0���p<a��ic�c��Ɇ+T:X$0b�Ă7'���%?a�̙5e�N]	4%�uYp��F�d�'��h�h�,�((�k��+�Y�O<���O_1OuST��2��=r2�DkC�ʫHS� �aH�6ufB䉢:��d �Lܾ3�G˄�o~㞌�aJ�W�S�!���"Zؖ��C/�� �C�ɼT��mZ���-%�v�J1�ܖ% B��* �L4��h�5���)H.bY�C�I%�U;�C�06�BЀ���`��C䉐BF�=5� pR q`"�B�ɭwn.�9��C�� �&��3:�C�Xrha&�P�@ָ�q�E��1�^C䉎7UF$٠��Nmܽ�TE:m"C�	�᪐�vO�G1�q���ڻ}�XC�I-,�D����P=x����F�c`.C�	"� dY���QxD%�E;�*C�	0H�,BTf�XN J ���C�	�
 ��`�,�L���N��22B�ɡt�c��� .J���-�&��B�&gtZ#cܾj�\ug._% ��B�	d��E� )�|-8v�����C䉓.�6a��ĒNS>�Ғ�]�`�C�ɥY|1��]�t��8�V�A;XNB�I&=24;��)S&�@��΀�D��B�#8 �cT�V�=���kp�@#D4\C��2@�r`�' �}Á�u��B�I&XS�41"��t̊&�"UTC�IdǒX��̖���r'�(C�- �Zt��Zx�I�(�o�0C�I�1`"̓�*1s���!0Y�Y�BC�	�e��xc��5{�б�C�0C�ɣq F�`rJ�\��A����X�B�ɬ�&t[vM�i�d�)�*r�JB�I	x|���0&X�[$�_>:B�1M�^T���;b<	�BG�DP*B�	l"z����{T�!Y����C�ɡ1�H�ÌV[��Q��K=-�C�ɐQ���1'��7�\����Rr�C�	�u��H'J5f�X�S�s��B�!������1޵	��]�w�C�Ɇd�L-���I�T��-��*.I�C䉷mFi{���Cа���G��r¤C�		�0죓G��;�����Ƅ8LzC�	'gj!���I�,�ՉֲN�VC�ɧL$U��f��;�d�BW��O��C��^�(�ٶ^q,�a���KT�C�/O�L��6�R�lD����N[�<��C�	�����dI؃p?J�)�
 ��B�>���;`�'P��Z�,��L�B�I��8�Ɂ������F�p=�B�	���B��ؐQ��-��$���2C�	'v�1	��Ej<��B�n� K�.C�	�mͨ ��<P��ũBJ ��B�ɥ^R.Y�+O�>���"�#�_^4C�I
.t�T�/U6�]j`�O�X��B�	w�v4獄�a�@�#a"-a��B�0:F�a�D�L
H�Tq84B�I��B�A�Q�Ū|q۵�6O��B�ɞ2�TX9e��J������fB�ɿn��Y���^����%왠9?�B��0'�E���86���X��Բ+�C䉐SK.���ѴY����Bo@*\zC�	#a���Y���펰#0i��F�pC�)� �㣌��|����ͩ

���"O*�V!UjG���r�?O�B�"d"OD��7��)C\��`蛃l�*살"O�X{%]�ȱ iT0R��p"O�H�"-�n&��Ӂ�'a��"�"O�� ��i9(}���N�y�Z"O:�����F�YCo͍4h�4�V"Om��n
��6���&9DiB�"OΠ��k��U�r8�@�9B/!(�"O�h�f��0�,��x9 *e"Oh�ʴ8	^T���� Q�&m�&"O�`cED�j�*�m�<���A�iH<!EG�G��0��1P>�����<ya�]E0�E33
C�I��,R��Hy�<�����C,�u�h|4H�(�jQZ�<��a��JNpk��c��Au΋V�<�V��W���7�_c� aѐ��S�<1*�{����zF]�� T�<���,]�B���K<czx!PO�Q�<�2�ؖ \2؀s��*���(NX�<�e�8}Y�~�pb��S�<�5˒�w����$��9Q�E
+H�<����� �Fɐ�d�d��`I'cC�<7cW�/�qڒ.UyZ���}�<9��PRC�"L�X+����!z�<YF�I�u�r�e�n�2 �� �s�<�1l�Z�i�k��f�T� F
�u�<A�%�,wꆀ���ތ�fՀ7fHt�<�d��9@	*$
�p�,��"H�K�<yp$A�1*�ys%���@F�<v�t�MT�W�oi&ؐ�/�\�<i%j_L�X,`���(_Gx��$��U�<ٰm\�j�F���ʈv4x���J�<c�&N���a�ɉb!��Q��H�<��΀3>�N8���RUR5T|�<qC-A7-8r�r``C̒5N�,��B��{bn�S��B�.=<�YBi�$~�B��9$j1(�%L�k�`�4y�B�	�	�D!j�e 
�4��"N�y�~B�I	k��Rу�+*!����P�2C䉗%h��pc�^	d t�̍�:QC�	\	Sd�����Nn��s�H0D�$�Q
�1~�K2 �.��ū�#-D�Љ���?@�����O,\���?D��Qt��x�L;�gT��`Ix��!D��ʓ��-�t�+A"��]���A��!D�`3,�<���ªE#G2�}I�?D���A�	��0���Aֈؕ�<D��KD���h�횈n9���5J D���Հ{U``׉��O�����L0D�,���F�Z�n�I���0>�$�*D��֧��ivep���0Y�P3�a'D� q�/��!RQ.W=O�l��&D�8���-L��1�R��x�#D�t�B��3[�HԱaE pOZ�;�%!D�PW��%�n��g,Ű.A��h4D���fR�!�de�����2D��K�G�m&؊��ͿS��%1D�P g���p��bֆV|���9D����Iìal�$��6�̥*T#7D��Gƚ�	��1V"I�Ρza�'D�p�+ǈ1 �R!�6+�b�h�h*D� 1!��W�R}:���+.b$be)D�dq	^�c֔X*���"0��Y�o%D�� ܸ�я^�̅�&,�n`,
"OB5゠�'H,��-{T�<�0"OX��6a��*���&/Ծz�f�Ȑ"O,��&9�YAH�3C��p*�"O�����d��pF�0X�{�"O�D���w��i�Kǿ[.z�!�"OR�a���V<h����.p�|���"O,R���Y��T�D�]2$�$@T"OD|��(x{(-��Z�R�L9���`�Рv���
�����3o+���B�.D��ǒoD֘r�ֿ=b^�AG�,D���#Y4RBB���!&RD�CN)D��"���hQ�PcQ��^��@e�&D�\⣊��x�@d*��\�
!,:q'#D��ؖl��D�����:��}��)!D�h0��[+q��u��$>��=��"D��!��6��i ���v��8��5D��86�׸H,H��e�
%�i�14D��i��
�7yqI#�I�zAZIt"2D�p��/o����q�F!/�pY0B(/D�Lx#᎛2�&�8u��&5f�µ� D��@�.�Lb��iwa��_�1��>D�\A�@�7Cv�Je�P(9�!�h?D����!���t9�� J�Ryö�8D�|j��R4L�tP��N�T�,j (4D��A���v�y��a@4q,II�D0D�조s$`�_0vQ�9D���g�/q��@��*qJDH�g+D�b���-Wfmr��ؾH^8p��'D��z�̓�Z�b-�dY�1$�i��"D�h��8v�D�VM܌>��5�s�"D���C[?$���ɛ,$f�0��L5D�l�)�F|��"i�-_����B1D��@	!WQ䀊���4^���[sn:D�̚�+2	&4p҇�=]}�UBa�=D�d��ø�=���E�<�9�,=D��n�\f���C69V ����(D�0��jį:�B�ې�J)��с&<D��0���iE@4ʊ$/�3am:D��jW�"c����'�|��	;�e�s�<���{!�x���6'`��S`�Z�<1��/��#�.ش*'&�����l�<�uIEO��t*�ă-
b���K�^�<)��@zZ=x����y�(`2��[�<�AQ%$H���-�QqHɶ'R�<�¦���4i�`"��|��@!j�d�<it�ӣ��q`1�������d�<)���u򔄸���f�h�
 G�b~��'0�u����q\��a!ʟ�D1ΐ�'�X�
��Cf<q���X�C0(��'2�ԹNP�M~��zq�Ŷ7���Hӓ��'��M� @?�[Y��G -S��'�} �gI��$�(�n$	6}[�'�<��&�#A�J���2�4r�'����c8\�R�0��=l����'tݫ&Ȃ�+E�\J�ϐ��,�	�'x�Eð�7{���F�΢==|8��'߈�:�m۶OTLr6�?�ht��'�:(c�O�j�P�cψ6`ġ��'��<C���9p'H��N�6(�X��'��Aӂ�&(p���X1Qܴ��'Dr� �C:\�L���"d�	J	�'��!R'!�@O��O'�D��'*����� ��q�hO�2����� 2zB�P*LX�KVu'ʽ�"O�DcMó�����P�"x��"O����[67���.֦~����"O�yq r���dg
�e	��)�'�`a�4aC'XVu)6O-}�x��'�x�ؒ�P8]4ţ�#{'�l��'v��RFϑc�R��q�I'kl|ٲ�']�pRp�[�&���!1`Pm@�'N� y1�����w(����X�<%n �"@R5 Ղ1K�yQ׏Q�<!���&HԃU�� Cir=�c�WL�<駅řN,� 5�S�^�H�EJ�<�U�Z$z��	��Yz�j2��Ї����@�9'�,�10��-ɮ$��vӖ�a�Î�@(yIg&W,L�.��;�p�@b��]��U�q/��f����g(lL�d�ӵmU�����yF���ȓV� �*BFP6@	b`���3(f�$����q7���2��zf��8ZQ<��{�>8Q���'���*@Jҵgi
5�ȓcA�JmI�	fVE"-R�	��Їȓ]�N�r�-Y��|��SM�.H¢Y�ȓN_����C�"�������2�5��X��R7l��(\K���A�Ȇ�}�(�� ҤK̠(`�D.Q=����^���g����KT�)&�	��wC@�гG��Q,*���L/z�\��w�r���1P;(Q�&dE��>�ȓ��æ��$-#4�Ә4�"e�ȓq��%�7�TZ�8�ޘ3G1��S~�B`�Uњ���E+@�p�ȓk;�YJtO?x� 0�B$GW`����o������,t%��b*�lF���ȓ"�Lr`J�f������GY*�ЇȓI(�c�<!|&����Y)}�BY�ȓF|�<sG�ڞU"�%�G�J+�n؇ȓ��)��HҜu�<u��b\15Z �ȓ&b����]3�9y�C�+,��ȓT%�j@t��$k f|t��>P����"�Xw�A�9Tцȓk X�FJH�O��a�vL��, �ȓRl�)������I��D�;
���+B&�S����/h���2�Ab~��*G�m�o6�D��N��̄ȓE�ḇ�Z�� �T��Y���v��U�ε<�F��Ɣ7⊍��;�<#�oZ�8��ħN�Zd���ȓT�*�;�O���D��	��(�4��m?2T�QbC�t���j�EA�F�i�ȓV�`� �C�`��Z��V�@��ȓi1� �KX+d2!�͆O��E�ȓ0����e��t���&SOm�M��)�PP0I��r����f,NZb݇�VW0 *�$
��F%����"9�l���O�*���)U�q�<UX�u�"O�y���1�\���+�\zP"O�Z�KV\�H��
:�t��"O.��,ؒ6 ЁW�f�f��"Or�[�#A~Z�8q�D�K���E"OZA�0�ڡy�>��c'+�2  "O�D�*�'_��Y�$'Pf�
�X�"O���C�H?7�
�S�K�p�R=ie"OH�IAHJ�'VXIE�C(f� s$"OZQ�r!ːI��������g��l$"O� �����7o��4fсZkB���"O�YS%^�e�����A�|�P {7"O��3��9�:�� +AL@I8$"O��K+	dh)�g%5MA���"O�3����J����n;��6"O0�S'�S2ND2|2%N�	2�d�"OZ�!�Qj(�PD�,t�h �"O�)���4�����aK!`[l=s "O"�	���jx��%\ FER@��"O���2��,m��X9�%�"h����"O|̃���*�vEJ��J	�"O�9����q�&f���L�!"O.�a��Z�����Tŕ-Y���#"O"I����I<I�V ����!"O���,ԂJ� @[ScN�i{Z%ȁ"O�-��B�o 4a���ԗu>�0�"O�����lM\���G�Ne�dW"O�����9'j�!�F9PXv�ʗ"O~�B�Nۜ-��Չ�=W��"O�\['�FȄ����P�kQ����"O(�0�D�q���te�(���yv"Oxm�Gϒu�T�eD�`�V9�R"O�t��U��%�^�,��r�g 	�y�M[�@��l�iă��@��y��Y7İ[R��7A� �	���y��1N�� 0��<'.�)��̳�yB��QR����c�.!V]�����y�g��h�z� �G��H��g>�y��$O��Yavb�9?0J�x2OQ��y��Ѓ0?Ȑ���*>G�qq�y��LZz�)k!ϔ52�B%����y�mW�����b�+�����		�y���c?���M6%��Ű���yBI�{��<�QǏ�?zy���y�UGz�����a'� 1�!�y­�8eq��q��Ѷ�W;�y�"[W�Y��jN�xjì*�y�Af����R�r�b���1�y�eXE�D1qN�Pb��K� ���y�#��9�Z<B�	�G�4���6�yҢF�_�eIу�R�h����y��	s�z��`�B
R�LH:��9�y���#ul4�ehK"[�!�'�E��yRBU�u��Q��X�_x���
��y�<�(��e�7\���[�EZ��yB��\ʱ�o+Wf���A�y"�ĖU��\��c�(Q��#&�^��y��2u+$��#"9�B�Ő��yr�)C�!��$���!��yBK[�'$Qr�hԖy�ε��ԧ�y�àG^)���U2y�P�xd�@��y�BS�b���*� ݛl��(�L�yb�C����$�5i�Rq��j��y�L.��Њ�f�eR�@� ��y�a�nN� "h@�?��D���yB�5�n-��E��.R ��V>�y"�S:sZ�������RU�<� �D�y�ZRbF%�IޮG��qQ �J��y���f�`�Ĉ��k�QB����y�
Ǥ7�m�t�G�:��g��:�y'�J����TJ��5h����y��ʶ2�X���jF��>�i����y��N�B��+�~,��٣OG$�y���H2Ptx'�Y5s��-���W��y
� 68b�G TBf�H1�bo�U�"O2��1�Ε\Z����Q��0�"O���l�,`�,��V�L�	V$��"Ofq;�"�&b��(鷅�8���Ѵ"OD��fIN5@�)�M!��<�"Oduz�<�����"ׅ��0	�"O@�@��G
���� �X�@�����"O���g��:�J�Jp@U6����"O�q�IV�p�:�Y�n��JN���q"OX��IA^W�`���R��I4"O4����ʃLK��S�!�r�iW"O�{�B�h��t�8�	��"O�cB�	�}�٢�c_%e��ำ"O�I��l��t�H�B]�$���"O����/P�R�0 s0B_����"O~�sH��x�8�jg�Wp`ȡ�"O�a*2΋%�����_k�ĉ�"O���a�E�jτ���Y��=��"O�}���
ixQxQ��W.���"O���a߻=ߒ�IsKB�I�|�r"OJX@��<�P����E��m"O���qI�:s'.�I[�D��"O�m��B��#U�Qȁ�. ���"O��H�%G�W[Ā�'D�c�dA�"OjE"ŞR39J$�ڡB����D"O�U@��֊0(HK5��	U
I8V"O^MH���$f�t���W�Vnh�x$"O�a��E�ȪР�@��Y3�"O�=J��A3_:ZA	`͐n��0��"O>py�M�9L�U��k����4"Ov�aB�O��R}��D1Z�+�"O��Дkި:�e@�����$m��"O,dc�NLS�|�c)Y;�@��D"OH��AGW�2�R�G��F�(�"O�A�'��&�@d'�6^���"O4���ؑo��`&[�R̈"Oȵ�U�O�@,:�c􄏆NF��i�"O��#��eM�����%�D�"!"O %�lNudB@˕�,J~���a"O�I�)̂e��8�bC,Y�0x"�"OP0�k�7-d�-)��I�l!��[���u�\E�l�Jtj
_!�D8\Jj��d�>:�&�3��W�Y@!�$Q�*:U�'��e�TD�򁀈,!�$���%D����a��Py���
A���N��	� B8�y�'ۨߒȂ��9V��Q�B�y�s�J튤eB0p�Љ�ς��y�k�A����Ǯ5,v*4Y�cF��y$@(k�t�E�G.:�=Z�O���yRh�	~�PZ2EV�0�*��I����=y�y�㋲-rT� �`V����y2��r���K� ��^)؄a�Y��y�&>�݃� 3^����$͞��y!:  I�3���AC���ToC��yr�ڦ$
6x@'B�569ڡRD���y�-�7pڨ4����+��Hk���y�ߴ"�p��_sz(Q����hO4��$A�`y�q0IC,����r%�#V�!��a����V�ɒj��ty�DA�*�'�ў�>�����mz~$����i�6���� <O��$6�I(m��*�e����RFV*�
B䉘n,�`+B8Kᰔ��-���C�	K&e�'�V��X)g�>l'�B�)� 0���z�手��� W@,����O����W�B�D�J@�]�B�x("e�3?!�dU> !�Cd���M֒%Z�B��&(!���Y�����(����¢A�`
�y�ɑsG�m�ŀV_~V�h�B$O�C�Ib�l�EKX�P�B�B����C䉷 ] ต�N�Y��$�_�yĬB�I���1D	N�FoJ����2�hB�ɺ
��A�g�h�6�2Tj\9bB�I�+h��h0�O��Ve�S��<
��B�-  �,놭�p�(	��,GC�I0?��Y�!d����L���V)L�B�	K��X҄O�v����N�1/�`C�� _0�q���(d�8��&U��`C�I�v�|\�Wk� {l� ��͹39BC�ɛ*�]� &A�-�, ��V��B�	~�����J�)`���a�h�/D��B��y�h��c�Ԭ �� bqd\�o~B��+Pǈ���"�:C�x�j�o�zB�ɟp��xa���R>	F�	�t;!�J�1|��h���&m�9��L3�!�d�K�R�K��Y�RX��0@E��!�$�/W�6i`wg[�|�P�7�U�D�!�
[䡺"n\><������	1�!�_./B�`��>�-@�(��5�!�d�/k`t�+�@Մ!c� �A��h���N��@�)F�H$�`(�K�+e:��+�g5D��ٵ�`��I +��C�X(�4D��0��\#{�>�ò,E�(���<�$�Ox���#B-�F�Q�����Ju�џ<D�䣅��DA��/wV%y�CЊ���;�Ovj�"�3j%j C!�Z�8��;%"O�X���G�>�A4�1^�N`�G"O���؅#�pY�F-��2���Ku"O�q��d�;��1�i��'d@\2T"Oج(nR"inޘ���ƟFPFP�p�|��'iў�ON��퓶n�4��¦G�i��`��ODQ�hڡV:� ��&.;��-J��Ik�OI
\�AD!�z,kB�.Ĝ�Y
�'����a FӀ��KW�^Ϭ��'M����L�3m�,[�.��D���
�'��ą�'�2�z�"U�Aq���	�'̖�)HI�!���W�3
Z�2�B�)�$k��Z���A|g�I��C���=)�y�X�PLRb�O�D�ɛ��hOt��Iׅ
dhp���B�8 Iq�̓,�!��Q5d�D11�~b��(AW �!򤏸A������>$=����\?/p!��AW�h�!���-A�rt05	�M�!��8q�l��fϘ'E��,�������	���?E�$I��c_v�P2?5Xts�C�<��O<#~r��̓B�։���L�j�x�R��~�<���]=���T�%��ȣ���v�<)A��U��1BZ0�� A�Xp�<iK����01�eN4@AX�ğh�<�$N��� a��ϔ�@{|�R���hh<I�o~xљF���u����'�ўX�'�~��Ө�3!�V
�R�L�(x���>�4����]=On���jЯp/�"OT�u�-
�"�R`��:p5r�"O���^!���;`n�?�����"O�k�ŵ{����$����hq"O&�ƥ� U��y��-, FН�7"O.�����0)�V�Зl�?)���J�"O� ��Y��5/�l�q��؍)$����"ON�����y�;�g�`n�*�"O��q!Ԡ`��@��
�0�̘�"O����g�s��q&ٻ ��0kG"O��:Щ���P���D����*D�X���^.n�x�!n��Gu��� L-<O�#<	�i�%]��(�&ɜ.,�k�N�L�<yb�	<5+!��*3�&iIDKOJ�<���
~m����
ӧ~���1#��F�<��-�/lP��O�"^QX\!�DJ�<��M�)�zt9��
s�ف��ZL�<W@|�$0������w�K�<�uF:�.�r�c\���4*�Fx�З'�>-���1���S��H���P�P���l=��X�hɭt��P�W�r�B�	2@��t
�h;��9���*��=�	çE�~p�&��% 2�h ��+3b�ȓwtX	��L�`�t�t� g��p��zk��r�F��O%he0���r���ʓE0�lj���x$� g��9���Dt��Ґa[[��`���8�((*I:D��E�a/�L��m�0_�$D��5D��X�- Q�J���:P20�*�f2D�dٕ�L&��BT2'_��IU�1D��A�̽&�)j�(�(����+.D���CN�)���!�0�Čpc`!D������ܨ��r�X�9G����� D�`�h�tE,| &`���tH�Q$<D��q&��3iﶭ���H�d���ҧ;D�����W$6�A�	#\�h�Bf;�$!�S�'x$����Hǆ0�i�FG���ȓY/x 蔣��h���`JI�.0�Ն�.Ap��l��9:�	t!FJntمȓ(- |B/V(R��!�� 3%@a��j�t�2���?{n%Rh`���Iq����l��M&<HTI�Dӱ��q�qC&D��&$ߙh��)03��4/B�}E�.�	e����3}���P�����3����B䉻J!����`W�f�`��a!OfVB��K���ҦH�.;��"ʕ	v�>B�T�fH"]v%� `�����B�I/#"} �&�����R�j�B�5H)��ǹ vaɴGQ��B�	1O/�iQ�ƃT��O[�~����0?����4�h���#HQА�%�R�<q�L�M�%�TK��RQ��/�x�<��l�~;t̙s�O�^�C�t�<y��̭fxH����u�=ʢ�E�<a�м2�6E�4{�UJb�Y�<I$eD;R��e��!>?���ύX�<�$�C�ڥ�a���W��!� .՟��IQ���QTkI�`�x����/NXT��-D�X
�PB�����R�1�D(�8D� ��L#oG� �f�U�6 ��5D��w]�̀�!��^6<{R�7D�d��Hꊱ�����75��s�0D���B��)F����B	Q6
���F-D�@�$F��^rU��<���D6D�졣.��D�Lm:Q��S\� �BH3D�8@2ŝe�tdJE�wd��!B/1D��!���1%H���(v�(-a�%5D��+5���8})r�G�Nˬ��5a5D�hpD��7n�2E녟u �D���1D�(�a=��8�OB�g�|x`,D�� ����\(+���#g���B��"O愸�.q�jy1��[S��d"O�=(aȌ$�Pl���B�[O�|q"OJD�"��2��b ���7���"OBAJt���[���IF�:��,�v"O��*U' &�R �I����d"O080AQ�c�͸I �J��5��"O( �SIɛko܉z�Dq�6=C�"O���/r?:Y����.�p���"O Q*dI�"}8g$L[�<��"OLh�'҅�,YՀ<H�Va#�"Oj�J��'|����B�n�4�"O��" Ȳm���+D�6��{�"O}��l�P:�Ap�� ���"O�I�M�%Ѯ �Qd�n��H�"O����7������~�t(�"Ol-1$L�z��#C�{�4�g"O�!¦V�B�\�[��őn�zL��"O��ɃK�������S�>e� "O�!����)b�;�g���\�"O����H͙����3gI+x���C�"O����ʕj� ����z��e��"OH��V�� �r�Qu�1�D0[�"OD���'ְ+�h|��bV n�T���"O(��)���J4raKF�դ)p"O�T��6I���3A�+u���Q�"O�`��eG:]�����d�,`"O���!Ѷ~yJ<�ꕼiH�-R�"O�����\���%+�6-b��t"O�;�@V�Y���VnV�{v�X0"OF0�ږ�&�:�Ĕ2I�d�"Op� ��(}�����g=��St"OvA���
x��ߚCL�C@"O6}е+��i=��Y�X<B1T h"O~��@	]3�b��d�)t�>�b�"Op s�j����R�З.q���"O��)#�
j����D�2�zp"O,�`�NB&:Й�CCp�|�6"O~}9ei�r���s&I�(
2��"O�p��$�¤�+��# ���T�'[�Ę�(o�5b#'G�#5Җ�x�ބ��'7���V�%j�r�ZT-�$lj`]��'��k��Ip5h��F*_|BM���D9�6��b�K%Be�a�Ns��	8Q"Od��L��d��#�����U�"OPP��=m:�����Jf�q�"O8�aQc9����w`P$BPu�&"Of�5��S8 Y�+O,!@�"O �c��3���`H �rp1S"O�\C��A�8��(�)��/ ��K��Ia>e�s����a�'F��g>��)��7D�س# 6a�J�y�g�0b�|=���?D�ę�j�m������R'_�����?D�����E.T�����d϶)2����1D��4�)0�H���B,;��y�pO+D�|�G���-�����J�0�i"�=D��j3��7��%�SG�K��Ƃ<��O�����G7tQi��hV`X��_�
^C�ɑ/���FL</ ��`��c�8C�	,D�,�`��Үj����―B=PB�	t��,+�J�2�j�2��H�*B�I/7t���ϝ>@�����[�CغB�I.?�V�)OV!
ܯ\
�C�I/[$81�Q��W�*9�p�#HB�)� ֭Z��@�q锘�V.�sL�ԙ�"O`�#��;��ajNۀH�^��"O��gi�(:��q��jF�^���P�"O��QvbE�l�D��=��Y�"O`!�e�5-d!C�?Z�D���"O�!�'��� EcR�A�@�tX��|��'[��ʣ��y��
�]�̀)�'0��d��L�F��ʘ,�¸8�'�pU#�X-@�tt�U-��m��'�R���FӪm6��:dg�*N}x�'(��rd^3��A��Bϓ{���"�'t$8�녾�N��򊏔x���3�'�F�0��|l�����_v]J>i�����&�������;|@����ڽ�!�z�̸b�	�6K"y26ŝ��!�$E�!0�j�j`��DN�x�!��H�mǂ����c�,��c�(~/!�DIl��9I@-�� ��ţ2h�2!�Բ������]ΤHyj�2���dB#`�`�Q�Y
�
��@���'�ў�>���A1�\�bJ�%B���&9D��Kd�A�t
,D���6)C>@��e5D�����r]p�0G���<�n�Y�C(D��H��!��;�B�=cX��b�9D�X#Ǩ 8f�1T(���2���4D��;�I�*aC,�&g�A�� �<D���U
в}��("0�\�)$�kp�:D�(��'�j�$)eb��Y �|�ao5D��U��+)� t�en�d�)5D�<�Q�<%Ȩ�"s!J���%D���Y,{p|�� �Q�h���a1D���c.�W��cu���F��|�Bl<D��խ�c��y"�{�b����:D�X��A.~�a n�z��%��"D��0Nˍ43�%y�NU���Pe�!D� ���F�-�2cT$����*D��k�!L�*3���ߏy�~�چC*D��aCb D�h��V'��T�A6�2D��Õ�����¡�"l	Rh�0D��ӵ�Y�f�0pG( �ܜ�e*,�On�ɂGh�h 4�(9�y�⠍"P�=�
�#������S�$�0���P<L8�Ն�\����&M��9���7d�8���_k�L��+Әau�y
��^0U6���/� ��S���;��l" �?��*�P��D�J3Q
̄����J��ȓoI"Iia�I�<Y� 1�	D���'	a~���9X�H�A��ߚ��լ��?ٌ�8�	м�A�(o��y��
n�|l�&�FE�<كD�8>�t��IU�b�4J�*�D�<�s��[7���`ᏜFt2/�|�<q�B޲X�BxrSi�Z��	�^�<y�ƙ���E1�]r������p�<a�Mǡ]&��R(�S���:UF�o�<�enH4�!	$D��ʌj���jy�W�D&�"|��غHR�	3!�AB���G���>y�O,tI�
mò�j���,\/�c�"OMPh/W���y��R�L/��A"O�H����֤@���W�>���"O���p�ʕ1��]�<Ĕ��"O�!�u�G9Bi+�oLc�>��A"O���3�B(�`T���HI��
V�|��)�B�Jѡ���Rp�	`$��B�$0|OD�Z��������0��8��}��S�?  ��6F��x�'_�~��"O�ю7(��pK�kb�
u"O��d�X�^�j �	D7X*13c"O��M"hX�	7*�r�ށ�b�Ix>J�-5���{C�!��3 E�O�=E���
�3c���t�Ԑ��2`̍�r�	i����i��"��\ x�����I�,5$.8��q �Zt �Q4��C'S��ȓ,ت��K/�h���Ȅ</:n����J���ˡ,�.|� @/S͚؄�n��m`�V�$�5�,d�fe��	d̓��ln���f5E+�!�x��	�<�?E��	�G� ���_s���Cτ�e��|"�'���4�\�cLb���#�[+����E7�y��E�d;VIz�˰q�4�t����yr�ZQӦ,S��S�s�6��㪌��yBjM9z(`	��� �v�B�Y����y�/�p*^�� �v��8�ugR�yR.Ƅ\c-D�w�����8�?����S��LyRs'�/��ܢ���ꘔ'��u�)ʧP��ӎ�,z%�0�%eG���ȓIt�����K�E]��q�E̞7����ȓ	���F� ��̇�5N�U(B"O�m��lX9{�؝HW
Pi�Ȗ"O�� ��0#4�m!%�&1=*ؚ�"O��p�Q,c�<�A��V'|86�
�"O��� �l�;�A�`y��!rW���'<�	o�3?��N�I�R4���95������۹�ybLU�1��T��.^�)���j#�y�O݋h���8#IE��D�3aF���yB [?*; `@ԨƸ(�9g���C�I�y����$��d�>(j���$>�C�I�T�%�Ԋ�+E���)�*V��C䉔v��XZ�l��P�y*ѫ��]�:�=�ÓCL�}��?`�СCh���!�ȓ]�hP �C��CBL��Ǌ��J��Q�
�+��0S�v�:w,��&��ȓ(���D*_9fB�!!�!M�4%���t~bʛ�ܔs�@�d�H��O��y�E���6QCkmxⅣ��y�Vg<���!e�����Fڏ�y�́�n�����9]��x+B�L"�y������ms�� P4�M���C��yr�Ħf(�"C��tꆴ� �X0�yb�>^=B-H4�D%Y�\���e��y�� ���V�W���u�Ķc݈4�.O �=E���"'�ju�Tb�=W�0�u�R�y�(\�VM���aH�&{~��3kͧ��'"���Ï��WK:xV�D���k-2D��)D�"�j0�䢃�x"	�`�2D��p�-��uH���5lA�_��y�
2D�d ,a��	�C
��Ie�(�G�.����`U�ʯ~_$�+V�Pg)��ӄ"Of� U��*&���bث��e(�"O�\Q�Q�b��jt+L(�6�P�|R�'��Oq��k��ұ8�5 �`j��t�r"O�4j�lE�y_\4#JH�aDt�p"O���U"´P!@�J0�V.H��	�"OJ�.��}�(�ᆀ	U��l�"O���'N i���DN�dՓd"O�]H0B�?KV%Aw`ݞ>�����"O��	�� �(�����aU.v��yc"O�Y���0QB�t���lؘKT"O[c��%�vP9e���-\T�("O� �<s�����t�U�F"?O~!��"O�a�t�U8@�z=AW�� <���"Ovu:�+˛85��x��	Ծ�13"Oݹ���jZnx�v�ӷ;�`���"OX)dƕF����D�[��)[�V�8��C�S�O���X!HM�[���X$�R�[�N8�
�'�x�JZ�5;0�!Tj�C�Z��
�'�RmRQ�[�L�r=���5����
�'#fd��Q�k���ɞ	*� ų�'SP�A�mM:kn�vꉽ.6�k�'tx��Q�-y� 5�hIP�}�<��BÌ����M�'T�A4��u�<��nE�$ne��CN��01�p�<I6�B+
N2�;�H_<T` ]�W�Xc�<�ĭ]�����"�[�_1��@Co`�<�1FR\�T��Q5\�ݡ��_�<Y�h�:lX��	hy�1s�%�`�<�6ɐ52G�%b��V���)�`[R�<IQ���J������^�^d�<9cB�{I�tc��D*4�Լ
��-T�����
��~�!�G��|d
,�p?D�\r���?�T��H���ٚE	=D�h��$H�E�h}� ��
ms.���D9D���	��F|Q���L>^D�b�6D��1�>S���Rf#�7	��E)D�\I��=P��������s+#D���e$�,4.>H����9^dص8��"D��Z��5HŠeI%��a� � D�8�7�ۓX
�r��ۓnXa��=D��8 M���}��ܐ{����u�:D�$�`L7)O�yC��\��^���-7D�c�/�w㘬c�f�Z���<ړ�0<	
��lɉŕ�fB�| 7�m�<y�c�LDD��P�-BV���!u�<1�U�R��E�ԓ8��d�CH�{�<Q$�?�u�c!�gA61��]�<9�� |��8�ŧA&�j(#�MJW�<�a�ܡB�4��ƙ��l�&_W�<�C�z�Zq��[�E ZUp�m�QyRY�8%��g�ę7GE+Ѧ�3�� �"#ըVF!�&V�@e	�e`���q�B��m'!򄅏i�~�3�	�]���֧܅f	!�ĮA����00O>t�&�ˏ	!��׼v����������:��չR�!��A�w�(��;d�p��ɒj&!��Ɓ�H8�Pn����,	@�O�Q!�\�p'��g�d �Ѳ���N��I{�IC
\��	i<�䦇6Q��Z P,�ְ�'%FZ�<�2̛2;���N_�RvȔ�t�T�<�bt@DM�P��G|�����j�<Y ���L��ȫu���d�d�2��Rj�<1s�� ��`th�=��ҧ.�[�<��Pcz����I6)~��i%�Mrh<1����YRL-dA.@(����?�	�'�~�v捒]����e�W��\4��'Uԡ8E��6~ID����Z�Di�'�$c@B�4!̔#�)Ӝx�l��'H�y���Nu^�Y�	l	�%y�'z>!���>PC@
�J	<f=�����<�*�����{(��k⨍�KR<lS��'1!��ͻc�fp��ְ�h��5#B�nJO��c�/�Zaj1��)��<��5�V"O8��Be\�)���
 �߄j ����"O�� ��K'c�����/9�x�"O� �aQ�HܥyN���FT�L�h�"OT�+7KN�"LP� M
�V���"O�����F�L�!����d���"O�b�(��)�\��[F��x�<��&͘Z=b	�g��GL����Z�<�U�(Gք�p �6
�p�IQ�<f��/(�\��i��P�!��X�<QcJ[7	��pٖωTRy�`�T�<!���%��:3aW�IGHd�V�Kv�<q��å(�:M��ЇC�L@����w�<��@�F��@pB�J�m�W�W�<	gd�-"�6e��7[J�aଞT�<� 뚭�<%	�!�6/`P٦��g�<I"T�t@��c҆N �%�p��d�<A� ܗUb �S@���J�`����U�<Ad�@(����6,�4�t\H�EP�<Dc@."�"�.T�0*�AxHUO�<���[5%���v1�#�kH�<	ѥ��^�,��e&�X@H�@�<kXT�IHO�<g��e	�\�<q�H�>b���r4�G 2W�)�dM�D�<��|Sµ1B��%`���� �LC�<�3��K�Q�#J8E�f��A�<)���4?1(�1���5Ն��'��t�<A��Z:D�y�@+2 />�1j�s�<!��M�)B��:��ޱ240��p�<Qk�=+�,�nʰ9��YpN�b�<�Sf&#��(�ߩް�����]�<�$�V�"߄�1�n�m(hq·�^�<q#��#:b-is*�8��jLc�<���W+�Z��Й�|���WG�<�N6C����b�;s�ji��@�<y�Fʅv+��zH>+�9h��@�<q��>M��*]�M�J�CGk�z�<!t���,�<p00N�SZ���҇Yt�<ّ�]��� 3���U�yKQ�Lq�<!�@�*Պ�G�8���E
�F�<��L�< ZI�9J�7!�w�<�@D/Q�P����M����ˆ|�<�w�-,��9ju��3���VK�x�<�@��"�*�9��#i>�]��N�r�<i!N�'I��i8�� �,;&���_S�<�fNK������OJ���w�ON�<e,J	&�pM�#��$a�)����P�<gDT%:�k��*Z����'�A�<��	�'�.m��#�$���`bJz�<QPcKִ��R.�d��ؒwR�<Ic@�k��x�̜�ePv��K�W�<��H�#:���&�X��Ej&�[V�<!n����3�#����N�P�<�c`ŋ3�8�@�R&6�P��#�F�<�TiL�(e�)��ʜ$Y�x���mTi�<�ӭ��YF�N��1`�Yy#b�<� ��*��Y9&���L�A�c�[�<��+�$$�n�z�MQ�;�Z�Hei�_�<AE�F�lL�dY�Jw X#L�t��y(Le@3�
>�-�7-pZ����J�6����񮁒�d�x���ȓ
g81ir��0Or��B(s1�Ԅȓ9lD�s�G�
{�	�B����0�Dx�#P��F�an��zH�ȓ }�	���+eq&�2gJ�k(���ȓ(*�h)C	·L��*��VT���F�Τ��i�:E�}b��ѬrΤ4��S�? �,����Ae�p�f�d��4"ORD�ǩܗV(Z�%$m�E "O�,1�(W,k*�XqaDI�`@a�"OpL "�32��u3�E4;�3'"O@$a�����	�1�HJ�2}C�"O6)pD��ʁ��/U�y���K&"O�Q�1W~���2��.�����"OL��@k%8dTS���e
�Uä"OĴ��� ��		A6{�"��'4@q����0�(y��H�u�#�'�s��0�Ay�Ŋ3?�&p"�'ע�i C]$bI*`)P	V�:.D�	�'�J�䫈�k\�P �A>8BnM3�'����
���y�D�#.(�H�'*4I�-[�h>0zgᙑ�����'����W`�{�=ӶH�\����'S� ���B}�|[�
�XtJ��
�'2z�GoQVY��Q� �5Q�^�b�'\�Q#�n:Cq����&H�5!8��'`�xѦlP#ڹ�@ӧ'n�%�'�>��M��If�qk1(O%w�h�'3F���F�D��k�CJ,���
�'�bm�� A�X̊EQq�В{c�P�'��5ã?I�D���
woZQB�'�{�l-� �V�Cި�	�'�`5)u゠ ����u�P�jZ���	�'��<��	�"h�1z
�f�6�K�'����.l9�p�vƖ�^،�[�'ŤQ���G�.t9�.+z�D��'���P�j��m(�[:!�N�q�'RZ�i�56@�uA3�[�/���
�'�����#G��\A��K�����
�'����B	@�Ln\�� �(�
�'b���6 e�}��IS�g��	�'>�����,���*�OL�1)�'�����G�̀��,��F]��	�'�2�3S�G�����W�'���A�'��yS4l*UNt(�i/��LX
�'q y�0oT�3�
9��R��0S�4D�`��/׏MmJMs�FL�Y;�rd&6D����BQz�0��uI^5N�%�"n8D��i�f� �6x�0)^?i�����4D�|�E��%��v�A��,�#�!�D��j�<��$�f����F%!�ď X�(u����
@�d ֩e$!��-H�[4b&n�F��.˾�!�$�[-P��Gɗ$���C�
�!�DV�U�@�$��Hi�+c�!�䝇�8�#eg�a�*Lے�r�!�D�c�Ha��R�8Ts���!�$|
U��n�\Κd��iܪJ�!�,�p"S/�]�`\��S�v3!�䗡k��ܸ�&72WM:%�ɫ�!�C(T���`K
_��!wj%�!�ě�z�8Q�䈑12�^Q�"#ՠ�!�$9���'�]mLųS���0�!�Ċ=�DH����5b9��� �L�!�$�U��bP|��DP1灠X�!��� [�|��Ʉb���s�
:~!򤈖?�̔�ql��
�X�i��#{!��1{r0���J�!�#�+7r!�!&�
	`b��{�<(!l�M7!�X~st4�$l�2B�d麡`E {!!�d/�`l��K?=����3��&`�!�� ����T%�u���h}��#"O�l�r���S&m;Q���5	�T��"O��8�c��-(:���"v ���"O6���0>H���*�\eb "O��)db���ppO�7;�"O&Q�wkHU���I�e��P"OИ��mȅT�
�q�� ��q�"O$\U�(ft88w`JI���CT"O��$c��|M:���.�&�j̀�"Od��dS�K���k&��:z<Y�"O.K�4A&ƀ����A��-6"Otm�QeȦlT\�d�}��i��"Ol|��KO�}"�* ��0*����"O�͒�
�
��+��ƙl��R�"O�Ր�G��r���B2�ːD�Iڶ"Oڝy H�����a����"O A�C�	X����ݨ;���"OƔ���m%�99S��@� e�r"OL�R�'ߖ7����C�21�*`�&"OD,3�χ)�����4+��a"O�~4HU��_!+� x�l��!��qJ|@�^�w��p�C��	�!�����Bt����ǎ��!:�"O~|���Ӵ��� �o�$K�>i��"O�E�V� =�ʭ;T�ٖM�$���"O�݈'Bʉ�٨�/ӫv L��'"O��X�└|�q�ș�����"O�i���?�V�#�f	<��� �"O�ذ�8fa֕�2嘨�|a0�"OX%���"+�4���^�l`�{�"Ov ��Ӛ�X-��Gʎ���`3"O<`���V�x-�AM���d8�R"O  4��g@� ���*��Ec "OzH�&���B<�H)"��"K��H��"O2d`C���v��1h�Q�o�Ҵj"O�a���+S�f=�2#�D@���"OR�#$:t^Tq;3"&@�Q"O>���B�G�F�ɐ�ǘce���"O��5�E�u�$\��xG�A e"O $�N&��RT��@��K�"O�9p�c�7|n�p �ȠW���"O&-:$a
�@/�:�h4�V�:"OL	�']a���8䈎-��
7"Of5
PnҴ)W�8	@gץp�� ��"O���P�-����EA�ph)��"O,Qe�a@1��R�fN1��"O���F��%
^�h���|�4��"O�3���.v��q9��Wm�pp�"OhL�d��������%�b	�"Ot ȃ�Yx@��7��4����"Ou�`�E.aKdaH��$@|5(�"O<@Q��]�!�"hB�|>��"OV���wX�q`��p:F��"O����m�8
whe���qDzт6"O9��f�~6�k3��h6N��Q"O`q�**u�H���֎]GM�!"O���b���|l��'ƍn���"O0���
�=6�����;ĞDA#"O֩p�	�>��:���-��I�0"O�I;5���y=da�K�7G��(��"Ol��7?H�<����"l��ٵ"O�h���&!C�,��T����D"OL$�%P�d4X���fr\|`p"O�`FF�+d�t�p%!V
��r"O� f�����bI��7c�88�%*"O<d � �  w*�@u,���c�"Or����!2l�P�J+P��i�"On��6.�4��}�fJؗ
�Ȍq�"O�����X�v%�D!�^�c�hp�Q"O���W�k���t���=b谅"O>�Y� m��aʃ�(��"O�$�� �+,�(DhCN)��hQC"O��K$��*2(]r%mۮn�y��"OIf*ǒ-���re����xQ"O�h"�b����a˔�*�d䨱"O�	�ue�l\D��g�MZQ"On���$mv`���ԝ ��]1�"O�}@��84�
��N�N��"O�d�ЯT���(b��%���P�"O��x$
�}�,Ӈ��>V�X���"O:����T-⴨�����;t"O�y0-A&� (�s��0R�K�"O� 3��U����wf��PSw"OX����>Q�s%�,*��PZ�"O>TAR�6�v�Z3�F�
�����"O��Q�C�kѸ�D�<r��U�D"O𹣗��������P���"O�آ�͊�,�<�kK?Iy��Qw"O=J%��b�����Rsd�8u"O�	�"ď�Ԋ]��
S�]4�*"O܀3��D���B5I*����"O��e�x�>��#BC,��p��"OZY��#��D��ٓGU�j0I�"Oȕ ��,�ȲUGS� �ju�"OrB &��#�P���I�t�B�)�"O<��ڟ$UԱ#�+Z�l�*�H�"O��6�p��I����	��i�"O�DH��ػ/�$2��n���;3"O���P�j��0c"�3�P4��"O�9 R����,@D��!^��z"O����o� x�H�K �9H@�"Ov�i��6n  r3`Z !X|�$"O�P5j�y���hVMՅB�n���"Oܨ��-�!�`9X�Ů���"!"O��@Ⴡ5 �@�V �{����"O���F��y9��[�n�"�n�(�"O��B38wN���m�G�0��"O�l�̎�Ƕ]�4�:<!ӳ"O �h���]���:v�4'��T"O�<�J��E-h=K5W�,)�"O�1Ҡl�r|�q㥫ȉ#��|ca"Oj<yђ}��!k�yՐ"OX�
��ȗWk:��&���~T,���"O�t�P�I�P�R�ݨm�va�"O�KQDЗ���y�"��v�,���"O����%?9(B4�V"�c�"OT���
��h����1"��Y��"O�胗�E�m/����	�;��i�"O^�r�J:A ���h�>!�pbB"OpU�t�N�:�d�"�I��|Ļ�"O���3�߆1h<��'� 8�2,�"O*Z��"!�D쏗|t����"O�����f>]��jȬ{�QP"O � /�zQz�"#�ĩ"�@-�"O~�zS!�.8�w�X MCr8W"O���G;Z뒘`ׇ�P0P=��"OT�J�I�+��}�b��1~ȁyP"O�s���&9�����)��t���"O� ���� �¤e�鍺i�d�*�"O���֜U��\��F�V�����"O�5�t��j���y���`� "O*9���O�|�j� �|q�C"OT�y󭍄[�R�iB��^
L9 "O�p��d��,e4Ei:/b���"O\����!��9��.{U�Ъ�"O^5����YL~�� A�QS*hy�"O�#4Ϙ1bzJ�� ���X8�q�"O�a2��#��eI��ס0+.���"O�h�g'��
i����Y�p�<,#q"O�Y��b����;�@��m�ze"O���)S��G��)$S�P�E"O��
d ),^��bOզ6��!"OܴY���$d��3$�J���"O��Cڈ�l�ע�C�Ic�"O�!�l�(Ϫ�id���Y���Z�"OHd�Ҁ�A
��;!�]@���"OJ�D�ƨg�s�Jۍo�6<;�"O�\#����s:Zl�
ϾU�`�3�"O2b�&�.��$��'�LyI�"O��;�G�:R�{��J�s�l��"O��(Ǐ	y��QsT$�� ;@��"OL��i�h�^Q��[�|!��"O"��'�0+������P$��P��"O��kcǓ4��#Ĥ�u{��[�"OX	��@�8'�\�!��S��$"O@�j�(}�(؉`��Zc�Lô"ODxˢ�6$������H".���"O�F��X��O΅�4Q��"O�x"r�A0��R	�>���h�"O�mz�	�:��Ԡ#ذ ��EA��0��a���H��U5I���ɬS�8La��9D�T"&ɛ�gڒ}iC�Bl%i��x���sӌ�qD�\�|K�5�t��3��	2�'R�O:��W�]#WHp�c�N!��ɩ"O���g����#�O�k�20��D �Şm"�����vd0���ëIǨ@��"���w��Y& �`,�p�H��'���q���S�`a(X�DJۊۨ)Q �R,�DC�ɔR��T��ϥb�`���\�QghɅȓ1��#�`�'<Y�H��@^& )�ȓ;X��IRB͹^�8�T�!RŇ�Q�H�aDg�"��]"�V%H��%�dD{����k��fh$?7���"�ٟ�y�h��`��C�$�/Ak�L�q�ۣ��	A?i�{���.	[�0�f٤Xhb��ŤN��B��|��i֜2�1xTG2c\�ɊbP�ad!�D�6@�d�ǯ��Z��u��#U�O��=%>! �
>hhT7�T0a�"�pu%D�,8�-��$�8]�2��%���8U�$���>I�y��TEN*���`���BDr��W����y�V�Q��, ��=���9S�I���'azb�F�j�e��34،ͻ�b���O����FڧJМAb���!��PЍ�<����DP�-�8@�D�]�q����	z��	A "��E���%̬)� K�Ji�C�`�:���j�Kfr�K�o�+���O�=�}� �kv��C�&x>l×�DU�<ɳ�k��]a�j��Ք��$�N�<���̐k�\diS*��#�6��Cb_G�<���	;�8<�B^��±�����<��e��@���j�B��ZA�Xb�L�<94�]H< ���#V����C�`�<� �����D�[��:D-��!����F�'9�*�5�+�6�2ݓ4�[���B�	�a]�y��ʴb�ĕ�'YwC�I�Z���!AA��ʕ`C��B�Ɍ���!�h��?PN�:%,T�WB���LU��ޜs�6�v�\� (�C��w��Jd%[�2��P�1�C�I20h�uc�ϛ�hy*�'����C�	6�����.M�$Zhp�֎��GT�C�I9m�(�9v"U�{�^@q�C�T��C�ɂO�Es�8���#EJ���C�I>qs� ��I$A�5�t`�?Mo�B�	?7��p'��p� i!��[��#=YǓm�d5�$��&t�*9��SII���ȓP����a�9���R/%f `�?�	��&�%��3�� ��W�i�,	�Ɠ^�x��	_�n���c��HS��ⵈ���'9�g�'`p���FgN���6��:?�>Q��ט'��K��M������Q=���O����N#�JUA���w����2�Џ(�!�CL�V5��4*�t����!���b���np�pϐ�c��	]��|!�eH'��Ι>K�؍YG�5���	�30<��N~a4�S�&ܵ(B#=��O`\uJs�á>_j)���P�+&���Rl`W!͙$�p9�+ fp�lZ_(<a2 ��b�j8(�G
�4왕�UQ����?����>[V��c�ʂ��%Z��FL�'��y�/ή�T�xT ; ��`Ȍ��y��':>�"F�6�<�W�Y�n������,d�D�@����(U�޿n�z�͓�0=�L<Ʉ�W>�F5�tǀlJ��3��Y��hd�x�͜4C�}S�jS(b���ʴ�ݛ�?9�'ұO?z�F�ʆ����\�y��iR�
H�'��':����H�
-���+C`X1:��@C����lZ^�tb��bMtd"s�a�̕) ���P��I�*F]%$�K�J��p��0<�L<g�±`|x\r7�Ȉx�6��$ZX~��'��ѡ�ꀔ]��P,C�Ry�x�
�~y$�Z��tPň�q�"�y@bD(rA����|<X��Vp`j5Q�&�#1��d��ɈZT�'��
q)(Nĩ����ĵ��Eè��IR����{���7A��w")��s)W��(O��=�Op�M��n^�:;���{
�'�����%M�Y�'��C��M�	�'�����nI,��/ �@Bl���'��zv�Εfʌ	p۸6�09���1�S��Þ0&,�UH�&m���,�)�yb�$oFT��δ��j�D6Ƣ=E���o�X���y'���ÆY,�^���H��$BƐC��Ӡ�N(eFP����hqaR �f(�h׌c?VQa�fX�p>�O<A��I5u��X���(�t)�C�<���(�~t�CAK���d�J�'H"=�OR�x��O
$4�-S��4f�H���V<"�P���tΌi# ?(��͆ȓl �)�Sn3lh(�I�kۺ���>	ߴ�hO�22�A�s�/|DR�Z'�^�L��C�	/0��)�]	�>)0a�J ���IC����V�K6,׃&S9#�HC5 7�]a "Oi��`�t	�W�)@�LŚ�"O�P�tUN	�e/ܚ,�TL{A�'��'}��R1�����V�l
H-�I��y�DE�֜���+a�@�x2��y
� �:��Βq��m�q��K��"O�<���ٲ:P> ����NH�S"ObY�N��)�j[���mږ"O�;�"��vLX����n�^��"O���kԱR�m�P.	�|��%�"OR����O��51��-!�9��"O&D��C�"�����b��*?ąr��Io�O�$L�/�	JWVx�K��t����'`�Q���S�ԐP���-iNd(e^��'"���3}2m�8@c\Đ&�7g�����#��y��W,(����`�
�d�����II��(O���Ą� pA�EYx������!�ArV<|�$�F
i�L�0h���^���/�2��K�'.z�ɲ`�b�4��ȓp����@�"�$h!t,[>4�݄ȓw�\�S�O����m_�ȉ�>��>�>Q�g�&б�`��8��ȓR��T�֦¿m�~l���
&���=9����D�+s���z�O���C�	��p=Y�}�	$<C��p��C*V��AU�?�	�'S��@DbS.~�6���.��l_�H2O��"�]i�S�'2�
-��(�
@�<qp牊e���ȓ7~��٣O��Z@� o��j��>A�ÁV}R�I�:����1_�ĳ'N?H�C�I�qb�h�0,Ѿ!bܥR�M]��"�'�\-�@A���y��.�� �V���'�2%䊃.pSa�� 1�'3�Y�An�>"�}KE*��tݢ
�'UL����-B�t&�"	F��K�'!��+���3L��$���-Ԩ��'H��B!���f�ش�� �<u��'�R(�$�.�Hx�ė�{N`��'[�D����v\0��lŬt�dP��'�v0�Ac�uZ�;�NT�j��0��'�`h�pbvL��*��6E.��'-(���'��un�
�lU�('
L��'�<aْL����|*A�ZL�n��
�'N6Ԙ�F�5�9
P�a��@
�'<ؔX��0?��q���4=�$T�	�'΄š�L�X!��{�M��Dt���'�ayS�ǨG�JA��DD L@�'�Ĭaq���G׬��w��#L���R
�'	h����]����ǰ�Z�	�'m�h�Ŝ�h8��c��6�`��'�Br���:���aV��$b�,� �',`�au釞
n�Zv��e����'�%W�D�H��q+��γFCD%��'^����ъ2 >�8�*p���k�'�����ş�j�L!�'P�r,��'z�#��H�MB��B�&�����'t��(�gJgL\8���-BZ��'?x,a���J|�EhGi�x����
�' ��9��B��0�V��#�y��'��h2i�-�2��gkI��`��',`����3#����(�). ��'��{sAӦM�~�j7�W6}�����',���2�!�.�1}�*��'�4$��Ռ(|��ɬ]�p y�'�d2a��	OD���U<Y���x	�'Ǯ����+ Ø��@N�S�R�p
�'��]�P-�2�>i��C���ǘ/�yRHu8<����� ��DQBi���y"'Hb�B���c�0@ "�.�y�o��$��N>d��0kG-��'��=H����q�(h��S�)�z�;�y
� P�T!�R�*y�FAN�+�H<�*O��i"#@�B����C;b��t��'-�*�#̇K+��`AK�"���'�4�@��F�d��0h@�ӑ�R�B�'P�I1��#e�䣒#��|�����'�ֽ9׫Et���²�\j�T��'li���ϗS(��c�ą�Yf
�+�'<�tB�D�-U��|�H�j� ܩ
�'����Y;!{�%�Cd��e �'D�IR�Q�$�S�ͽ6<��	�'}�mp�������#Ԥ"|���'Bb�s�,�7IA���e
�#�8 �'�8��֡Z�]�C���'�^
�'����¢�c:F�3��F;�)�'���&�7i������4< }�
�'�v��V��%�h��A�YC
�'�z�@�o�,;S  bT��*a�4<*	�'ĶY�6� !� 0P���-����'yJaX�R���Wh�)$ܰ�K�'J8daǌ^�H�X�X �U��6�c
�'��¶N�P�B�0���
���a
�'O��r��V%id:a���x�%D��I��)�\�x`�;V��U�4D��S'��L¼#��M�҉a�b4D���mU�a��h���0�dp�c�>D� s��U!�6T��� !��CR�<D�x$Ǚ%@B�s��&WÄ��r.D��e�;<�j�k�W���1l/D��Q���"�0s���o�����+D��;�M�m���8[<*xY"+D��k����ms\�!@����(g&D��c	4�ze��K�SǨ�I��%D�x2�oٵm8��c2b�#`?���P� D��h�����-�gGװ����:D�h��F>(�)(e� J��qb�n,D�0��"V/2�V�C`�"�Љ��"&D���֪'��U07�ɫ eTMM�<Iâ{N�(�E^&CKD@���H�<�R���^8 ���� �qmUQ�<y�1P�&�
E��5'5.Ȋb��N�<��g~f�pZ��U7N���R��b�<A ����n�'aW��&$�b�F��L�5l�˰\�'�r{R�[�\5��9�/��`5�	��'!D�0�E�(&غ]��@-7h��ʎy� �5m���V�L�O���(�Ǜ!\L��ܬ8YxS�"OpD� mH5	,�X'&Q��2�bFՊ@��Q���J�|�g����>�0�t�ϴEf����Bס�$.��ER j�=#!�P�ïؼ=Ub���i�& ���Rb-�O.�8��C�~|��.I��I��'�t`�Ae�-O��a�:ON�"c��U��	�1. xb"OZ��
�6��%��MPb 4�0�|��g*�j��Ę=�?Q;#@
�x��4���R�k,D��9�#��ML}�d]�(�@�53:Ё���<!� ����m�&�J�b���RB�G<8�B�I����k$�H�9{X�@e�؝3'ب����C�����N���&��(}�xb��#D�h�l)<O�pJ��E� C�@�Li��Q�i�D�~���f�L���ac@%D�ܐ��'Y���${����&�Iz ���GD�h�Q?�vΈ�K��ʓ�߄{�t9�VE#D�D��fC�0�qs���)� �z�H�{o2��H>q� �gyBW	8^n|�Ef�o�V�z D6�y"��	�T<`l��T��$CH2�yR�I�aB� �Ԏ�
c����˱�yB���|���R��t�X��y
� �a��/e�4A��)t�BX�U"O^jB����<�:�l^4=7f��"O��9t��QnЙr�<8U�2"Or�{b$.ELt��798���"OX-).	&^y���ΫU�c`"OLa �m�`[*I��':�$]�"OV��i¾p�t�Q�*r�nYb�"OB�e
�f�| t����J�"O�%t�?��T#��X�J�S&"O�t��c�A��%h��ƛP!���e"O@�AD�bTt䳧B܀�u"O^�S��W�b-dDsBQ?�\�9��>��f����S@)�82���aM��ˆBΞ)��"O*����3|��b��ưg�V�8��Nnb˓���rc\K�g�$�|E8G�QH�B2��gѴ=���#%�pY���P3�`�e���T����ǫ�m��19E�N\�a}���C����Ɗ�>nq6��dܭ��O
�fǚ)_����В����'l�zh�����,9�Хl5!�dP�~H�Lޏ.�V�C�4C�	�{8�;�N���!��S)�6aQeԟDXA#��.|C�I�.����!�!��eI��/`.��@"ͮ�~(,N^MQ����{2aؠq�=y5�O��0 Sc����?�g�X�w.غ��6Aa�`dfG*Zs��ˆ`��A+D��Gdr���{��i�>C��J���G���᧪����$ήV�c���+Ԃv�q����������1A��
?.�ܣd��&�س$�P���c>c���?R%�%�1�M+!���a��<�� ��6���Sk�l��	6<h�Aԟ��w����'n��Y'T��4p��`5lX@y�ד[n�0m{�N�)�5E�d�vJAd� #A�!-���Rv�(*����T��k��(9X�H�8��Ԡ{d�C���⌠���d�A�0�{RA�"l�ix��۸p�:]ðH�B!��ᙅr۶�4	�lp�'��R�d6§1H���SҲ]���!0@/J�����;�6���Oa��ѲČL���I"���Po�AA�MB({P~���'�` �I�F�0��ǥ�{F{�Y"�� ;��0[�H��m�>�ēf����V�[^�����]C`�����_��f��6p�ey��Y�>����fkKi
��B#�'�j}��'66}�'�ę���6�݄�XTa##3}��D�;����'L��x���X�F�o�0]���/~;F���G�YŀEpH��>�p��D��}1^H��ӨM~h�1B/҆R0�r�m��(��D�ם&�,qeCA��M�o�&S����D\� `��pbl� Q��h�c(Z�џ�QÃ�2~PR���$ə hp�����&]:u�s+�J�2��$�j=b�&?��	�$�	�{s\�)@-^|�
fύK\��P�P�1��?2*ӧ�ԊX9<:Y�c�o�:1�AaI4�����1��U��&/�xb�n!�q��A�8&ʄ95B��'�$����uk�`Y��D������!�l��$�ΞK���BKur��W�#�b�C�	8
���2�ڇz�LI�!��w�\�� 
�8��'�Z����i�Zh!g���x�&a�=CO�rÓ+\؈�@���h��8�&��gq4� M�"�ʼ�ȓX ;d�x��m�Ө�p#$��On˖�љ����O�Z�HTh٭C(6�5��/R(��'~ 5p �N�LI*�p�/đR���	�'u��� �%�p�!A���#�
1	�'�^`Se�˵a9�m�'�ۊ,7�@��S�,�d�V�B��q��=�V��ȓP�С{�aF� Ī�Տ�2H%�(�ȓ欪�.TQ�	kC�D�)O��Dy�$��	�F��H�6���sS�c�2�O��yr��O\BlƧ��D|1T�P�[�4Xє�ė`}ɧ���DY�P�M���&_n��[��(-�!�d�?lD~��6l��rTƎ"�R�W8h�ؽ� ʐk؞�!a�Ć@o\Q�"аu�ٱ��5lO�	:v��0>\,��c�i��Pj��K_�УtC�gZܫ)O,y�S�����=�GL�K�H2A͒�:R@ؒ�/Sܓ)"fQ�7?d��I�O�Њ�Oۓy�Е�䄌:(�b���V^�i�r�L�<	GB�y�`Ly�i�,l�;�*�t.��I��d�Wr���=K3���,�XUЙw ,�97�H�"�0��R&�h������� .QQ"�Ʋ���S�$�5���$�R�%pt�@OY;"JnPS�J�.YyR�Ǳ��������^�qC�(@�P��f��D��Z<�
��� `6mŎN}�{6�G:d�~9:¡̋l���Ot���p��^.DB0�a��'݀󒯙�o2�x��X/��-��{bW�[��v�ؖ}���#>�vu��o ��?�e/��" ����s/P�Kb�ͽ\�����F �	��ɯ@���F��>!��+$AS�����'�;"�:�?AAII.B����'R���/~f��p7��W����ߑp��C� -��h����x����7bV��h��p�p���H͜C#8jƕ�-��P�iz����cy�]�]Z<)�M@	W>4�BM5Ȱ=!ac�$�X��i��<�HE�Ht�[��Ĭi�*u蔴~�L��'$��S#^�Ҧ�ɭP�L�?����!I�رP(Z�0'�3���Pyr�¡i7Ƙ8'�Ȏ2A|�����6q&��̋vȔ�H��)z���V�1? �b!p���%R����f�'�O��5����q��.�-����Y���fi�9A1����N$>5t�	�`��i�(�#$��;G���4��pa�%�%ق���JӰs�<���ܦMx�x�O��z� Ţ$/ 6^�̰�c��n����ѯL�H���
:�2��/��	�(<z�'ʊ��į�.��ԉU(+����䘨N�.P `�0��d@�g�"��,�)0�굠 ���9�4���� �h�B��	Ĵ�cJB�C�FR��6;���g#ٻp�{P�1�~�W<��h�c^CyB�^�f,c� �~�h6�M�iq�A�F�b�6�q��ɛQ�wը���c��3�Ѱ3�Z���L��<�Fd�'e6�ڥ�uv���� M8}�P *&��*]�Uq7g�����n��Ԙ�O�S��I���_�p?��'��OdN0	��"��b�-��3p�غ��� A�
lk�u��!#'�-[J:TI �<@E �'����an�����p�g�'V�8R�����|����8(Pv�H�"�qC�i�V��=G��/�^�+�.�=Ѭ���ɜv�>equ,/�,Y��_�r\��ɫb�T�@���-��Sr�	.�8����O�}��=� d�.)/�0�2$�p���E+X��Px��׵w0��zwT�w&,+���h�Xpd�V
;Z��6�ǻ[����S�V��'^H�9�Ѥ�E� C �%}�<���	*_J�1�®ܮL���{�.�u_jd�$G�(�����ؾQ�v�r�U��G���;q��x���'��-�I�1oH��ȓM#��9A'̟u���P�3.����'}��k�3 Ȱ(��	�'ĬM�ְ�����Lx����*N~�mA"l�0��\�@¸����)3�K	�'��:�"�7�����N>"C���X�WB^��3��`�r�P6�Y�a.f�C��ծN>fC�ɱ( ���t�C_�nj�l� �ɦb.�d��ӸK
�$`�ķF���0�,�1$������y	`n݊e (HTƚ�!�
(%6������_�B$R�F�D2!�d���B�m��B���pe.�#!�$A6�杸t����)y��X?{!��D][�E��J�J���'�!��t+䖄`�+Ƒb��[����!��Ҭ>l��"`�3|��)x��ڠH�!��$w��i���)���A�ȝ:V!�dK9W�` #2OMڴ�@�A�EZ!����X�I@+�V���A$����!������SoGI�z��Q��u��'f�� cK�_+*�ɀ�S!�4���'���;AX)
�^�р�ۻ!΀���'&N�bq(�<1�ԅ�mS	r%����'PL��b%�9\�,4��jRs�4�9�'��
VK��|x��u�U/hz�a��'��1��$(���
n>0 q�'"9��-Ԟg%�0�B���
wi�i�<�eЮ5̆�c�&��}]N\�E"h�<��b�. G�Jlʔbй���g�<rH�]9�D���B(/Ќ����\�<��bA7�Dl�-�'IS�y'��_�<�e�<ܒ5U8�,9w��r�<ѓ+� �5P	�?�B#�o�<�@�I�P�J�*&��ɑ+�k�<y�fN>Ĭ$��a]Ȑ�f�d�<�� >y`��Dm�.�P%!"�`�<� ���pm�J���iJ�OK�U�V"O��3#n�25��	O�E:Z�0�"O~9�Ц^�:ۘ]���9���v"O(iY�.%4���钌_bl�g"O(��W�A''\� wG�7iV�!"OJ��#���1��<R�FֆHdP��"O��@�Y�|�ޥ��lB/(�^iP�"O� q�o��<b:�R��9YB���"O�H� Ri��hC1LJ�G�t��"O!��#M�dih��d��"O�X�R"O�Q�i�S���K�	X�2�.az�"O�D*p��g.4�g�2�D5�!"OB=�¡ѧ]�zLr��)q��`K�"O��j��c�H�@�%ؑ-�"O`s��b�(d;a��̴Ua�"O�0�vl՛	� $RdL�=KE�m��"O ���d�8��%?�@�"OʔjE�PD0���і7����T"OL���#�${�DH�Ph�:}���@0"OLlu�O}�4��w	�Of(��"O�Q�Ĕ�"�kƏ�;��`�"O�4�P��Xj�q�J�xۣ"O����OG��0"�L��~T�Xғ"OFhQE��Y�8��fi_�1~t;�"O������[�"@��häU'"\i"O��YAH0E��9� �8U�l�"�"O��c��V{�EJC-ԇ(&���"OTՑB �$u���3L0X�S�"O��Ud�/t�XI�kCW&&m#�"O\��܏ˈ��iX.J�AI6"O��֣�1jPH�Tm���"�2&"O�ؓ
�R�%�W�����t"ODm��m̕<�e��oT#r�P��"OЀd#�#zt��R��<����'шa�'��\��tqDh�Um��'�pQ���Q;e8�@H8FîA�' ���e�.>&6�����?�� ��';�(Y��˘G���r�H�FV�	2	�'�0HUL@f��%��W
���	�'=�= �g[dnX)�I�C�#�'A�r���^t�%@�T;�lP�'C��83�
 ��i:�G*I�h��'9��a���n�0�A��L�@��'����1N��U88���BM#:����'\�La��-��<��DY_PL�	�'yt�ҵ �<MH`��L�n��i�דZ00b�?����"WǤE+EBS�dS�m����3,�!�$��[`��*$Kҋ @�����s�1O��ȧ���q�j�����I����B$M.uO��"T Htr!�$wJ�HyR��	_��9���jLMI��ȕ&4�IY�:���OJ��f�TX�@���%K����O($ㆦ��.8pWb�@p� ���H3m`�U`��t!���� I����2x�}��E�!~9�y2)3}�M�'A�|;��@ [�t@��olmH#f�C�N���ȓ[�)��5X���9���	�\$�������B$����[�O����D¬5�>y��/�px@��'b�ph�έYt$Aok~�"�&� ��Ȋ-O��a�9�3}�k�^D�@*�m �l�rXvK��x�K��-�]��N�y����*�{���2aZ7�$E�G�'�ޭC�R=f�H)�R�2@�ϓf�P�_Q�8H��'�*�뎱�x�p��G@ɉ�'��yQ��v#�tk0�P�8R�q��y"�P:W�e�v.P�O�(��'�)5�q��i�g���'�p�z@�'����әs5.]�uN���.�O,U���Y�� ,����_'0�Ԝ�(ԧk�&�JG"O
�bF�׬'}��K�%C7ߤM�`"O1��	�W� #�D�zV�E�$"O�\�rm/����$�$Lx�"O�])��<=���`���z?��0�"O��"�nj��v�������Sf�<���.S���NJ�P�S'��I�<��Q�N$����\1m������K�<��P�ZCZ�{��vU�I�g�Ql�<��ώk��)�՛QK&��`�<A-͊
�� �Ο/V��ٴɌI�<A�	�y������
�@tH���J�<�w�Q3F\V}�1ٍF8���A�B�<9�Y"Y�x=z�kEY}�9���~�<���U#:��q�v�Xq6h|f�v�<�s�q�x����ڈA�J�8�Eo����l�(Q���0|Ғa	��BɅ3��D  �j�<9��^�4��=�1�L��$����,aI�@+OL�T�O5D�1�1OPd�bɐ)��s𬃩u�����'�Tp��^=�� �1.	��J@���/Q2��s���1斄����9Ny�T���~�^u���I�ͬ�?��R�7��F�y�%ɱS?�UH��a�r�֬ܯI��)�o2D��3D�T���*TI�vz��	�<PK�'_$��᳌ɤO�#"�dy
FF�*��YwgF�<9�C����A4�.`� !���*T2���@�Or㥈�;LH��qO�)��.�JUQ�I��L��pIf�'��5��� �,g�4 ��V�]u�Lhh�=U0��J E�b��u'N�7�qOVb?yX��[ޔ�R���
#��2T�>��o|X���3 �k���~*��Ow���"kOP-��!����P/�	�KB�g�1��,8��2d{�lI&��=�8��'ʔ����Y<�v���
q�O�� �à�Xxl . ���礝U�>��IP[}h��IZ�⩚@e�,e��e���N��n�j}���3ǔh�O�\U���EͲa�O�y�N
U
�i��֗0 <���(?�O�m ��y�驅��7��Ssi���
�s�������4� �3Ӊ����a�O��]��/:H*T�T�4���Vd�h��I,��'l��q�n��.�h�q0)E��b���'��9�"���F��inF{,^P�6�r�)��/�
��$N	��'+ �J$��9���?5�S�?!�����$B���+H?�z�yC�7A�|B*A;�?�!�=1����J�����IZ%l�&>���4L�8��g�PpL)� �s�6@�69�6�(G�*}EP�@6j��rΨ�'�'�<�x���d��+���8l> u{��_0M���r�*�ݷ��%q�xӸy& ��<1Ǡ+�\�bG�$D
��]�'"��#�k�vVd$>ٙ1	��-����f$�1)2ޭ�7��ݟ���-�>hM�1�RC�+}���E�(D> ���dj��j@0��F� 2���(	�1�dB[����?	��ڛ2�Ǐ6fT�J�A� ���YA�V-��<dVC���-r�ys�$��q��k��+Δ��J��1�J�6k_�-)��ζlk�O�c�wcT��?7�ΑS҂*���	�a^�;�\�K�L�
BB�6���2!3��Պ���"'�c�ܒT�4���&Z+T�nx`0��5�>�Q��0OX��%cC�3n�c�H�6��	c�~�B.�ԣ�"O4u6&�/��qW�����2c�>��B9]!D��?% W �"��Ȑ���P��1ӆ@=D��U��[��9 �R�v�J��G�<D� �u#ν<<�뤆�6yW|U�:D�H��@D�#i@E���6D�ܪ��ۨO���
�-�Qs�5D�nm�6��|k��ȓ|jt�p�/D���P���#�����M�,�x��-�ܨ�p� �'4y2͒̒<��jwF nr��ȓ�r���î:���It� =`��ñ���E2�K>E��'X�9�d�"j.�YSd�;{��}��'����u�ĸ�t��Ճ#@,�I�_�B�CQ�Ǎ_?����Fa���G@�<ɨ������l؞�YM�0<����kӀ�1�E��{Dx�1K��BDZDH�"O� ��"�{��y�����<���d��UR%�Wg��Z9�"}Z#�΄N��J�iVY����(A�<�R��o����'�em&�rLP>.O����ώ)Lx�I1C�Q>�BlM#C-X�	�\��� "�F��ȓ P��)�2%��=ذ�	�p .�k ����3��a{R.V�u,�<`���0�s�X"�p=�_
���sH\��Mk�I���^%�J�8n��9��u�<�Q%��.:ܵ9R�|@F�
��s�!�B-��N�)_F|ى���	b�Z(�򊅞k���J3)��$!��EUj	
�c��t�2���n�6l@����:��l�>�|�'�5
hpx�
?u�ui�'xd����"v��i���j�B`��g-HR=Zǩ��0>��F�f�$��-͢0k���N`؞�ITƍ�c�����Ua���jXt��d�5H�,Y,���3�����[�WG��*��H(�}�'�Z���X:#�\l@׉LE�O�ey���|�@�̖�I0p�	�'CV�+�l�PɁ�ǭk!Z�zI<���WY�J��Ǔz�D��@�H�uG� ��6GL0,��I�*��V)�'�;-�N��"�֞sDLA�Ot٘�f �a�P�`vMRxU���	�;mhH�
�d�1���D�:)�ly#nFE�D"O!�5/�-V���sC2*���d�O�x���5�E�H�b>��D㑂^�j=8����c�b�'�]�@�A0�"Oh��W�muP[�&����Q �k��Q�b��D��D?��$��S�MиهL�J��"H��0\<��dL�_N!Ca�jFl��#,*���0��(T�FdF/>�ܸ�Q�!}r�ӵ~�����&]����"e�tE}r��"�I�e@J�'}!"���2Wd�"aK��T�'D�Da0�
�)�~\��II�&��
��^ (Η�)<0��0V�� �R� 0q��S��gTlP��I�0�,5Pt���cI1h�##O%{�#��8L���`6�3�ēi�`�#6#��q�9+���2D�O�	V5����Aڸ�NE��U��2K�4�jؠG
�I�Ɓ��ߗ{�q1��js������U��u�O?Ź'@R�#� ��d�N%�t|�a�Pk�<15�E�¥itC��V �+�J�my�&Q%$NM��/DjX�����֘3d��JY�����h5�O����U;lLd%@��W��i�,�R�^��c܂��x���Aa�13��Ϗ]k��+��¦��O��Ce�L>d�?�ӄ@�YB
�K'��@?�q&�*D� Q�Kr:�ДK�$e��K�̫�X��i�-YqO�>��lλAd�Lx �ϑ|�l5b��2D�X�V ��K[�}�Ӂ�>X����3D� ��#!�\2l�$,�B�Zf�:D���v�^�N@P�پ1tp��@7D���KZ7-8YaCԎ-�~|A� D�Dj���K�Qc��U��A�1�3D��X`MK	F�(� �)$\�i��1D��0���Oy�Xا-U2�f�as�,D�@IIʩ>b0	A ��B=�	+D�z$�^��	Ҫw�Ƒp�<D�!���&B���T��
p�e�4D�ѷa'N��Ԑ�Q�[炠��C2D���1c�w�����&�-b�iYF�2D�\1���i��4�r#�X�S�0D�@���N�R�n�4̉)@_� @�1D��{�o��"4<(����<������:D�d��[�S�8ze���Ylڭ@"�'D� ������ݪ'�ĥD��}�'�6D�H�2��(�81����#8�Yc�3D�IQǉ&X��)�lA��dm��#0D�`Z�M�f�ư�I=�D�Zv�/D�`QfM�k���1g�ڑ�J�s�.'D��c�l�8I�v(\�P�m)D���d����1�C\�.�ڀz2":D�� "��P��aF0(7���]v�B�"O�a��J�R^��K�C�F�c�"O�Q�
�?L�Ԉ��^�/M�a"O�2�,��\:�5������x�"O���'�Á��b`L	b�L���"O40�`J�*���a��� ����"O�Rf� :cM|�#�#�-I�@9A"O�]2׃_H� Hq��B���%�d�9E���� �T�n�u���1O�
gC*N�0��J�/�  ��"O��y�O��H|ekr#�u�Hq@V"O^��		o�Q9�b��� e�R"O��TFP��rT�}�"<q�"OAH��+���'/�]9J(H�"O�u���\Љb��T5dY�E"OȝX�֨>ҼE�c�V�1��4�&"O��u�Ͳ�J�;�萑E{"iq"O�;v
��tf����c�s�"O�S!?��W��+PV�D"�"ON�ɑNÙ(����>c�"d�"O�qJ�T*zY6- ���,a�z�(��'.�*׹i�h�a�	��&n@Q `A�	?�>�Ӌ{2��z��O�OĒ���n�S���Ӏ�t�%ǁ���3q�
�}���F�,.I2Wǁ 
.����3o�����Фst�'���I3,�`��!I;Q&F���ҜD\v5ˢ*V:��$\�Kru����l5��+�$�$�Q�j�2<��Q^�̚`fI*A���
ç.>"�r�܈
^��q�� ��=��mO���'W*���K��Q9U]�����]]LeY�Y���Sť��t�r
��u�dMc�OԨ��`���7Á/*�P;�a�j~�Oƃ_U2ĩf�Oj~m���L�7S��c�#H��f��(O�H�&�� �X��!��b>W�O��:K�e.`� #A+H�� G�'�V(Y&�B�	3�ڐd�>E��C��2����Ƅh�M7Ş��M@ƞ8Ԝ�M1	��{v�� 2$����D x6�u�Vi�R�\=M���I�!�gRR�̓����Oaz�]�{z@����^�p��$�	�'8�E�2$�#ۺa���d���	�'V$m؄i�A�衡�R�D�\���'&�E	V�悝����@!�P�'s@�C�Ή�s5"E!��	 k����'���)�끁lc~L�2��(j��i!�'4d9��K�e�iu��_h�	�'s���AL<�Z!��-�7J\���'��k��A�7*�M�ÁY �J�2	�'O�p���4F\$i!�E߰^�ε��'�����9>!��D��V���'O0�����!t$���]z �A�'�.e� .%1���'q
~E��'bl�`� �=�B\k��Z�!�{�'-\8x6M��(,���I1���)�'�LL��
�;���O��N���'՞9�	տ��̑��J9=m0��
����,	�%��K��_�44
NZ�yr�V����mƫB�RP�,A��yb.�+�0��4C
�8���	R���y�(J	m���S�\#'�6%1�*ϛ�y��9$�"���]�&Y�YQ���y.S+z�xq��#r�H2j���y�R-$LLxڅ`��f���$I$�y2�&Y�
-��R�\���Q��y�0m�v�`/cI�G`�)t�xy�ȓ:�l�)V��1V���딭ؤz��t�ȓa䰓�fF�k�����J����ȓP�*ܰ�Hϖ$�5dN�/Ҩ4�ȓb�Ē&#�EÜ��2FL�]]@���l���@��3Vh�[e�Z�>��?�@8е�oѲL��.S�e��S�? �@h�BT�pz5@�aN�KpH��"O�ic�iF�{KF��Q #s��C�"O�4�"���U-��rR쀃�"O�D��,��)u���.��c"O��P��O�UɺLq�GO's��'"O|�0�Q�M��u �e�]�h�� "Oʝ��4�n8U$ǣ[�ɫ "O�`�@U��n�2�bP���P�"Oڀ�Q��/��U��2<����Q"O�|jQG�!1~*��A[��V��"O��R�J�/ ���#!�Ry��"O�P1# ֍�3�1�(�`"Oе+Qx��Ҧ�V����"O4q�bT:
(1��� /�n\i&"O �J�bY�a�<S� I�J�4�"Oh��b^�A�(ha �{�=#�"O k�o˒SD�#�dO�T��@v"O�#��=@�m�De�"0PH:&*OȰZ�BD���Q�R���	�'��	�\�w�!�n��b%�@r
�'��p��O��m��`񩀆\%n��
�'���K$��$.�*��l� \����
�'��ũ��Ըp���`�܆A%l��'�\�`���&I�p��?*����'a��2G�طiQ�l��+�,p0X�3�'S����㖡t1��̎ur����'�fAi�����,ġg%
y��'����6L�p�ҥ�M5�R�'�ȝ��j0�2A�eE��
��'��<��f��+�B]�da�'yHX"�'
P2d�Y��C�,Y{)R�A�'=�����D�>�A��Pz� �
�'�ͺ�*ܟOg֭��;D�N̲	�'׌�X M���@ZQ�@*?�J0c	�'��
Ηa�h1�󡖊0���J
�'x���� E(�@�&@�� â1a�'�D��n1 ��a��� \-J�'�"�Ò�_��>	��/l�<�
�'�ʰ����jz�yƬ7"��'����L]-�j� ��©��<h�'�q2�)ا|�E
4F�g> 1c�'C�I��c؀��i�[�q�
l��'h��7�Q;HQ�a�˜Y�Rx��'�@�q���c9�b��]�"Ƹk�'�aY#�ġ/xd�"A̭+;0 ��' 6�Чg�8K4�t���)r@ɪ�'���#��̷��݃G�@�J�'d֝�a�V�"S���f ԾY���a	�'�:�f�.�0I�ŏ�P���	�'O���࢚8Ǆu ����wq��'8ԉPV<\�r�#Z�D�L��'],`�Ɖ�d�me͝�9D^���'�", �ԷYUT5qg�Z�/:�1`�'6��gׅII����뒑Bf�
�'��uI98Np��s���!Ep��
�'�H�1�1Z�����̘�c|F�
�'S��&ed������/^��R�'�H�B��:�ԨSm�%&�����'��� #�M�5���HR�Ƕy��'�^�#���!%Z�x��.�JH�J
�'[H�(G#בh�:��W"y�H0�',y;�C�%~��uh"�hT	p�'���!��C)z��J��+]�0��'�69�f���=��I�ǝPꐘ��S�? 2铤�'ʢ�ȵ��� �<�I%"O(h@ �ՠ �Τ�A��J���0"Ō
$�X�I�!&B~Gj�"O����Ή9�t��"J�T�A��"O�8Ʌ�I�<���!ćE,�Cw"O6�	p�^�x�ִ���L71�l§"OR��Gf�
k�̬��hT7d�
�C"O�pQ��\��l{���2O��̣�"O�cU��,�S����.Xx�"O�|��jD� �r���`)k�tyi"O�@����5f�y�S/���a�"O`I��l�(NS�E�
(2T�@"O|�! ��i�eQu!X�	ܨk�"O�^r�Pѣ\6b2�H��!�D�Z>m��Oơ�2����$!�d��F�ig��#c�5��"�K�!�!��\z$��>g҈9�q�é1�!�dޖnH�@AK7W#�p���^�!�
��̩�	΋nZE2�	*w�!�Dң,�P)i�eX��-���J']�!��;>��I
u
��{��#F��E�!�;4G�PQ�C�\`
�$�72�!�S6\|\�x�#"� ad-4V�!��ߐ2mFAbgĊ �v��FMM03T!�䂿X���8p��,k\�pa͉!E!�dЗX;��q� �;L��E
�&#!�dHB��Hyw�� �i���;a!�:oKT�`�@�G�a0�ȉ�cI!���h.���D��M+����a�D2!�dG�r{2�蔩ޓ*��0�֟|*!��-$~���펇&��q��͗.!�D�1S�8y`�
��L�r�_�]f!�Dx����/�T��1Ü� !�da�P��v��2�z"L8b�!�dZ�N��U���V�%+S�T6Y�!��Ƞ���hY�g�eCP̔�(�!��̋s,��z��K�M�@��F��PyҮȊO��1�c,�+4m괂��y����PĜ��V��-n��ԡ��yb X",��a�u����a�%L��yR�*C,�{AI�)p@���;�y2D���1Ӣ�՞4�Ʊ��(�#�y�� :¸�ԭ�ΐ�C,L6�y��);�񫡢�{~�0����yrHC�5 �r3�A�`��1���y˔����uMX��٠�y"�hpl�ː��a!؂F�>�y�I] *l�AC,Ə\ V 
��P��y���"��(r��׵Y�⨙��� �y��¢)��Po�Y�0B�̝3�y�ۮBs�kA��y\n�dDL�yb.@�Z����vfV�q��]��a �y���9e�T�I�d�v����6MЦ�y2%-d~ꨂ��L1Pd���۫�yb@
�T��`+dC�xߔi��e���y�
!Ԛ��uk�&s�TM[c�*�y�Om�P�(� ۬!�V�yA���y��W�c�j���%�E�.���oM(�y"dģ+dr��aÁ�̄c�I��y�eA�/��<�Vc�'�hY�]��y2b��!��T���	�xh�������y��&c�NE8�@ �r��U{�B˳�y�O֫D8�A�íkc>�Ɂ�D��yR�Ro']�&�D�rV�31��y
� $0v�@�T���SA.]C/Й��"O-c�6i�Jջĭ[(5�H��"OR����ϘQ�r�ѫ�6�D�F"O���4�K�k`����S1S����"O�`[f�C�?�@�	�,$����"OH�p�����(��a��J&"O��(���(B���t'@�EW�I�"O$��.@r���� �B���5"O���u��x�m�3D�[�"O�$"�a� jC����o�-\$X�"OĀ�tIT�Cv������`���"O�I��>4Jb�` ��m�|���"O��G@�r[|���	���y�"O8���Y�P���2 �_�*���"OT���D�QB�9�O,Os�"O�ȗ�V)Y�](�D�Y�Mj�"O�|�����Rp�)rS��WMır�"O� AVF 8�V��l?Z���"O�P2�ǌ'�6����'%�Q�"O�ɺ$�� 9�l@���D	��y�"On�!�O��^n<��f��=M��V"O�x��΄�Gǖ�!@�d��=Q"OؠYC�4F�v�#�dN?���0F"O��`�'U�N���ㆡ�@eb�"O2�Z������a��Ce�j�J2"O���+��j�By���,`�bp{�"O�C��e3��aw�%X�V	JR�6D��*4��z���IS�0�X�F4D�̰U.�*HNt���ܖ'��$�1D�li�l�)�$L���V�E>8�UA;D������]#>Lё+�,t��`�e-D��*bO�� ]�R�P�?H� c�(D��3�N߮���Q�2	�!6�!D��"��Q}��q3�p��|`P�<D��S���u4�Qa�"Gx����#9D�\�҅S�[���,*6n��T$8D��[�Э
d�z��Æp!h6�5D��0�N   ��   �  W  �  �  �)  $5  K@  7K  �V  b  ;m  >t  P}  y�  ��  �  V�  ��  ܣ  $�  u�  Ŷ  .�  ��  ��  Z�  ��  *�  m�  ��  1�  �  `�  g 8 
 , C% �, :3 }9 �? uA  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e�!�S�)�Z%����� �Z��I`n!�ͷ�JP)���4�H���,\��Z��(�*�-�pZ��N���V��YQ!򤈧6��r�7Lޘ�զ�]�$�O(L��fÇ�0�˴E>]��(�q"OR��х�=~�6l�F���
ٚ�"Ö��hY)F^L��!I�l�H��'G�����MP��SR&K!J� �L4D��xÊU�l���ᠪ�D�2�ے�2D���J�p=����ސ!�&���#=D��I�b�".ū掛�6�b�kf�r�����d�%��$h&��n˰E+��/�!�d�K�"H�&�%���s�'\q!�DؙX�^,p*��y�V��Şo!��0��(g�̏R�j�y�JA�e?!�D�-Qv��o=u*@�#�\�m>���)��Y9�һ/�����>ސ�a�;D���rfʣv6<X0�ڏZ�z�B͹<���2Z���y��ӂ+X�2������0HX���$��}it�u�$��TAζI�!���!����?@�hLB����2f!��7/���O
�/nZ�:e,L+�!򄎺o�~}��	=\G��aB�!�d��=SdIH!/M�E2ne��@�2�!��
�Aj�dqE���p=na!�b�#Z!�D���pu�$*L@�� #Y!�D��b����#21v �6���?�!��A Q~�y���*"�<����� �!�ʒr�X�Q����0�_�:�!�Ē<_����eb�
1�L� #�ׄ{�!�dTJ�D�٢5�y�ī��!�$�@h����*ZQ�s�ǩ>p!�$Y2:�~���Mf�W*�3_!�d��7VB�7�ݾ�*4��)�K]!�� v��d	�A� X�������"O���!H_!5�*�j���2��PKv"O�D���C�C�~,H�k"H]p�"Oܥ�Fe؋�P$`ū�	*��1"O�xX����J�I$	�"O"�ғ%�tQ�����mt"O~�4FO8P�=��@��l�Z@"O ��҃_	2fD	����������"O>�%*��TD�٘AiN9Hy\Ŋt"O���S��� {��H����"O���!!E�U�E��lΤ��"O�})uaZv�����y��8"O����!?��fO���1�"O����W�8����
���0"O�`A��Ch��#gk�:k���R"OFԑ���l7����CŪa�Pې"OF�I����B/�aZa�R����s�"O���eN@��U;�Mi �;V"O�eσrf�Y��"�	��E"Oȹz�m_�c,�����v���"OL�e�R.��Xa��a��M�s"OصJa��4xa�H1U�uj""OT[�d�ڈy�'�L�е"OZ=�Ҭ�kz�׻8J��#�ŞH�Q�0 �6\0J�{��݁gC剷!���;0mH�P��9�T�v�C��.nڨ)�K�'6��	B��ހp��C�ɳRox��ᐝL4�)���[pO�B�I�JK&a�[q�8�h��U�C�B�ɘY�$��o���=�����Pi�C䉢t��Е�]Gv��G��&w�C�I�P�\�cG�<'"���Q��
%�`B䉥9M$ Cb���}��D��^�%�$B䉪s�y�1
Ǫz$�aE�δ�B�I!�lP8�(
2~�e�&!�'gNB�q�>�@�@�:��������-��C�I9;)�Lq6�&( �4����9`�B�ɳ>������"^��(sLA��C�ɍl(�MyG�AA��"� �,®C�	
�8�ka[2la0�0PA�C�	q仂��;�J��E�A(�4B�Im�v���(���9)��ս-5hC�	-`��j����P$O�w���7"OB�:m�n�
7m�E�~�V"OVcv��+��
s�U�/��� "O�[mS=$6N��Ӏy����"O4HI�_4��i���Z�5�"OB5	�D<Y�~�+1bP)'P�y��"O��;�@�g�I���2c4~�p�"O؅�%i�_ΰe&�Kw���"O���� �f ���e�4�h �"O��2�ݼvW��bqEF^�>U"q"O�� *��q������uF"���"O�ay�Ӓ%�z]���ָ<@�0�b"OdE�*�q��5�.��A����"O^�r�JT��Dؘ�F
s���"O$��̩U5�p���`ihm�&"ON���ǅ�gV�1�C�E�8�2��`"OH��e��?���Zf�� _�p0�"Ov����->Jq�&,|��{�"O~��h~>}�&f��?���J�"O�I��\�"z�%����0����"O�������|�&��d1�A"O���F�`K��S��u�ٻ"O� �`�@dO�n���sȬX�ԥ)�"O���Ejɩ�9�@̇�*�(��""O��ZLƜg3x4a$�.*�Di2"OFu��Ü0�����k�h����"OHq�q!2�� 	q��K�V�[b�'���'��'a�'�R�'���'�������$e�� r����"R�'D��'|��'"�'s�'���'J�8
I��H�Q������P&�'���'R��'���'���'���'��Y�mֽN^zE�!n[IL��Y��'���'�B�'���'HB�'F"�'�����ث�ByT�]q��P�'1"�'�R�'�B�'�2�'Z��'?�a��m�&9H���"b�*��V�'��'���'"�'���'���'ʈCV
S!� ղ��F3��e�1�'�B�'Z��'��'�R�'���'���r�K] ~oxH�������E�'�"�'pb�'�R�'y��'���'���9%�#I=��R�&U�\��T�'��'���'��'���'���'�h�`Ŏ*=[IҴ<'�F\h��'Ob�'0R�'���'M��'�R�'A.�R
�-nt�ٱJGy��Q�'���'���'���'%��'s��'��e;�`���^����]�(9��'�'���'OR�'���'"�'Xh�^�E�h�#	�9y����'��'�R�'x��'R�"uӀ���O�̂�h3��J��
'|��X��Iy��'*�)�3?��i;`�5g��Hr��� S7���e����������?��<�����wə,#��i��@�������?��K��M��O����:H?qk䈟m ��s�$Dw� �6�Iş$�'�>��`[�w��^�h0;����M+6�YC̓��OQ�7=��X�u�X;b"`���՝�ݣg�O��`��է�O#�@�iN󄃡P�4]��A��bEP���JO��r� ��U	�=ͧ�?�Q��A�P�P���J����@�<,O(�Or9oڡ,�b����+I6^��`��m��8~���By�;~�I�`���<�Oh�J�D�� �-�����>���擟��	�hD �+�- �8hE�-@�|c�m�`��xQb��o�}���wy�S�x�)��<�W��">h|p�b
�=0�`�GA�<9B�i�Ը��O�po�Q��|a�6eg�d�`$�8~=T-yW���<Q��?I�v*��sش���|>j��;�Z�"AI�*��ñ-�%Z:Y�Q�5��<�'�?Y��?����?��	ҹu��;��0C��M�G�]��Ц9X�I�����	ş&?����_K�y���T;p(\�xd��X�K�m}��'���|�����:{e���ӂ2*�QH�q�����iK�	!Y|�I��OX�O�ʓK$�)p�^�c�0Q�s�����K����������˟��Ry�`a�����e�ON���))�2y$�ݡq�dH����Oεnf�Iɟ�!�O�D�O�B7I�t��_�b�@c��p�n���Fy�>�;,v�#��l��M~��;2U4�����i+� �[1z���?���?����?�����O9��[���
�ҹ��L�]|�1�S�p��.�M3�c��|B����&�|��4%G�E�a$U.���c)
=��'Nb���ë+i�֓�p�H�.x���fY	 ?�M�G�Ӭj�����'b��$�������'��',��k�
�\!�L�.A*���'O�^�@ �4r�R�a*O��D�|�2 �L��`2���hڑ���m~���>���?�L>�Oۆp��S��hň %T�+Ӝ��m��8Vp�q�i.�i>a��O��Oެ�愞�N�ܜ����-����O����OJ��O1�2˓*G�Ɓ�^�*��V��wQ�m��$]��X���'�r}�"�h	�O(�D�Y�L�d���O�ZXxQ`Y������O0E2e�c�t�W�ZY���3�5{N�J� w&d�Cׄ@�?Z��	iyR�'s�'�r�'��Q>���C��w�J9����~q�}z��3�M��n)�?����?�O~��ƛ�wJ��@H��_`��̑�/���'$B�|��$���.7�>O"<�c��#V-Ĺqq�\�Q�@�6O�8���ޛ�?��*�ľ<ͧ�?�al�=t}�Bc�N�$Z<���ē�?����?����XԦ�	�֟��	ǟ$��i�4ڴgT=��eYG�@�b��	՟4�ID�	)	�¤W�!e��!�o�<L��C��9�FK^��M+��4�V|?)��D��T!ļpS�Ć�s$X�a i�-�?����?����?�����O�|�SoN!����#(ŵs�bAy(�O��m��?X��	�@�ܴ���y�Ć�Yy��4�2�vi��� �y��'s��'��p��i��	��e�sП|�c�6�t�Ə
R�8'�>���<����?����?q��?���S�~y~X�JC���a+���$��P6J�ßT����8'?Q�	�+�j@ )R(գ�lW� �U�O���OړO1�
h�E��=d|�z�Ô~��YZ���L�^7m+?Qg��?'R6��o�	Ry��H�6-b'(��_"�,Z ��n`�'�2�'��O��I�M�	7�?AU���5�}`$)�-\e^�3��,�?�ųi��O^��'�b�'����1��b N4SdQ8�A֬L_�h�i3�	Y�2}�`�O�q�(�� �\�WOL4.����k�s�]�=O��$�O<���O��D�O��?�x�C���̠%`ҡ�Α�Cf̟@��ϟ�Z�4v�@�ϧ�?qջi��'���P+R(����jN4�9ן|�'.�O��p�i��i��� RTȰt�%_�j�2�Q��Z$y�Ʌ?�'�IƟH�	ܟ��Iw��x*�(2f��q� ��JV.����H�'�r7��{gN˓�?9/���$X�"y~��%ĪS��Q3T���Z�O��(�)R"O�o)����S:s&�V�%����L�*BO !q/O�I��?���4�dڷ%r����.`.����G������O��$�O��ɬ<I7�i��XB�˒f N1��F�[%ҙ� J��44�'�~6m$�����O��o�M�R���H-o�R1@V��O��d��)�63?�;`�z���'j��˓,�"X��(
7E��`mI-J�������O���OP�D�O���|
U� �,�#��L, @  ��Mi���L%p�����&?��I��M�;/��
F���d`
8��2xy����?	N>�|R'I(�M�'ԱH2��;�n\�'a��*�Ƀ�'��ٻ��e?N>q-O�	�OL��ͺb�fiR(�%E(1���O��D�O��D�<yr�ij��!��'�2�'=��gԅ\H,� �O��i�A�Fw}�'���|�dW�~�H�gY�
*����T���$ϲX�z �7�1��Z��2���Ė�m ��[��]犖�c�d��'Y��'uB�'��>���+&��#Sd�/m'���2DC8����7�M�4�¹�?���E�f�4����Z�_�Q���BNa��;O,���O8���J�d6� ?�U ���Ov��gHZ� �E�c�L�Ka� DJ�	]y�O���'E��'�d�0PF4��I 0�^mZ�L�A�I0�M� ��:�?1��?�O~��p��(��,h�m�W		 ��!�CY������$�b>�ӇD@x�T�#U��R����L<\�amZ��䐖_`����'��'��|#PP���$�X�����7���	П���ڟ��i>%�'Qj6�9�b��V�q��QE�+���p��=-�h�Ē����?Yp_���	���I�N�T��0�J%9;��!�T�\��FR妡�'Pz�p叓�?%�}��;lqT���) ���j2�Z��` ϓ�?���?���?q����O��鰤ԧW�]���Ť|U �@�'��'�6���3��O �o�h�I�5�~yZ�N���a� �-Q32]&�`�	����EnZx~Bi��_�h���ć�0�Ma��S�L���#A�VH?�K>�,O����O$�d�O
��n�GC�@q��ϔC���CԠ�Op��<��i�PM ��'�'��S~m�r�Qޅ;0�$�"@�>?!T[���I�$��'w�r����3A&:]�t�	wa`8bo�/4Cf����4����N�<�O�ԫ��1*�}��cV���jQ�O���O$���O1�fʓ%ٛf��:jx5iU�I"j�L�����<�n躁�'��eӺ㟜3�O\����R�} .ԼC�z%�%a\,<����O��J���Z�q���%O�r�OCr�1�A� }���m�n�D���'8���L��ǟ��IȟT�	`�Dj�w����'fǮ`R�ic��);��6M��b���$�O4�4�ӂ�Mϻw���b�ʥ2m|���+�4y��?9K>�|���'�M��'���8G�(O����K�ZF��'q4���N^?�J>Q/O����O�4!L�f�8Da��˿P�X���O��$�O����<�iqlH�e�'c2�'��@9�I^�'Tv�)���*W��A���B@}��'�|rML�&s���aJ�&I�ԑ��ȁ���䔦Z�����y��c>���O���B,'��5��±3V
C`�h���O����Op�d%�'�?��
T;qjR�ڱbR����aB��?�f�iD-�s�'A¨tӰ��]�y��ucE�Ȃd���-5?~��Iߟ���ӟ�p�.Uܦ��'O��K���?j��3��xrI��d�p����'��i>�I����I͟���"o��1M���m����~h�)�'a6�J��O���+�)�O���Q!�7��e�u��9��]��ꓼ?����Şg������:/l��ADF/*��<@1���M��O�t��@� �~�|rR�ȓ'FT4X��տ4æ �F�H��`����Ɵ��sy��OM:r�'ȶ��P�2-i�q3�"�w=�m���'tr6m,�I:����O����O�$`�@�%\�:����bI
=�Ph��&H7�4?!�dK!;P�Su���ߕ3v�T�{Av�	�fٰ#TXP��.p���	ߟ�����h����P�:�ʃ�0ɺ���`���a��?����?���'A���'�?Q��i3�'��œ&�-0]��`a��4u"�8�|b�'5�O�>����i$�I�q��p�:Fh"8-��W@h=����1<�$)��<A���?����?�!��Qjؑ��E�7K��$��?9���d�㦱�"M�����؟ �Ow$x���M(X�ՊŎ��(��Ou�'�r�';ɧ�)۲2�F��a^%���k����-�a�*Iv��<�'i��D	(��b�����̟�Sp��0��`v1���?����?��Ş����%RJ�c�t��Ć8%�d��c@�g�x�	���4��'���?هG�D�d����[�(�Z�ٷ���?Y��+2����4����е�M��N̙-O� ͸���,q� E97�Z�C�<Y('6O�˓�?���?)���?�����i1r��88r�V/��x��mE8梠o�)`���''����'��7=�Z���jT�/��k� W6=ˬ�j���O���/���M�P�86m~�����\s���òv�b�J�v�X�5c���<��<	��?Y�U�	X���F���eY���F�ɔ�?����?!�����ݦ�R�c�������x�G
����G�x� �W��֟4��O���O��O�Y�����RƋSJ��ɢ���K�ז\DtS3�FA�Ӓ]C��ӟ\R1OĶU*�ɚ��,i����Sc:D�5�X�d7���0-Q�]�ˏJ��DK��݁t	Q��I&�M���w�&<���f�H��"�7v��i�'qb�'*螓sz�星�!v����S�X�Ze	��Y&���F�ZT�����|�T�����p��Ɵ��	���Z�
�L�e�_#+F,aS�Ŗuy��qӚep��O����O�������;P��)��
�Dqɕ'^����'�"�'�ɧ�O��y�W�ƩRN�c�%F�6a���!��: j��dP��F�G�rJ�S�Ey�R	6|Jl�gD�.��qر!�����'"�'B�OU�	"�M�1痀�?y��P��>��0�m��$pcN9�?�e�i�OH|�':2^�������HvB6�eR��[
 ���l�_~�IE+o�F0�S* ��O��Ѷ$�� �"a�N��@��j��y��'&��'�B�'����A�R'P��cጀW&j�ڶo(B���O��d妝;�gh>�����M{H>�!dT$���d�D?+,d�d�[���?���|��Θ��M�Oj)ŉ.X�v�IS犱\ui�(��S���'V�'A�i>9��֟�I�A~$��ӧ<(��B�+�	ˈ�����4�'~6�9���$�O@����)ϫH+WoWl����gѕHN�D�O�y�'��'ɧ���'T�(h3�+A8�{������&�6t���i����?-�1�O��Ov�9�(��{��0�@��&R���Oqm�.�P9�%_�O[pu�&�?z�	`-�ҟ��	�Mӊ-�>��	W�{��J��,�Cၙ �"Ț���?I��J�M��OX��� P+���P����!�" 2h��F������j�,�'���'t��'���';�S)n ���'ҧ_Ĝ�A�)
>8iX|�ߴ$�J@���?���䧵?)���y'%�(�	���"S��qe-��'�ɧ�O�\�Q�i�DO!~�J013�B�r=lU�f�H2�$380�'��'�i>����9~�̙�O�O�y(��%v@���IΟ��	՟�'�7�X���D�OB扝*�dƄ�blD~^�,��OX���O�Oİ�c�>0���$1OcT�
q��(x��/B���J�(�؟�{V��D>��H6S|aS�L]��H��ğD�I�$G���'�&$�`�*""��6bUE�VU�#�'�7M��N�D�O�hlk�Ӽ[�c�0:�
&�A�onJ��c��<	����DV�]1~6�8?��f�u8��>N��1���,6��r�҂ig(̫N>�*O����O��D�O����O�љF�%a:)*��9c� �	Cc�<9e�iop��W�'�b�'��O�r���W��`X�'_;�B�h7b�$^�(꓌?Y����Şm�����̖�4U$@"p'B�^�D�#��(�M+R���#Z�1`�-�Ĭ<1�
�E�e�R�s����W$�?����o�d�i>�'�j7-D�_��V/(R��Û��L۠�|f����u�?a\�d��iy�����H��H\
F$��i6霻^�n����il���s�zI�g�O�'?q��'t@��FP>�:��;�z�I���X������W��X�~%�6Aܻ$�bu�g��(nsl0����?!�fZ�ƨ�����Z��'�쓄o�=>e>� r� > �lt�D D~�	���i>��ƎWߦ��u'jU�?2�i�.��6����uPJ �#�'��M%�$�'RB�'AB�'Ϩ�:3D��\���K��Z\P����'^R]��!�43������?������4e��aQ� ���d����������Oj�0��?�)!eH%Z�*�)(��e,ٝ|�d��O֦���T�s?)M>)�Iڟ(
�İ��F�go�2��ά�?���?���?�|�.O~�n� �� �.�p�� ���._�}
v�_ɟ��I��MӍ�>�����R�� k�q��"\�4~B�/O�����aӬ�ө�#JҌ��t!�2x֠�{3蒛y�X���_��^�Ixyr�'���'���'_"[>1�"�J(y� ��Ҍ+?2�$�=�M�\ �?A��?qN~J�Jꛞwn �sCcR<���9,�ұ����>H�B���=|F7�u�ĐhZD9���É�EK�e�w%n��A��p:�dd�	Xy�'a��G
!h`���0�4��g�߾- r�'@��']�I�M�0�Ў�?����?�7�B-V�d�Ǎ�u@6՛�ٹ��'����?	����j�=iAdΆ?�X
��E'P���'}�����t��֙�����īF�'�����΀b˪ĳ�G�����''2�'?��'��>A�I�SJDQ��D�N��(BI��<r���B�iU�����'q��u�\�杧	�}J�%^#C�"��,U�$����O�ʓ�>@cش��$����-q�'d�� �$�#�Y�NI�����##�2�°i ���<���?���?i���?���A�>-�	��O��1�B����dӦ=c��	ן���ݟ��z�9W�x��b�ۦv�P��5�IIH�������m�)�(ߚuJe�Ry@�j�ǖ�K�*���E�'{.��� \v?IJ>I(O�B�#\�T&��ꢪɉ�@
@�'w6�3��DL�0P"4��G�T��E� P���$Q���?�@Y��������	�e�d�#���-��9��O�u�~�����ڦ��'�%�EMYf�O~*��K0��cIù|�$����P�6�~���?����?i��?����Oj�J]�x��N�7D	r&��������4	�j�Χ�?Ѥ�i+�'�:(�S�K�L�I��փv���d�|��'l�OwF�Ʌ�iv�I�
����/�9��v��z���Z&�=���)�ļ<y��?���?Q�d�U7*�� �PzȐrBo��?�������z2F	��l�	͟�OF�=�ש��x+1X�@/�m�O��'�b�'�ɧ��2�`��,V.d=j"���Xq�ѫ2d9��2����d��*�l�1�@�P�Wݞ*p:ä�;���'Br�'���Q��zڴX^��[��@6�N
�6Pi�&��?i�/ڛ6�d�t}��'�`�S���6c���D��/	W*���'�bj
\��֒��W�X#(�q������0q;NuBw�C�	 �@��1O<ʓ�?���?����?�����;9j$8��,١??$\{pʁN8o�f.�-�	ğ�	k�SğL��������Z�"�"C��y�B,5��?����S�'|�@�޴�y"��(	 �qeC�8}{g��y��h����O�=�K>-O��O�a����"%2���%E�X�x���O��$�O��<Q��iݘ���'r�'�,��r�\ؚ�;�bL�kȫU��^C}r�'�R�|$Z7ܪ��!�< ���0b���d=x2TC� h��c>Q���O��$B�0�e��5��x���0����O,���O��S�O�
`�r�H���tY2(��&� r �r�dp:�n�O��$Vۦa�?�;p�����^e�����)Ul�a��?Q��?�b$�:�M��O `ʗ�F��GDK ^�0E���05��L�,\�cȶ�O���|���?���?��/��ã��\�=+A�&F���2(O�mZ��2!�������O����b��&���b1A�
8��F* �����Op�b>I�&�͗�`}P�!�&C"���'�	���hQ��Uyb�_�D(X�	�G�'-�ɧU%,���Ը���`g�4X���	ǟ��	��i>�'2�7m��?�4�DI�)H�H�s��pң�\���������?	�P����韐��!D_fq��@��F��x��HN[�
 8�J�ަ��'l�*0)�V2M~"�;*��1�4�^,��L�?1��͓�?a���?����?�����O�)�+J��p#���p��{�Q�D��5�M��H��|���#���|rM��+��E
� **l�x��γ��'��]������ͦ��'�T��!��Y����r�E69�2d!Q�y���	?/��'x���� �IП�	����@IY�ͨ�k�&Ү9�P���p�'��6�#���O��$�|���V�4%�'��� h�E���p~�f�>����?yH>�O�f1�bHܿg��E�_U1�um�*���U�i��i>�z��Oj�On����W&P볮s�.Q�+�O`���OH��O1�˓)��C�8D> ��爬e�z���R`h؝J��'svӠ�O��DPo}��'���B�(Y��x���@?����'�ҧލr:�����ݦ�|��@w�I�{�j�����+;A;2��j��My�'yB�'s��'�W>�y�D�"]r$��^z���ޒ�M[un�?����?�K~��[v��wqpU�_�$+.�/vfl���'�|����i�4O�1:����Z�?����~��?����'y�'��	ޟ���|���v1j%�ʍ�j��Yv�'7��'�R_�4`�4�2����?���f@��f Ih�å�:�ڡB�R��>���?�K>9��IT�ܳD�K������A~B��l�D͓ƣ� ��O�F��	f��z��DRb+:h��]"�)��y"%�h!g��+`=�pI��%H-bs�LLP,�O���W�M�?�;
D8��h("q���~�Γ�?!��?YV�A��Ms�O��
��p��A���Z%��w���䑢y� �K>�)O����Or���OH�D�O��H��OA�Q�H�A}���g�<���i��t��]���	`�ßX���?.�v�Zw�'��D��̂��$�On�$;��)ͭȳ\H9���p+Ph"�-�y� n�f~��ļ0y�]���䓽�D`���h&aD*+��*FZ�Q-`�$�O����O�4���"�����<��e:|�X,�ҏ(�6�ă)w[2�d��㟸b�O����O����Gm�	8�ȋ�����RN���؇Bu�*�J}��#b���>��ݸe�<�[�B�%�e0��L%��	�����ȟ��I�����E�'s�U��ND ��3b)�%�����?�:�������T�'6�/���>�8��
p����-^��p�O��$�O�I� U��7�)?�ab�O�? ��V�M�����^��  ��~��|BX��ӟ ���\��ܥ�R if`L�8��|�f�@����YyRb�Y(c��O����O$�'6~��@�+Јr>8���e�ځ�'x,��?a���S�D��>=���%uX�Ðʔ�E�0E�c plq�Q�擉|Wb�ZV���(a�N>q�u�1]�}���Iܟ��I��)�Ty-a�t�@��1����Kv&%�SNC�i ���O�eme��2P���� j�Ϗ��QW�w���FPy�e��{<�������"�3p�D�@by��ٳ5��$�ufA[���+���yb_�H�	����	���	����O�0J�`ܞk��H�i�36$,J!kdӚ�[a��O:�D�O��8�d�Ʀ�{
�k����8�\�o��8�F �I�h'�b>�˷�ɦq�A6��R�G����q�P�/�d�d�hP�dK�O��J>�,O�i�OҌY2��'u�u
�%#b�L0A0C�O��$�O���<!�i1� �B\������(�2��X�B�H(4׭$J��?QT���IZ��>� �����=%t��r�S�ڴY�'zJ0A�
hV�}KU����N˟hK��'�v���?>���G�FL=D�u�' ��'���'��>��	=6U�p���>"����UKܨ|��		�M��얾�?	��4e�f�4�� q%��Xۋ� ��)�e��y��'�"�'"��ʠ�io�ɼxR�YQ �O�pj�HB�G��;�E�~%���FKg��Ty�O���'J��'�jՠ ���(1c�)[��a�D$(��I��M�бM��㟀��N��\b0C[5 5j(:`�Ԓ	���������D�O�$/��IED��a���&����Rc�1ː�jq�j�'��Y�E�N?aL>�*O�m� 'ٗ�����d	9�Z$����O��$�O
�$�O��<���i��HHd�'�Rq�УI�,E)"�UL �`f�'��6�"�I���D�OX���Ot�F��
��щ��&~R���8+4&6-'?A���.���Sr���a�``��n�r���C�8s.P+�$w�<�I��T��័�I������<�q�`D?���2EH��?����?aB�i�H�O~�)`ӈ�OV��Q��h�轂!P=A�@ta�d4�$�O@�4���klp�\�U~���@�u��P���	}u�p�H	�Kl�$�����4�����Ol����m�$,�:rr��*�d�O�˓fl�VF���2�'��_>	 b��Zd|��QL�A^d��D;?IeS����h�S�	Y�E�DjEjhy6����_<���+�)[�v�yS�擭%��^�I,Z�Q£��d�z�Pw�7�����`��՟��i>Q�ɮ���'�07m[�2��i�ILqM��S&��]^�M����O��d�Φ���py2�'�r꓁?Q��=BVqaD�\*&D����?���z$iٴ�y��'��H�Z���	z~R��9�~I���' l���!t��'i��'l��'���'3���L賋��Y̎KrDV�c�. ٴu�u����?	���'�?���y��ÈIp	C�9c2���K8��'4ɧ�O􂐐R�i��DV4�,q0 �-�@ī��kR}h�A�H�OX�S��AX�z� �$�p�A�)ʣ�0<���i*�pyP�'�b�'��(�$S*�4E���ĄLr�x t��]R}�'M��|��s 8c�NG1k*����'��D��B֌!(��|�"I%?YK�O6�dZ�w0:�(��2�Tӳ�hv!�DK�v��`��� q���K����.|���ͦ]r`
������1�M��wӈ�ɀdďPc�l�3ΐ>n��
�'�2�'���V�x��f���(z�����8�hRB��c����!ӵ��bu�|�Q�Gr�H���Y��7��0�σ��d��{0����I��:�U+0�j���T�bW��ӣ+W.]D�I���	^�)��(��CBK���b�*�uKt�� *OR�����~��|�\�����T���ԻeS(6���e6�O6Io�<d���5^y�H�(�4q	j�6�:�:]�I$�M��� �>��?��~CE:�-���4�GDT�@)��M�O��]����o"�)��2���o��P�����	�0M ԪQ1O��dZ�\QXE2�oE�Z�|���E�Ic����ON���̦�GK,��i<�'B�7jH�>�2�C�O��sn=��|��'3�O��l�ӽi��	�PF���f� c_"0Xq��. ���:Ld��(��<!��/;ڂ�!�k�/k�@�[��O�oڪ/�2x�I�IL�ԫ��^��#�Ȱ3Pr�E�����S}B�'=�|ʟ��B�ɂ�@`�ٰ��>���AL,i���(`��.e���|�CC�O���I>1�*T��\�"lY!��T�ס�X<�4�i���2�/�e"�����W����2ҧs�2�'-�7�5�	,��d�O��Q��J	�J̳ǫM��������O���(F��7�5?�RN����fy�&BAb601F=[Y��R�=�yrV�`��I(9�XX%��f��{"�ʞQ*>m��4�J����?����O�T7=�޴zDd�4o�����{��u�$��Ov�D;��ɔ)]��6�w�� �#'�HH^�p�ȋB7��@�=O�T��e��~�|�Y����ӟ8���F^��$IA�
��\�P�o韈��؟<�I@y�r�VљSE�<A�V��ex�Q2L��[�h�P�y��d�>y��?�K>�����6	�;E~Y���F�U~b��%%��40Եik.��*9I�'^�ҁ�����]�^-p���)	��'�2�'�R�ҟV47 �����-� �x���+C���OP@:��'m"-s�T��]�8�n��1��8xxT�P Jk����O����OڜɃ�r�d�� �D�?!���F$��|" ���sGLP�IPy�'�B�'��'�K��
Ja[P�O:�ljQ�ŵ1��ɏ�M���?���?H~���"� r�惦z�I:g&B�)�´�6\����ٟD%�b>a�p^?/�F�Rp�MR�������ަqR/O���E�E �~2�|�R�0����,�Kge�}�<�*������	��`�	��Vy"�z�0)З�O�A��ΞV'X���)���%�O��m�k�={��՟��i�UA�ɓ;w�!�pnJ��r����t%�mo~�F\0.A�y���A �OQ�O)6xq��'4$��y�r�J��y��'0b�'��'W��I�k<,*V�I�&,) �X<ڔ���O����ɦAz�c{>U��0�McM>����I�T4���3�<��������?���|�'�L��M�O���^�X|B$�H�6��e�֮ײ)FyhEi�O��"I>I-OJ���OB���O�E���O�de����.تB� 0ʔ��Ob��<��i�>�qS�'r��'��*wx�2K˿t��Ӱ�FP��ӟ��O��d�O��O���� ��D�0=���IV�·3
�Z�B��!ѓhLy�OlX�u�M�K>��_5%���'�X�U�q�G�Q"�?!��?����?�|�/O�o�X<Y��OQ9*7B�r��I'$%�@����䟼�	��M�L>!�[��	� �tz��JÇ��z�4��ȟ(�	4S���o�T~�D��}�������$_" ���@��vPV!!���� ,�k��9[�)���h��hCԴUBhSTB��bx&�����<$|=+�DN#h�UKE"ՒnF�ysA��.W�b<����:J$�!�G��p=!���WwTq���%s�tYfF�*���5���v�'ϕ�VL>��i�C_��p�+o��˅eA�>���C��(XQ2 �϶2 �!q�'�d1��"�<�C�C{������ �r��ʸ.8fD��-�4��3*���ݺ:��U�ſD't���� ^̛�'��8O�D�>�-O���K�m�Vɠ5d 0ur���S/�¦Y�����D%�����e"�Lr7��)2�A��r$X<Y�i�r�')�D�'�����O@��7 9xAJD�)-~x��ZB�1�B���n禒O����O>��;����"�`��r�Ja��l��<1F����D�<������#ե�0�쵣t'LO��b��b}�Y�
iR����ٟD�IHyR ���b��!R]$B���C�534�0�aC�>	)Oj��"���Oh�d�2vz	�0�fp��h�$R�A0��Orʓ�?9���?�)Ou�3���|�4��4�T�s�C�\���W����͗'�2�|R�'��'N�z�bjډx��1S%H�h�|Q�/W�����?���?I-O�8�M�Q���'��j"hF�A�vc�����b'$h��$>�d�O�d
4���t�˕3\�0}� dΪ5H�c�Ge� ���O��ed���Z?���<��'W��w��5�4,�RG���P
J<Q��?1�M��?	L>��Oj�m��
ۑN�@p�/�{
�H��4��d V�\�o���x���<������<u��H���8���2?O���װi���'�"\���#�S��,tZu/C8k��`���ƘE�7��g�~hl�(���<��y�\�x����	d�(��0���`1f�:�M#��A��'���$U}V�{1��&\񦱢��
����n�ş����<1�%����<����~�C�Tʝ#Q�D�G&�{�gX��' �Aw�|��'��'TR�R�J
�H::��Mіii ����g�P�ɴ__"$�'�����$�֘�K�~$p���k(�[���8]� �IptxK>a��?�����V;K~l5r��ͅ����U*[�֕��ǋc�꟬�IW��jyZw�H1��(��rqa��O$܁�4�?	.O��d�O���<��DȄO���J81�$yr�k<}�Ɛ�n,�������~�ky�Ot�d�Y#����dٲ�c���O��$�<�Ee��(+���"rb�a*T-z��$��[��Im|��?�/Oz�	�x�A/�Tqauc�=�B\����M����?�+O���2��A�՟��s�]`����)=,̐1�׳\���A�(�D�<����?�H~�Ӻ3%�>h�D`��5!��
u�@t}2�'��!�'42�'4�Os�i��S��0=�8�QE��N�(�!�w� ��<!�&p��ħI�D9�5��d��33
�X��n&.�����4�?	���?��X����ц�hdJ�,JC�3�G�x�@7�O���O��O�3?AEcU�m���� ��K�����j׃vi���'�R�'f�s�^��'��Ɏ�����(j�M�LC�-<ӎ�\X�'�?��'�X1�FI5Q�`�cB�-~��M�ߴ�?)�C_���$|�D��_��L�$��4 �K�,ݼT��H'��`�&�I���'u"	!� �(���z<�y# �W��{AL�"���OZ��-�	럼��v�F��0{�P��B�d�dun����?���?q)OT�)I��|򡈛�G�u���ɰm�佐�)�f}"�'�|2]���ݟ��A͊�'�����@�e�����*϶���?�(O��$*!�ʧ�?�D v�z��O�Y�T�0��K7!����d�OX�&(�0'�|���8���'�� �J�t���D�<�� ?.pP.���$�O����Z����'2��æb�qhdUkךx��'��I3Z��"<�;"�p����P*V�C���/N��m�zy��f�6��\�t�'���a+?��N�b�� ���s�����_צѕ'v��'Ӻ�쒟���N;l�E26�
iW�I���M�� 
:ś�'S�'����8�4��a��P[.|��!R:��%)���Ϧm�IΟ��I{�)�'��@���.բm#��e�$ӥ�c�����OR�d�@�v�S�$�>�%�̳uh6��w(�.c>�*��=&m��HH|���?��3�r���Ėr�����fJ2�u�i"�i&P��O��O��OB����,7Q0��6�U�y� (Зp������'���'��S�|�-�d����2mJ�/dy@��;�`PN<���?9H>�(O�W�Z�����F�#�8B���e���'��'�2\���	�|,�'J��9)�P�bB�E���\�v�oZ� ��a���?9,O�%X��iw24�d�=`�T�5�هj �B�O����O��d�<і�Ő^����0�D�d�(`g��O�I��$ũ�M+����d�OL���O��C�1O�ʧ޵˕`z6)�f	J�`]�H��i���'��	(M��EQ�����O��)U�{B�`5��1�\3&@�klB��'42�'��#����D�<�O�:\)�g�S��8�&������4���%(��o��x�I���������2�A�(n�����2�i5��'�<�'ErS���}ґ�T�f�����;�Dpc�C�cQ��%�M���?����r�^���'p��Vi̵}��]SǊ@갍ٰ�q�q�p<O���O&��2������K��1llIЄ瑥��[��M��Mk��?��x��Q�H�'w�^���ҎW�$�~�1p@�:M�pX��i\�'��ġ�����O��d�O��##PfOB Ŏ�/�m0�Ʀ�I�Y�8*�On��?�,Ol���B�*��R
'��A�D�_ ��S�U� ��w���'���'n�[�Th�B�4Ad�����@5��d:�#Vf��O�˓�?�)O���O�����ԅhP�H�u�,D��R�w|$��;O���?����?y*O�������|�ƣ�0t����3���D��˦�'m�Q��	ݟ��I�u��I�a�4U�'O�4s�(is�I�2|���O����O2�$�<3��Qn�S�P�W�X�X��䈗/K�cORl�BOܪ�Mc���D�OT���O�1�5O2�'���HՂ�4@ȶU��EU�~|�ݴ�?I����J3[ך��O�'��T#>l�<[3/KQt� o�IcP��?����?��N�<�/���?EAC�^�Kt�5��~� uӊ�6�d��i��'��O�~�Ӻ��aדaJظ�왡ۼ��P�����I۟8b� s�,'�0�}�C
ˠCʸ8��!̎�0 -�E�����M���?������R��'`a���R
	*��s�Ύf]>l�u&{����4O �O��?y�	K5�U7��0bs\9�→M� `x�4�?Q���?��Pp,��py2�'��d�/N�L�7.U�=��c&��-�	~yb]#��4�0�$�O ���%�|T�#C�d�<�`m�k�H�o�ϟh�P(�����<������Ok�L���I�,�&^7N�hE��U���6<������ǟ�����8�'��u���_�)8���G��-�vp25�4O�����D�O@˓�?y���?�0���3,&�s3+J�?�Լi��	�0�r��'}B�'H��'o�I�,%:�O����4lA��8�jU;]!��ܴ��d�O���?a��?9�J��<��IH����h���U����%/x���'�"�'�U�tA�·����O|�BbD�j��Y`3�U�N[ �y�ڦ	�	{y�')2�'��z���4.�"Q��׃M�tq�M�x�}m�<��nyҀEHy.��?����
DI�^Zr��a"яw=�Q�����R��ϟ��I֟p���`���y"ӟ~iÃ%�FX�+�2?6轒��iy�ɱ E���ٴ�?����?��'+6�i��FfY
~D= ��G*`|�r�e�����O���4O,���y���ճ+�r,IR���"���Ta�?Z-���%�L7m�O(���O�	Li}�Y��aԠ)6��8�t$ˋ>��(@KS��M+����<9��D�'�ؼ8�ḍXj�ij�C�S�е�"e���d�Or�ė�P���$������$��V,�HҒ,�,k`�Б�C �Al�Y�CIt�H|
���?y�1��|�*w�<�R��C*v����Y�rM�4^�OF���O�Ok�
,(��#$��*�B�@�E\j-��"lG���{yR�'�B�'��	��pIq��$By`9�����
��W+���ē�?q�����?y�5��h��T��U��,ŋ]y�ES�.� ���?����?I-O&]�M��|�T�һO,�%H��6^)Tp9&�s}��'��|��'B@ӹ�y"�݃�BE�0�)ʄ5I�ˀd����?���?,O�q3EDp�өЀ �X�i�:"�fmѰ)L> N�}�r�i�R�|R�'�b��y�>��$כj����1Gˠ=��1��
�������l�'&�K�-�)�O��)՛m}*ɱ��Թf��ˍW}�%��IןQA��埔&���4�:�pa�r�� �ta�>vogy��6s66��q���'��#?�	�B]��¢[>
 ��s#Ħ��	؟ȋ b�&�d�}�Ă�E�r��[F�!ꄅ���ና�%�M���?���bs�$��p����S�	�h�f�ͷUf8oڣ?�0�IU�[�'�?��C��m��a�U�vCX� �
58ϛf�'!��'�髆�9�Iڟd�,׮ٻr	N�;&�X �ے@��AnZu��P�H��L|����?��k�����
]= ���a�
4c���%�i2���]�0b���Ie�i�]�ԋ�6�� ��˴0@�V���D�����d�<����?���'WZ�H�rⲹR�����D���a쓁?�M>���?g�R�&&��@Ί��"��M�Y�fϓ����O����O8���O���-�O����ŞY��(!�X�l�`y�@��	֟��	G�I֟��'�v���4}Xr�q&/ܡz��,��/ɜZ�fP�'���'`"S�$;4�(��	�Op����E�U���Rum|�EO_<����'���$�OL��pAgʎw�&QVk�3��K��w�d�D�Oh�d�O�U(���O��$�O��$��LY�	�>[�$A '$��y�,[pK�Q�	쟰�'�$����Z@xq��Qb6�R�B�*e��Q�\���I�imT�	ɟ��I�$�S埔�'Oh:�	��V�G� 	xejM�k-�Hn�Ж'�������D��E+rQ%ăi�f�I��ϼ�M[�>!��'s"�'c�DH$�� E�Y�Ӯ�	�R	uiS�6[�=�	��?�2�2	]�Pt��6��x��_�?���'���'����qh!�$�O������cFD5Dt�J3f�I�hYA�%�I�4�Zc�d�	ʟ��I����VN$t�cd�. �^��ش�?I���. ���^y��'��ޟ�X�yt� �$L��t�\SA)J H���%݈ϓ�?I��?i��?�,O�I�-;_�� ���uyR���4��}K�^���'�W����ӟ$�I&KE��80�ͥ.����h�)�7f �IП��IߟX�'��s$�>�`�M��̙X�N߳��ř��}Ӷ��?y/O����O��4g?�P䐥`�1Q�ԳƁY�y��aoZʟ���՟$��uy2�V(����?�1눴��E�S`� ��)@B�nZɟ��'��'$��>�yB^�i%�K)ԑ@��� ��$W��M[��?�)OV����Te���'m2�O^,łS@�,˄��l�+�,y1dD�>Q���?���M1>�͓��9O���C{�(��3N���T Q<_#�6M�<9Fꖦe��V�'r�'�4�>�;DݬE�T�o\����	G�l�������%��	���9O�>���&?'��[�	D�Fb<@���c�Ω��OЦ}��ڟ����?I�O��+YEr��W�8�(�U�Z�%-���i�����'���ߟ4�����H×l�5[9��PT�
>al&��D�i���'���26l.���d�O��	\�����R��)���$�d7��O��d�O��ɰ4O�S���	���{6�Z"M����,
%�^�i��4�?�%�F$��Ty��'[��ԟ��}j$��/���)/v7��O��a�4OP���O(,��L����'5\ ��-��pb�����.��1 �"OX�3Ŧ�""���3RHZ���#��I�Sn<
�Ȋ�'�����ѻJ�~���'S�3�VЉ��:7LhDX&gռ�J5�2��~���ӃD�knn��q*V�ڙ�"��O����g��a��,�Vcź)7�A�%B���<�e/�d�ȉ{3��B�)���V��h�F
��n1$���C���Zӆ�$`�ak����P��|** �@�֜"7���X�3��9� �d�O����W*-� ȏ�P�<C�`ت$`�O<��*W��5��隷��U���R���U0?UzD+�$��
Y�T&y���LA��%DeC�B� 6(4�V�8�>�`#���ԟT�:��4�����0HN !xq'T�<Q��>��r#��4?ˠ���3����I��ēt)rx���56���p������Y�6!J,j�S���i�D���2�'���La�hA�J2c���Ӷ�R%Zl�em�
d�H�[L�e}*�\c>��� r�'��<,װ4�elM)4�^Lb ܺL�P£)�����O�U��O�o{���Ӭ�{���M�/д���O��S��~�hђ���ҥ-�1�4E�fC�I t)�1;�m�e��i�PCP#<���)zFA�&z��L�I��=�]�?���j�������?1���?)�I!�n�Ol��!�aR�e��"ʜ"�D����gӐ�Q!��
�0pk������۞~�A����.:�
}3�=5fq�	0}��P��L]� �U2�՟ў|I���&B�I�q�fZ��q*��,	�L�O���!���d�D�ݣt��Hc�a�k/!�䇣�^p� �Q�F��\j��Ӓ#F��Ezʟ,������i9��m��@3dh�%J$��'�B�'�R�=�'$r(K
9�T0�3��� ��qG��I�*[.��Q�
�O�ĤRf�?M�(� �tXg��Oef����$^�~��T�!�O&����'�ԩ>�
��:#r �M!V��'��'��'�OD���D�Pw� �p�0XZ9{�'�h�J����%�@dS�*�',=��И'�6��O�˓ S���?������84V��4#׊W�\�A�(>�J�G��Oh���O̣0kv�$��'i����_�_@��a���>�f�DyRj�.L�ʄ��:kp0��,������
���<�AI������̟��	A��# >Vxm@ H�E�8��ԅQ5v'���s��`c(u�ڬ�RKOY^� {��5�O�5%��‌�,��P��E�6��gs�$��cI%���O�'RH	���?���V<,�Dd�g��'l�b�.����w0�EЃ �g�T>5�|�	�?f,1*^/�i#@IA�c�Paq�Ky�DوA�2}���'���P$?i���`�
�K@�A	�!O���'�"�'?��:򺨸�G��={v壧GX�>���O���$��)�BB��er�<0�_�+2�P��D�|�����T��#� ۞�`�����x�m��,!��cHۀo�ؽ��(��yRi���N�i*EXt��!Ő�y"���"ڀ���H	z�H	��KX&�yr	��H�:�;3�֡i�|�3tώ3�yr��%[�5���4e���Ώ��ybK�.L0����e��-nD@��'g\�(7�U;=��-���v�x���'�P�*�(G�hXp�k���+|�Lmh�'����D��]��«�ڦm�'XnPم(4gIJ�b��H�Gk���'�nQ8a̕BHi�/��-"�'O���h	VlT�����=(�����'N9Sb��Q�j����6�`9[�'c�u���%��=*��^�3,���'��q4�5dV��ᘟ&��8�'u���47Mt�2���05��1�'QHAiF!��$�h-*�`B�4��� 
�'�@}3�m�(f�>�C�рC�DA�'A�@�C�
z���r��
J��m��'W*`j���	CWe߯G�N�X	�'��eH$�Di����կդB���8�'�4IQFMQ#b���B�3'xUY
�'�6DK�-�4
x-��NN�Bݰ�y�͈�y�4����Z{��y���-INH�5|�<�+P��,�y�`�0GT	R1�>x�(a���	�yBfX�S���a��[}���Wk	��y2ԥ1 �bPI�<ZҰłG�9�y��*��$#� VrAAv��#�y"�O�����]G9be���Ӱ�y"� J#\m��/ŗ<��U8�F�yr��A*(��U·�T��׈4�y2���4�,�c!/��!���?�yb(.g���Ua�ud���Z��yA�j�p�9�
��� Ү�y�31M+�N�x��vᑎ�y�����(Y!F̕�8z�n	��y�!C�!=(Q"\!w:V��i���y2 �'|b�i�� �(LԢUi��y�(1A���㈚��q3u.���y�'ↄ 4�ߔ���*4
��y�/ï3��YrWL�9x�yj � ��y�p�Ȕ��i��C�! �F%�y�HզR���4J3K��0�6���yB*���C%�	2״�����'x��A+7᲼����mpD�K�'0*�����Hz�;!��=_���Z�'��T�0�j.����yE�0�F"O� �1
Ys5V�`�@] B�=�"O:�Y�]�^��(���)I'L}`�"O��[��,�t��$ћ
}H�"O8"�`�^��9(�	]�Mr�)�2"O�0Ydk�>�*���(Afl�1V"O���$FX4iy�upua�C��`
F"Oz SQnҒ��83�`���kP"O�t�����s(�Aч`�PTܢ�"O�Mi�'�#�H8�QܛO �ak�"O�d�DH��8T��	Ge�(�"ONs��+F~BA�_�1Jh��c"O���YKp����&�"0>���"Or�тOӟRE PFa����"O�=X���u�.	�W��l�$���"OnYi�CA�ܰx�M� (oNh�g"O���b�EZ��9`MS<TJ8T"O2X�g��,2�h�J�%3�b��"O*H
w����@�Cʟ a��q�"O�ؙq�}L��ˆB�&q�Ĳ�"O(��Í�٨%`���&xD�h"OH��5\�n)�E��^8%��"O��Hת=2&���aT�d�Dw"O@�R����
}����2u�́�"O�f��B�p`�A�q�,���'�P�E�Z��i�CQ\�p���=l�JB�	=�8�3�	ޒ2���2�B^�AM�c��rpB_p}B靋J����~�����@8�x�a��B��)�`XD�<�eH�N�葡)اg�̭9���D�I�.�޴g6J�F��O��4gT;I���甔_ɨ�{a�'�~$�敉ca�S��]�C�`Es�ӎkZ1��F�!J�{�Fg :�������<1�n�*[�XD��,�4���7hK�'~`e�͎6:���@ ̼)��O$�H7�K�R H=��_�(���c�A��p���k��Ձ�p>Q���x�@)eZ�4R�N %�z�����1.�� )W(�S�2N x	c�A+aR�N ¼{t/@ <�vu#�]R]��s"�{�<�ī��^�,��M� j�jDh2d��+|JY�7l� �D-���_�B����D�����O�(��Ѡa��nD��$��C�
-{����a|R`�3]������1ے)
(Kf-r
� [�����IQ2�1�h�g���
�-̎uBH0ؔ%�O�9��M�"u��Ҧ�x���	/u"L1���%�1�@��-ɨ�S%F�'�T" ��U�$P��BŷE�@�H%OM��N�&D���د`�*��ӨZ< `ȸ@�[7ny����[E*����k�<t����� F*��נJ8(p����Z5jq�T�s�q!�i�;y�T�G�_�.c!�$��wzJY�r"��#���)͉/��Y{���<�4��T�>Q���V��Ja��	��@�'zf�j� ��(>��QAo=A����'��l"�/X5{��3� �et��R�Ǎb�"$��K��5"b�R@˓E���+R'R�-<��X�B����	G�Q����dߊ(Rց�<��lϪh�ր�%,Z88�5�@�*�v�'���抛�a���2Q)�%
�[�l(<q6l�v#�L�XJ*p��E�\b�9�h�QĦi������>�'b9�qͻ$�1##ܛg�`L��B�\Q�ȓ=����e�PѢ���	7n	�?!$��!��PE�(q �Da�Y��Y�y�y����Y&�𺷡Z({�z2`��a<�l��'�f�sWM�+^q�1O�jhH:�C87U��V�'[sੂn��s�����$^�u��0iv<���_%�qO��ç� ! �!�f�ì`���J��|䔽Q�MX���]�X BՍ[�N؅�A�LHsTs	� ;��
;G�����ۤt�@d3���C���q �?�C�w��Di�a��cb �B5�Zh5<� �'�^`Rd�ʁp��0�&&'0Q����d]z�Na�4>��X;��X�1O�,�BMѹO��*�Ȏ�WP�h5�'��5���W�)�p��,�/<��HX�HI�uo��1 �PN���gb����X�H[��͆�	�5����u���p5pǉd��#<����� a��aj�(4�M~�fB��B����:R�6E+ 	��c�&��'�VI��LM��T���V�
$�S�`�?���� �\%[�ht�TH�����9�(%�@d]/aE�HA"b'u)�t��"OZd��MZ4���1Isj��Q�Ux_qO��*�OR2��Q�X�	"��Q�_��P�>Wp +������pQ�8�O,�h��U�#�$U�� �s��O�o3�H��A�j5"��'���2+��I��@�R+�-�p<�wČ�yzMs6�Q�=�2͢�H�'�ڀ�s̜�A�zLq2�A�}2̠/O�\@&�ݔd�@�q5���9x�
<4�T��#����pG'��sӖ(c�m�v�`t*�Wn�e2wf�C�,��&e�>�}�1 q�v��:"`�GJ]�E��5��y_J�� O�b�RH�Ɵ��ऒ�d�����\���S^J�T�Njܓ����N�ΐP3�������I(#}��
��N1V�xZw�ֆv���3ψ#A�|a#��5W�~��,�X�Ih�y:�����	 ��Գ�'�8y�F�N��A����G�	&���"��� �H� F�\��!��Y�m�����jT\A#l��Z���� \u UѤ�8%�|�������z��'$�
!�M9�<)d��S�jB�	�� �Щ_�S&�0 F朾:��94(�K��	rg��+ ݁a�]D}��_�I:����.��~^yt"��p<I�Ǜ�,Rj�~�Lc&��k�pGD���ZL��q�b8�B'�O�9Q�S�(�� 0 �"+��
g�x�@E+@^�O��8Ȑ��Ou��7�W�Y,�L�0 �bhb�
�'�h�a�4p�<h�%���U�
�'ІP2�J�V pA	t��D�h�#	�'ߔl����N��h��L(?d(��'��19@�"�J��qƔ16�4]��'@��� n�)X2�	�mD�d�`�'�����I^�/�,��W#�U�XD��'U��a��{)*%@�Ē.zy#�'�0`⣤� �~Y�F��e���b
�'�6��k�	{FH�kȿ9��	�'�d�:5�2�|9x���wW@�9	�'P*�*�� /�1��Ԫ&6�I��'i�T8G��-q��Ri ��@��'��4S��\�y�тȞ��Lz�'��S�#�g���9�$+Gԍc�'�hS�]=4DɖJ\�vY��'�j$�p�A+ �hM8�gD#g���'u��!�O�f��]�u��V�$��'�R��ҊD��X!qEꐆ:,���'���!��6.�R�3U)
�섡�'xp��d^�	���jt�˵.p�q�'����7-0B�N��C:~w�`k�'B���%�D'��q�)ʛzʾ�*�'�:)Cc�ɰ�"H�i�&'�|0�'�\�s%U%[а���
�!*�a	�'�8��b͜	l�%�T9Ĵ��'������P������<w@�9�'�!�L]�BƄ�)��Lw��(��'�� CG4W�,p *D�a�	�'9�Q�N���,���ǮEah�y�'Č�xshALl��-�8P�|	��'���Hֹq��$Hǯ�H"
�3�'ܪ�"c �m~��B+�y	�'�fY��+��R��vt�8��'l2�##%\0��E�PM}EDD��'���H�ϔ`�����K�fR �H�'P:�y�E�>m����6�v8��'�Z<*lE(1el�#�S<-Ob9��'�n�9Ъ��+,q��T�n���'��a�.��s!l�@ƫ®l_�YI�'�:I�$�Z�*(�hEnF�`��hB�'̎]�`�)?b�D�1c.\z�'1PJ��܆�<́��Fqk���'T�0�O,w�1	�!��f���'b�\��� 4@�rKE+V�ƀS�'<����;
aF|I���<���'�D�X��|h��a���-�^`j	�'����FU1G ��I--`~`0��� �A��[�8@f���)8.*���a"Od�0�@2\F��He�)^	�<Ҕ"O9ЉԳUUP%X��C�KXb�0�"O����Mśk"�YХ� Q��X1�"O�ɱ��N�)݄@� �3f�]�"O �B�;@���]'GRJi{E"OFq�aX�0��
�+or�yC"O�����2�T�zl,Uv$�f"O���d�X;�5�fϏ47j�0�"OJ���)ϐ!G��;�$�$p||�"O���	�t�P��&v��qZ�"O����cP�-�0F�B��\��"O
�QDHnu¹V�W�*ڬ��Q"O4�����>�`�)��|q�"Oq"��	0d�		���,oɞ�Q@"O~����I[X1s��S�E�U��"OU	��R�@z����שmV�:#"O��A�h��d
g�M2�@�"O�A�ra��Z�*�Ŗ�K��y
t"O�|��W�g�p����27�"i�"O8��ό�;�He��u�P� "O^�8��ղ8􀣤��1a
��W"O ��[��AyQBW�V�uT"OV���旣�Ҁ[����)h�z2"Of���o	/jx��c&G_t8�"O�I��W�9��%��x)�s"O&hy��-�*Ղ��2she� "O�a�&�)���PtC �
��1��"O�z��=g���6��Ab���y�G�3�����l�,z�@:a�d���Ri@���`G�4��D1uc����ȓN�FQ�dU��⹪�n�^FdT�ȓ82(�@ʜ����U�P�&��__�i���6���%Ŗ1�Ѕ�0Z�5��:�v�d�R�pRd�ȓaW�u�eCҔp�k'C��A�`̅�; ������v�,����d"�	�ȓM�$T�g��t�����-~lلȓDݨ̰1��3I�.��B�I9�I��-���5�&��!�r�Ԅ�C������!9yH�c?9�"U��Isv�c'I�k?�ԫ��eꝄȓư�V�O-`-�a�i��}��m�ȓN���˿a�tE�rd�7�Շȓl5��� �}�.�:�+ʻ<��!�ȓb^hd�CKA��ԥR�Y�B�&`��uw��y4�],�Z�B�耞&<݄ȓQ����hʱ.z���sQ�Մ�s+�9���i6t��>h�`��ȓZz�y8D��1r)*��v�Z�-��Y�ȓ �=�DY���7k��LŇȓt?�(v�J�Z�f�����$ �ćȓC���+��O ��q��$j6�q�ȓY�5��⍆\��u�da��`oXa��\�9��Xtf��+��A�������),]��򈕶Q�ȓ'
�����b����AY~���/�Z�Q�K\�^����	T��@�����(��z#x���v����:E��9�Š~Ĵ� �ܝg��ه�L�� �N
I��`�4�E�%��l�ȓvʒ�;�M�;l���s"�le��J�n�0���+E�������B���g�0� �H3E@>%��O3':@��S�? ��	�!j�t �F�O�^�� #a"O^�T+�$S�B�0��I�e6�R"O����iU�4���h���W�R\��"O6��ri�2��A r�9?�Ͱ!"On��TÜ79�č�K�Q+�d��"O$��a��A�����&&�z�"Od����EI+D�%b[/fm-��"OtX�JP������o��EZ�q�t"O,����_�]�p���+��_:�� "O���fU��\v�U�(%$)�"O�r�A!CD�ҧ�!���8�"O`K�@���Ʃ����H��@��"O�e���̭�2%�hҎۡ"O�8yp&��:���%8�z9��"O�=�FԖU�x�k��ɨ0�)y�"O|ȹf��7�|c �O��"<{4"O8�0���H,^�2a��*0�.� �"O�Cv�U�W�\�ꢌ�N�,��"OjةS�A�'r�	�L�Tr,=0�"O�4��n׉Z/Vq@a��ThD#�"OȨ�͇}lt,{��Ԗ�*��"O�!�d�%;f�P��F�E�p�R�"O�l�o�"7Dn-Q+Wv�d�b"O$�3����?l�� 
�2��,@�"O�K ���!�]Q�e�"Oi*c�Օ.�h,+� �$�ְ�u"Oh�it̙;x�����W���:"OH�U߽(�e��̊H#�hR"O���!�ɯA��ʳj�pn�q1"O�j ���Lz ��j���	�"O~鞴����" D�cG��h�!�Ęc��M+eK]�z� LHUn�%&�!��l�� �PW�� TgPk!�D�$��%*#� 0,��v%��c�!��/ ��I���4^�����e�>j�!�[�B(�mI��-<��3�U�Z�!�Dt#F8A�Q�+����b�q�!�	<��p{�-�8q,��0�@\!�FI
M��㝤|;��he�!*�O��=%>AKuF�/:]��Q��C /WN�V�%D����P%5|6EK�#�����8�f>D��b	L ���Z�z�F�g=D�HC���6�T�2��<]�"k:D�h�1*��F���YQ�Tv�	)D��>���铉n�r�X�-��6$��9d�C�I�#	(i�P�����I��	�~��C�ɒ}�y����-Taʘ�d�D;61�C�I�_�僢�T8��pz��ÙK0C�IH��S�$ŉ%$� ��C �<B�	6*�lq�ؙ5��10d�NLB䉍z�E��i�+C����H'F۔��hOQ>�z�&�9<��51 b�	k�Dl �$D����`�7���
���7~}�\�$D��ǂߗ9і�GU�V�萂�N/D�,��۵��WY�*
���Ms�<a��	X�v��Aѹ6��- �e�<�I��h�60z�Ew��[��e�<��GH�h�nl�R��w�4��HDa�<ч��{���:��W/c����'Q_�<��m:���Ma���e�<�㣜�:ߖ�!�m�N�R4����k�<����A!�� %�B0�IHG�Ne�<yQ�	N_��³/WR�(�P��^�<!��èR�����Ѝ$M
X�	�r�<� *=�0A�VOn���� ��9��"O))��	�7l`T�']2D�0@�w"O`US�m�7g�D��J��5�g"O�H+n/�LXx�P$�j�"On���)�=>�� qаBA"O"��J�0{R}�ǚ$!���pc"O���i��!�ؘ�`+
� Dq"O�`�E�E�c�HTk"I�,Z����"O��p5��17��21�9c&��w"O�T8#�ڞfo�(�"�TN���"O����Z��rF�*n6ͲR"Oj�pփM�������.�N�� "Oެ{�(f���]����(O(y@!�V@ʞУ�lHn�za��
J!�d·�&�#e
P��$�T(a!��M8&�
�tIe��q
��%����S����(�
\
�	����: G6�ȓ_��v�K=m~������Thri��<��X �;0�EA�/=VGBa���~ *A�_�h:ɨ뎵]��ȓ\��AQ-V��A�6��.sW
��ȓ[B2��NS<I*�0�]1&� ��Y���s�AW;Ty4���)��@�ȓtH���?R����g��\�=�ȓ}����FdT
0�"�:$��py�ʓ|b�7��(-X�fI6��C�I3S�Y�p��kS!�DF�,(g�C䉸A7~ �r��H�)ҤA��C�M��q�!O�j�@�O�_9�#>ɉ�iOW
jհ���iv�Ej��ѧr�!��5J�������O����Q��!�dĠ�D)	&*ѐ`X�xR��!���A��2��t7�$S"�-�!���X� K�a �8T�:��� M�!��P�D;fT�F�L�*��?�!�d�~���%�)a$��N���B�.ғʈOf%��'�kh,@�5�����h�"O�M�0aP9|�H[WBQ o��x��"O�M3"ț��N)�a٪�T�"O���+]�_�(��/P�@�J�P"O�ł�D�@X
D獑�
�l�B "O��B�R�`��Ƞ�/W���x"O�@�e"5���I��r�����"Ob��C�U.T���(�X��|ˢ"O�գdl�g@��q�C?��a8 "OJ��)^� Vr�t&��L���"OBMAB9�1�fG�4:ɛ�"O<����k�HX��
	>�� �"O�}�qT)����3�K;H�.܋�"O^ثeJT����I��mH�I��"O8]2�
��w�(�`�g_ e�x�"Op�[���0-x�+!Y#�l�W"Od4���hTL�F"ԣs��"O=��5��Y�#!�6mT�ܙg"Oд�-�9��@�e6�\�E"O���g�^g�Θ�3��'��c�"O,��SGW�.��6f�R�8�P"O�1�"E�=�l(�WB߀%��*c"OfuV ��(�ҭ '��,-Z�yD"O����*LT�qe�y78�"O�m�%0aNt�(4E� ���V"O�t��m�$��\CW��mX:�"OdA3&� 9cz���M�\�Z�`�"ONєo\�X0��;���"O� �9���d?���Ak|�p`�d"O:�c��КJzi�I7$�@���"O���E@��n@�Rȓ�?�έç"O`����Nx��J�G�!Yn��"O�1jtNH�+汱-�O��9b�"O.D�&�C�Sӈ<�CKC�0�"O��ST��?���e(F�Lw����"O���2D^9ou��-BYR��"O�E��N�^��DB�ǌXV�Hr"O���B̒,n	����+�X9�I�"O�9vHR�`��]Kp�-G1d�z"O A �X˞eS�ˊ@Gr��`"O���C[�0���HS*jǪp�"O�s`�_op�]�կ��*�Hж"O�dpT��wj���O�;H�0ö"O�� '�G:/6vT��H�Ka�1"O�d �m�
pe��YcD�w-,Y�e"O�U�m�h0�毑�rLpc"O~(��
�E��EOfD�cV"O:�Ib/�&Lh���6�]�L@ġ{v"O���~�x��M^��vl��"O�U{tn�j�6���T�$t��{�"O�D��h�M�H�z�E�9c��"O09"�EK&$��k7��c^��"O�Ew�i��qo=%*l�"O����ʂ,�@���_�R8�c"Ol��'��4:��t�Ի�`��7"O��	���Z��U�31���"O���d��"*�T�Fe-%P�Y�"O���#�+PN���dD~A�̨�"O.K1�R���s��pE�!��"O�]3�K½T(�`R⠂�~&L�;`"O���eV�t4��R�An�xQ"O�Q�b&N)r������'?�Ij4"O� 1��Q1$�VÙ
����a"O����;��q��3?M�$�7"O-����<�i�0Ԍ&'t�8#"O��P�iM�AM>-��lO�o�=�t"O�@9��]�n� x��)���$!�"OJ�C��8,�4*�`��=r'"O��A�S<N�I�JV�]��Yj�"O��(3�@�bj_�A�����"O�� FX�3��LR�Ȅ9SP8%��"O���R��m����p�*0G�H�"O�]�)Ţe�X���.0 �*�"OZ PD}��Aq@E� Ĩ�"O��ra�ʍ�(u�P�=x�Z'"O�H�5(�;7�4!�eIq���Rp"O���BX�Fv:��ѡՁ1���ˆ"O��Vh�>�.�!c�0�.�j�"O0����.(Ș$y�$K6&���"Oj`���&L{$�^�4�#q"O�d���`�Q�*��m�a"O`�"�%��I��o�-m��˗"O�,K��N��@2`a	?J�j̸$"O8���`Ꭴ��m�7m�&�x"On|{�է�X/�~~����"O�|ز��9J���QP����J*)�!�VX�ԉ"4�B�j�,�)&,�]�!�G�:�h���\˄��`j�>v�!�߀a�P�5n��T��-��FO7<.!�D�<R�P)Р�+�V���`
�*!!�d9(:Dd�D!�!`�!��yQ�qj i��Cv����GM�!�� .!t�*7<j�kGF�:����"O�x�aG�>;�j��C�?$b"O��)A�\6�B��a�9h�58�"O���s�M�/��bG`��5Or���"O�TJR��* ,#Q�;v��(h"OD�e,�g� ذ�0L�8@��"OޅxI�N�Ԍ�UfQe���p�"O�%!�/�r"�"��X��ЕAb"O\@b�Mϭc�~�(�`ٺ|<Ll3"OFE�M�}[蠸p���?8�P�$"O�qS�U�0LZp�K���"OL�Zƥ�,,N)(g�T���e#a"O \s�M�|(x���昗S�9$"O�0D_$$ʬ0!qd�~���{�"O��zb�ғ5��Q���@�*(�"O�<"F���'B���Weޚ
w�qj "O(���^�X��XG���G7ֹ�4"Ob����a�Na��O�Z��k�"O�@�B�M�4��ba��A�"O^Uх��RĔ�;s`ۥu^��"O��2���1\�e��mͫ��*E"OpI��o�q�P!�vC�>8��<ɀ"O����'�<�vH��!��V�s#"O����b�^���s  G�t���H�"O.�Q�L�{�}����l�l!"OL��B���a�Ơz%ό�U]0ؒ�"O� B,F�2hLh�[9@郇"O*�b��o(>�b��.e�� �E"OF�+P��7����S���7M���"O4U2�I�>f�$��6�"O8ģ�e�d��(I�1�L�0"O�8"��E�c5fL�q�'ZM�L��"O�qS*Z�X����� v2���"O�@U�?��c�y� Y�"O�:�Xa��th�烀[;��1P"O�dԈ�D�С��z�yJ�"O��NQL>N�+q�'\� ��"O��P-K�r�t��< � �iV"O�Hȑ�K3[�v��3`��8�"O`JA�M/Y�� �3OަYip3"O�0�1eS�`�j�s��_R쀔"O���
EZdEk�R/�:�"O����ށj[(�#�އE��s�"O��C�I�<6�FHVoE�]�L�"O�ٳQG�y~�TdLH�;;P�Rd"O��b��+%�n��Q�F�!6���""O��;��[���H�1+�$ &����"O�R3��r���0�R
"y!"O��!'��dB%x&a��l�Tyv"OW	vU��,Ƕ
��o�*c�!��^�/�}�b���K�+��O�!�d�U�v��b��S�"�3JʼF�!�ڍ\��D����
�z�Q�i�!�~I��NW��t��ӄ4�8;�'m�A��뛜+��1F�/���;�'O҉+�^<87`�a�P�J5��'���J�%P�����@��J�$x�'�&�X�$�U�nt�p�ƼU����'V�X�T�^-(�0���V��"�'|а: Dב!��hR�`�)[�ʑ��'�z���tN�}����P�9�'�v�9��A$�����B��1��'��{b��w2	[�DB-��@�'�6=�΋�^�đ	E�U�dթ��� �`�)J`�b�K��ΓH�r�	`"O����`�/*����]������"O. �nV�Z LUJ����P%��"O�D��)31��X��"��U=L�	�"O���D�Y
Z9t�T}Av�z�"O�d���"�����Daij�"Ou%�Ϲj�̩�@g2�Sv"O���D�m�<cs���0��`"OL!��`	Z4�X�k�GyH�S�"Om #Ņ7^�(�M[*����"O�}�H��:�l0�T�MyiS"O\�)�=�2(q+L:x����"O����\�F�mѠ��Qa�m0�"O�iw�L���Z`�ݓsxt{�"O%�s��g�Е�$㔀l�`��P"Ol�b��+i�وu�I6��uI�"O�dz���(-w���pF��C���;A"O !�uH�GR��{�e��^�0W"OĨ��j%SЄ����G�VP��"O�9�����Ȁ�;i�{�"OH�#��+.����K	^P,Z�"O����gI?5�z�ʡ(M4�b#�"O�%ٱjK16�(����?�8�0�"OZ���cZ5p��S +z�SS"OR�{`)���@��G�Hq.M��"O��0��5��=���нF\~]s"O:���C�5L��2�.�'
���"O̸CS�E+RJ�%r��Y#W�DR�"O�ݐ�
܁TE�@�^(D����"O��J��I���3���j�T<Y�"O������nY��$�P�'eD"O�]p�I�@7�̊��Z�@�@��"ONtq�n�|Ɲ�чX�
���"Oz ��ڵ<�8�hD�U�<�l�"O�Y�2k��B���p�ܬ*;
 HS"O�$�Bi�z�r �ץ�@8��*�"O¨B���1R���'�ʉ|��P��"O^QQ&�ܮy�z�vI܋�z���U��Y�KҤIQ�i�ǁҤ{����h,D�4��=��т
:Yˬ���F'D���d��5v���,Ŋyvt���i&D�<��c��H=�LX�ǔv�@�#�#D�`#��ܪ?������ ~�����>D��&F�G���׭#'1ig-:D����S���9TaH���pC�#5D����.K������m�ά�* D�l�%hD�R�0����7^���sN<D�����M�<�m�P��9D��8&͛7H:�QdYXH�`¥g;D��1�D� u>��B U�&O�<#�:D�H���WfV��MѥAtا�9D�LeiU1"�l����(_��E�j8D����Qx���'R%7���7�4D���a� W�9�$�PC���O3D�l�%m�#(3l��`a�n��@���$D��P�j�a���A@?:�p9e+8D��;�X��j8�p��&T�2����!D�Q*]�\����>����F:D�����k̴�q�5<{����C3D�d�ª��9 R�Y�c��)eb��F2D�x�D�6�^�KK<g���G�+D�����F�q䤑X�o�Y���1"<D�X�$k^�nc֡�f�$��"�;D���C,�̬ܲ�Ɲ���2��&D�� >P�%�O78���qG
�0���H�"Oj�K���+O���T'��R��U��"OD�KŐ�h���#�f�F�H���"OjPB6c�I�@CT�y�D�"O��)T�U4 ���
{�i;�"OFh��R�M(������؋E"O�����I4 jD4Ȃd[A��(B"OR�sFFU.y����unP%OZ937"Oq��Lߍe�(A�gĹR
����"O�� �(W# �
(�Q�JS��w"O�}�D�Ԩ
m2����O,9l�q"O<����[�$�4Pa祏6~��,�!��Ǎ6d@�U"�,m�)k�3�!��43����0Y1�P�C��&(�!򤌙.������r�D�(Q��!�d
>!�V,��#C	��	t�&`�!�$L6�"���HvL(�4�I�}�!�dMS/�����%���a�:!�$=j2phcv.�9��rc!�dK�������~�ly�A��(!�$�r����'卄g�ziaa�tX!�Һ~g �q#ʷI��<H���sU!�D]�u��9�b��#��щA���.)!�$@
|�F�R��ŤL����D W?!��ǵ8�B\�E�`n
�вυ6#!��[4�p3��u� �0�!�J�41%��/�5Ƀ�V�l�!�ɤl�T����Qhڞ`�F�U
�!����+�����Am�j�*�ńS�!�U3/�.0Q����f�{Tş#z!�ć�"�D�;D��c�>"��y�!�D������D�w���Ӎw�!�dQx"KαMZv]pO�b��9�'����qA�p��} �	;X���
�'��P`b��OWf}rǋȒT�E�	�'Ŋ���QZ���X���	�DX���'q$(�D*ۚLT�p�J��u��p��'��Wi�t�HH��o�3|��I�'�`̛EʄM���0� ��� �'�r���႗;�z��0L�}�>�(�'����؂lފe)�Cm�0Y��'M����M+.I^E��J�k�F�+�'�ڬpPf�(H��MC���`ܲ���'�f!y�c�Rna��=�HQ����x��E�l��w�DS�R0;�X4�y'K#Y���Q��5 �"�'�$�y���!���J����p�)���y�&����cj�4�{�!ϼ�y�M� 5���e3!��y��%$�8D�"��P�Չ^��y��)?B��Qjd���`�̀�y���0��٨�U[�2��vhP��y����B�KLH�Eg(�+_�>���r���F)L�2����b��-�@�ȓP\�<y��܍[�F��"��'H�����Zq�#� 9,Y��ژ���ȓ\��y�I�TAذHP�Ja��t�?�
�
Ĭ�*��RuZ����u�x�ȓ�6���V�JU�A����V��ȓ���&ìIq�ț����>D.T�ȓiHv�󵋊� �L�C�K�5�0Єȓn�`t���X�D-~��p��AB���P� H����*�c�Bs||�ȓt8��ba��U�^<���p֔��?���0<� J�*��7)[�x �f�w����"O��3�E��"99֦�2X��"O>�#&J�m8���4H��=��"OPA���5:�<\PA��:/�l��A"O$(�Q
�!�USMޣAb����"O��3�$ʙ
��;5�.̺"O88�R�~��Y0��ˑ8� ��"Oʩ�B�iz⅃G��X�Vٓ"O�=@��>�<R���@2"O��1���@��vN�X����"ON#��D"V�R��p�Vk�"O0����i�XBٔ=��eC�"OP��@��076bP"��%"�f�D"O�Z⊘O90���)ɉ���"O*�E�^J� �H]�|<j�iG"O� Ab��������?R:�5!P"O`���S�&�t�L8���²"O��ӂbΔTT�5����/
y�"Or�`Ԏ�1r��	��K��4��f"O��fo���N���%b"OR��tI��@`F�����,W|y[�U�DE{���K>���k��,�QŊ�J�!�L \���2���,E��#��C7p�!�D�N��C¤Jm�5�SC���!�dC@,���e� ������i�!�$(u�ЌYRᆏ~�ȉ���,KX!�$MGJF���I�1a�P9B$�C�DF!�D�o���\3�6m(s���.!�䂘6����U�G4�pT�Qş�)�!���om�9x�-�����#�7>Z!�dY6 Z��7瘮-��� �� L(!���0F��d0�	�^��ɗAU�w!��Y�!2��P�0��`6@!�䏠
��H��[��(j�E�D�!�$َ~8��dI�0J5�TI��!���O">����T�|j��F(n�!�$ <Z�lo�? t��!c�I!�d9g����!N�)��u�h�T�!�$�<D�<<X��	U��q�AGR��!�d���R��` ��c�� �׈ٍl�!��Y x4&� �c�;�GH�^!���Mh���1�L�q!B=�6G��!�
�'��{���psd���2y!�dA�u���yW͖/�7D��7r!�d� f�@2��'���Q#{;!���w[ i:b���2�h�����Q+!�ā-fn-�4NW����i��T"!�0h�����[�ā�Hʺ
!�D�$)_L 4Nِ��aJW��%Grў$���0�u��̪ )-��`," �B�&>���XT.Ƈ~Ԫ��Ԁ���B�I
 "�X�E�k���A����C�	=T��d�Y�������=a�B�I�j�tl�0�0/�j�b�A8��C�	�_o<�a���.`��B#d�fB�I:����%��P ��MAf�B䉪G">1���9$��睰E��B�	�6�&�`���
a���؜!	�C�	�V�F�(�(j�����\)X�~��	�'��U��L��Gr	QbPy����'�L��Z��$U�Ț08-v��'�詹�%�9�h��_0�hZ�'��,�O�)mŌ��� Ձ������)�tI��a��b҉ǚ5��x�%���y
� 0�� ZR��;�i��� "OJ�y&���h �ڬU����q�'y�'��)�'���T�U�[�`+��ιk60�x�'��kG�6�0i�Ӎ^�e6\m�	�'��@)&*Z.��R���_��(�'M�mxP��S�����:S1a �'=�A����0]�F�%P�DµJ�'�j,"c�v�,+�C%=�P, �'�:�4�&!c���,1F@;�B�)���5��m���ܬ_(��k�@X�yҥ_*{x�����=W㞔#�C
�y��T�̸�/
�Țy;����y��\gZ�(V���P\ѳ��_9�yR�
X<�q�5�9;Kx�i��C3�y���'2��	 �2-5"�K�����ybO�4�|͈�O�'�8sd�_�y�ɑ8�y��A�u,��0gީ�yZ����H׼k��0�DۉsV�)��'��	P�D5$^�H���̈@��H�'�\�K�#�4k��Hd����O���!A�5>�"Ă�._ġ)�"O~�ƣ�?h=2r���<r�D��q"O2���E-|c4���s��"T4!�J�����CS�(ȧ�W:!��)D?P��F�����t,�+U|!򄊁o�pJ�ԪdtJ�v�> o!�D�({e��1!Öj��p��,t_!�������
�^X2h��.�!�Ğ�IpP(r�k^�\��1t擦s!�Nz|Y���T��p�A�R0	!򤚩':�;7%G=����V@� �R�'3��'O�0�@�Gn<b<I��� �m;�'� 1���A���p�Q&q�]3�'�Z<��Mĭ}�5�qfAfi��'��T/��.gx ����+Q�X��'2��*Au�+�A	0Y
�E��'PR �pއM�>� F��e�~�*
�'�,h��]�l�����F�K� ݐ���xB�2ĜM�&$�%)�q��yr�� 8��D��ɘ�&g�հ���yR� T�J��f
��ӈ�
�hO ���JW�ՔN�D��ĖJ ���"O�	(��4�b����
�#�Z�c�"O( Y2!�0��is�K 4�%
&"O2xp�OHg,�Q ��z�����'�2�'`a|���)A@�1H[�'O܀�7���y��G0|�����jM<A���,�yBb�{A2�ӣ���R�v�[�$<�y��Ȕ���pW���G���J�����y�ˋ�W���K%.B8n���È�&�y�
�! <@PBl0o�"�nל��>��OƜ�p!6I'΍�$��+���bd"O�!'L�2)X�x�%~rJ2"O�I�0b��-[��uL�J��"O2m�w@�!=�aaD�_��1��"O�J4�I
'�t5�@���b4���"O�ഥ�O�(��pL�,Q��"O9j6�V�#�B��i�kBU�"O"�R�O�' �	���iL��"OP�B��i�4�:a�	9LU:R"O��T��;R!h(�LZ.LH��E"O��s��A���AQEۖjD���"Oj��PN�1�2D�B$++<r'"O����7Fx�E�N�)Y�u3�"O� ��Y6N�'^*4��G�-2K���"O&(��=I��E`��[� a���"ON� j�Z����Ƈ+DP��"Oz�Fۧ��XK�Y]��ku"OX}	S��5_�P����ф0KP-jqO�4��-��bB}��3+s\��t� D�����1S��&	F�6�AYщ?D� )��.V����ĭ�UQ��=D�P���{�����ï*L�����7D�ܡ��[�F���qc.��*nx4���1D� �Q���t��,��I(MI�(�$+D�� e֛H9��Z�G�'���yC*D���S��(���A��EF���5D�A7J�<cBX��jV�Z6Ĺ⧠3D��"�ڊ.��4d&�{�%3��/D��A�+�k,	���S	m2���gA�O<B�Ɇ8R��ʆ�MSy6�8@LvtB��C ���T'&�p���Rm�C�I��>�P�dC_��a�K��eo�C��(f #�X��� J�
�m�nC䉘��l�'���r����$�LC䉺I���j �S�~@�����'�6C�	8 �dh(5�׊h��	3)B�O�FB��36�<c�.�,Gy(#,@.e;B�Ij0�t@�A�X�q����= ��C�Ɉ(7�����0N�Ƹr�o��C�I��P��ћN�J9ѿR7�ʓ�0?���8��e��Ɗ,��0I�W�<�p���|�1/�<�쪵��R�<�� ��'���5O�0�4���e�<!�k!|R`{!�����!��e�<iS���dP��X'%ތQ�|A���b�<�fF�*4�{C`̡VG��s)�J�<qq�߳?�*��`�ɡq�0���n�<Y��ǿwm�-	���o��f��q�<���'$h�� �6b��6e�j�<A�MX�4���R4E]#��p���e�<��O\V��Y!D*�D鸙�c�<	���
�b ���	[�lEB�Bd�<!���^6����n^��xi��\c����<�W%�/��DK�C�+�8=&+�s�<)�l�,8���dA
�!,y�<IRKZ�;sҝ��.ڡ?mF�c7(q�<1!�3z)�g��Ha�){DdXa�<��W�DUP0��[0:4�!Ǆu�<S[���Po*?C>�۶�p�<����,Q���M��5Q�\{�GEB�<3�BT��ɡW�Wq�Jẵf�v�'��x2!ӷ���g"A�@���a�w�<��HZ9=�0���*/�Z�Gn�<!s�ƧR�v,ԯ�~��Q���c���?YÓcƁ+��\-l�8X����j��<��^$�T�	�/l�;��i2F�ȓ2�tp'�>���҇�0sw$���#����!?R�$��eF�=֩E{��'��f%0�\���\6(�<�r	�'� 8`@�G�WYF���H�7w�����?9�����+NejJ$oX�Uv�� �F���(�d#���(�8,Z��H*	�<�!!D��إ, )hP�4i��{��9�0�?D���@fT-J>XiB��8o��Q��B8D���E��'zt"�y��;8;>��fn5�O�bb��VgO�U��'`ӿI,̇�VĪ�΋��x8��d�b��S�? .��K%|�,��s�)M��t���@�����p�X�
�Y��Pk#,*D�T��b_�e&�b�m˻��,@b,)D����l�45Ff!K��)���I%D�L���ѻl<n�ɵL�.^��bG$D�D�dG��N�f=���[z��aP6D��p���:}�ͺ���
E���2D��hg���J-����a��yNu�A%D�r��.��`˰,��c<YZt�-D��N�A��f���h��DF+D����L��O3������g�sFJ(D� ��M0\ю�$Ë/$t�Q�d-%D�Ļp�( ��%�w��}�Ht�M=D�x�f`���7��,J~d��F<D��zl�3{t}c�*�� ��bE0D�� �(J�o<� ���ɳ�A3D��Au&�'.��І�DW�t��/D�@�#��,h":]��۸�J:ړ�0|����,쬬���#Uh�����E��d�|'/�W��]9W��hpr�,6D�0AW�	�Y�A��# m`�G�2D�hۄ�]84@��쐳X3�8i��<D�Ԋ�A^�n��H�6}��� &'=D�|��."�p�BS�N�g���Cf8D�\SvȓE;�
Ё�2��݁��6D����y J���K� d�5��4�*�O��BD�˯>5JP�
�+ݰ���"O���#A#N����Z�r�<�T"O���r��;^L�W�R�n���S�"O��(Äd�dM��@��@xi�"O`�`A�%~��%3`�^#:y:��$"O�A��KQ���Pi��ᢀ��yB�׆�P��6�ӅA��m����y�F;�ݳT%[9A�fh� I��y�c���t�C� �9	�x�,��y2��2��]��&@�.��8�$(�$��'�azRM��v�d�&ϐ�sҕѱ�S�y��ɻ��������?mX�؇�y�b�9GXٰ�̾3�� �`X��y"�Ԇ'v���� *�("0C�yR@ ��Ѫ�BҖKcRYK�N��y��ߋ$�ZIk�bKCo�L�fW+�y�&��O4I"��VA�`R��[>�hO����^SFP�Fm�9._�M�L6N)!��KL㲀���\Q��c�B�"!��:F"n�A�!˷Iz�r�ʈ�1W!��۶nl���C�W�%9\E��)22�!򄒝g� I��F13��!���2�!�2S�(m�v�,w�@����J}!�
�(,NزF��5>�{��I�$Z!�$
h��P{qDƲ@8�V��BE!�$фF$�<�4��4�b�8�e��!�D
�6�>-��kG�|n�x��D/!���"��Kѥ��p^ؤڱ�{d!򤎯7�.���UgMbAۓ�$K!�L�S�:�x�eZ�IA^hbNȡ�!��#%��ze�Դ}.d!��{�!��=��*V�:l�����aP!�7zp���$h�UK:���@��e�!�d���:@��-:,��� ���D�Q���ȋ-Nл�D*K_�C�	8��$��h�l�Q��G�k@�C�vBL�2D��U�d���0�|C�I�j�{���,�T�B�=�LC�)� �X	�"�4(���%F��y�^,��"O��B���7������	x���g"O^袆��p�Z�yd A� ����R"O����n�	\���2��]:e����	a�Ot��+Ư�0@���GI�5���#�'�|�Y�H)c&x9�5h1�����'`���J�(C"����V-b8���'�Z�HQ�F)`��#H�s��@�'��I�p��
���#
f�]0	�'��Ȱl��>��s���e ��"
�'n�݈�F����P�s$�+j,A���D;�A����ף��hS"..H�ȓ[���xa�@�+�䕘.<B4�ȓP(0;���
��$ҋ�<���E{B�'G����VP��rRc��~ �
�'�f|
�(��Q�I�J16%D�h��E
f��5��V�r��i�g�?D��"�$�c|F4Xs�V	'�� YE	?D��KQ�Ľ6=}�F�����(aH:D��1�O��0�Hic�ϖ`|��(�j2D�����0Ytk��
��,��B$D�0��!_�Z�j1@O�Y�lÔe4D�Xc�Dt�Br"	�
%VD�ׯ>D��y��!*g\�b�f�cYX��(D��ᅃ�/�8XFh\;n͞��O��=E���O#6����Rը5�t_-M�!�dK�-�Ҥ��X&W�:����k�!�䈿c�t���DV����S�e�!�d�GMz=$�$�������!��_�;ˌ8�2g��o�6��FL�i�!�A�Z��m��0�� �.e�!�G7|�p!	2�ș*%�Mh� �%U��O�1�A�R僰.7N����"O��[���*&jȑ�N�)F~dq��"O�(�&ʐ�"2`�A�t���f"O�!�pG��V@@����[z4	�"O��J+=4!m�mX�@U�y��"O҃C�@�v���l˕Hk
q�B"O��듆zʌ�Fօ1,��cW"OzL�0�V��l��ώ�l�;v"O�!s�,��p��I��$�~�sF"OfРâG8ms���Q�4@�>�hF�|b�'���KX
�|PN9El��
�'?��+��־Bf�e!R=AV�	
�'^��[!H�z}��5��5�~u�	�']��B�	�<�b�+W�����x"�օT�q3֢�*J�����B��Py��ˏO�`RЋС3L`J�+�XyY�PG{J?}s�$�?Eȁk�� w���5D�(+b �& s�;�٫4ɞT�w�5D��(�Ǒ8U�r�F	�X�TLI��'D���h�7T��q����~�,0�Ul+D��j�a��?�f̈p�%���;�K'D�+�L�0�L���+��/�V}�t$�O��O|�=)�O�A����Q����RI��qx̻0�|�h̓@q.�y�(ëZ��$t��,g��'�Ą��l��%r�%G�RN����D�hC�	�XI.����7p�:|	�O�5G�JC�	Ol�Ix��˜:ԑ�&Ƞ[LFC�ɢ~�N�6I۞;�@D:fˀ�b�6C��&s��5�P�ΊT>*#@�2��%D�<�q�o�1����v`"�0CL1D�$�	�9&\4�cȞ[FH�P�4D������kx�E��^1|�6Eqs�=D�� :�����R��ag`гu�\%�e"Odpr	W,P�$����Ѥ�*`�r"O��3�!m�@�zE��2��s�D5LO�` � ���l�q��7I���H�"O�(R�ʻ<ݚx���Q��Ts�"O�S��/b�ma���r9�$"O��X!hkt��#.ʈ*��I��"Ob�$mǅZ�z�����'K�<h�"O�u�E�C.㮀Ȧ��1�]�$"OL��A  ��B�"X��q�"O` ѐG/n��%��Ѣ&"O.��@\ D�������1|nB`"O�D�a�	��٣��'��F"O2���B[�,v�l�-��!�.ez�"O֐8�.�k�Ԛ��Z;^���K"O�	�c�	\�гpJ]2T�lm��"O�"BW�U�	B@�Jm��˃"O^�XU�}���� [����'��sl� _f�����	>���kr�8��0|b�Me���!(�e�J���l�<12�n��W"�ܡ�E�H����~&l�k�o�=	�����Y='��хȓ\��	u���ht�;�)���ن��I~(R�\|C@#ϼB}�%���J�hO���DRmb�R+�FKܨ�d
�!�DЪfUXܪ���l1J��t����O^�����\Y6M����y���@d"O��nۣ;�2�����^ոIY�"O�Q��C�  @��#)V�:=�"O�@��̖�����""��dT��3"O
lҴ&��Q�ݑ Lu�XaP�|�)��3��=��B��`���:��D�C�		�>�iFM?"��l��B�&�P��I���d�w�ih��A{�<2"O̰��W�0|h�!g�?c\�q�6"O)Ä�/G�8Yh ��=MZP�""OԀ�A���X*��� �Òv��,�0"O�Qa眽\���d�KBa�v"O����k���Q��J�^����"O�a�o��Qc�����|����"OX�'�ɠp��}a�BY�����"OFd�a�X�lR�8i�>	�Ty�"O�t�%`�9yF��ubD�5��YB"O�k &l@l ��9��1"OjI�4��N}�<�
�xF%��"O�q�d	��^[�hɅ�E�Ѐ�@"O��m�5y� "f6R��P�u"O���g��n�5�6�ņq�V�q�"Op4#�KE���t�0e%Jt}�c"O�0��C��2lI���V�nxp""O$��G��Lw��s�L�r'"�9�"Opt��R�`�~���:)p���"Ol�y�EV7��a�D`^�
���"O|h�ė�=��ЉF�^�V(����'�1O�Z`�Z�\^�( R�Z��Jc"O~*�8~:���P�,�� ��"O��;��G�0�����cHp���a�"Ox,��F�>bB^���������"O�<���`6���<A���je"O y�E�Ҡ
0I�FI����0�s�'p�|!C�bvbYi0lP�H�~z��O��=���	� ,h��R?��3�8b5�	m��Q�H�N��U�O��v��K&D� A2�?z�tQ��̓R}��ʁ�%D��  5!%�"`2T��1��#@"౺5"O��bE�б;zy
s"ȴ]*4̛�"O� B��@�Zʡ Z��j1�'��58#��S��H0ܮl���_�ͦB�ɐs����A0]Լ��f��V3�C�ɝK�`�Z�"q5���%�2-/�C�I�Vx�@I�e�;񶈺�	�%znC�ɁV*�ct��%�d�V��#�8C�I��|d��&]��JQ��,��B� "������4��e0D���#����<1�O9#`(ͻ8-᠃M�"(!��+P"O�䉷g�8C�a�T��z�p"O\�a� c|�TZ���/�@i`v"O	`�C t(.�;�,��}}�E��"O���fDӱtN�m3��J�.Nf"On4��]O�d)�+O�zƜ@��"O�U��RsÈhhB���2�	n>a)��+p��a��/&=F����)D�TcP'[
ʘ�g��%`.<u���*D��zm
�6p�����}��B�-D��`��ݡK*A���L��$���)D��	�'E�r?d����f��RG'D����n�y=L���g�6<�V����#D� ��8T(D�Ҍ�I]>4ʴ��O��=�O��I��񊓈'%ѩ!�ɊK���#�Q�<&�>C�ܐ$�ל�
D`�Dy��'?�Ĩ��$^��H"`̊A��9�'�B���7P��b����J���'��;&nL�b6�I�!I�z���'��1���ͿQr�i2D�u�d�H	�'t� ���%2��Tؓ�\.X�>���'T����}.��)cȣ~�2x�'(C4���@Iڵ�ǰv?L�s��?y	�M���+��P����w( �
�1�ȓdF)`�ƞ�%����GC�p=��n&�� 0g���ų!e�Y��Ň��"�ۥ��*����1�QK�x=��5���Z�'�72�c\�}���'�ў�|Z����H@��P9������L�<�dm�siF\�!�S8r�n�  �\�<�R-��M����4m2����HM�<)񍅥RL�}I�/O�1�J ���a�<���3~�$[p����	�,Pt�<%�H,Y�C@�/\�P��p�<y�n��J_:�1փ�%C�6��#Cf�<1C�o�f����5',�pӂPj�<Q��L�{��Xjd�˝�©[ �e�<Yw˖)<6d���G�i����b�<i`-X�P�bs�Ēv1X�a�Ly�<�B"A �<��eL�S
,�`��v�<�A� �f~�B�l
�{Z28$.�q�<i�a�)�8�"��z[�b���v�<�B��|�X����sa�XcE�}�<&jɥ,M��!��#is�r&{�<9�mA����CE픫E����HM�<9tlP�Y�"�h.�+:"�mQ�k�J�<�U�
��(��͂�"J�,���F�<��m�G�|����Xo1b܀SWK�<Q4E�Pd"�q�n8��H�<����-k��s-�o|�⅙C�<ٲ��i ����a���$�XB�<��K�8'�h�
��j���z�<�u�G�ܨ�n�@|L�Jq�x�<i�ِ_���s�CY�4�@�
�r�<� p%bՏ�y�����!D9�#"O�ڷ�� &k���`N��6rp"O����AX%����%`b0x3�"O�#��ΐ�<L;eoO�/�FcR"O�q���@	%)��"I
8T��A"O�u�W�д34X=x�m�U"O�ͱ�,�T`@�R7A���59t"O�9�r��lrр��̭
@ଊ�"OX�j��R�s�@��E��"�*�ҁ"O,=fgB��B�= ��(S�"O�pÚ�Lej����I�0�aI@"O�mB�l$ yZDlڴޖ%�d"O( SC)ܶ&H�a��!X�%��dJB"O�0;�*�^4a��Wr�����"O(]�$�[g��ч�L���g"O ���f��x�ΤK$��[�^)8F"O�P��̟�rʜ�ᆎ$s�",��"Ov�)�+����R��`�z�$"O��K�!ԇCC&0�P-"���"O�{tC�'z/�2�WF/x�2"O��1Tg Y4���g7t'*��V"O�0:!�\� ~p�+6�k�آ�"O|�$�{��p�g�#i`��"O^���� �z���Y��-�S"O�	@<X�8(2��%)��S"O�e�E���u��_���{�"OhyB�X���9��80�)�"Od��JؖB������%�T�T"O����A' "}�ӄ�K �K�"O(��R�,�#�
\+�"OA�"х^p�#D�&���!"Ox��)U'U;�-��ZE�i�"O�y�5 Z�vǎ�q��1����"OHe�攂[�C�`�>�@T�"O���ډl�
T0`��Drbɲ"O �BA��~��$�e�T�x::s"O�k��݊ ��:D��'�65�E"OlMY���8Gf�j[	e��a[�"O�� #�V��4��h��V��x��"Od���!�r�d̃��Zf��|!e"O�"3EO AT��gݳO�I��"Oz��Gȝk�T��"G0`%�u�"OFe)Z�t���� ��� �'�Q�!�L>2(~�:���$P����w�U6v:!�>
̭z��R����W���|!��Gt N�pvKP28������n�!�d�) w�`DoE�	ۘ�!-�Q>!�D�j"D	�W�]4g�U0�5#N!�dY]�,5��b#[��R��m8!�䖫ksj\jTiK�n-��,A"!�dS�{��9�Pg��Lz�D��$K�!�d1���q$J�!�r��M Z�!�DD���6,CU�n�+V+ �!�d�{K�HS�(����L�����bt!򤄁l��9��Õ
MVG���pe!�$^Ȣ�hV�Ϯ H|�� ��\C!�dB�E1ʀi���iGԘro	'4!���
�2aDa�308���[-!�Dl��zQ��pM�$�6I� !�D��܀q��DE޵��H��M!���5����e�O0Hm�!i!��z�A֜NT�-��"ܝ!R���"O��c�+�! J`/��m��"Ov�q��8F�ݳ�$��G��ʁ"O� �i9��Y@��2�:�Ʃ��"O�%
�#�CeO��F���"O��%��7�B}ѕ���?���"O����j]$&G�XxJ�����e"O|!P����x4(�
#���U� ��"O��%.�-0���R�(>a��0�"O��u�T9t����7,U�Yt��Q"O �s1�̒;�L@6"łw�d8�A"O��2��:f���76m�Ȃ"Os�'մ>zNL1���N!�5%,@|b`�H��ؘ�ԭ�=!�B}"@�qn\���Kg�I�(�!�䕒D�H�+#���%I`ˠ�!�$�N�����Ŵm�ޱ�׃��!�'�L�*���d���¨�`�<�T8(�(YSƠ2\�W��v�<A�M�k ���!o_��Ţ�Z�<y�I���m��3`��j�fPW�<Q�� �a5����I�u����e�S�<��Ōd7&���͖�l�0psaK�<�⭌�f�-z&�_�+���`��G{�<�d�@�6`9˲*\�0l���m�<�QcA�k�dyQ5g���s��h�<Qv�ҭ3N�	��N�E���b-�j�<��)έ�(�i��P�s�l9�P��h�<��1@/��y��2�N�����]�<i�.�)���x���q�  XB�E�<	 (R�-�욒ǎG��x���u�<�֭�O��t���	�+d�A�D�Mt�<9���*[���Xg��T�q'�p�<9gdB=��� Ŧ�C>X��k�<���o�v4YE�gk��J��f�<I�k�<X.�)X`铈t̺�h�cTd�<)#�љ:r!tm	����ed�<�7�����Z�8�t��U�G�Fk!��$}�N-H�	�5(|��@꙼%j!��j|��(W�@p���J2$i!�$ѓZ�҉��e͑W�kI�4ic���vz��� pv]��Ĉ�y��ܜ{7�A�1)��f�J�uΘ��y2�،�쑻%�3ZÈ��
�y�l�$4h�*�L� ������y��K0" ���E��Dyr��tD�)�yB��'}��(P��Gf9��H;�ybIJ�vI���5n�B4 ec��Y��yB�Р�����mS2@Z`�K��@��y�N/6ǎ�@�B�2@�D�b��y�D��xjr��X�.h6�hR�E=�Py"N��>��Jd���o6m�)�|�<�0	�&HY`M%J��Tc�HR�<���S��,�DZ�!%�ȩ�#�v�<�@�I�[��( ��7^���yB�]�<9�Ѽ~��"�߯���q��]�<��X��4m���]p��Р�A�<I��B�cxDaD"�Q��d�f��c�<�r%�$8h>�h��@.)ҬZk�<��a�"o�6-���#�b���ɚj�<!D���!2@Ջ�G�\XJ�����~�<��!Ԡ5�u���4z��|
֬�e�<�qdQ,��S�'1(�f�k�,MG�<�E/��VW��qХ�MVPz2�QX�<�V�B��)�6��
}�����&�z�<��]�r�lX31)��H��e��p�<9�ӗK��<��	?g�j)	�M�c�<� �*G�G���2�-_5-n��U"Oƥ�T�\�a`N�e�Ͳ(����"O�a���M�g���#曬X�0�"O�U��a��Hu%E7MG��3�"O�|��i]+\�z������� NRe�<a�(ʰ,����$h�{�&�a�<��k˺_���1"d$j��x�<iFo��4��x"��x����At�<��$ܴX2TtB��<��E�<��!5��]�m�����ƌ[�<�b!B�Ø�у��g�x����[�<�A�_:r.���aL����a�U�<�u`��M���/��+�!����f�<�3*\�+�v��פ�D�2�h��a�<!R�5W�%�7"��񞄐�E�F�<�CN�5+���z���C�D,���|�<Yq�|C6�i���@�ě��^�<a�g)an)3�ɑe`l��-�]�<��G��v��-J�m5g�,!��EC[�<�0^�t����o��P���p�<��a�J�Υ؁�DǮ���KCE�<Qg�q��	G�O�x;p��@�<	g,�6��K�ۦ:�2c�}X�o~}�O��\���P�		J��aխġ�yR�¡2a��j1av	ZE���rf�	G{��O����S�F{b���.��=�9��'gFH��"���c�ǜ�];$�'�6��W�`bQ(���PS��c�'�hqq��"P�D�vi��I����'pd�2��8W�0��V��8�'w�l²��N�y�ea[���'�����UW��jU�Ֆ|^�qy�y"�)�S��p`�2�љ ]�G\	.�C䉑l��Ѧ�L�����>l�#<�ϓba��ID�Ņ&,�������� �D ��ϓ1k��@gݖ��\�ȓ,������
��H�`�˞e�ȓG��q��B/:l�P��m[�f��чȓ=�^X!s�Ζ{���{"dU�jr༇ȓ[�6���l^>T��W�1y�ŅȓN�vu*t�7�x�3�M# T���s<���.M�5��!�t	Cs�6���)�t��NH,����I�0����%i8��SU��ʼ+ L��k�a�ȓ,9 ��@&�{���T�l�ȓ�jP�fРB���U���[~���ȓr?BY�aE�(;t1p���� Y�ȓn�rJ�����0p ���y`�����L�����ŨI:�y����B������b�<�p� �>�k��;+�DrW�BW�<a��׋����D�=,8,�R+O�<Q�l��R�*�c���?\��<��C�<Q�"�0! �;s��=�&��oR{�<I�-�� �P@y��Bf��p���=Q3�	 �Z��Aa��;�AG�<)aH�
 Ѭy�`=��ȃR��By�'_ uC6�Ӂ>;vL��C&͖T��O���ǔ&֘d��NN	8D���n =�axbP�X�>��%\�$1	�,�� ��m�4�_j��0}��"�'��,:�k΁4ul�s���5=h���ē�4T���04\��R��݄U�LP0U)IQH<�'M@���r�aH�6^E5,��<A��4�>1�>��G��4\4C���`�Hԁ�.�?��x� q� s֪
&Hx*���:}���_�� :�T���f��d.ѽD�vT{7"O��bL�6b��Da��9�Q�A"OH��!㗸Q����-����g"O�E!�j��R�ѓg�ѭ2��� &0Oz���
�=�Y4�3 �6�S�fB�	L.$ᡡ$]�w��	&��V�C�IY������*-���Y�A��	T�@���.�m�ԍp���`"��#��bH<ф K� �BX�`ҶX5|�8rI�'=N���<��M���s��d]biڀ��"]@���	Dyr:O�7�:o JU)�@4]\�σ��c�<�dAH�f�x���Q�6�[��t�'Y�?�j�ɒ �����|ږ	�D�6D��c#�'	6a�����H��%5<O�#<I�k�.�"�1���%�n٫0)[}�<	a��qgFq��	�pH¦A}�<�b&�Uǲ�1���K��)�f_v���'g��^��F
�����``׵vwB�b�84�4Qf��;3��0��ܜ9޼�u�:�	�<��}Zw(�	Z�!�o�+*|ءA@�4[�rC�	!jk�	ݻ1�U�t�� )sr#<�A�Uy2�I�ʌ���:H�(9)ы���y��KX��S$��Bx��@�)��dB�	�9D�L��iۂ��C߳�B�ɬGЪ��`�W>9������*�6B�	�n-r�[�f<0�����L��}}*B�ɴZ�@�c�Vl�x�(d��~T�B�ox���xw4h��`,���d�<ѰA�e�b��ՠӉR�V4b1`R�<�����NϾ�bGÂq����CO�'z�E�tO�%��EY׏��F�|��.G���<���K�Zֺ�;D��v��֤�%[�TF{���'oM��*=Y�X�hB�+���N��xp�6�S�'}�TR��`od|��ĻDn����?)E�2O���c�03<�#P+	nܓ�ў�OeY!�"�VL�S�>;�0���
O�p  �L�-Z%#�G�	��y"I�9H��@�cK��4X�vF7�y��"`����L ve�8�š�%�ybJ��A7�����i�2ȡ����y2���f���e�|�c���ymT?*þ|x�n��Vζ�S5)���'nў� q� C��SL�����քC�D�2"O,��p�L).��10Zx�����O����!��\B��E5Mw���ԡ��!�G(x����e�����PCC�<�̃��)����2Z`�����L�D�"p�C'D�`s磋�Ip�Q�
��<�yBf��t���ZxνC�h�^8��*�+ݼA�pM̓�hO��+���vE���bK34p.!Ȗ�P��C�I�(�a5m�O�<���g��q��C��<c�*x'kS�o:���bZ���C�I�b��;Vf�nCũF(٣b@�����1,O$�y@n��w[�a�S�S3be҇�	K�����s�!w`@�9�"���U!���v� 4�R�o��P�s-	����,�O�Z����CF�s�F �%,�={FOh��+��w���LQ�Х��� q��ć'Ӓp1(����P˝��yBl�(�	�.M�.�
D�w�%�y�B�GFU9�(=z�q(G�^���O�~2���D��,qB��>:8V��l�<1ŋQ�;Jv�BNRG�iy�-Bj}��)ҧ�u9uI	�"	��bT�q�����S�? ����"\$2�,�"S���7L��"O�DI�	�&8�K�㋝a�ld�s"OjX��A�bR�@r�A�w��j%"OT����T\�#Ce��J�!e"O���Q��Oa�8��D�/U���&"O<e��C�M�@���J�3-:#D6O��=E�$�D ,Z��	\�v`� ���y�fJ�����Ҋh]���S��?�J�0�O���8�t�@�˄���Bp�Ș_ ��ȓP���� �ɚ�JVmX!�ȓvǈ��OU'Z���t(���ȓsƦ9��هn�ld�Y�Dk��ȓZn^��"=��u�0�P�Z�p�ȓrM����Ԍ*���)��c"4�ȓg��@�Ht�8�V�0:�.Ԅȓp��8�����mb���|�ȓ�x�IBJ��P��hB� �&b�V��$êI� 'd^��� 9���:(d84����-2�-4>��ȓq��K�$"ΠL�	�1���ȓ���2w���9����Tgt��f�����j'�آ�2ߌ,��,y8��FZX�Q�w�[19q����ox�C���mœ�O+*M�Y�ȓ
�0��N?`<s�D_�P3��ȓZ|i4c�v�@�������tUP�����Ւ=���Y&6y��SN�6	�_8�x�%i�{+j݅ȓ`��)b�˂?�J��f^�T�L4��$�@}xg/�\�`�Yv�\�:0��ȓX�m��,ro܁!���2#r���ȓF�����f�ƌCE�(Vf(Y�ȓe��A�K[��$�C�.`!�ȓ�A�c��J��rS����B��ȓ",�Db�Ɩ7E ����H�7Fa��{2DA��ϛ4K@��G�Y")�-��;9^A[��>G��à��V���ȓdVn�	�n�$ �$�V�R�8ܜ��6'�2�#�u����W��.C�d��0�����1p���GK*_,�ȓsP�g�+|�)�<�du�ȓ�؅��s紴����$�P<��=�6M�� �3 r�1�v�Q��by�ȓ"訛 R�	X��!��ߪHB�bO9�>	����A.���&晉$#`�����=
rB�ɂGX=��h�	Nv��+P���X��C䉉"�]�bƒ75$�]s�&�#I%FC�ɔO
m�Q�:�="���.C�I"?<9J2/����s�BcC�I<��0 ��"Y%�(*V�.��B�I#,����ѭA��({��NhC�I�SxfU���(.:p,9�!�ZilC�I?PniB�� �4P1Æ[�B�+,���6A�F
���ebbB��:`s����]F��q��'^�st�C��>cQ��ӕ�{~�QpL�
פB�	"����D cp�����0 ��B�	�G
N���딨��%2�A��5�B�I4]�P J=F���àL	�`��B䉝�\Q��7,�(�KڊhNC��� �`wC��c�tX0O�n�XC�	!�f�0�B~�����A���C�(ސ�!JQ�9�xp�@�Л�C䉑o�PEq���g�L��eBحvLB�)� x���E߆r"��B�d����"Ov�rU(ckv�����k�i�R"OFYzTM"(;v��3�(j���@"O(6I�/d�n��G�R Fc-D� H��R�p�ڄ+�(}�:��4D�d3�C<���G���/U��fn0D�
���i�ʌ�aM!ZH�ҁH5D�0�^�@�ӏφ�<���C>�2C䉡mD��G��0oJ��� U�.��C�	�g�qs��\h]�$9��Y�̈C��iL�p��lp�*�3����z�jC�	�t�qs�L�V8�ۑ�> C䉆?5iw�	9_�ᲂ�ɸE�C�I�=���b���(c���ڤ��/k�B��H�E�rC�Ѥ+��{j�C��"D��"5�ϓ}U�k�,�W �C�ɞ5:ʜ%�A�U�>ܙ�@Ji�~C�I*`�fD�L���%/��^<<C�əg��
����r�`ܚ�E�g��C�!7+��{�K�o¦H�f@'�C�	�,�u��h_�k��D���Z	h��C�	[Z�Mk�3f��������C�i�����pǤ�x�C�	��x��k�h��[��(>��C�	+Y�IGmδ���"�m�]�~C䉘{�hˢL��t����VjC�I/
V��Q:>�}���X")�B�ɓ`�����B�J�d�PA�6CTC�	M�d�'bC�Z�^)���b�B�V��ܨ��Ǐk��p��I�bC�	�'Y|q�� �!��8H�Fܩ	�VC�	k�Z��Ʈ�,J(�AQsH[:R"C�ɖN�N�ō�AB	��v�C䉙v���a��8l�8��A�{RB�	C�H�0�i� jZ�d!�*�,3B�Xt(��̝���<�D��)�B�ɝt�Թ#�P'6�D��n��� B�I+�t�'AS�Q�$9��Pi�B�ɹx�}R�F5HZ,a�6���3��C�I�.DͰ/k!eώ*H�K��=��ΪH�C�{���g�8(�D�( �q˷O���y�g� >=t�'�Y�"�,0�G�̟_z��K�\p���>�q��'X��
Ҡ�/R�8��/�9�)��_Y���Һ0����BA�\�SӃI�%�$�+CHN�.�1��;4?�����z4j��EA�����;;��$���Q�O+H�#B�T,�8��JA�~�VI`��H�(�`H#��Л"S2���-�D(<	p�Q+g�%�W%�V��XcƔK}�MY�(����5$��3�T�HU2pڜ�2+)�S�.q���o��+1,҄ Y�T�B�I-9 �J��4U�����"Zz���c O�7dŁ�9H6�%�>��ʂ�w�6d�'8nlY�:�YzA��He�IA�bQ����e��49-j2���8V:�"�̈́;.�3���"���%B-4�T����;O$�)#̓�~ep1���]O�(���8Fj�A�Q-	%�1	�t�Ǧ@nZ!Q#:�%;��AhD2��5�dȗgM
�L�Q��Y��j�0��k�Q���P�.[j(�|�7�L �T�iEL��Q�ҟ.@@��IaL%F�<`�Xx�"Odu��? ���c�Y�`�\	�Cȗ�8��鳡��8y�z�Ԃ<�ne�8����3'Y�e�D=��8��P�'�4KK�A���%���#�'ф��8 zD��)ET��(d�;J[x@ړ�F�z���$�GȠ��%��<,fx�wk+AS�O�s���?Wײ� �a�@��`��	�b�<��G�[�" ����.����Γ
���T����]*�KZ`���K�/E�<y:�n^e����B��U��9�N�I���a��@%��f
ޭ� D[�jV��n�T��	1& ��M�V���e�A�M��|��!$$A!�m�y�<��=3��C�O_5e9��!`\�48�cC�?D��IV�^��%{�aR��J�'�h�H��x޽:!Œ �Z�zG��Du	2&6�O���Uj���� �-hcmW�
%^���K#.M���Dڂ5�|�����-C��I&���&k̇��O�p
VAG�-��1�dL��|-D���ɯ}#�x"&F�+������z!P��72���j��]���pQ�εZ��6�i��K�@@2(bՅ�h���;v)��^���8�J&8K.���<a��x��IP�zH�Cd�k���'EE`�n�';N*����z}4i��E��R�����^].C䉽��aر�ǅa�X��V�>W�>��0��Xt@ �,mr��{5�Ӽ
��i���<�o�9̿S�^�,b��:�!�>�^]h�Z���=!�.Շsq�����.F`yD�
fz|аW�P.U90Б6$��E>ލ0&��D�.�x����ûS��sca¨�nH �(a��O`�:�l��q���&BS��HP���S�Z瓕��Dx��T�(�d�V�I�tC�I�&�=�/�*OVaQ�I@$$,Qs���/�<�rP$V�
l±�6#��?Qλy�Dxk�*��|��A�w���V��X�ȓy�"���{�Z����g9tOQ>d��M����>E'h�A@��i]&o�X"<y��/7�>XH2n��?���R��_�����,L�*?z�)dၬq�Z`�3��Y��i�Ή�DnFJ'��=��q��kOQ���u�֊=d̐�*Ǒ~��Q��1�I�9�,��+�w4��Q'� �"-��NA�|�W�/fʒA���,�]
E+�_�<����-w �!�EEE�&�p�y��țt�ZW��]^@�:�߆���'�缃4Jۉ)ԉ�s^�_�Z%�TjS�<�� Zr�Z����lˆ�� 8�!0��Ÿ^�THq����j�'�HOލq��=Y��k�	1Y�D�d�'��#CJ��@��-�-d��<�G����:ᡎJЎ�R��#C�_�T� 1eC�QZtEr,� [hd�Q�ŗjLU�O���h�-[_�0B�"
�lJ
�'w�xk5�ƨ!�����&%�A�)O��F��.��8�͆��ȟh4�`D=$���C�"<�Mp"O
�2�+M�Jz�T�����'m�2!*v��|�]&�d a�����g�)����Q'C�%^&����\K�|���)���Y��V&&,J���� ��'�088�bC��a}2F��άp���
Oㆥ�O���p<1��M�L-2�#������P�b��ӡ=.x$.Ѩp�!�DԈ�9� ��j<��Q���1O>��h��F����TJ�ޤQ+C>d���ǩ�s�<�`�ր+��=��n_�zk�����׶tl	�=i�+;�gyb�
"M ç�	`4�㲠��y�S�:FX���,�3e��c�L'�y�,d6xtnǏ NN�� B7�y2n���ST/�9sf�Q#��7�y2�Ǟn���Gn�8�bh��yd��[TiSካ[!�I�D��,�d��m�3����@�`Ь��ȓu����B��B�qA�G������]0 ��ӏ#�"|y��6}����:�,�rG��q�9�4�S6�j�Ey"�;�(�F��N�-+�V��c�r�	uoA:�y�T�EtF��!'�~ Aũ�� �J�p��8nyzϧ>E��'�qS�HxO��ۆ ��ō"D�HIS�_Q%�p��P"x��aI�Ozx�uE���d�	ۓ:�m颠޶i���
EN�&Rd�R�4Dr�`��8��6f˧jԄd8d�%�2�kD��ZC�$[HQk��Tf@PQ�L㟐�!�!5D������i�@	���F���K'L�'@�B�ɔkw%��)�1�
�P�
��k,�X����/�lE	K��E��'�f��F��4��6�U�H�@��
�'�ry��	i�\0��Y�5�4ٳ�h����VJ��{����
�gP�b�P�E�8�tbĈ;/�{2�2M-R������)ŀ��qhh0{����BV��)s" D���퉀X�ؼb��
v�Q�
<�	=KpN��#)� ��>�P�a�G<H��R=]�!r"0D� ���&z���eꇴSۂ�x�O0m��I�HN�)��<aV�	&��B���%�8����T�<Q�#֥\Ru"�c�>�P۱ DV?����2���U?8�h�(���,_�h�Puo^"^!��5]������pC&L���nn!�� ���r���enur���&c��U	��	�A}���b�S�J|�@���=;�-�5�Ȅ6�C䉆vA����-�13�	�F�Z~�mxW�˘�%�"~�6Ј�H#���8�|��$�k���ȓp�9Ӵ�P(&�ܤ÷N�a'���3L��ZR	;}�a{򨈁xV�P{��4a��ccK���=QSƏ�5<�d���hӎ�+v��D�>����1�h�t"O ��GOX�`iP�@��X=�&��W*ќp8oޱ�H���L��=*�z�E�*R�z�"O@L�-92�Z�#M�pz��S��t�ܠs��`��-�g?r(5J�6�ҥG��C���Ch�Q�<���vN���0G�d�t�`��䟈H�ۋ0�h��'V���MF'xZ���_+�%Bߓ���P�^ GR�6�V��
�%ģhEpw#� �!�26���Ɉ<5��0b��Z]�O��!K˚fj40Y�����aϺTJ�`CFV�!�ď�I�� R�M�<<Ԅ<蒀�;�� �t�O!wچ�O?�I�4�r8J_�0Jd�pj_8EUrC�	>
�D��L�C��U�p.۬V��	�g���U�'����˪_��]���*c�N��'��S
�!_�8b��\=o��@��'1h�B��_	 ��Ξ�K��
�'�X��աȹ�x阄�L�Mu,�S�'�j(tc�8n�@�nK�F��'�<P�ʕ�Y)��])-�P��'ܐa��cm�U��oc44"W"O�ᚣ�jn
E V$�%yfpYbQ"O�d�,R�WW���ΣI?��K�"O��P�A�y�P�bs�SR��q"Ox��Nԡ*D����J�̨�F"OV��'�K����ٔ	Z^|&�W"O>|�Ah�5S"�s�BB�1���"OR����I�Zq���[�r͔1E"OTeQ��L�Zl�aPvb��J���"O���Jވ90��GꙂ�VX�"O���6� �ej�d��"�"O�1�HM��޹B/ (J�*G"O�����"V0�"@�T;�ɢ"O��)d���O����c)"sr��"O�Ԙ��ͱA�h9(S��e��"O����$��2��Q3W�[�Ra�"O��3��os��u��U\��"O���q�ƼvPP��t�I? V�S"O��2�y�8��Ά$N0"O�]qF�F# �-��A� 'X8Ja"Of������2��(zp��"O�������Y2�����-�L��"Oj���b�3
��I�kG?|�V���"O�<J�j�Ac��St'�v���#"OnP�Ed�;��ঢ়��"O]���+8�^���4}�t"f"O��P�K�yx8�TfŮ$��$��"O���>0D��&ѺXl0�cf"O&�!\�h�p��.U�P��"Oq!l��K��� ��$"�5�v"O�Q;D� h��B�B-,���"O0�K�̂y��|�
�#E����"OX�Ӆ�
2"-0��&xp�
b"O�BuOE�'���T�R=e�p�"O�,�b���A<S*��"OT���"i+� (�&5:���"O�j�®g��TˇA@�Xٹ�"O��{R��n9�n�"0!���"O�e�@�ՏvFDm��$N��0"O� ����㑩 h	���?BF��q"O���#��W�������M���T"O��K��`P�Fϋ'm'K�"O�lx���i�ɫ��%y�"OQ����6�ba���Ȣ"*���B"O}�5�ͭQt4=��*�\f�$��"O^�jd�ʞ	 �0
wX��!�"O���S��S\:�wj�&_G&��"O�E��G�i�4�C��+B (�Y�"O�C̈�^��1���cq"<��"O�P*3��<q  �R�Xau&8b�"O�X!)�(o���`��}a,M�q"O�aj�.��6��N�B���Z�"OȸA��]"e����-.S~)��"O��k���!��lKEJ��2`"O��C��Z�P�4�÷1\�5�W"Ol�J�	T%\�s�Q�mI�D
�"O*���O�F�hL@������U�"O�� �'��P����aU"�*p"O��*�]-v�P�������"O�9�MX�D���;� ��vz�:q"O�lJ�Ε�!��a��P�T�1�"O���O�7Xz�j NHGܐ,��"O�X`B�U�;�`E��dхg����"O��3�c��?{��{�eP��8�CV"O 0���A�/��U3�U�n��A��"ON��ख़3F�ȱ�j�'{O���"O@Da�/IT�"�1A���"O0����"gO��q�	�`n�PF"O��uNǟgF~q���k�:D�"O"���$��Dܰ�C�$�xF"O�������)c=�&�~��eZ�"O<�jF�Ό!��P�@&"���z"O>���&��T�l��#K,`�z�"O̥�r�^2�1���^ Y  �"O 02M& )�\@�a
 *`�+"O�8I",#e&`����Vd���4"O�,��.ҧ<tM���e�P��y�J*J�\b5�ο�N��7���y"��z)6�p@�Y����qW`L�yB�ƌ
MD����ƚX|f�
��ި�y�F�.^[l�-Ƃ$X�� �y���/`c8��U�=h�	!n��y�(M�b��p,4U�8������y����1�`�+Vʅ�A[�A0M��y�iĴ{f8	;���:m��b����y�o�E�|#FÎ-��@��Ƅ)�y�A�8T��C`��-C4)4����>pY�xr(V[X�h:&L�9�f�b�+5���f�<�O`h�co|z"a�1�hu��W�Wl����NG �Px"��%W�2��wĔ�#�Aᕯ��hO���)�/O"���(��:<PUya ��DF:��D�ׅ2�B䉩mg��2E�҅G<j��8'U��$�(P:u(D ��E�l�S�OS����ڄ-���Y�oVD��<j%"O(����"7#6d��dϹ%�$iU�����א;���ԥ�T����c�U��P%�L�����A`+�O������j7.xyÃܚk�l�cva
�e�a!��49�C��&-�Ț7N�)o||�w�"R�r�=��`ɉ6����䉊^�UЄ��l:`曈6X�@`DJ�`�����&�V�<��׷W@*�Lͪ'	�1"@.�̟t;Ł�W���*Ҡ}���1��.��IU��(�O�0+H:��8v(P9i�1�'3b8Hb��rV.TeB_�J����ɋ�(�B$�S#�ɂ�	��B�����o�sW�i�l��&�^$+�/ø=x*�r��D}"��q�.L�b̛�v�f17�� $�T0S��\��t�B�J�HGdi3�'I7�,��Պ˅)L����S�? N�h���Ze�Q�M��}�x��O����-iZ����΀2#F�b�J߭3۪��V��=� �Q�OL�<`�R ��T�Uh� ��Y��'�HDR�$��s--|��p�6�K�rG.}cAB�18����
O5n�T874���Ur�Mϻdb�:�f���`ĩ���S��a���#d�~��5
N��D���ÿN	�8�VZ�,N�m3*�˴P� ���I�f}6p�q�'$�m:��N�f���Dd�,QJQ���D��%#�]Ze�d��҄$�SH�	��m�Р�Q�Ry����77ћ�A��@j6��\���RG��9G��:xjqA�J=H��B ܸE��9�'�g�j��4�ݮv��<��8cUc���`��;���s#���e��I�/�T�!��G4+���HŮD�r�H@CI �jt�i�U�D�GHĵG�<��LG5*���x�^�\�����u�G�!p��ɂ6� z�9:Ǧ?�O<�ː�P;3�6��sC��v7� 35NA�p�:�Xe!��︌k��2W� �;W�#?�n�d�ң<I���?n�:��	�dǲI���,�(���Rj��|ږi�E*S�U�­Q���Tc�*�F��``�t��[� ]��y�kS9jM�10F	�&���@gS�S�8��&���`�dE�!��7z.�I�8��O��nՃVe|�;4N�"4��B�%�!�DZ�=�0�s��
�r⭃�������� �ґy0�+!�.�@�O�:�#��ɆX��ݱ�틘i�.$�u��"7�����B�Z/l "��_�^��5�C���4'��B��A�ଢV(�1:���B˒*�����C�&�	Q��-�Y6,x�O�9����0�Pe:�"�,0�c@�2nZ��S+E~Je�r�ɵku�Qȕ!h�B�	��H�YGaųe������A�@��-�wZ��O�~g�2����Q>睰D���q�R���pf�o:C�uXU�ЊƘ@��蕻 �pDL�v
R]���F�A���5�M���F�'�f���U�H��]{s�� _�0���| �B%E�'(K��6eE87r$[`$ ve�L�D��oU^����%)(�9���ݜgx�؉�a�~�z�?��q�����b��'r���֥C�jg$i����-s����ȓ����)L�s0N�R�L.<��|�'7��xU
ܖ6��	�|�O�>�8@��&K-�I�g�C�P�����'��A�V��?��x�!�ۓO�r�h*�m��	Hْ`���Fp�3��0$��0��ǭi��$	F4C��0%���yN���i�.h��L���@�����(��>ɇ�YM�i�%��:@ʝ�$\y8�0	��ׁ=M�'��H}�b�)7�E�Ӂ�!_�(��1�yB�g�f�SKԷ'�6Ku��ݘ'�2c%���\5�?9QC��J^�SD$�;XP��q�!D���f	bP����ƕY�er�@ Hi�➼`��<�u�ځ5*RjHy\]C�E�{�<�CϭWX&{b�9/s�L8!��x�<Y�i���@�	qA$|���!�t�<��
�e��d!�
U�2�1C��]�<	�`I�J~2TRc�_ 41�T�K�X�<iƍ�	#��1 o�Y�@ ��U�<�V�@&p�Bg�=@��!�k�<Q���9�X`��3T�pt�D��i�<���x�`�1%��@F��Z���e�<1e�A�n��0��Ǻ5���J�E�'��Y E�i�O��[3�#ZM~�s��FTd��'cT4I5Cu󚌹v)�3�Z� EV6��@'�|��9Ov��q�,{�l��m��U2Z(j"O�e;T�C߀E��� 'p��P�'D<�q��(�
t��	�Ri�U�C�Ԃ�Xy!���7���ĕQ�,Uq���M�PE;`϶ q�F�{��M(c�XN�<��Ë9`1!k�!%]��׉�J���4�8�ǚ
v"}Js�P�zG��`עQ���k�N�z�<�E,��o�)��*N�.�0�C�,��_���0�X����h��d�5rA�dO4rjУA�݊N!�D<uъ�`N�kgND���2�2��<��F�d؞��v$�4H����=�B�@Q5|ODp�j�
�\���4|����'�%c�xM@`[�i�����؈$q��9;���e�
2��?Q���0�	a�$0�'a��;fm��0,L���Q�"�ل�$V,��v.��4"C�P<X�z�KBE�n��1�J>E���� �zP愱;���s��1h� �`S"O��{t�Q�UM�I)��x�ڬ#�Oإz��9�0>����X���f��@1F[�E�W�<�q��	x�Dtꀩ�4�B-K ��P�<�bg�4�\Ͱb,Ü5�f({p�T�'6I�B'[J�OOdh#�%��qZ3�A�!��
�'t8E��ݻc���b&�W�t18R�S��ԭ+֘|��9O�P!mؔ��|c��'3� ���"O���0(�y�*���(f�D���'����O�)LZ���I:��HD��Ze�2E˗V�F���U�([�T9u�D;�M���+R"����	$�
d�&�N~�<��'Q�!E��z VdQ+�}��M'dMۧ�� F�"}���S;}Y��޻%�U�B��z�<�M���	��)��R4*�f��P,��Y)�铐h����:y�ѱ�C�5@2vI�w@��5%!�D��~<��aT>�Y�7�6C2I�>^� �#U؞�°}~ݒ�b��"e:�Y�,3|OB���R�0�>��4\��t�e(̪V$��P5_;DB���s �yD�s�f�pt�N�F@�?a� W���(ҧD*D�y�	D�T��!�sh�u� ��w���!��z��4BӮL�j���{�����2�O>E��'`Te0ӏX�n�<X�IX Z���'�f�9�"(R}됾�e�7!b?	���U�8��$<nc��2�_6��-�"� �>p!�d�)�0H �����	���֑e!�J"��)���H�V=��� x@!���xI�@���/Aod�Q�л!!�D	�`����(!E^y�Z(z�!�D[�o���(wht=B��J
��!���K����f�~Ml!�d�!򤌲B��,D���^>�)��@= �!�D q�|Q���C���rA  !�DQ#�6��A�)/�tB�a@�uk!���:Of��Ģ��u�&9�!�+6�!򄃊h�2���< ������!�`n���%E�wzd�z��ӷ\9!�$`� ͘���.Q�D҅�|�!��K�t�½sB'�2g�zde�((�!�$��&셛��R4l��`e�E�!��8�*w���rD^�[��ߎ�!�V	}�hQAGM���tx��a�9o!�]L����%.�*�DJR�#v!��P��L�|"h�P�Y�t
!��,����P��%�F�@L��i
!��F�a&�i%�Ź���+%,_��
�'�e2V�U2p?�����Ɲ``j�
�'��	գ�����1�ѤâP��'�đP�/�)�z8p�eH)j��Q)�'O���Vm��&1�e� ��#k�V��'�8Ar���6�y� eJ���']fp�`۫x�<|�f���"dL��'��y�'t�����@<"�x��6�
�b%=c��FdВ���*�~)�ȓs���֨I�e��S�j�@Vȓ|,��$A�&'z��bo�G��ņ�z�~*���C��TB��K�<�ȓ$BƑ�1m� �� N��{-P@�ȓD���I���>"¦U�,�;|�F5�ȓ9�|�C�]E:�i��\ɲ���9ћv�<��q�Dʖ�����a͋��ɭ*811!�ڗ-����3�'n�T(8V*J�%�1��.
�GCb�'��@R�Qp$�`>=CTk��3��!㢀G9�x�ãóD��}1C�^�.��y���<E���Oz&y�C��.X���i֬ć��l��Gҷ>U:튵�f�H6�\���? ԩ� Y�N���!!+�q~d|�b�*n�a�ܴ7%f�I%��L>� �H@����HA�պw�	fD(H�̈́T���	-{����qf�4,��?�'p���e��A�𐚥
��)#Z�
�?On�d.O)Y����"��l�O��@�����X���]�d���ZufՀ4^̈��M�N��!@���.�?E��43��$��� :hJM���k�\�Rn� ,����h��	P�L>�'L�T!�A��O��T ��%-,��DkUB�I1%,.����~�u �
� E`� '�
�j��JG�<��@�[�"�{���&w�����đ@�<9��z������E�s���4
Cy�<�n��a����Ak"�7��y�ˀ=�"�����*�����ŉ�y"�O���F%ԝL��uSLĳ�y��ݬ]b>C���=�d�a�Z��y�D�.)Va;�P<���Fn�-�yR�R6Z��G 83-�)B�'��yR� ��ȠE�(� \:�Ώ3�y��H�w���sfh+J�����N���ybC� s��!1�_�:l>����:�y�$� TX��?:O� QC>�y�B. S��z��_��9J�d�$�y�gr��4!#�֢^7�`BX�yb�G%#,�u�J	�[��yP�����y�˖�g-�L�7-�Li��P�JL��y2��{�[S�E?	X9�D�(�yB,ȇ"�:��`ȯ>�����>�y2�ןc��]h���g���'r� 0��ӓ
G�麳�M=b3�Pq	�'��H����sjDs�E��*����'��{5��_d(��1xA\M�	�'�4E�5k��x&�QT/Z�B�Z1�'��,0r�Rش�$��IO]��'y����k�4�d�2��[*0O"A"�'~ �2)Q,�Qꑪ*�"գ�'���
�
�/k��Jw+A %D��'��@�"V0y����`����Q�'A��`��[����&��z1$��'����Ғ0�v���n��uƖQ�	�'�U��C���r���<���'%tL��� }O��)!�2�f��'�!S�nׯ���+u�_%&�vu�'Mh��3�ҿ��H���r�Z�I�'�����;��JDOl�r���'�r!�	�#���aGMk-��a�'�T� 3���vvpP���dM���'�zh;��ޱn�� p�	]]����'�\u��,���0��!�On��'q��A��մ9S@1�a�F�(�a��'.��S�1w�0��n��V��'����2��&we4��6�^3Ֆ��'
ʀK@n"g{.@`�ȝ�8R���'�֝�'	�����w�ʔ�D���'\�4��ҁU��I&�M5(ul�S�'� �4��OL2�#Sb݀$ծ%�	�'�hh���9b!s�N	'!�|�	�'1b,#�Ɲ�'q(��T�Ų���2�'�vTbe^�h�hԋL��-��'����ǕX( ���^�z~���'
�㥙�,���'�V��Xih�'p8,*���jԘy�!9����'���4���A�ҁ��\�z�T��'�ȠR/��[�V�����)�$�)�'Ml�)w�Gr�.��b�W(��'�� V�;VLƙ�h���Lђ�'�Bp�(cP���m[|�"�P�'���A�*Y�C��l� -Q_c@���� *�zR잙���j
ë�2��"O>��1���SZ |�eHZ�6��X�"Ot�����WZ�Z�a�Mα�"Oq�&E�kdJ �^� s"Opyؗ�T�S��%oJ"=�"OR��/��[AFI��N͡~��2"Oh�Ƃ�.l1L|�ƌ�!$� �p"O}���UC�R5�cK��Ұ]�"O>� d`ĩ4�X��`+MY @��%"O�tyuό+c�^����݁R�"O�i2'
/1�}�Ňȣ;@��"O�!�և���p�9)o
�r�"O�h��B���ڳg�<,(���"O6�	��W�q3R&���Q��"O p�peK� {�	�ޖ�(�~S'"O�d�'�ԎK����i�<��0Z"O��KH�?��K�H
�9
D@�"Oެ��`�=tԠ8EB�x�h��"O��
�m�"g��!�u�C3u����"O�H��g��1뤄�:��R�"O�HZk�	tdcv�X=���b�"OYb`B:��:P�v��`"ObicRaE�y�.!1�iY�b��%��"O����GÐ}���'�-ږ��a"O�i��Ƅw��@�de�5c�vը�"O���0��{����$�7�<*�"OP]p&+m:��jWCC0�$8�"O0��`�<�J�=�tEK�F΋�y��:beD��g�� W���M˳�yb)�ۄM@AM�zp�3gO[�ybh��x�a1��eP��r���y"�ț!��u�aF�23<}Q��y,/F�4�� �ʴ5��H[s���y�P�96dr�g�h�Hs�Г�y���H�X:�IP���i"�[�y��>'	�e[�H�s8 :a����yr�����I.�.E0ZJԭ�yB�ـ[B��!�͗r)D��`o�2�yb�F4[id0��K+d���Wi���ybNZ�Fd~�����VXp�3�2�y"��49�xl#.[;P�"����X�y��+{�H ��C�� KC�
��yr�V-1��[f��>�΍�u���yB
�"kX�QI˲2��Mqf��*�y��ؽ>���W���$ɪd;Ƈ�y���&WDt�@E�&g�H��#�y2b^
h6f��u&N4u rU��y�+�L��iy��D"�d��$�R.�y��4]eb,A�A�L�^}� ���y�!f�
U@Pc��/G.�9J��yR%U�l��U�-<�0Y�׀�y���^�]��Ť7B̭�a�-�yr9�� $!ް�	��y�Ҭ�&�	��a0��y�W���x��ֺJ�М��h*�y�V$��5i���<ۼ%�����yRRc�l ��kI�:�X%RTս�y"E���H����}]DA��kO��y2�-E���s%«} #3�œ�y�f]"?�°X�R�y��M�� V;�y"�͌F�^�J�
L�d��pAZ�y���}���>f�@x ��!�yBIU?���*���	cp(٧����yҥ��x����'EՌ[��i1@�і�y
� &I� '!-�� �j�� Xl��"O.Q"�&��OfpL���� <�r��4"O�����,Y$�	�Gir�"O\�ʗ�B�����!�.M��`;�"O�`qd�mk\)��K�p�j�hQ"O�x�aC�7��:2J��}8�H�"O�A��&�̲��Ӊ_-b���U"O� Ĥ� aC�� �bҏ �ؓ�"OR)�E�_��u����8"|�ay�"ONhp���8a]��r4`��7�@�!"O�P��+YE�68�w׋6��aqp"O���$�8g���0�Z g'�\f"O�-���)�-�n�X�e;t"O��x��ë?=0}!���&咅"O,\ȁn\0]l�Rf��5L\�[�"O�A�T=Yd�0��k��W"O 쩢��_`�a��'��=Jb"O�L�b	���UJKnuHD!e"O�If�<���È�m �pT"OXX�� ��y\��I�4_:��a"O$@:�!�4a���@�(Ǌk��@J�"O[A�ܝu��,�g�!g�B���"O��xbG�"�����w�u��*O�Q�����r1
�+�"-a�'؍Hc� aڄ� 񌔂 �RX	�'L؍�� �X�p�!��.�����'���Ч�� ���bOP�u~ `�';�O�A8Z�x�i������'0��*�oR�/�8���犹H(��s�';&9�.�0Z4��h��Rl:j�"�'�2�6n@	S�@(;aNeg$|��'�>(А߃EJ ѡj�0��!�' Ȉ3*��t\lh;��͓*�"�'��9�'nŝ)��l���S�����'@���b�-<`��H3O_>�(�	�'�~�: �Ֆ(ؒ��r���m��{�'���6�	3����b"�Ps�',u�mǡ ��!*���S�:8B�'I�)�f�ߢ����p$��K�����'���:�$=�j���̜�s��0�'��(ց�7Si��@���f���k�'yq��!����Θ�,=��'�p�8��B8#<΍��@ye�	�'8�p��"w3��2�ƚu"���',p�2%h�(s�i�nx1�'xV}��
��C���	��Xp��'°cԉ� dx��a鐨>�"8��'��5Kș/4,t���	F��'�^����G�.F(P�KK;J��x�'>VT{�$��x���g��� ���
�'�&��`2}�-�L.�u+�'��Z��XJ$r,*��@�?r$0�
�'��Li�O:/���1& �==%R�'���j�k[�G"ΐXuj?0e��
�'�މ"u�H3>4U�d�K=`R`i
�'t��1)�������P<�d�x
�'�n ��J��
9�YY���A(�A�'R8��g'ǭu��`�Ԡ>x��'�T��*�Ӡ4�&��7�����'�IV�"$<��lP>5����'yR����,CV��h�9&Hnqk�'�RQ�)�4)���[�̍u�"�#�'A���Q��*��xY%�#�(@r�':����	) ,����&69{��� �F�U�J�B�L�9"OX��)� �4���H�"2�0�KE"OD�1����ʂ%�W��Cx�;"O����  �#\��v�8lBp;"O�}k���2i�RA�V�Ӈ9�Ĩ��"O=�b�����`�N�f����"O��sS.'��Y�T�EE�BR"O�Z��_�`�L�ȅ� �E����"O~��E��n~�8r-A�9.��cc"O�����ڵQ�>x��KI��B"O�����QvT`H��<SϠU��"OxLbcCN�F�.�3��n�J���"O4"��&�F@K�Z�`��c`"O�Q�Y�H�ƌ����?�֨�"O
-#"'^:o����`e� �"O�ho�q��M�9�L��4"Ob�Z"�>�	�a/�X���F"O| ӆ   ���M)99d����'!���"O8l���ٔz����WÁ����"O� ��H�~��!ϻj�"��"O�c�̓�h�T-c�&H�|o ��"O��g�ܷK�� �&˦0f�5yw"O��S�Oײ0Ӡ�I6&�(�z�pB"O�jaL�^U��@�|*ƨ9�"OnȨ�;]�:�2 *X����K "O���İe8��� J��M�Vli�"O��{W
��Jz:���6)p`��3"O����O�m`�,�,s>ҥ�%"O��	�-A�x�vX��S=���*OI�D�X%V���C��*1!	�'����b�^5�d��W�iޠ���'��\�  ���   �  O  �  �  f*  �5  ?A  �L  �X  �c  ,o  �w  |~  0�  Ύ  �  `�  ��  �  7�  ��  "�  r�  ��  ��  ��  1�  t�  ��  ��  ��  f�  � � � � q! �) �1 �8 =? �E *I  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy�"Ob\B��;h�`��Ɇ*���S"O�h�T�ÕZ(jܫ� ��+�Ƚa""O�A���I�{"��qReM.v�\�J"O�I��cR�G�Fm+De����(��I|�O���#�H�R!��њ]��p��'_��uʆ�vӲ�R�c�*m�'�*L��܉�` ��ڭ\�����$֮w4I�1O�,��g�W�b-h4��Ӽ9�HMB�tX���;%�2���IЦ�Fx��2R^zmC`� �p��#�ȵ�yRO����!�L�q�tR� K��$"% �"|���6U3��B0)зez��%�~�<)0��.)�#U��4��뵥�T�<��۞@J9������
�ĥ�F�<���R�}��%�	2a ��`j�<�d��W��aP��ۆ&Z<�j�g���'o(�TA0g�]j�ȺS�����'���G U*=�~@�g��J��p`�'X���	B�z��X3'�R�m�4u�	�':��D�K���@ W/�S<������ �\q�C1������h=�A�#"O8��N� Gv����^�g �<#��>���tl@aM�/Dc��2X���ȓp_�B�"'���BQ �萄��N5[�œ�J�lU���V ��-D}�����Q��*�	��ȴ�� �C�I�qv�d��+̅Z�����슃'�B䉌�����"� TU��gɭ 6#>��C?�'w�6��![�.v���a(3�i��j�X��`	O̙K�aX���YΓ�hO?!F��*e�@y�FP�@�XɫA0D��:4��(N���q�S�/�����,D��z�K��U�TǄ�'TI�9�+$��g0��9�� �:�����o ����9P�M���4t\�\����ayR�O֒O�0���xb�Ӷ���V�{�"OQ4�B�|;z��&T���S�pG{��	�d�\@A �K���)��/�!��>P� L"��"GBi��&K/}�ttFz��9O�I��rL,y`��hX�xp��'��+K�Q�����T��������1��]m��<)�]~��ʆ�&O`�3�X'>��1��	k}�K>!B�;q@ηn��l����yRaA�90�����Zcz����Y���OL�~:��N�8aޜ�A($}�q��a�c�<��R;/xВ��E-�:ѡf�c�<Y�Y0�����j��u�C��i�<��#=uL-R��	�+($Q�E�]�<񳋟�%D��O�g��,P�I[�<��g�&�:�r&l��G�.a��&A@�<6��_N^�R��:���� �y�<�w�ґH�yz �3�`��� �j�<i7�}�2٣QO�p����2��q�<�5�̏�xq��T,�s�F�<�#��![����UN�t˞�b!W�<��k���≨��Q &Р��|�<�ƤS��ڑ�UF�JIj3�Mq�<���ߣ��� �M�1vN�Y©v�<�q#����g�)��!��v�<ag��R�F�� �>���Вd�V�<�����Ttހ	�[\��,3aL�i�<�a�C�2��-�I��T��x���F�<q3 �jT�㶦ւa�j0I�~�<a��WB�<�S�	?sC����j�o�<�"��P�:���=bJ��&��n�<�/�"��ړş6K2zD��c m�<�6�P�*���^�B�ވ��ŋ}�<I���1�0��#�3c�R͒��LS�<�$o�^ľQ�ԀR;1�:�Ns�<�d�)0��f�g�����/DG�<i���B���UB_�&���SFG�<i���b��C�Hܭc�����<�k��FWL�#�M�%j(X�FE�<�ä���8�d��&J ��DoV�<s�T�\���9�2M���Q�<��/	�P�RfD�<��l�F��e�<���G�#�H�1�K(v�d�4By�<qB�"J14Y��͏%�B���t�<�PHZ�:0v�a�U�E��!Y��p�<A&	�W�� ���~tb|��o�j�<Y@��.k�:��m�9pt
Q�5%f�<Q�4F�(�3�����k�'�F�<����r��t��v�J�{F�{�<!ݚa��	���.����d.�z�<� v�B_�0�q�� �f�2���"O�}p�4�V%Y7b��i�!("O(h�`�lB���5�B�	��""OJ5�f炖l��1��Åw ��Ҵ"O�IȒ��&$.i�Vo>)#�ı�'M2�'�B�']b�'V��'P��':L�Ye	�#?�T�*�j����ͻF�'���'���'N��'���'���'��q��(�.mZ���x��1r��'�R�'���'SR�'.��'���'�:�`I޽f��PmK;�8h�t�'�b�'�"�'?��'b�'���'���# ��4a�R�QB�Ɣ�f�'}��'���'q��'�r�'���'s.�[ukF<7aq����`%6���'���'2�'��'w��'/B�'��p�D܊o6~Z3�E$#d����'���'b�'-B�'��'�"�'�8}�#ެN:�J�MI�?	����'Q�'��'��'b��'7��'B���
I�s�t���ع5sx����'�B�'"�';��'/R�'�b�' ��J]�<�K��ӧc%tQq��'��'0�'�"�'*��'/�'�b,!a� YH�,ܲ4��>�?����?���?)��?����?���?���� #�d���B ;�
1�A��?���?i���?1��?y��?A���?�r+�
�\��,O=4���+� W�?Q��?���?����?9��k��V�'���Y�i�"qR�)�	�~��5ET�3����?�)O1��I��M#E��(���h⦇Vvb�S�"��'��6�.�i>�	ݟ*� *���	%K�*$*)�u�����~ �pn�j~�6�D��SI����#�l��"�D.B�"����1O��$�<����F$xg.����,$Ft,PnƗ}�oځY��c����S��yWl�#��XbO� ],��I=���'��>�|j�kݯ�M+�'>���1�G��T�P�2Gz(9��'����$s��i>��I�dpi3פ�+�PEZ+6]���vyb�|�v�m�r�$D�H���rωD���d�����v}��'�6O��'��P�ԖqfD�F-NC�H�'����p���i����Dş�i��'x0�&(d�s#��c��u�QQ���'���9O 4�7��*K7�8��F�.�  "�?O,�o�3���%כv�4�>�(q#{����́7���ڴ;O<�$�O����V�6#?��O�4��ĉ*h6�Hc��qJ�x2�F�@&>͢J>Q*O��OF���O��$�O���C�K�8��E�@K��v�H��	�<)�i�t���'r�'��O�	Z9R���Jf�D�S8Cה�@V�fE�O:O1�0�0q�Av����+S-#�н���{H
�W��<a���!y���]������>׀���_~�rуr%�.C����O��D�Ol�4���p���b�!d�!	1]�:4x�L4ځq����y��`Ӻ�L�O(�o���M뀴i��*�J�3�(��LR�4�n�ɶc�V�����p��,[�C�������*0�v�����1���[b�]�3O��$�O����O^�$�O��?�[��##6iB��7F�pT0����\���H�޴z��'�?�&�i��'Ύ,��9,�T�r� D��,b�(��F���c��|1�ƃ�M�O��FoJ7 6��J��f[L�Q׌��>��|;�s;R�O���|���?���k�@-h�� (��E�#�^8l�X`���?�+O$�n�)f�`�	ܟ���w��)^���!�힝$�,8��;��$R{}�B~�b�nZ���S���%;~��

���F�օj*��s��"V֠p��O��-�?A�c!�D��6�.��P.Ta��Ѩq&՞��D�Ol�D�Oh��<A��i���b���*��'�n>)�uEO�RN���'�7�(������1Ғj]�e�I��j�_�46���MK��iJP���ih�Ie1�5�OK�'u�@;�ֺL��Q�k��%Cp��'���'�b�'���'��d��u�N	P��ȫw��pg�TQڴ�d�9���?������<��yw皥hGj�"��F�&���@D(��7���I<�|JB����M��'���	7��?�6IZc%�� 1i�'g�<�sO�����|_������r�d�2�{��	>F_T��6��\������	gy�s��E*�d�O2�D�O`)Q���?��k�d�1$%�D�7�	�����O~��.���An8Y��b	.��E�I��v��I\ZX	��>g��c>I�Q�'��Q�	��i��M�i��.����Ο(��Ο�IS�Ok���Q$JA[q,�++/�Q�󬞝9���~�.�Pv��<!Ŀin�O�C�2��j�۹
�6�Rb����(ߴO���؊��&��leϚ�&$���:]ĬXć+9������L�T��u%�������'�R�'���'��e�2Zp�&��u�&�D���$
��Q�G��vy��'�OB�ܣ\����ϒ�p~Xr�f�r���?���3:���O�t��MB�N�^����;��x�i[.kU$x�O41*�"Q6�?�$j>�D�<9fϘ���Y����I�T�v�̙�?��?����?ͧ��_���v��ă��m�t,�~0Ij�H� 3,������M#�Bg�>����?��i{8��ۑm!�IZ$�ɻ^�\i�OXD�F��\Ҡ�	���	��� �t`+T`K$|���R7>�ҹ��=OF��O����O���O��?A��l_h��a#�B,\�&�(���ԟ �Iڟ�Cߴ7'\y̧�?ya�i��'~Z۔ K�/�.p;Ô/�Z�c�%�$���c��|��L	�M��O��شII 2�&H�oѨ+MR�q�4i��s����<�*O�)�O����OY�Bi�3`s�`���ѕ�:���O���<q�i�(���'*�'��mK��x�,�U5F��r��_~����	Ο@�	��S��.���d��GI�h�>��N��r�i��E��p�O�)͙�?A��O��	ƞ%�˙
7���fC�=Mb1Q���?���?��S�'���妕����=
�4gK/>��9��*E-N��u����3�4��'��ꓺ?)1�ڦ1���@�\�Ђ�ۂ�?Y��i�(|*f�i?�	U�Lp�v�O��'���[1��p� )�8|)>����$�Oz�D�O����O���|���5�ؕ�D�& =$s��������,z"�'�����Ԧ睐\�,H@��p�X�@���	����PyI<�|��Ϟ6�M��'�(��2��1�ƌZ���e�R8��'�XYR�.�韨Qf�|�^������! �§4Jx|�7ǋq�^��fKP՟h��ٟ��Qy)g�dhj��O����O6�d̅5�H���s�����3�I�����O���c�	�P�� h�D$�X� �Ww�H�<y���$���|��l�O���BvN�bL
�[�P!A���-�}���?���?���h����<}p�&���Z%�T�>|>|�˦�A���ޟ��ɟ�M���wH���a�7(�8�� i�;*C�ت�'Zҹi��6�/{h6�0?���+f���.DG�Y�Q .T$x�A�R)$�HL>a)O�I�O�D�O<���O� b] �,�RP�V\긐X��<�2�i��[�U����G�Sޟpq�!����A�ìQbx��U����Ob�Vl�)��<[��a#D����9�cf{\Ms#j�09<�-�B�2Ʀ�Olx�N>9.O|�Z��К����Oo��)ie�O���O����O�<IQ�i�ZL���'��
; 9�t��Ð�HZ�؊��'�t7m'�	)����Ot����ųT�[	0x={g�
`G
���	n�`~2�M)�(��SMܧ��+�c׼��-r*��kB2�c��<��?����?���?!���hQu�@�s� �E"Ri����'B&Ӱ��d1��D�ئ�%�r�)N(mWz���ObB0�a�N�#�ē\ƛ��i���K�	�@7-(?��E�v^6�H�I�$�D((��[�%"Ų�%�O��@J>�/O�)�O���O*� �/�b���	�/I7��9��O����<��i�h�g�'�R�'���<o�� �b�GN��0`eJ`���	+�M�ýi��O����5���=�}sg�0�z<z`�Z�w�b����:?�'���5��4�4���<TjmJv#��Kb������?���?�S�'��d�Ц�c����|���-MtxL�#g���:���'�"�d�����O,}lnb��x$��	Ar�H�p@����4��6�3g������hd�N��4�~�vݔ3GT��(�,h$m`q��<)+O���O��$�O����Opʧ/��(�P��:U�W�Z\� �iT��c�'��'W�O�bh��.�
D��y�O�AP�m(Ф�A��lZ�M��x��D��	[�V2O�UP�C�6q�����mm\30n��<���
�2`����$�����d�'V�U�Ba��@��۶1����''��'BQ��Y�4M��D	��?��<G��S"�O�p�Ѣ!��~T�T؋r˩>����?���xR�D�H\F���!=<��d��D�B�P��)�!#1��X��&#��$^�B�Y�� $#�$��-�2���n���'Z��'��>����M<!��͍�j�DU�$���;�B�	��M3p��(�?9�%�&�4��I�w�#_��:�.�IRY��0O����O��nZ5>��oz~",V2�(q�ӽkZ�噧�ǘD�윒V�F3y�����|bR�������ğ��۟��r���ԙ��@�Ya�b�{y�cp��0�P��O��d�O�������>$B0\x�OC?��� P��PѺ��'���'H�O1�f蓗��
~�b�a�b����ؓ ќ�����i�I��&FB!H~�	tyoڀ0n��VAΉUs��8Gld�2�'2�'��OI�I�M���C��?��H
}
щ�	����bO�<�r�i+�O0��'s�'v�W�"�X@�NS1}V��"lJ� I&X�i��	�)���Oq�&�NܦV zM�k�)&��� u/��OD�D�O��$�O��/�]R�g��.�H"��qN���	͟|����M##��|������|�A��8pE����h=sd�S�(O��n�9�Mϧ(X��4���n⤚�)�w?���!��j�b]0CM��?���9��<ͧ�?Y��?��L*5^�V̒7ņ��6�A��?A������Ħ�z�)�ʟ8��؟d�O���	��&j���;s���,�(K�O�}�'Mr�i'*�O��3MϾ}�֎J��c��#0hPq0E��=�:ܸ�%�>��i>���'h�%���p@����ՒܒO��x�䉈���������ɟb>�'��6�O+�h�I�K˓���9d���V`�)3r��O��$�ަ��?�V�,o��DX�9#dT=V/���QHE�x����ٴ4e��M�|O�V���)#aT8W*��~� l ��J�>Y�:�Zv�>T��1O�˓�?����?i��?������ҙE)f�k�.�=8:H%k`fF�X��l�#@�	�����Ie�������Sg�?;�,`Pf/�XZa�Q<�?��a􉧘O�bl@�i��V�9�~�i%X�<��q�CǛ�N��ןP�M���?t��O���|j��X|p���-J(��q�U���[��?q��?�(O��n����9�	Ɵ ���36��Д�ڽ|�Z8@�(�?�P��ܴk���x�)�37"���gW�幒I�0���ϮJ���4ƕ�f��������a�0�䘪V�g��`���c��	���D�O��D�OV��?�'�?��I6<N����+O�t�c���?ѱ�i-�YS"U��)�4���y�EE�B\�@J�c�&V��y�jdӨ������j٦��'�a7���?�P� 
�>�X*L�/�v�y�m�1��'��I⟔�����	������ߤ|�@��4M��yZ�/5���'r6� ��b�d�O��d)��9:�9��;L�jt��$� Opf��)O4���O8�O�OHLaQ�ٞk����5���|�������AwX��Rsɂ�~���s�pyr�F09��ոD�A]��N�\���������iy�z��	11��O+K��)k�Qt�ԥt�`={�$^�<��i��O���'I�7�	Ӧ�JشK2�݀���7��A��h��\N\�b��]�M#�Oz9�p+ь���D�wJ\%��E�	B�@-���2IJ�pq�']"�'U�'PrT�b>93��(�*w���)���%�_�x���`شX�D��O��7�;�䛎%iV�C�-�/Bt�A4�K$v���$������ӊ6j��nO~�MG�4ζ�d���R��%bX���lYX��ȯ����4�
�D�O��ē�w�Ж��=�F����D�u��$�O��6E����/
jr�'/BR>�2c�<4B(�x�N�W���:��/?ASS������KK>�O���ZՃ�v�(�R�J(+K�P;���U��t�B���4��!��YU>�OX9����Hs�%H2d����@#$��O����O ��O1�>�sޛ�H�	�Be0��]�o��a�FCL�ى��'^��r����k�O����7�0Ԑ�*��Hߞq�s���e��ͦ�%`���!�'h�QU��?�����X��OUdp���J��!�±�;O�ʓ�?i��?���?����򩅑V,,$�sj��YØ�YIY��X�ɕ�2��O��$%�9O �lz��h���%n�|�Q�Ռ_qZ�F�����v�)�>mw��nZ�<��ϟ�J�~�8`i�*H�ܔ�e��<���͊
����L�䓉�4�d�D\�
�ء+��2x�B�*�$�;U��$�O����O�ʓE�����.Kb�'�bJ��B.uQ
I�IN�}ð.�"��OB�'��'J�'��	Bg�}�*AGJG�����O���Vb_�e�Xy��i�?� �O�]sp�O�4cJ�B�6�zá�OX���O����O�}R�6��L��*.�E����K�Dl ��p��V�K&H�剉�M[��wռ��a&��c/�Q(Q�B!����'��7�����4OǼ5�ܴ�����nB��C��2x8I��	j���%hւA������O����4�����O���O����ݰ��I.�f�0�.��.z���6&��wB�'����d�'�D��c�s�a{3�ƌB���S��>����?I0�x��$��F�r2�ț��X�+��hR� ��(�����W"T�K����|bT���8�9A�O�$S=jA@0�G�\��؟�Iϟ�Ny��~�
�1ţ�O��f�D�1y���=D���1O�%l�y��O��1�Ms�i�
6M�<��Lr��<rr��#�b}a��M��O���Ӈ��҉�4�w�^�P�ML4�*dy���'>��#�'��'���'�b�'��<�7Ɛrذ��Ԙ
����ƥ�<��v3��.���t�'�D7M=�䕀2��5�&�T6y��W,��6$N$�0�I���0���o�Q~�J@M��xy��D�i
�b���%>��R��֟����|r[�����I��:��K����DJ�x�d8��R�(��ByBtӺ���O���O
�'u�z�Jୃ93�i�'��/܂��',<��?Q����S��E�6�6�����9���׾}^t�`�BG:��O���?�'�dԹF��1����!@���*֐v��d�O�d�O��ɪ<Iw�i|3���"g9I��4!�R��3I��5�M��҉�>)�1`!Rǀ/@h�!��	]	�$���?!@NF��M[�O����R��2J?�� ���81~�D�s	� &m�`�'��'���'���'p����E�=³oR����i��+�6- by����O*�D0�9O��oz�EAubZ]��W�ū/�fEK�F̟�	A�)�ӄ�]n��<AU�� \ˠ�Ȕ��N�lRam_�<ѵ��E���˦����4���D� 8BU0V��[��h3h�.F$��O����O(�UE�V��H'2�'�o�i��A��\�B�l��FO���OV��'�'��'=RM�r	�8�#���98�L��O&��DN��'z��f���(�?�f��O�J"�?I��x��.8F�Yw�O��d�O��$�O£}��'P1{��Ȥ��) qC�m &�Z� ��ʘ�'��'jz6� �i��/ٔ\�2�0Y6�X3�����	Ԧ�۴,�z|��4��$ǘ�R�1��z�� �dsU"��2.��7��*!��x�/�$�<ͧ�?���?����?���ـi�	z���yTIЂ-��\��M h�ן0�	ğ�&?9�Ir����vE0+Ȑs��� j��\�/Ol���O��O�O0`��p��� �d˥��"Ur�(g�L)$���_�D�e�\�1���Om��Cy�-��2ɐk�T��&�@����'���'W�O/�	�M�wcP��?f�ǸZ(�Hqf�ߵ�����i��?�'�i��Or��'�¹i�6mT�����A	tшU#�)tR�t�e�f�"���U����>��]D���s��_%�n��PjU�t������	ğ`�Iğ�Il��z����/d�E�����
\>�����?!��Lz��nN8��IP�m&�ܢKұ}d���EN,h�p�A��/���?���|JA����M��OdQ" ��>�Rԁ�Z������VQ��O*�OZ��|���?���fU��V�%�Fݹ4��z�P����?A+O��l��(��ڟl��A�h�&	�I�U,͋6QVp��e������\}��'�Ґ|ʟve�Bd"�:Ys��F�F�P�r'W6 D$`,�5R��i>	"��'���$��a�E�X�Dt��iWa��|��ן��Iϟ��I�b>��'6x6��+V��qЊ]�e�x�3�䀨Wz<M�q��<��i�O`��'~"6m]�*�x�6Ȑf��@8�lmLlZ��MK�+�M{�O�|`3Ë���J?!J� E��p�z��[6Bs,�ɥ�x�P�'�b�'���'�b�'t�S�Z
�<�㇆ �����%��_�\=(ߴk��0��?������?�R��y��Qe $�FH=�쵊�'�(SqN7��ğ %�b>���R̦eΓ(S,I�r���V�����H�.�t$�,�ݒ%��O���H>�-O*�$�Oƍtj؇�
պ��X�J�	j��O����O��$�<	��if��i��'�B�'3�q��"T-04,i��)�0�!#�Đ`}��'���|���n��d�T�[�\d1!㛜��D� �� ���7<`1�8��9`��d��d�(��-��(>)xcAK�CMD���O����O��D �'�?��Ȕ�?Z&��M:_���˲fX��?���iU��J��'X�r�j�杈*�B՛���_Zp!�I^1%��Iş`�	��MS���M��O��(&/�	�b��f��IC���7m�D�[�O&j��ON��|r��?1���?��]̸��.�km��Ī�.j�le�,O8�lھ[tA�	���It�'�X�u���s	��K��حqebi3^��Zشdhr�x��ă��`UHs��+LSh�dK�Wz��Yv�+�� ,!^��B�'��&���'�j�@",��'l���ßA��y+��'���'@"���dX�(p�4w��I�7�V���FD,����6��`��)v��$[}2�m��u��������V-p��J<{i�y�"&N�*n�o�A~Z���c��?�Q����wN���%� �	�l$(��Ƹ���'���'�"�'a2�'��ѓĊ�m_D����[,�c���<I��xț���9��D�'�t6M?����) 2LHDN�	ReN1�S�M20���$�r�4:˛��O��-R�iZ���O�����Vh�ur�G2�%:�`�%%D���'�ޓOH��?���?!�������!f��Ux��˼^������?a/O�n�>��������Il�c�'�}5�W(�#4�ҝ��$�E}2�'�2�|ʟ�e�pOI6a�&���L�;z�5��[&!�F��C��?��i>���'u�M&��z�Ξ-yD�i`��޷<�ڼ+���P�Iɟ�I�b>��'�~6-�zZPM`U(��Eߖ�a�9	2��E�<i��i��O���'Y�N����K�]Q�P��+'F/B�'T�jt�ii��9��H�O��++�p@ͅ� e*�&�� �������O<�d�O��d�O����|�2&�
;e0xK����8$�2�K�
3��dהokB�'jR���',�7=�T2%��T�Ԅ��_�A��2�e�O���-��IF�Iq6�l��q��� x-1�J�,l�� ��m�h�W�3�A��Wy�O]���%/�v����-�D��⎪#"��'���'7�I��M��g���?���?�!R-��lѡH<0uBB.��'���?����.A���L:yռ����1����'�9�R�Kc����$՟���'�
x�a�Ɗ,+�|���CC�(Y��'�r�'E��'��>I���h�!Z�
$@ !J'Ob.(�ɰ�MCa��?��&˛&�4��{�L�fA1 C�4M��1O��d�O" nZ�<�zToZ}~"Ќ&�`�(eՒ$��O-��ه���/E�SE�|�Q���̟�	ȟ������!�J����jP��+1�����$GSy��k�L�Yפ�O����Oj�����_�F�,�:Ʈ�f��q���B<eh��'��'�O1�jx���\=S$�a)�8Z��,����~�K����YVB�$bj�x�	ey2KR<���Td��7���R��B�s�B�'vr�'J�O$�I��M�L���?9�(]1R0�I
$�JRzr\����<��i��OP��'��'��Ά���{c�+�8�#��!{�X���iP�	/�[�1�O�q�����MΤ��K����P5b��d�O���O~���O��$>�Ӧ@s�UQAfA�B8p���p��`�	՟��	�M#�@�|����F�|��_�=D�Ь�xb��ïN��O�0lZ(�Mϧs�.��4�����6� J�a�iښv"0�DϜgN؈pf��?�'"���<�'�?y��?�򏙖7�����m�
G�|�n�(�?�����D즙�&C�ԟh������O�L��Q!U�bSJy���>*����O2��'��7�ɦuXM<�O� �c�oٌ\B8t[�]�!Yx�J��F��t��C2��4��a���nB�O8ѳ.P�!�.f�ǃfqP�$�O����Oh��	�<a�iۂ��D��%q��D��y÷N'^Ir�'�x63�	=��d�ܦ5g�Щ x2���A&U>� �_�M{5�i���ˁ�i ���!�2��F�OA�eЄ��H��>X���Aa4�ϓ����O��D�O����O��d�|2rOM�1Z�����
a�<���F�(��6g��]�R�'����t�'��6=��q�RKX5	�P�K�{��C�'������4@`���O2|����iC��+4O8�8U�ݜb��i�@��	�$ӌ	5��y�����O���|B�d~9�c2Z=� ���),�:�j���?9���?a+O��m�-����ڟ�I�E�d@���8ؤ ���F0@I�?qvY������ K<��0U��<U+F�k����i~�V�$�b�T\�͘O�f�	�MzҬ&b���3���VbY�V%Հ�"�'B�'z���4b�F�s�X=�G�ޤ�៼�ݴy�����?9f�i,�O�I�m����D��/F"��B�^
r����O��$�������˦m�'�%  nE�?y#�`>��r���!R���yw��\�'��i>Y��˟��������o��H����\e	���)Ȯܕ' �6�۹ �ʓ�?YJ~��;��ʃ��.Uz�&�+<g���Q������)K<�|2Q E-6u0�a�r�fU��ϧ��kPg�l~�ЋO$*����Y<�'!�� t��@j&f�:4�����H�������I����i>��'��6M��a��3a�a�$ڬ��G��&t�d�$��Q�?Y�]�;�4��ieb��B�\}A"�³:���c�D8�v���Cg�B���Gr�S���:����U֜{ +Z�@���S�Ns�<�����	럠�����Z&✕���ف��v���P�̞�?����?e�iD(г\��ش���Z�Iq�X�`��L�c%^����0�x2�j�)lz>�
P͈覱�'�E�s�$H'L�{�ق�x1#H�(=�i�	�G^�'9�i>��ɟ�͓DI%`��=Ev�@�<a ����֟��'�$7M>���d�O���|B�����8�#Վ*WF�V*}~r	�>�B�i\7-Gd�)����&6H:s�źS&��tI�4nn�m��+Q��tP���W����f�|�M�>�Z���E�)7V�iC�F�8��'�' ��tP�\�4��%3#�͒%4��K��6��q���2��香�?��[�xjߴn+�y�7
�_?�1xA�*u�飲i�D7 tT6�2?�'��P>���6�d.�"�,pcP�S�h$�C�ߛ�y�X�X�Iڟt����������O�� �n�:=�|�G��4Ir$$b�X$ٵ��O��d�O��������9w�`*�$S�=�V-�a�
)1��	ޟ�K<�|��ך�M#�'��y˷��	W��T�5��Y��'�
�Pd��lC��|2T��S����B�(Q؂/�:�h��e�ӟ���ן���jy�CiӞ���OR�Dh��z�d�-MN�P� tG�@�F&�	���d�O� ��I���Y�6�y�#��{�I)㈹aaΈw��b>�i1�'��4�I�NSJM�vmT{z���ǨlrT��	۟$�������w�O���N>���)lVX��$*�D���`Ӣ	���O��d�ۦ��?ͻ)j:Dɴ#D�Sv69r�n
��"M̓l9�v�nӌ�o�h30�l�[~2��9t0�m�S�(����ba��*��ey�oB	 j���w�|�_���͟�����@��韴3��	g��!-�?0.T��F]ty��l�nE����O���>����t�'��%c����UN����]�r��<!���M��|J~��K�v�Ԡ9�k�m�Xh Ā�9 t�����U~�9i����+��'k�ɶ5�<����W����L+'���������l�i>=�'�P6m�pO��D+im|�p�O�~����3��Ȧ��?��S����ܦp�4=�>�y����y��1z��E��t����Mk�OF�b���
����w|Y#jL�.����ś5�T��'���'B�'F�'o��:U�>_�2=�w��	3K�q����OT�D�O��m��=�����L�ܴ��[��}��#��LXi� ֆK��e���x��'7�O�8��Ƿii�I�F��A�$K�)n2�X�b O0#�o�O��&�I�	Qy�O1��'u��^���4ժBDԄ�0l/!�B�'��I��M�B
�?���?9.��(��ԛ<��zGS!�X��V��8�O����OH�O�S!z1r��b@UFǺ\�����`���&Wb��u`�L,?ͧ+������X��RT�S�3�Ș����9z���?���?q�Ş��D�צ��EjR5���Y�'kU|}#�&��4�$��'ؘ7�:��$��D�O9`O��Q����"Ş*g��f�O����8z673?�"h��wc���8�d*C,J�+@j�#=ʌA5k��y�R�����h����`�Iğ<�O&�Xf��|�;�U���Y�dx�l@��@�O:�$�O����צ�ݻ0y��(��]C��cE��X�J���蟤$�b>9����i�S�? ��8�h�$C��ե�@����q7O�Lr2��?Y�*�$�<ͧ�?���O�$<S+I
'��5���?���?)����_���H5EXyR�'۬܉PM�#Xؘ�9��� �2���F}Rce�p4�IM�I�s�2 �`���x:
6r��7:r�Ǐ��[�,��H~�o�O2���\(ڂ噱G���WA�y�`���?���?����h�~��V6JV�XQ"Ȃ�Ne� k׭
�x����Q�������I��M���w���0��!-�J1:�N'N�JY@�'s:6-�韠oZ.21f�m�I~�N�@e��NV�(uI�|�P�Zpϝ�GB�js�|"_��I�`�	��,�	˟��6D<df�ЁP��#G�&�H�Nzy�h�\H�$i�O��d�O꒟��&ąP�ڇ�(��T{�|��'4<6���%�b>���� 'ҬS��V�pP�YڲNE�CNɱ���hy"i�60��	+��'4�	 u*�z����ln�a��LA|NLI�	�L��ٟ��i>}�',
6�E2X�^�$)B�����%8¨�K��R�./�����	�?q�Z�����3ݴ/'��	e��&� Z�J�k �Hf�V��M+�O�1 ����:����w�N��E'�,aSJ�D�TvPM�'u��'X��'���'o��Y��2`����Ԩ~��"�O4���O��oZ O�@�����4��J�
�K���n��sd���3��D�|B�'˛�O�$�0жi��I$c1��Cm�L\�ȃ"a[�b�䩃��\�<����|��wy�O��'��/�!2�=H�������=���'X��%�MS�����D�O�˧\��	*��plf| ����x�6��'���8����w��q%��H��P0�eY#]�Dq����IL��$k�|C��r���x~�O�|���q��'�Ƽ��KI��&n4�X��'�"�'R���ON�ɴ�M��)	�'-�J&��`g�#���<G�Xtk*O�m�`��fg����M;R�D�\d���G܆{���J�O�3��+a�l9�Fp� �\	�z�G����O2�ū��w��@rP�A�JC��О'��	�����ܟ��I�����@��$ �u2���%@C�x���)4h��h�6M.E� ���O�$)�9O��nz�Ah�P�`2ȝb#���\���,�M�i��O1�x9�&|�2扒,;�P"���-�(3E�0!\0�	$e��P�'D�'�������'�06n�|�<uH"m�%όEi1�'���'��X��[�wx�@��㟼�Il�&�3�Ölf��d��N8���?�qX��	۴m<��b2��I7
(=ٗŔ*89 |Jq�<% ��(U�r$�f� y^~b>M���'J~<�	�@4�k��O�VT(F`X�5n8�I��X�	ʟ\�I\�OI"�=a�Y��N����b啢)�48�I
�Mk�����ަ��?�;:k@�A�V:>���E%LR��Û�!r�2`m��|c�1l�P~��?J�� ��>� �SA	?5��\�B_�kv�|�X��Sş8�������Xɷ��$7D4��E���T���UZyrlh�j�	���O����O����@b��
K�>&�A�vE�+�Z��'��6�F���N<�|� A��>���覣N�w+,�Ps(Q�APH�"�kB~��P�&�����5��'��	�|�F�cW��?
@:b�B�^�:a����	��T�i>��'�.6� �D���d��3t�S &X�\�&ē���e`���5�?��^����ঝ��41LHi{�,׾p�V�2⍥<�z�A���M#�O��$�O�j��$FF6S|�%0�JM1ܔ�y2ēuNj%��[��DS ό�1wT��&'Q�bTԅpQIJ?��H��Ɩaf:����P!��{Əda�I���8Q�:��]�{˔��'E�(gL����"O��̓Ģ͏(�FX�!#؇f�0�!e�S"F0�(�>ڭȇ��L@��E�ȁ4�6�#� ߍr�`a�V4jhR�y! D�@��ղ�,�+_5�m���x���h[&}�ZlR��	q�d�:�A�\��5r7/�!K�Ͱ��55D@���&� H�x�a�7��A��������I�Γ"`���	Ο��O���Op�W
�, *�dZ$��sn�t%�H�$�
�ꃚ���'B�'�J�j��ٴ@s85 ���5Ď![#�h��I�}�R���O��O��|����}쾙cq�	�N�Hl2&������J�2d��Y���t��ǟ����h���-0jt	��T�d�֍X�D�[hK�;c5�ʓ�?1���?�J>9��?Anv�������Y�	1C�A,��ɘ0��d~�'��'x"�'���'�Hk7�X�~��p�L�9-�����wӎ���OP�:���OR����mت i!�i2���qge�,�kU�X�&(f\��O����O��Ģ<���ߥ���ğă�'��E��%��J���#޼�M�����?��-����{�菧v-�� &��FB�����MS��?9+O���ǎ{�4�'t"�O�ڱ��,�k?�Y�KP
8��u�-��Or���[ݚ㟐�'6鄴�kQ�
 S�e��*�Lm�Py��Z�-�:7-�O��D�O@���g}Zc9��A�M*C�T!d�ڴ�?A��q[��A�����'�q�rQ�n	�,Y�D�#8�r�(w�i�Ah��v����O���&��'q�I�v[pX9�U=b�P��1�,zNM��4#@Z�FxR�i�O������Z�ɗ��r��ţG��M�I����	�p�
0��O ʓ�?y�'�Z�8'�T�So2aQ���~��|ݴkz`�'��aas�'(�ڟd�I֘͟�nRP�$�ڳB`*��إa>7��O��B�L}"Q�,�Ij�i���� -�.h�3ND*&�8ЁϿ>A1J����?Q��?�-O�T� (�S�/_9S+`q� B�\�P�'��81���JyR�'A�'�B�'��h`L�H���`��
S�`��FP����/�yB�'n��'H�	1���OV���q��)'�0j��ś�6A��4���O��O*���O�5�Gj���ȕ)�!�����ıT�T����>I���?����$З3~��O�)Ɍ{U�qs�,��H��׈ޟ�M������?���44x���@��,�'Dq)�BH,h,�%�Ф��L%"۴�?q���$$�h��O�R�'9�ħL
 ��iQ$C�H4l|k��dy|Oj���O&@)tG$��^�s ٲx^Rm����?t-n� dȒ��%�'���bf����OP����p�ԧ5&F�p�x���=`��0IV�@�M���?�����'�q��%��h�;PP��ؖa� Q��i�2�qljӆ�d�O���@�'��I�D�h����5p��(�m��-�J�4G&H���i�N��'+���$v0���K�?��E��Ł�Z�>	lɟ`����X��NՕ����<���~R��l`��΃K�������'�P ��|��'���'.h@�h[dx�%�ҍ+$�(��}� �L6)W*��'��I��ؔ'����m��i�P8w�U���[���}���%�d�	ğ���Uy��(.!��;�	;'��8 e
@8q���l(��Ob�D9���<��gʁ�R�R|ր�;6��X��n����'��'��[����N�����L{p�C��98	jl�4	������ON�3���<�'�?`�C�LhRp�0׉~\ ����F�J��IƟ,�IӟP�'(�3Q�+�	d�f� t��ӌ��h	B(Nyn�ܟ�'�������'`�{�4(i�f�a�1�%��i�0�m�����`y��K�k����$��k����P�MªOAڙ[���e��'��	�|�Ih�s�֝- �j8I��Οc�q�v��D��?�/�6�?����?����-O�NƴZ��6>cJP�d��>	���'5�	��f#<%>�؄�D	_s\��䯊�9r����`ӰYA���O���O��럎�S����h��W	�?w���*�iV�J���5 DDx����%�h��ֈ2�~� a�.+���oZ���˟�A�APyʟt�'�����#N� �RQ���	j"i��@$r˱���d���-6u5������9f343�$tӼ��֏�p�(��}��m�<�`�K.bX
$�qے7肍���x�	ژ'��_���	�I��M�g�̩*�,H����]����#ΚDy��'"�d�O��ɰ4�J�������<a�GU?6��6튶c ��ޟ��Iڟ�'H:�j��n>�I�b��?��	����J�bA2��>���?�L>�)O��O �Y�J�9�|�,��HQ�R}r�'���'\����HL|�F��/-I>�c�C�1Ll䝢`CK�c9���'n�Y���F�D�'?�'T���@ѹ#r��ŏ?��l����'.�H����ȟ����?�l"�X��B\Y����uc��}[JO���Oz��1��4�1O��9>[r`���#4<�G�]�/ 6M�<�ѢZ�F�f�~Z��*Ӟ�8��Dx���@�I2�b�qӖʓJgJ`���%��O��M+��޶1�I�E�R[����a�ަ�@�"P�t������	�?���޶,�H%Q2�u��s�"M
)oq���T�?�)�'EI*`���ĬF���3�H
q5H��W�i�r�'�"�H:��)I�\E�G!�2IX' Ѱ9������:��'�>�-3�	�O����O����c��D6Bx'�q��T��&����I�T���K<ͧ�?�O>��J�����MQ�ac�ܩ��R��ɖ	���	^��şԖ'��-��3��@`b'�;a���#Q;%~^�3�_���Iʟ��?A��?����g��Ae���q:~�zW(܂!*����`~R�'g��'��ɇ��J�O�q{e�K�vNr��e.ǼI�LLٴ����O���?���?��T�<����?��Yci�	L�����H��z���'�����'�B_�13�����OklA=�P`���Ѻ���w'�r~�v�'��I�����џP9�y����y?��P��T<H",¡R�Ȁ�pM�ئ��	ğ@�'��tc�F�~����?��'HYZhh6D�`�҅lW�k�s�T������2L�:��Iy򍒬����?U<�c��>T�����K�l��W�����/�M��?-�M���#_�i��v	��h��H�u��YT�$s%{�,��On�;O����<!����a�܈��j��>�m	���M��LЛt��6�'S"�'a���>�*O ��ɕv�^�
t�W	�(����:тt��&�,���6W�s�]<l��nM��l��iAR�';��d���D�O��	�\���#�/_�}z�)�dXJ득��� ��i>���۟��ɾ��b�B�^����7��7O���ߴ�?)%�Y�%��	OyB�'X�Iϟ��N�\��PǑ���;�ƌ9+���X�̓�?A���?���?a+O�tk��Ẍ́e QfC�ڸ�3e�<V�VU�'�����'��'�"n�&��g.
����ɋN�-��'q��'�dA3�'YW�|�uo�;���8�ČK�H߿ꤴ��鈭�MS/O<�ħ<Y��?���(����t��G�Z*Yfl���~:�`�i���'��' � ��⯟��U�? �H�q�I
%L�\�WO$0���(e�iU�U���	�P�ɴ\����Y��*��a ��A7T5��JB�I8���'�"X��qJ�4��I�O��D��T4*��[�es��h�h�4"�r�е��M}��'���'�����'���eE���FG����6��+�!��@��n�`y�)�8U26��O���O^���F}ZwN�-K�OߞM]:M�uU��3�4�?���N�lΓ�?A.O �>��b��!w�}�'���@�\p3ƆjӾl�L���������?aR�O��G�VeB�,1fd
 *��S�@��@�i���b�O ˓��O���[�r���T>.��ܪ�/C�e#t6-�O��d�O�X�l[N}�^���	r?a .PHxjt��.Ҍ7+��*�i�Ǧ&��A�.~���?������S�8@���8̰h	Ë��Mc�^HX]�0S���'��P���i��m�N��؊��	!���� &�>�E	E�<���?���?q���$�>"P�A/��� H�f��8�Z�I1b�E���0��z����4��VtL����A�l��⁋��AR�q��'+�'�RT����mѣ����*��`�`�ԽȜYsw�0����O,��8���O.���/���GURm@�I�%-�};�+�5g���'�B�'��_�HJ��B�ħVFL2F��ifH �����6|Ȳ1�i�"�|r�'����<�y��>��'�}]����Ҧ)! LF��Y����t�'��i9���O��)�%��=:�	�#0 Y����2=��'��I��)��q��$���'J�>��3�
O�4�@`j�-G	��n�gyrE�S{j7��n�D�'�4�6?9&k��0�Xs��	}��"����I˟ps�����&�$�}�dD9'��5D�?d�4���RȦ�ѣ��M���?����֘xB�''��a�͋#Z1�����/�|�$�`Ӣm��O��O>��"/ ��Ӄ�*����cq��ܴ�?	���?A��D�h��'��'��$��y�@��f��� �öE�2,��|� ���yʟ:�D�O��D^�gK��a����S��\ CS"e��d�96qz|�>����K�W1,(ՈX�,[����l�_}���/�y�U��������VyR��A�H���)>s ժ�Sy�t�4��O0��&�$�O2��M7!z�����4�6y�g�ԗ}C
A �'��O&���O��/l	i31��%�`B�*&�V8��ӄ;;��՟x"�'f�'M2�'��=@��'LL(�Ƿ6������I�\���K�>9���?����$�_�5%>�a���l���Hpg�!��x2��˕�M{����?q��?�~�s����	���9(����cL��'�D� �J7��O����<q!�'߉OCb�O�������1��U+F-�$'�2�4H4��O���̼K��>�D�?=�b-S�(ntJ�$ܺM>� �jpӮ�Z�Li*װi��'�?a�����D4�H�A��?����f�ߔ��6��O*��J1_��d0�$6�S0�v��Ɵ�(��@ge�6�ZtP�oZ� �	ٟ����'�v,��*/=�(�`�ϣ�8��i�P�۵5OҒO\�?��I�hs�!���ۊ3F�l pL 8"Vq�4�?Q��?���*@�O����� pDL���4����۩O���� fӎ�O�-��HAL��ڟ��֟��[
<�4�x���'�~�X'h���Mk�e�bp9��x��'�b�|Zc��CE��zC ��%�[<2� �O��*�>O�ʓ�?����'2�ƴD�Ռ'�,I�,Hen�iЦ�r�}��'i�'��'E��F(_�!����S��>+fÆ
{�b\���	ܟ���qy�
A1��擌SP���ҷ�����C�%�2��?	����?�x�j5�+(P� DO$��lI;oX5	_�0�I˟(�	`y"��?��( I�/67��qm	�?Z��E����D{�':�D�'�����R��w"݋vH��U�qӬ�D�OLʓu���[�����'�\c `�gO�l�8\{F�5X^�Lڈ}r�'������'Q>04�X�F���{RjؠU
BI��bgӤ�����'�inv�'�?��'
����&5�\X�@�	cJ�8$�E�=�>��?����?�N>�~�F*�	=��y�@e)]��XǦ�ň���������?ɗ'�S�r��8G#�99'ѣ��J���ߴ����[_�S�OEr�\&ac�0$N.c�����#$��7��O��D�O8�R�d�w}2^>q�	؟��ë�3mo HPVn�+3~� I l���'�aQ�yr�'�R�'δ�7E�f8�%k"Ӵe�t�wӢ�)�@˓��ٟ�&�Hіi,7���Q�/� UV��1� ���ޯ;��UI���$������IXy&L�A�9�sM��U��4���nRtI��>A,Of���<I���?��,�*e�0*�W�¹���>Y�.�@�,��⟜��П��'b���.q>A���;E� U��h?��i�e�nӊʓ�?�-O����O����k���(m����`����� �%5��oZ՟��iyo�����';�mط��~��*:J�HA������t�e��iHbQ���	Ɵ$��l_6�K�䙁x��$�Q�=�~ à5!����'��W� R"�@��)�O2�����#@� q�j�J�/��}�����G�m}B�'�b�'̈́�i˟�IJ2'��#�&	sP&�ܰa���妝�'�.��ak�,���O$���aէu� Bl(���_�<%�b&q%�M���i���'ڔ��'�b^���}�U���%��i�`TP���[��ۦQ��V��M���?a��ʦ]�З'���ѫ�x���۲��� �ȝc�`kӨ`i�8Op��<��T�'�
�£�A"Rr��F�
=!����Hl�$�$�O���,|�u'�>�*O����� A�f��V�:�3��'�"i�n����<�KM�<�O�R�'��	X�$Q��:B�->r6X�O�ag���'�^t�E(�>Y.O,��<Q��sv)O=s�����"a,^��bGY}�JU�y��':�'���'+�I*}b9� ���~�S&՟~ hL�1������<������O��d�O����)��u��4SK��y�L��!
.���O �$B�AdR6���$��=��O�O��,���A�L���J�(nT�EK�'�<�s�m�;��M��Z7`1l)��{���0��ՠg��k����M@���Y3�jZ
t�AP�JȂp����7m�@ff	�C��|����vǾ������kr��'LŘD�`ʴj�|���p�w�|�1�F4��� O���0��fȖ�6YD#`(J�l9K���!\���� �ʬ&�T���i, ��5wb�?閯U+X�@dr��N��8&�I�?��?�*T�㘧�Т� �  �N��ӡ*F��!F<}2L{���O���"$C �x�"�(�<R�ҝ�O��E*�O��9�)1���9O�����#j�`d�I�6X�1Oh��3<O,��D�V��,�W)P?$�^L	�'KT#=I�OZ�s j�c"nʶR:")��֖uy�Iן��I�F*� ������I��iޑb��|��L�KY6(������P#]���N��[\�c>�O"��o:֫��)Z.�cH��d��`��>Q���t�L�>�O�(0��Z���Ӷ�O7Vz�Aiq�O��m���i>AG{Re�7�p�ӗ���E��$��A[	�yR��}�7N۰E'�D�V#S� � �'t�#=�OX��3f�(��$�X�:�*��W�9[1�AaA��C߈��	���	П��Xw���'��k���QD��;/P�hE:F�Ĵ�v)�*�����H�F_���$ȁ2ξLY�	݄qHh9���.�� q
F�U�͐AɎ"N��䆏U඄� s��[aiݛ!;0��W�'
r�IP��r�2Q�b��c����c�Dr�:�ȓ=�xUIg��%g¥�	��16�e�<�2V���'1�XB�El���d�O���R�X�=9��W�T�	e2)(K�O�����V���Od擆	V�1Jq��o�I�oS�i8Ag�5����@�̞d� ��z��k�-�$Řp^=S��
�}�&$�"�.#��x�lճ�?���?A��0�d��ׄL#���A2�P�L�*+OP��*�)§Dk��Y�iUa�fs ��H-����;�����?���S��0�q����y��)�'D��(k���<:N�R�cɏ:��ȓw6D�1F��?�z&B��sjͅ�8�� �����V����!��:<�4�g��[�b$��L��o�!�ĕ@`$�
��	+y�j��e.��!��X�l h�]	����2��6�!���2*����ţd��(7'�!�A�}n�a4~-j���/:$�!�evИ*����]����.x�!��"F\�s��~�<ui�P&�!��e+�dy3�4-��0�CC�!�$Fb��`#gW S�I�1#�2y�!��fb�H#�D�&3��k�ۚZv!�dG&M
�A��
V���ic�惙4v!�
��B�p�Փ}���B����z�!�D�J	�D�A` w�v�To@��!�d�$\L��'�6+�<ˁo�9U!��1sH)@� O)���
���xQ!�$�+����C=�|i���!�!򄏋"���OV�4���&�X�!��!DD�1Iέi�b��D���p�!�D�4n�8�"�K���0����a�!�D�� /������c��liV�I�!����y`�R*�vla��	w�!�d/}�4U3E��Y��LA� @�!�#a84��@��xpp`C̗f�!��5)�2%K��M8j���boY�#�!��J����ZEL\��l�sҧe�!�� ��� �Z44=� 偞,�,8
�"OX��BIv�m�4�ɷZn��R�"O,��b��b��#��Jl�y�"O|����R�hiI;q�O9���sc"O�}�,ˀ$E����K~�Y�"Oh(�4��7#yz1��>`x�-9a"O�1���>�EZ���6f
��"OD���kW�GI�h��C���$	�"O�9/�;���6āDm�L�"O(��j��\�$�Z ��[Jl1 "O�qc��r����!ڷV��� "O6��V�D�.k�#�Q}�zhg"Ot���LP�RKN}a���	�x��"Oyq�0�����G�	ʞԈ"O�I��f��,y�	�	X+Z�D��B"O:��Fo��.�
�X�ɂ-��9Jw"ORi��oP�`�H�s�Ŋ+�T8"OZd{�������W*�>���!d"O�A
�#�j|��V�y	3"O0�� ��Zq�U����I=�T;D"O.4�`�ew6���- ?>�"O\ܱf�5Y1V��j�:H)��*E"Oj �S%)WԐ`��P�!����O&��TO�O���䃄rzP��O�.�Ƞ�	�'
�\��hY=7��#�k�({>ൢ$�ʧn��O8�}������t��4U�Աt�]7a���ȓKF]Y�dK!"�P�5e��!�
�ɗqD��Q
�t���ȕ�Y��s�1)�J݇�4_�0�*O�I��D0s�(���Q!����"Or|(�� kP1�݈qN`�@V��.���D����&M�:���8��(z��ɀ�y�Ҋyn6`ˑ���A���`��%l�:��g�:�g?�v#�j�P��M�z��u�q�Rj�<A�� �})V�#p�
�U�P��t$��<�b?/a}���,z�N�H��EpNXXe�U�y2���H\dff�?D�@2���yB�R�Ob29[��YwǠ)�Y�U�ȓE����̑>:����b�ҵ��%��r�x�a�6�Vę�
�1y�=�ȓ_�F�c��jR����ჺ:��h��YJ$�v�]�+���e�A5b����J�7*�3b�Y��"�P@�ȓm5%Q�'��AG�'.����ȓ?X�X�DA�5��ei��D�76�ȓ(��A��L�HG��dl;�����f ���/�Q�d�w%E�zf���P�BT��"�g1̸p��J�7�J��Or�1a�*lO����gÍ#���s��	�8��d�'�.9�V�i�P�!�t���G����q
�'x��W�% :��C7�X������$��x=�"}�#I�L��L(+�pA��お�k�<'Eո�nl�wM�	N��%g?��c½���h���X�hR4{�f�bQ�.f��e�B"O Q:��Q;���g��\�܌jp�>I��:�=���ƌod�a�� ߅H]ңFVK�<9�A��6�vUC�Jv��9�� \�<���@� ��0IFOR?h��PgmQW�<Qt ��>�\���[=��9�͌T�<)���?e`�C�n��(k�T���R�<��(M�?yl���)B���R�ER�<Q�+5���''�g�=X���P�<7�H$u�Xx��k��=�T�#���g�<٠k�p�"��dO�H���0S+�x�<���9EB����ȺfR47��u�<� �XYU�̞(�<�J%����(Bd"O���o�f�Y�j �s�"O���+�D$<t��N;ZT�m�"O��ac�1q�䔳A(�sAʉ��"O�@z�d�yX4�`�11࠻"ObЪ���%��4��8*��4"O���	?uf�Hp������'<
5��V��QE	"]
n�+�φ�R��q�'D�����7E�.�#�m�/Bg陵�#�}3�tRA/�']?�|	f�D*L�R���E�#4���ȓ]�j�`U�Q�+�Lb�x�D`ٱ�F.%�"~ΓU�h�`-ٕA)�ē�/��v_�i�ȓf�@(� �˦/�`H�r��1k���N �m�66�O�I���H�(@4 )��@
I$`��'J���I&Z����7@6�����%̊A��F"(�!�D�8s�8QꉳM���de݉) �O X[sj Y��ͻ��	E�z s��f2��T�ȧ@�!�$�I�R���6x��pC�V.F2��P'�>�M��B=��h�͸|Z���Ś<�~���o� ���:�a}2�H�1�z���njPB��f9��s����#BG�(����\�����۫n��a�UH�A�D�B��xRf�D��H���j$�!c&��'a^�j
pҠ�d� �%h"�����yh��A�JEYH���YhƌG�MӰ@O�l����KM���&	�0�|�����Á�ïH�k��Gm�@����Q�R�Z�L���!��,�6��U%%l��EI�Ʌ��r���`j�d%Zj��(�SRǑI1ZKA8d�ڄ����4@�K��=�&mk�j�%"ȭ��B�sbX �f6(�X ��:N{�{�%�&�H�Į��O��,8�,Ɋ�HOV���O��0�m �DÇ"��A�� ��'2/�����
�� Jң��Y�X��
v~m��.Y"*	�U��h�mڏi��i�IU;�aPƫq���ئ�s�)�g�+,��#�Y�t~p�� D�`@��O+x�
Po�c�d	/bD��:�h�H�g�!'st(�$�|���d�K<A�lp��a�6a~�G��	�Xb� F/2�(5�Q�
�$���O�	nl6�U�X%f0(�bľ��5fӵ�ʱ� ��5r����'8�^��'�O�1�2���OQR�ʒZ�}
	�2"O��
R�S8fh�D��2�qX6��NK�YS���54J!�8<� y@Hӿ����$��b�O������J
�"���=�uoN�_�x��{��9OX���T�+�(�
Ңυ*٦�1Đ�P��U��ا����3kYo�h)'N�d�8,1�5O�dr�.���p>����&Aj.p�����!Y�U�N���l���kz*�n�\3
�kO|�ȟ�DĬ�Th��+=� �{��~��NQ3v�x�l��U��u�ݣWy��(7B��N�y�U-����<x��Z�(�3�I�Qb�i�
üM�gӮq��܈OÂN�Q�Щ4�˔9�0��Gޭ(p4-�e�O�h�qkԋi��Ѻ����>2b��'SV���+\EyBN�#^MGy�J��	Ò�E���bJ֘�&b��~���Z]�Q���Q�yH!Fߤ�ēm*���O@~����/��UV�Q�v L�Й'J�����OE8��&�6~8�j�-=09�\�A�T�(�Ni�k�@�I�,��I�?�;B�е:5�v5 �t�ذI�iF�'��P"�M�Z)8����xBz�j�$ήVHΓ�`��%��y̓1;���#�ǉV���h���8���b��O�>�8&-��E�� ��A@�'��	� リ#R�[���! k��Z�N�����w2��P�;�b��'�l��' ��r�٢��;���S��I��m�j�S7/�_D���b���}�'a� �o�5k�y�D�˖7�ʨ��O*-�&�Ƈ/�e&�(U~�(��%��.�J��5�H:1���Q��	��X�ߓZ;���@��1MjN�:pƎ9�"���kڿJ$�Ѡ^�����ξI���id@��3����`qH�e[�)2��5@��@ �4�O@bu@�����[�焔�>�
��vU��s��5>�Hx雾Pa��?��wJ�#(t�	E��j�t�:�o�,2�n�Ѥl�$Y��x�N��P�џ��%O��Ud�H4��-FB�X'�ܙ&c�ɱBK��6�y!eEVL$�����hj�'2�d�c�Hڹf�jȲDG����'
��%`�>����g�n��M���G�(��k���������	�G��<y,�2��Abc40� -N�r* ��$��3�E#2NOR���D�2H�$<�'�F�I�l��BT�HR�'ɖM�JM�,��-��Fړ��%��'*zd�&�O��Y��[
U��jQ���x�'b�� ec���KR���?W&��R$@�(m�"�� i>���w]���D��4�O�b�������;��S�dC(i�N��!A���p<��L\�	��c���s-K*F5U���O�o��i�	=?��E�j_j(�2l�^��dK��A�'����K�iFh�.� ��M<IP
&!T1O�%
�
��XR���#i]�%{^��殇�{0:C�I+n��"AǱ�8]���6���pAh�g�S�-�~��L��l���"��C�Ɇ`8l�@r�H��Ȅ����!�(B�I;,�@�:��DvYB��ڗv}BC�I�@�����Q�f�z�����C�5�L���+��7O��������B�I$"V2m�v���Ʉ�Z�&C�I3	��ٰ�HU�s�|4�����VB�	GT�)b�'�!�" [�C��0��B�ɸ	v䁑�&T�i^N�[��O�`�C�ɤa����BH�|���c�M�U�B�I�;�z�JƇ
�=y�Z'�<W��B�	�<�D�u+X%p��ٔ�[4tC�I�}��{2��/6A����v >C�I�3��y���?J�J��޺o�C�I�|�d��g��i�
l�� ��,B�I�t��<T!7���y".[��6B䉯, ������+*)���JC�	�c@�8�%ܯW��l��.H�3�B䉛Kl����'�h�����&O^B��6}�M�R
jVr����0XLB�ɂpl!�$JǊ{����"dC�	�?1.-���֣Sg��Se�M�5�C�I06p�Ch�7[X<�rE^�7�VC�	B���䏼�� [5�q��B䉂��l*�"�z���X�_�B�	.Wbh�@�B��<Y!BxTB剟,d89zGQ3p4:D���E'2(!��L-�R�
q��{2� �C�-!�䘹ݸH�W��ܲ��&!�[N�xJ�)	~�v���ף�!�Ҫ�h�mͨ|�$Y�Γ�$�!�$[�NL���V�D׼|Q5��!�D�|TC`.��3HU�W�1'!�D[�V!��f1���W�!򤉴5}�!+"��9ON��äˡ�!��5^r8�q�'�7&r  B�/��چ�.����8Y2�C��z�	�g�$60�H8T��E�xC�I�eⰚ��AtΎ���Q#U�B�	�_��!&M��0J�i�ώ+�TC�ɨE
�q�3i��V8���>(j>C�	�h��)�B��N�(C�߯XCC�I9G;:(q�H@�>\�p�ܲ:9�B��CU$-�'��/m.1���N�tB�Ʌl�J�Fٿ5�,�Ѵ �3PTC�	)$w��"�!��# i^7��B��$uԄb�A��(�xb��U xC�I�{�L	 0&Rs�UX�l���VC�<'F$��ҳ!��%�Al�pHC��Xj��sଖ:9Q����٠��C��*jn�jq$�2~ikb�VvݢC�rq���m�W�X�a��c�C�	�UCd1S���b�NU��Λ9l�C� =\D��d�\u��6,T�D�C�����#��1Y�꓆^|C�ɒBC<p��2g�a[�լ`xC�I��Z�Kr'ʥEd)��bS�=�NC�ɐK�\p��@ \p��y
�B��B�)� �43�+םz(�3�̓�,?�E�e"O��W$	�v���`�D�v❻�"O0�e�Ŭd-�y��B��b���"O��Bw�U(Y�ؕh��R���:7"OQ��[�,�HW�
t��Z�"O�S#�\�x$�@�O��R��"OD:%��:���{$`U6O4@�4"O���w�B?C�����B��T"Ox��Ŵnv�-��O�}p�Q"O2��F<,Ld�9��(E�b){�"O�� �n�I
�́/l$�(�"O�������|
�$��jP#vf�a+7f`H<Q�Q�QD`�ۭA�<I�M�<a��+���$Q�fvX1)XO�<!�HѢO*��*R�	&!R �Jd�<aCl��a���sA�u��D����]�<i�#W�b)K4�V�~����E�\�<)���`��RQ$�CŸ�c���r�<I!���l�� �uy�{C�Yl�<!��$ǆ�z�b|*P˧G�r�<Y5i��S�b,������DW%�z�<�'�#����!YT )�@�M�<9t�R�R�B�c�����jPr���F�<A�ӊ\�J=��T=q-��� �w�<�`�{�BHX�ҹ~�pa+�/u�<�FlA֞�O[ �B����j�<Q�ʚ5�h	� ��=i0݁0�e�<�$A�c�p�	A޶HF��ӵe�h�<i��Q�f4�AX,2"�s��Nf�<�d���>)� �4u8�IdIBc�<a�e��M�.�2��?|:`R���`�<)�cRgk�ʣ-��3_H��� �g�<�T� G�4�0 �֎��*Ig�<�ъө+��K��If�t���Q]�<��-S>̴��n\>r|]� �]o�<�a���}�d��
�JPQrv@ G�<�mV�f($��c(�7)~ls��C�<��06�h��,�)#2ţ�#]i�<����G���c��	��1ӧN�M�<1#O��m��h�W�R���d�B�<a�E��^��!�Gƹ@�(Q�%!D��*�5�b�q���8��[WE=D�� ��:.�$��G?[��)&D�����'+��)׈��D����&D��
uj�o��.y*��#'7D��/K�R"8`ȡo�^@��.)D�t�E�ŝfTA�����].�e�wM'D�0����f��5�v#0]���j#D��spJ���lP�[z4���'D���s�ό*���GOO8�
�`d#D� 0��_�.�$�ӐL%.2��?D����6W�Z�C���phY�%=D��*����`�\-�����#����CB9D�ԙAn��$,�th���D 2��æ6D�B�B���(T���*e�9D��z��U�O�|چ�A� �
E��9D� ���	�XqP���#U�,�ڔb�7D��8���'U&|G��� ���C2�:D�X��Q�,\"c���0s�b7D�����U��ZÃF�Q���E4D�����ϖ.��A��:Ą��3D�ܑ劒~�l�LC7M�h�a�%D��C��մZ֬x�`͞�%�xt��B$D���D�G�@���'_��@�G!D�� xA��R�TVj5���"`��I�"O�Us�nm�8�dF�.t!�H�"O6��'KƥL6`�@�"�v�H�"O��;7eǍiP"E���U:�>A�g"O,�Q��TQ�E6M��A1@"O�B���4uӊ%r"��e� %*3"O^���?@��P"ӳw�z�R"O���S����r�(��`�Q�M!򄉻{j2�r�I)3�v�D�A
<ў���ɧS�@��2�T,K�)8����I�C�	+�x����H�<xBj� [�~C�Ɏ��CRbY);������ 4\C�Ʉ+��x6,���d���z�"C�5�|�.M=� @B�Ⱦb��;�"ORm�@��
GP����d'a&20�"O�9zu �1�qAF�57�	z�"O�)b�P¶�i�%K�A�ƅ�"O� (`�D�B����%C�9�:���"O�����W�D�c�ɱ;�pH�"O�H�����H)0��<*C"O�9��)�G��D�g
M��"O��a���6|��q�͗ 0@�au"O�1R��?��H#��(�Q�"O�4x�ɜw�2U	�)�&T�F])�"O���1�E�[�@ȳ�.����f"O��A3��):F�p��Wx.��3q"O��H�_bcX%"6Nи  �A"O�34�Y$�����:=�x�r"Od�r�-��<\�a��� �ڔȃ"O��7�~7xt�a��<����#"O<Ђ�ңw�d��R�Ź#i��� "Ol�H�h9\�`�¬iX���"O&�AB;l��y ֦TZ��`"O6i��H�OSܨ�G%�|5.�Cu"O�`��"[p�9VC��"�5�'"O����+�W�`�bF�+@���""O4���ɧ ^��wAA�4��"O0�"V��wZ���R@M�*֨�XS"O�9��2ZY0]j��-tD��"O�0F-�?��)2Ə��P|�7"O�$9B�N�j"�=���E�����"O ��u偦9�RÍ[��b�)�"OU�`*T�!/�h��S� ���ʁ"O��;���;D+�,���2\;�h��"Ov4��	�z�$Hb7
T�FN`�9"O�XK1j/J-Z6iۅf٨� #"O
���X��� ���T��3&"OѺB@�{lw�R������8���k�Y3�$�-y�q�u��,)z�C��'I�|��R�%"v�z��D4TU�C䉰1�~�T�]$�p���-W-,���.���)��!��H��2׊�
Q���Z_�C�(Pb�A U�FTLt��(х2�fC�ɍ����4.0���\�A*C�\�1�-�2,�VpD��-i�B䉣D��m��K855^��1� 9 �B�	�L٨��"�[a�!���bY�B�I8�l9���43k�BD�w%�B�I�C4 ���̍/�i�j͸2��C�I7��T��e*��z���]�C�	$d��Q�n���%I.TzC�ɪ<�: ��[�>�SbbE>^ZC�	�\l:�Jdf�P�FtP��A���C䉧%�LUY�b�^sz�hR)��C�)� 
�!��K�V@��`[��[g"O4�3�i�.��!��̎2�<��"O�1�2����]�s�ە[�N���"O6H��++丩�c�To0��K�"O�	�$L�(IU�1�H�;(Ű$"O9��)�(�h�ьB8	��F"O(((po�'��H����n�,rp"O<t�h_�#����k��8�`��"OTH��+N�ukr$����@ؤ�`�"O����J�9yS�y�c�W�\��"Oxp��ɗ#6�a
��w㲉���#D��"���(3���5�D!�F���"D�XJ&`�*385*$� /x��bej?D�@ZTI����:f)���(��A<D���$;����_�8�;a�9D������r{����!'dwJ���k8D������'䬘v)Q�@o& ��7D��������8�Ȑ�T�H)�Vh3D��:�W�Ar9�h�"l�ca"3D�  �`��sd�8$���{Nyt$2D�$j!o�BUܹ#1�͚T2)�1D�(�4�@�ᄐ>!��`�Tm*D���C��^{. &Y�̍0U�&D�0Ѣ�4��:'뇟��a�Vc"D�h�H�@�T(��D�.ds2�;D��-�$O��� S�Ц+�<�[�;D��iQeU�x:�
�o��V&"����9D���A�c.� c�$�Uk�6D�4x$n_12�<
cD�́*�:D��)��	(D�¹�P�Jez���a�+D�`Unev��Q��J<HШ��(D��@�D1^�tE@����T))D���.V+}����CeE���t')D�\���ڞ'4��q/Ņw���cu-;D��S@�T<��(�@�"7�J��;D��� ��88I�������P�5D��2�,�TTL	����bd.Aj�4D���nU:�`� �JM�r���!-=D�0z�N�&Qjx!{UG9'�Ƞ37�9D���� 0�Vmȳ	x�����5D�tR�o��U�lk��/^�E�q�4D�ة�L'�N�QgpWsY�@q�'�Z��A�C	#	��s��>n*@i�'��P/X![��!�" ��O/>,�'i�i������R�Ep���!�'ќ�����
A��qI�Jȼ� i
�'�2G�M%)3�pA��	�}�,9@
�'$�y�T�v��a �k�9%����	�'D�D��-L=�6dZ�$@�K	�'��M�����`��;��G��$���'����&B�.��s��#����'�¬�R���_�^�ċ�/9w�40�'�t�B$��):2��xec�"0���	�''���'�NGt�p�*���}b	�'�P��Q�l?T	2��;�,��'Ԟ!@תUD��9$+�)er�)�'���v�[��p`A&����Ѡ
�'p*�چ���Ix�������Uj�'XXpwAZM�p�ҰH�4{�'p�sC�@]�>L��D�������'��yYv���o.����( ��
�'�~Y#!(�y��-Y2�	3m���	�'z� c/�@3>qc��)]��k	�'�Vu��@*1��C��7��	��� ��ϝ6}�h��Z�'X��"O\���&�,ڢ]�C�����@F"O4X� �.
@��6�?�~��B"O�y���X�`+�-zw�A�"O��enYg{n�3p܉I`P�"E"On�1b��.���(��H�f�7"OHI�`k�3�8T�"�I8f-�j "OzJk˞d]0WC** �"Or�2�G?`���B��-S��}s�"O�-�ׄ�+0�����`Ҝc�,YA4"O�	y�Đ���m`��$!���r"OZ\�d�8k d�v�յ?r�M� "O���F�
;xR��I�SJ:\��"O����a\�J���`[�Z��}"O�H��	6�0R��������"O�@����@PUʔ�G/	�H��"O����o�(B"Kgf��K�Lj�"OR�@/D/D��FB�Fr���R"O�Hb�+�<X	,�i�d�}@�kB"O�|
�O�|&��Р㏼J��y"O���b�%+����+I�u��15"O��b�y�J�R�(�\�
T��"O�,��ʉ�H�XL�A'�E��P�"O�@c]�;WH��GoA:*�j|�c"O�<�0MxB�`�� 5��9�F"O��hB���f>	����?Ң��t�<)q�R�n�� @��q �"v!�a�<���_�[��e`�d��m֩r���Z�<9���OP���VU'�)��R�<�箃2��q�	�+�TD
Ţ�C�<��]�n/��a'���}�Ѣ��<N�9��a��*�f����~�<�kP�0�l���F�K�X�y��@A�<��l+~���f�5�ܻB~�<�s��1}�5h��@(=CRI�Qm�v�<aЈWt�TE�'U�A@@hv�<	c��>��0(C#`�p�[%�u�<Q��1fУ� �R�3n�t�<�W&R�q(<� ��M�XM���n�<�q�J�ˊ͊C�O]~����t�<�bN�0cl�e�e .-H�F�<�� �p���K�޵��g�<9`'�6��9
���7�b�@��x�<�5�_r��J�ʌ\�*���Gq�<��A�K�m���IP���Za�<�T�`52���N��c$$�@F�<Y&,�2>� ��		���Q��x�<�v�@�aH��k��·q^�����_�<����=H��b7$Dr0F^q�<1�H�&�2E�#��0"��Snp�<1�+�7F��6H_�#G��c�)���y��c�l1qE/"'l�����y���	�X��ܷj���M�y����>1+�����e䌋�y ��,8���PL9$nPIu�Ȑ�y��C"_qD���JA�ml$W(B���z�*$ b��wв	3���+b h��ȓlXM;`a?k�݂Sܑy~����Jy�40�D]&���B�-ƒɆȓ1�<��� dZ�L��ȇ_ԩ�ȓ1��]3�^�FY��UCs�n�ȓ����J�oX�)��<#
��ȓtg���"Qg\�0�n��#�Ƅ�ȓ~	��`L�R6�Hx�JZ�z��S�? 0@��#~��lh#O�F��("Ozx�Ď�C�l ���.{r��a"OVR�G�5#?��j��j"OB)B���5�)(���1J�5�P"O���'Hw���Pʓ!e���"O����T�X�aiU�4�K ��y�-ɞ%���S�_:z����L�9�yr�Z:d\A��1v��Y�gcW��y���pe�Ԧ�zL,$��&D6�y�B��m� c��hKȍ�U�B!�y�,�<G�(�weՓ]�\�S5�_?�yBdU�B����
&X�vc��y�������uc��� �5����yoCn5jG��).P#�"�>�y�#~h��w�~)P�C�0�y�_\��-�4E�>}�|h�Raы�yRJ��<m��Sx����F�_�yBa�D���� �Ԥ쒖�A��y��*&��q�C6���!�l@�y�aЎmM0͙���9,F�	V�U��y�lL#4���皨b������y2��B���9��	%@��W��y��"�Μ��@� ��BW��y"nܧ"��L�e�%�1�L��y"�M
�J)[g��z�x���f	��y�̓F�̃�"{���x��"�yl� *�84�4�E�;���p��7�y�aՊ$�ND�"ꜥ-� ��wH8�y�W�a�H��&�) �L�)f%އ�y��
u��C���vo�5�y�<^t8D��D�� �֥� C��yҡх~j��A�:f�,E �:�y��u����v�(P�@�R��y"O��ay`��A' Y�IT��y�kQ<0`�Ȝ�0�Q!p.�y�DǬa�� �3#ړ*�ԑ �h���y��F�o]�SAEP?3B�"�֐�yB&هǨ҃�� �hI/���Pyb��.Q�%{�CR��)�	�x�<7F�V <2�cE�O�͙�k�k�<��\�py9�c�V�����HS�<��.o�T�1�k��1E��x�<��GO
���b��|R�x��Pw�<��	K�S[�bb� �,1�H�o�s�<)�،=�l,�&��224��6�Cl�<q���9U���B�M3n!�kLi�<�vQi3hy*��"^�|�S @�<	���84d�:3�"T=��co�c�<�a�+�0Y`1�ƚ'c�)Q��`�<Ar�\�o9�� Q�M-%�i�fK
^�<i�`��(�X|a� (Ÿ�O�~��8�<����-������D�W���c��~�<YB�қ{�$����<�@Y3 j�v�<�RAVVO��`솠h.�@Cu	u�<�Bɔ�NDp�� �-���XG�<�'"˅Jm.�9�\&#&��R�OD�<qbɄ�Xp]��̊���'�w�<��A�*X�E  �'n��u�§R}�'�ax@�i4i�p��Kf�;WC��y�ɟ�uH��@A� �1r�� ���hOq���"���0U�Ӣ�G(eP$Q���'R�D�
�Jdӥ�¸,�+d!�J�!�D�5@�~�q� ,:�� �*�!� J�tu�$�' ۢ���I�x�!�� 8|ٶΝ�rܤ��G9C,I�����O���D�P[��B�nJ�[�|	do�'d!�$C�om����X�<M(d�dH��)b!���e6�����+8\��i��qQ�y��ɍ=!��th��9O����Pi�8C�"q��͡���P?j�s��VU@B�m��ayG�t�u�"���z$B�	7�8����1*�d-�q'ѿo�B�ɥM���@�h4"X�Wě\��C�	�|���!N�N]A�kF
z��C�I�u0�|��.��t4u	���)U�C�	>�8,/�j����	A�C�,7���N�4J�>���@�B��C�	�k��AK"o�qv	�WQ*	}�C�ɫ	�$�)�t�r*'�Ӳ)*�C�I��P\��i�({���H���N<zC䉞!uz� d^z$�:�(ɢW�B��	#s�|(GN��\��ت��*t�B�ɦn�\����O�yl����Y%>�|B�	�^��d0�o��q:ř?aQxB�ɐ	J0�,H�q���֩D*=�8B�ɘC�I�	\���8�D�+"B�	#D�`��ȢZGd��� 4B�	��d��Ҋv�6D�c�`�\C�I�=J��@�����X�(-ΔB�I 6`�2�GCq���p�F �b��0?��k�Q������L��ayN�J�<�#�*H%���T�Z� �x�g
�Q�<)�N cPv �蝆D�a��CJ��̟���	9,��La�$�#oB�z���#'b�?	��I	�O1n\a�d�Tl��x��R��I\�������4��PK�g��F���"�B3D��s��Y�"��'��t~���tN/D��[0C��m�la���'>�d�Ǉ,D��0'
q�h5Z��垠q��+D��`�`~��[��T�np�-���+�$�O��=��D�I�	�Kޔ���&Q6��S���<)��1[�N�h��� kP<��"K+џ0F�,�{i��b�l�)wh	:��*�y�B��[5K�,���%���i�d����D�Y�{!n�"�K(w�9��a�k��\�a�4��+Ρk�hL��7`&D"��ُM��A���&_g�	�?����~��%�/Ӓ�s��W��0B�Jx��D�<��ㅍhRb�:�!��|���)�P�'_a��O��&]�����[2�����	��y���nB����m2*�.qC��y��.Hܙ�D�@okr���	�0�y��F�l�F��C�-i����X�y"�_MH�$�	��6��43���D�?E����r�Xq����6$���G;��Ox#~�υ� �������`�ѵ�G�<QB���f|�mb�셒5?�İ��j�<��	�C6�����FI; ��ύj�<Y �"XD I��ͮ-/��Ic�d�<����1�;���H������eh<YE�U����4�S*P18�� ���'ў��'V����$@iG�ꘈ!���?����!MCz���e�԰2����"O�i!wJ�_k*��A��?+I�c�<�k�=U�ҀRă��&�&�I�<y5�W�n<�33Oͽ7U|3!�Im�<Q���*�%��g�5h�)k��j�<QҤ�H8�Q�`���b�
�EIe�<� ����D�+R����(j���i�"OJ�X�/��m��+c� �!�<1��"O@�3w�ٰZ;$��W�ݍ{��i "O���l�!z�h�#�e^ez"O���F�u��7`����W��y�@˖L�,�)S&�T w$���<Y��D���X"��[A<M3�M�S�!�D3R�*�)BCj`�rA�u�!��N�,v�)�H��Kl<����!�q��Q���B�d�B� �yT!���1V�� %��I�0�� _*sr!���<�ڂ����P�.t��"O<�R�M�smRڴLڢr�Zh�E�'��ɯNZ�H ��"(��B5��
͞�'�a~"�ԕ<;Fdx��U�
����"B��y��9*[�n\%?~��d-���hO�����E�Hqb�i��"�W$�!򄈈(y4���@�T�����!��P5m�Z��r䏾�L-���[�!򄁀u�0'�X-�f�Ad K
?���>O�\�7ː	[W���b뀪H�>��"O��)1#��@�yD��<��[�"OZ�26 �;5.�;��Ӱ$J(��"OB���Ԋ5��B��٧r< �v"O��2.@1i�aJ��H!�y"O`���E�;DDn�!e��Z:�x�"O숈v�F�]���ؓ*�(-3���c"Op���.O�vpRJ�L1Ȭ�1"O� ��̌D��XCS�2)��P�"O��OC q�t4"�A�H#!��|��)�!?�����^�tX�I��<�C��	<�T1&�Qy�8�TK�*N6B�ɡ|9
}!C�HVJ�a���*2�B�ɱ]EB�"�W W��b�`û-g�C�ɺY�`-i����.P� �U�j�d8�S�O����@�!|��AK�U�"O:�3�퓞:���8eɀ�����0��;�S���7��t��W�T����1 v!�$ �z��lc�IԜIqD)��،Du!�F�R�9�r���Z����ž(
!���A�&8y`��\<
��ҏ��,!�_.^�H�4��4.'�	@��"�!�S)FV�Y2��;���7n�f#!�-\��8��� e��%:�I4e��Iq���ÀgAab���`��m�y�L;D�pH�
ί_��ȳ	֘&q�a#��8D�(�3�1Oi���U5yy��c�6D��1gN�;�P�S��]FUz��'8D�| B�qΦ��D�G�y�dQCP
!D�|�W�F��d0"1#^�&�De<D�0;��<A�l�!���,p�����O�D;�O�P�͝%	ZH�� Y�VK~��U"O�щ�� Q��V��3=@%0�"O�5qS�4q��eC{ `X[�"O))�Ζ�r�Y$��s|�<J�"O2	���ľ9Xvy�΍>H���ɡ"OƱ�����x����lЭ��"O�r��'Q<��%��	xT��2"O�\31H�"GFC�G�jV��"Of�HP�� ������MĬ@�"O�L�	Xd����$�� P� �"O�a�1�ې/��0s�)�S�f�;�"OX�	4@J�y+�59vI��v�X5"O���K�/z���SW*�9)��=�T"O� �k���M�|!�R
ʽ+��5�W"O��@E�C.�tٸ��}}x�p"O�T��l�Q�vR1��Qs����"O��qv@�1x����(CV.��s"O�X��F�ž|�%'��j!ji�s"O^�3�.��+�m[���L����"O�8kĬ���p7�39��h��"O�XxT���t����g��E���d"O��Sq�\�,9�%�
HzVP��"O���rC��n��%�c㓔jy~y��"O\ݐ���%�x���ۑge�E��"O���K7	����0VbE
V"Ot4��$Ğ�$l�A��3��a	b"O�ieꟈ?���E�Ƶi.���"OجU�I2a�`	���.�� G"Oҙr�h��F��玀�����"O�����\�l�2P�ly*�"O�0�E�r�2Pc؂�ꤊ3"O:ȠW�Ko�l؂gh�����"O*AUD�i����Q�����p�"O�q�b鑃8@B-��)�+0	$"O�����P���(�N\$�1�c"O��R��<)MHЃ�H6R�x�"O��:#���g�FQ��G\�v0��
�"O�0���	�� 놦�,'��;0*O��� HE)\](�;¢[6[|��@
�'Ќ�B��[�"޹����Z�8)H�'}�T(`o�u�Q�����
�'��m@��'7P�������0
�'� 0���ٛ`���$�t�b��'�*��g-�,	�VI��a��[A���'� Њuj��*b2h"TΗY.���'Ԁ�FMȌ*�m����KcvIR�'��P�&�%wB��Q�ɫm�%��'�D4���V# �����˓Q%����'법X���&O�\ �F\5>˦p	
�'1X"a�MKh�r��^�?W"��	�'��L�S�[/Da�)�4!]��	�'����@+ɩO�}Y�oD�ȁ"�'��8rP��U�p]a�nA���X�	���yrJO"%`��W�=�ƌ��O��y��ƙG������%
vI��yR��	jƺP�$��(+��pQ/���hO@���� �j�s&�$�r��G#]-�1"�'���{f�Y�2/�ay�+h�\���'�Ң��`�&X)�Gݎ_
���'�V����/{�^��c�Y4���	�'�~��Rk�YU�UrS��T���'S�1���A��;C�T�M���A�'�r�*���D���U�u��Y���.��L9�F�'͐h/�0xr"OdD��dN�?�u9#GĞw���$"O�ж�B�j�b]y��O����P�"O�d��'�VM9���'
�@�"O^�`0�0EN����:f�0�j�"OZ%�% ��y���[��3����"O����Q?��z�ϔ�qB�4�$$�S��J�'@l+��+��!�p�!���09M�yd-��l�F����14�!�Ǵwڬ�iS��w�5�@=�!��Ob̠��tjS�7��K�JV�!����69	T�R/J
����-��!!�L-y��q��i�<�����T�:g!�d̃e�Q���)Wy�pp3L�!�� b1�cB�* �VL����[��YY�"Or�k���2�LI�1h�!��1�"O�Cc'	ָ�0���8� �*�"O.@�l�Uނ0!��=#spu�u"O����M�q� ��e�OgEĔC�*O*e+��^.t�vI�����,'�HH>�	�;�5� 6�tX�/ǐ`���ȓ\5�) ��(�XX��rjƕ�ȓmg����*�@���gLp:]��Z��;Q�V#~�hQ�c1�R��ȓ=b���铼v��@�e�H��0�ȓt�`lS�y����f6�\�ȓh7�C�R,#Xb$B�@�\�(�$�G{��d��&,��N�/߬U�Rƍ/�y��&7$U
	<+��q�Q1�y*!3^�p�%A�⦭y�I%�y""Ԣ0�L�4�X�n`��ӫ�y�
{Eb�٦N�j���-ذ�y���5��1�@�I�%��%)�E���>�O0�Y�@�>m�\݈��ă;���B�|r�)��8i�q�e��mà��"�y��B�ɀ�H5y�᝝9~f8"��"L��B�	!	�l�����ry����#��B��&$U�D4C͌Xh�"[C�I��T+B�W��|�&�H ��B䉪L��	p� ;_�yh��Y��B��|����τr�5�L�Pp~B�Ƀ4{���iV�;�9iw����B�	�7 �3����^=�sN�Kv�C�I��m#�c��B�\H�)Ә/��C�	��L��Ş-I���ЁoU5i��C�	�*�X�jǙ�,��逌6�fC�I�$t�u@��%G���v,�0&>C�	.u�p2,�"Ȃ1�f�4$��B��?�8`b
�T�~ib(E�-��C�I�TD����c?V50�� H [~XB��
_�`3]Y�,�X�B�@�*��A��-��<���ч,��C��Y��̲�k�ja��2����B�ɩ= 2���Ҁ5ِ� 7��f����f���V˧z�P4�Bd�Y%J�gF(��0<�!!��h ��`Z�bf
`�<�U�	\vh<�#ϒeXm�a��C�<�g΂DQ�آR,�W�tb�WJ�<��$�y��8��_�K��� �d�A�<Ѣ�V��f��`��Ԓ��,�T�<a�*I06MrI�lZ�`�My"�'Ƹ�4�L���R�͢r��V���F{��$i�9�T��3��&�ǯo�aa��!D���w�����sdF�-Ђ�Q 5D��X�\$\�Z��&�D�D|pU	rF?D���agP�>�p�R���,�
��o;D��(��J�1���;!m�V�6�k8D�<ᦔ*`��4BC+y&6�"D2D���&�[%���3 <���QpH�<1*O��O>��Vd�
)���d�B�܈{�L�^x���'�؉A�V?߂��P	gw�x�'8
�������扭v]�������y�J�#������̱Z��Ԁ�y��Z�'����ǘ<�6ԀƏƉ�y��'+9����܇{����L��y�ƏJ@:�0U� {�6�F�ތ���hOq����	�3AL$12�r�x@	"�'��{���0Q�⟶W�nJr�X��&(D�� �Ig��,���	4!ԟEXL���"O�Q��	�7N$��QMҔP<�E�5"OBiQW`?}��(:�,��.扚"O\P)X!m��aT�Y*�U����b>��߮X�*)[��[�CW�8i�O �=E��/J�VIBܲ��kz]cD/���F�� �exR���؁ŌM�d
�L�扄�N��]+5$�P��٥�	)�%���Tp�0eQ�)����Ƌ		x�L��D���'-L�(Z�PG�O���`��U\;����I�"0�!@�$����	H̓
KN,�q$]���@AN%]j�1�	�@�?E����"pF:���n*>���*�+cZ2�|b�'?2�4��`�èV=G��Uk�kخ�)Ǩ<D���G��֑�B&ʗ^���r /D�@���� cF@x���D��,D��Y��ו:��E&��D�v��T=D��B"���Q^p]�k�l��%?D�� 恝�C2Ғ��Q,l�sD�Ol�=E��N�2N
0�(��I�Nd!�N��_��Ity��|���K'���C��(V�0�e�!�$�
���s�Ri�L9�N֮�!�˖1�h��(����@�K�z�!��[8!x�	��$d��`���[�!���7�v���J7I��	�j	�!�Tf�$B�=�qu*�/�!�	w�,��F�؊6.��9�L���ry�X�T&?�xϮ��%�K�`7�)���]��R���'%t�Hf���
�:����r���'Y=ptoJ\R5��:w(ȡX�'�ba���<x�����=!8!0�'aP`@%JT�;�<�E��`�F�b�'{��q� �;6�p����,	*���'(�A���Z�8󆔀���$/Ox�{t�ű�� ��G�(�̔��"O� ;� ����El�6���a#"Oش�D̐J�(H��%��W�V��E"O�9jRZ�܊�C��L�p��'����ta��{G I���U�ON�tB�Ɉ~��=CQO�L���C5�M3JB�	�JG���5���
-p&V�T4B�I$�H�ˢm�tт�2?B�	{D�e)t"ְl1����"<��C�	h�<(��[�"
��vDЮA�C�Io� ���D�<C���� �ي
]�B�I+��U�@�E45��L�ub�h|��hOQ>� ��U�?O>�s$�ɹm>�� D�(KRiD���ƃȉvuQ{�6�I��G��'�>	D�_�*(�&��F\~9[�'@`_2����� 2��T�<a�+pF6���O�
��i"DEXS�<a��ѓ)�^�{�� z9��{��Q�'?�%Nļ/~���g+��� �4D��hf�\+@��E�#�9؎)ya?D�г��!-�U��Y[�d�+6�>���O���>鉦��'k�r�G��6�0�@�'D���Fl�,R=l	�@,,&� ��#D���O�$ �dSTKS�D^�A?D�0�N]�PFL�3vU?=
�S�9D� u V�te]�SK7��1��M8D�XDjݰR?�]�FJ��+]�QI��8D���gɭ!ڰP�pa�H��#�&9D����X�S�d�X̓cޘ[��6D��W*�%�, ��P�k	��`�� D�� �A�ֵ#��S��Ư=2�j�"O��DA�{ST���W9l,���"O�аFH�Hv�5p�A��a)t�x "O�X��<T���e`݀49���b"O�|!����lpK��
�y7�BGT����n�S�OlH@b%@ךY|ڀBWhH"̒�	�'��8��l0�x��Je����'8P �l�+�F,�rh@/<cʗ@�<Y7��r�&�8F	��P��V��S�<)�I�6^����ઓ�y#��Aw��M�<�3{^�[�Mݼ	��ə1��G�<!���i����d:Gu�}���C�<����7ScVqq��+��J���|�<iwB��>G.TIfJHUz�`"���\�<����|����6H�f�*J0@�c�<�7���͖��h��;M�D3�FI�<1Ʀ�1?��Ī��*dI� &OB�<��%����P�У3�B��ɐB�<����� �-ᓏ�<�%Ci~�<��B�
D�1r
Z�b��2%�J|�<yw���vЦ8IS�})�ͺ�j�^�<��4�0��ȎFr̴���AY�<�G���"Gʂ%92��[�<�l��Q'p�p"�̲a�ԵI�.�m�<--Ƭ2���P.Z��BJP�B�I��<(�`�-��} ���B�I�;H麂��	G���j��FK��C�	-t�va���B�^�#��D�EnC�ɆE��ehK<LF�i@.65^C�1|:�`�-�-JM���D1D�.C�ɠx���E�XGb�@���0B�ɶ(�,8���4.�&����[)y �=Q	�m#2X�BL�
m�����<����Vn���d�.%�6� E�A2m���ȓ����;c����O�+vZR���0�^͢�
F�Y���O�+��Ԅ�x��|[��!�\P $m�a��8��a�&���W��Hey�l�Y��B�	�%a*����;/������R<c�j˓��9��?�'܈Mɗ%V�	�jDˢGB
G~B���'����5��<tf��-Ժ
UJ@x�'Q�D*6���4���D5�qx�'�|<!�L�B(��@���d?��	�'�4��7,�;H��S��O���M��'f\ۤgP�,��(5��
���8�'�(�񗮄$����m�y���1��?�|8�/ǘe��C��4�E*�O�C�I?#Җ��5�-�R�X��hl�C�ə/f`�3 -��>��d��hC�n���BT8W����f�,�B�*o4UYPN�8[�qQ'g��B�	�� �"[z�Dy�
��\�VB䉄]AJ=�3��T������C�*.'
49��78��� t,���<�	W<�K���UQ@H�N�������a�<�e玙;�ޥ{E-	u���3�PD�<q��̸@R�dbŭ��?���l�E�<��HP"~͐�%ϊ#@���B�D�<	G�@>R鈡�q�լW<.�3�[U�'a�����D& ����E�_Fv]KƠE��?��'�8ؠfX4���e�CH��I���xm�O�.dЗ����6 ��(/�y���!�tY����ՀQ��DC�y�&S�}��i����"Ψ�`�΂�y
� �L���� Q�G!ϪF�d8��"ONдܰw�x�� N�B1w"O6@#��D�o� }����r�ޠq�"O�$��$��u�Ա��I�O�TE��"O �31(�W�&�p��6�T41 "O T�!�*K~�hR �6bb��w"ORm�'��`;ʠ ç�tG��p6"Opu�E8?���FI>t�Q�"ONQ�����0��C>�T  g"O�H�Ȱ>�P��%������1"O���Ƥ��$� $��@��"O8	�¯8��q
��P ��;�"O*C���!?wr���Y��*M��"O�(����@O������~�i"O�ؓ`��I� �����9�J���"O��d�6FW�I(��|�bA��!�$J.�~)���G��TCa��C�!��M�y^�Ĳ�Nݶ>� u:�`H=3!�dڶ$��t�Z!zl	���ݚ$!��2S,�h{i~;7�S�!�$%��EF�6Xc*jS��%�!�d�]v�����]sd��B��"s!�d+]h�1B��WE��P��j�!�DQ�#BBL+@Ġl��A+��_�!��%��;�N�0*Ī@��P!@�!�dG8_��s�N4Eт,�ũ���!�����h�e� ��x���t!�$-��AV��/��広'\uu!�$�/_�l���P�J��T��E�^~!�Dݻu4���'\�O���!n �KI!���.Mٔ�b�
B�N}R�I.շE9!���TBl��흊 `� ��ݛP�!�^�S��m��ɚ[#�M85B6@!�$���M�y�����P�!�d�P9�d�����"�ܕr���>�!�$	uR�<�fJK�&�4���(x�!�$Ƿo�>�Jת��+����M<�!���,bP���R+�D[$d�w�!�d�o��403���3� q��^-!�!�Ğ�r���AT�69�|D�4��!�;f�1ƪ�g���Pd"� $�!���?���c����a��{D���'��h�HO~�l� �AM�^�l�'Wryu�Z�{�&�P���41U@�y�'

}jW!��#�f��F>�����'���Ӗ��zUڢ�(5>i
�'�Ε�v�Qpt4��Ưyz��H
�'	L�ak���d���y�h�;
�'\��ŭ:T�<m�4�N�p��i��'��4��]Fu~�����ve���'"�u+A��zXV���Ǟ�Wy����'?��&�A8	�`����L���'J��'KT<T�T1�'G,jP�@�
�'�TDl�+7�q�1��go���
�']��� �8+�0�R`�;tQ�$�	�'���K�Eүe�h@�祋�vRy��'���x�"B�{�F�I���k5zmx�'��0���� J6P�S@R`��(��'<�4 �iӵ{ܜ#)�W;^u��'Ѳh�U
�L��@h��W� �~Y��'/>�;B�1+gr��!��(��'~\Y��C�Xz�L_�[8H��'(���+i�`d�u䇟:�B��'�0��#��:B`��DDC6+�k��� �D�7`X�PZ��@7�ӋpY^�w"O:�q��̩(%��"��� 4j"OnHA��Ę��-0C!�5�H��"O�]����{N"-@���1`'�iqq"O�9S�e��t!�Ī��D�ĸL�@"O* 2��a�j(Cq��+G�&��"O,��6�ߛJ��Q&��=��, "O.D���Fe�-��`]�Xx�"O\5+�㗟fl`h�5l� �"O$���g������`G=.R4%"O�ŀ�-ʗT
��ʁ �7��`-�yr�V�b�4I���L,ygN��6Eä�y�"�>i&�IP�G�D��j�؅�yR��e��	�<J*h���K��y��'���%��8.mb�a�IS%�y��Z���K�]K84�����yrK�TF\��6g�7R���
�M;�y�@	~�,�� �E0,	��ʁ��y�5wk���ED/H���r�ΐ��yrf��H�0�ě�<V�!�l[��yb��m��T���58�ސbSe�3�yr�����gD�1|�b ϙ�y�a��P�^�)z�а����y��bW�I	�GU:1�PT��ǣ�ybE� ��Q��	+�YRF�	�yB(��A���J@Q��6-��`���y⭎B>��C����jiT ��yE`��K�@6@|��/д�y��+�\�c܌Y���	s� �y�L�Ci�@�B��>�
`j�����y���J��]�m'��Bȥ�y� G	o	�T�BnT�`�@��+�y�%�`�ycP"@�
h+�i��y�^	��A�!_@=ʈh��R�y�&��TJ�9p�ʋApP�{�̝��y��E���`JÁ&"���R��yb��ǀ!�FF�G���3�Q�y���E4�k�d>�)��D�(�yB�(lܹ����`���	�y��Zd�})��\U�$��щ�y�'Q�]bs6lDӀL�&����y��تCR�T(�A�Wf��f��;�yr	�D�s�8{s���;�yb�3_�&a� Nۢx:5�%]��y���$-+j�4g�0r�V4�BJP�y�)��'b4�PƉ�3i��=�E� �y�9=�4	(�*
j�9 D���y�Ӥ`�����0V��x�"& �y���-�8�怌�ݪ�b�7�y��-J���+�[�'&� Q�2�y'Y=i�Z�͋�a�(��K��y��	�E=�� ֿ��y�`L�y��Z@�~�q�dW96!B��+�-�y�
�5��A-��5u���4Ɵ��y�E���T��@ڼ1����s�J(�y�O��YN�1x��aB�W��y2'��r�$�ߒiٚ���B#�yr+ɏ���2E.�3g���P���yB��	�8i���^��Ԩ�dܑ�yRȓ� �� `ҶN��U
�#T��y��}���Q�L'�a@7��y�Q�F�h����)A���0gOA?�yn[��Ppɀ(2\���R��y�aR1��	��&�(A����c$_	�y
� �}�v)H�N��3��#Fy(m��"O���v� ���i���O�p�.ၤ"O ��]>�MZ`%0Z�d��"O�6l_)��L�F)/}�)"O ����5��UA��E>x�zx��"Or��0Ċ;/f*}�&�@�[�V�b�"Oxk���2�X�׌�o�<�F"O��@����h�z�KׄK L!�"O� �Ʉ�r+�|K��߀6�Ν0B"Oj4Zd�9x��L"R�`@F"O�	�$�L�#zh���L�VD�X��"O�aY��K`<��k1�_�0*8(� "O����%OUf)���/-!\�@�"Oj��k��xC�-s�8��"O�<�r�
^�(1��b�1�84{W"O-9$�_�>�h�Q��w���A"O������T��W�[?Z�Zju"O�)����n���R`ߎh��EI�"O�1��C�:��h�`F
IIpq��"O�	
c/�? #��1⎛�i��iCS"Otˆ�Ѩ:rT�MZ	aq��V"O��#�m��-y�)��kp6lID"Ou���P��U �	�� gn ��"O�a���t�P���B�9�,e"O��$.X��XR���B'���"O �'5w�\�ȓ@ق"O�%@B��}.����I&���C"Oh�+&#J�T��	�Q�,�h�"O�4�#CPn�<V�$(��Y""O���"��f�p$�W tBP�3�"O����,aC�h�Q��
H�|2""O��s&��O�II�A��}vT�"Oꄑ2�6 -CѡN���=�"O�i���9������5�MQ�"ORI:���9|�ܵF�W}2*��E"O
!���/$��#w`�&T�LT�"O�!(�\�	"L�BΉ�*��M�&"O���O��I!����MZ�|�$h�"O$��0F��c/Ѱs�	�ab�0#�"O`e�rdБ�41�a��]z�	$"O�ds�IȂn������B+M?���"OR��IM�^(2��A�%�:\�"O���\bZ�lX���2�B�0�"O��PŎC�;�bc�ҫ��
�"O�a&�$md��;�DW�z��U"O"Q�#�ϓKV8�`@c�+<��r"Ot� c�T?=��q���B?.	P�hb"Ol�rǉ��#���!���I�hճB"O�(��x�a
G�(@���"O��s�ŵz��=q�/�6<�Z�"Oj)����% ��c#� ,��""O�Y��k�;d;j���ȣt�B�6"O~Q�V��Z�l�ab皲g�d��c"O��ϣ���	�H���E3"O�8h�g2Il�4?����J$D�t�5iF R2�(���<K\�	��7D���$.�&�D�s)_�F-��h�8D�Dsg��L͋��J���h��:D� �PL,�Y��&^jd����7D� YGɖ 1RTT�"	�g::���K4D� q�ˎ],��""�[ac��3D�,
t���\ȲQ�<GcH��N3D����=y�ri�kM3�o1D�x��C;{R��2�&���4���k/D�� `\1��ެa�blHv��^0����"On<��DL@���*46e�w"O�=�U%I�{�Z��v(�4x��X�"O~ ��A�r��ʞ;��t��"O"�mޠ>�<$Sc��?:9�p�2D���F#	�e�!���`�@���,4D�DIp  ~��H�`��E{�� 2D�A�N�h+}�D�^�0��c%D��b遲B۶ыũV4
*��f8D��BAҋ;���gh��Hh����5D�D�c.K�G3��k��:Y��up��1D�И��c��С� ! ��"d0D� �V��-�V] 1.]1%�ɛ�.D��V��*����ڐ{ް��m0D�@c�&�����W�T����`.D�,�������m�f.�A@*+D�d!q�B�qDT��֫Ɨ��Īł5D�ܐ�C7�5���H14*���%&D�d+0)m�
Ԛ���$���IЪ9D�`����I/�X!�nS�K'-$@7D�Йf�� �<1����&��K�/D��P�G2���vL�ӦL3��,D���!%��&4��,;�ܙ�i8D�l��Gɧ�����ǅ���Aҷ.7D�Ѕ�F�L�Ђ ��f�X(�S�5D��w��)�X� �����z��Q��yҫH9:1�g++�@������y2�I-C�
 �#2n �b)ȫ�yBb �c��I����.�(���@��yҨN�o$>	�`W�#t ��#��y�	�*h���1Tȩ%/�9�y�A�*�a��%'o?�L��h�8�y�mP�j�ͭ2r����`�\f�C�I��:�엠u��ʲbț+}�C�ɹHp�$���"np��ʑ8��C�ɍ:�����  S܊��#�T#P�C�ɗ�����2���燘A�C�	"p��iI����}�, 䌆�G�LC�	�@�����&�4�,�t�O=�DC�	�W�H��A�b�0��D!P�.C�	4Z^�����ծY�H�
I�!S�B��&q�j=�d��
��k�C�p��C�	0O��H��Ey[:�*¢ ;�fC�$,�ܘ��M�8�$|�EɈ>7��C�I��n�b�fN�Z���X�D�p,C�I�@"9'�լ���$��*: C䉉'�·�6��4P���(��B�	#<����M�A[�(Bg� #�B�I�nt}����Ѯ�0U��0f��B��(Rn����� I<RвR��O�.B�ɏ��IF.֣B'F 3�&�0.B�ɓrL>���?)�0:��%E!B��$ÐᲨ�u[�P�& �K��C�	�#톉���8z(#e	<2�C�)e�>	��12�iIF�R�^B�I3f���qn�Y$��@���NC䉋�Rl:Ri' -�VG7q��B�#_v�u�B�3)�Ui #��avB�	$� �
�Z �n�I6���%��B䉟�|RuE	b���#��>h$�B䉠o�1&!W�@I)u��#�B��+Dj����W<"<qh�f� 	ҐB�	�b�v�!˃qLX�H �LB�	�,<�}�U�ϳm�"�4�#iLB�)� حM�2,��@�f��9�"O�d$��c|��ő	�	T"O�8� �	W�.��)�s}:mi�"O�Tc��	��T�2*X�D@i+�"O�e҂^ H�2��)!Ό���"O�L ��L62$�#� �p�d"Of�Tl4~8a�ud�7(�b<�$"O&�pW�ko��
4� �8�"Oh�x��H9`�ikf����0S"O��F�%nn�����3��Б�"O`h+��ϙyv!��� ���0�"Obd����G;��"A�3j���b"OV�
5Ûq��qڅk��	<�3"O��y1�Y��eK_?G$��iw"O�@S��!�	��̟4W�)0""O��h�:V���*t*ƹ�	{�"O��vNE3�!�"Muή��"OD��U�^��$=�U�\��v�+$"O���bV�x��;F,�)T�40J6"Ol�q��CSѐ��!.ݒ�B"O��KA@ O���Q��P8�Ȁ1"O�D`�1��
%�0�"O������<�P��W灚:��Q�&"O�E�gAL府b7e��*�:R"OBX�F�K�y!��gƙ�[�I	"O��#���J\l|�Ҏ�YI����"O�U�f�L�%N ̛A�596�"O(�b�X#� �U�߼E5��0S"O�ը���G�*�gi��a*l��"O����'��5��[7�¹X�Ӏ"O�%P�	G,>.���@(S����6"O�]�!I��t� �8@�Z�p��i�s�0��`���
�͛:8�Bڵ-f��`F�6D�!$�ڲc�ȁ�e�Z9$�� �gӸ�=E�ܴ6����5�'��(���a����c��|tVx`O3�(9h�;2@ʸ�ȓm<���AoҤp�4Ac��J�A��U�<�����Z��� e�U
��	9F4�!�ċ�z�,�b �K�h�&l��d�� ��IP~2�)���^�th �v���B~vP��EZ���x�
גM	�A��M�D~~�3�єo�!�d�.D��cv]�Pp$�&���/�!�E=alh�c���Ā(g��4H�!�$�>F�FT��L� ��x�M���'�ў�>)#��&~�� e
�I��r %D�L
�m�Z����!L�;}�y�1o0}��Or���>�"fF�hy9�l��5T~�J��h�'��|&�$�}�Q�ֱ]�Ȥ<𜔢�ǇO�<2*ƩU\�kgKϽ��R��H쓍hO�O�b�+5/$_�L�tcņ?o0tb�'\Z�I��B��T�R�4�Lu�H>�O�b��>�Q���6Y����o�����[�?D��sƯ�F�(<�B����
�#8��Y���kč4���d��3x$��EE6�����ƔK�x�KP �n<��=O^��������)��j��B�
R�&�a|"�|B�Q7�	s��#��d�Q�Қ�yr��2�<3$�N�	�\!����
���hOq�ִ�W�E��PY@��!<p�0"O��Z��	�d���ś�0� h�"O�e��YA��;:`����!��\/*���06�ϓ=�d�%h�5uA!���F�t��� �F٨�l�6�!���0��h��א[ʦ�a"
3�!�� Jeh�I��?5��8 ��Z�A��'I�ɯ,�0A�Q#Jz8��SA4=$�C�	��ް0�׾w�E�-_X��B�	5'�RѸ�M�<��4�q"���B��uv(5��F�b?py@��dS4C�	����f���zc�9Q�B�hWC�Ig��!�R8)RP0q�Z��B�	�y X`�F΃BӀ��ɀ&�B�	�����,܁�ve��F��v�B�ɣ8t҉������U�����Y,�C�ɪ_ �D�V�D�tT��$Y6o��B䉩;�^��g��7^�^�3AC�FC�.?���Ku�
r^n��n�7.V"=��t@RY���*B$�Ӣ(F� b����e��L9��Y� �y*�  5s���?�
ӓ{��IW
�i6��D[$��Ɠ �aI�� I��q��/x�G�?�Qs�y���F}c�2>�I@t�ѯ��L���ʹ��=�y��N�%�|�b恉�tS@���oK ���8�Oh�+�),J`�Tc�>4?�UQ`"O.4�#��.'���9DLpW><�e"OapD��3��|`�%�9q�Ah�U����ɹl6���^%r�xB�͉:@C����Tz���2�D�Lư8���w�?��p<��G�f�f��$�@F��d�Zz�<	g\�� �����1K��!�ѦE��8u�h`��ʻ<���K��I����ID�J��8pf��
��s*�^��!Gx��'4
���
)Gw�` ���:�d�'�"��N8���G��9m�<%�S��0>�H>iI'2�Lm��עC��A2$�O�<�	ӓ�ēM��UJ��02���yA�8��IL�'�X;C �#��EPcǥ0������yR���'j\�� �A�8�3хOP�NDyxR�i�E4#tbЭ��E8qe��uY�I�����IO�b��B�V��Y��^(M���I\؟\S�S�8c�,�V&�`���T@%?iÓ�ē{b��я?N�����Ɔ�AHd�'��}RBJ=��Q��GϝQ����/�!��>���>����.0� ��uB'Mzt*FKPm�<	AŃ ͈����7�"��k���j'��n��J����3�.4駌L�5�f��N�ȥO�ϸ'��諴��>cWu��Ѱ'�F�1��:�S�d�@�&�dxy��;}{遑-H>�y"H�g����`)q��%Х�E�y�4͘��e��o��=+���y"+O@b�����f��im����TG{ʟ�9���q�����$ȵc�C"OЍB�HA�I���H�f_<xC�`��
�}�������8r��"juc�Pc�!�$H��f� E]�j�f�rD	XJ�$LY؟@b�i��#.<��٦Wa0�+�'2�O�O,aq�F4q��:d�^@z���"O�)�R��R�D�+��AQ]���'�	
�HO�~��I�$�uF�p��*	�E�����2�ě�$����GbC�ԛP��$,�!�[�
݉a�	�X8��EC�)��O7$�S��N$@*����߀�8�:�� ��y�i
*�(|�S���|�8��'���y��)�'x�F]!�M�,݆�G��53���U� ȓ�&�'>�2����]2��ȓ
?�b0��X[����@��	�<9H����dW<䈌@��1	��A%I0D��!���	:_�=[�)��H��;G<D�� �lac�@��j�ɇ�f>��"O`���-^%�� E���� "O���� (�, /�Z��"O�9G���Xl�=��4Jx(!`D"Omc3(U'r�Nd��i_�uʲ��"O���̎�w� ���_�k]����"O�iwJf��8� �]�g]>p����Y�O��=�Q���D�Y�L"*��	�':2h�rLԆ7�Ăs���Z�
�O����S��>Y`�؅$EvPr�#�2xtp.a@B䉖��x���OKpy2g+�!m��<)˓x�!"��Z/9�r��L�#޶�ēU�l����T8"OFiJp�c�x�b�"Ob,(UfX�a
UB���E�!��"OX�+�:�Z� r�=%t�<��"O�i��D�ުq��FN����0��,\O��b�T vz�+�.��\wxy{�"O��2f�ǇE�qHPL�4��LIs��+�S�S6oH�
�mE<<���$�XRj���$�ɡ|VP%8$�O�	�u�3ώA���=��0s�_
A�`S�-@>c�� "}�|��O�a�c�V������7qu0m:t"O�y�����|p���S�̋���<��IJ�'	Re��/�#0HQQD!�Y�#�'�����̙�� �>�B�=D�P���.p�ư��Q�M�!f8D��H��Y�-FܔБ*7)�&i�N,D�h�E�,=��)�𣎁[]Ɓ�n)D�\y��_�Y��i����i^�E���%D��B��V�tHlۧ�n��b$D��z�`��]@�
��ڥa)����/D���3�p�:���dI�U��C)D�B���V��G��:� ��
ahB�I���@�/MTt��It�RB䉣$(ՂGb˒�r|�A�|mB�.jQ8أD`LZl�2@Ř3�B�	0Fs��Y�ئA�n��7�֦<�bC�	�}��1�d`��!Q
�y ���v�B䉏'0�,�MJ<�0ۅBӝ�rB䉊 �pxccf�,S|��2���B�ɲ�����W.!�>�s G�I�B�I�,�^�`76�<��၅4,DC�	�Itt��%G��Nq��D�qy!�̄*����e�" ~j�f�I��!�A{�Ɯ[SG.oUp�D�6!�ؑ��"�N�AixI0�D۳*!�ǵ؁��@!��ɠ��s!���fV֐"�)�d�� ��pj!�ē&p�B�p��	��\sF�G]!�dے(q��b6̓(@���7&�H!����g:1�dˊ�:j¸��J��I!�7
XAk��:,m�cH�>L!�D��{���2�j�{����烘!��ފs~�)�Cm�2}�9��Կf�!�$�#j�r݇�@��fH\�b|!��Зeg�p�%H�)%:!,x!� �Px��gn�)�a3a!�R�|�ꕓÖ�H���z!��O������G݀!nŐOd!�$
^&��!��,SԂ  �)U!��4�F����,�4UB��G�ME!��K�h-鄥���<�� �4-!��</�,upb�D/]��1PiE,O!�ϲU`�x�J�x��$"c�K4`�1O�Z���g��#��N�f��X�7�� �Tj4OD	s�0z��Č,���Ӄ"O�7/�Q�R����,odIs&,"D��X၃��r��sd�1�\bf5D�D�3j�H#$��I�,�.I��3D�h��Q�������/k��Fk0D�8ՀB�~h.{�hX	U<�9hbF8D�hJ��ԝg_�px��̃7�`|���4D�P�&��%�N`��*t*��@�0D��h�
��=EБ[b��&����N:D�\P��D�d�� �Ę,��ESЄ9D�x��Qi5�56-ƙ/^<�g�9D�L�%��,2@R��F�p�&H�!i7D�|�EM�`�a8�ıe��7 /D�c��i*��� �4�0#,D������ �0��FL?��T�6D��r�e�t�����k�k<�ar"2D�p�uC��?�)���[�$N?D�X�Xn�|50`L\P�X!�3D�P� �ZOZ�zD*Q�*ʶh���3D�T�`��"]d���#K>4e)��.D��c�� =��9���Jl{̄ХD/D�� �h�3:aH]7� ڒ�,D��q��`��uX���:�$�:�N(D�h�R%E�pL��(g�ܴ8�)D��B�ǌ2�@�ɗ�u{��ڧ�$D�l�#��>^<�����M��h�E�6D���!�E���ы���V}���È.D�pXt�	9\�H�٫&�i��;D��x!�
@%���ؠ {�	��%D�:��_�8�$��L� \��!� D� �E �-D���AA�^��8p*O�����j���#���&p��\�#"Ozc�ʏ9P�)��L�� �1"O��ɱMްa�Z��FnK%4�����"O��1/ M��s�DT'"�~��"OJEyqk� &���;qe��8� t�r"O�m�DV?Zw���$�o�BeC"Ohd��îG�lEY��=rtl�R"O杩��n �����IbH<a""O\���@�Mvi��H<sl��5"O����\%��KT�A���0�"O&�Pt&�i�Ⱥ��$�����'�*M�EI&: �ɖoP��Y� �"�@��BgQ!\zB��2g�`�ӥ�]�~peE�*$>&b�`.O�&;,<c����k�,$�@H��7�H�FO�O�C䉟@����KHE�A�}��1�O�0�ʓ=��!���L�(�G S27�r�q�)� ^���Q�$4�h�dbϐ[��)�$�l���(�M �$�MP�JzȆ�	�@"ൢt�׺c�Dy�A64�B��ė;`�\IÁ���7�F�0���8 �D�UQ��mJ
B�I�Š�3�O�6b��Qs#�+��O��iӣU-�� L:�Q�fHc��@+S������CLƵ�ȓW�xȅgR��p�ߣ�D��O��Y/栕'�X�B���>I�q�v@ C�����5RǇ�Kh<����!�t�1x?�A��	Vy2J�Vv��`��d����rC���j�c���L:����ɚ �f�[�DܔO?���	0�T�A(�*�Z��i�W�8���U�����8�`&�@@��<�@�LBE��q� ���s��JL����+)^X�ȓ?�|y K�;-�A���n%h铍Ǒ��'$lE�,OT����as�t�Ɩ�8�A"O���֡�=>{�09D% 6U���"O���U�b���,e_4�7I�A�<Qs��<Uz���J�{� `7��E�<� Tu��l�����'��>d��"O,p�u�Y�=��೧��f��"O�Q�2��v���h��*=�����"Or]�P��!�D
���Xq>8"ON\�Q% ��9��Q.t�����"O�p��b���%˕g0`x�i�"O�|:W�
�8`S�C�Ev�A"OT8Q�U=Jzk4�چ�05��"O��S+��b�K���(G"O�x�F�·\~ʕ��J�1'��p�%"O�%�3"T.,Aٷh�\$���#"O�<b#�&��,�fĞs'��05�>Q2�=4�J0�AJ6�>�+u��4zC"љQ�ׇQఊ�"O��k��Y�0�*�oOs�6]Yb������=s�Y�$��L�g�dö�
Ѕ�L�@W'J'vH���	eƺ���B\ÜY�(�6I|� @�'<-(��E�4	�a}"����s+�<o���J�@H��O��
N�Q��A�����ÿ Y����O��−�m�!�DE0 ����:�5�U	6�剄xH��r$V&N�(hz1�.�ʅٶǹW��t���3npC�	)/��m�I��$��	)�O��⪙��~R�aĖHz ���{b�S�2�� ���Q�q�`�kG�'��?�6ӱ4�:��V�mܨy��?��C�.Rax}Q���v<��ˉ{��	A�Z�ȁxR��fh��2Aܨ4�џpg��'*���q�ʅ<r���*P�"��8pŞ�2#�f� �%���r�]d�$b>c��f
�*h�dQ����y#��<���پoz�ʗm؊rè�|
7�+�����O1&�`+�A��f��+�`Z�;����Ą3��r4��MpX�+`X�F<aC�>���^����Z��_@J�
�$:���'3*-�u�lb��=U�و�'� 1ڵbb�&��Ԡ?k�3���0/��Pp�B<B�s��2vOR�O"|2 �G/�Pa�����N8x�T�o�'��E%�s]0�$>m�� ٕ`�>�s��D�z%�л�钷�?�m�9]N���"ʾ� �3����wa�0d�ҕJ�(4v9�'���[��V)��ؤO�	����𕨀�~M\��D��}c��݆0�6�i�g��U�ԅ�	�3ezU��_0n�x ��_�S���(K��`��=:��5�F�-���[f${�v�=�y' &Ni�f�����.̚��?�q�� �T���2xV5� �e��J��
�%���'���r�Lq��A�D�W[��<Q7��#�P�8N��+���U�B�'����A;�@$>-��.J����A��5( �ҟ\���ς�
1� 4�-E"��[-L�����^�Ӏ�I
���C(4��C����?5S%¬##.!%�; wR�[D�.��My�jRS+\�P%���O�'��A�Ɖ��$BF�S�-�,��qO��2'J
XG���B2�Ե�y�RL�h�ؠJ�=v
ԥ�E���?� i҉O"t@���E�6,��><V�<
��B'}.Eq�)#�Ɇ&y(#|n��@YZ����Tlx�1,��J���$<=]��B�8��<\pjt� &WlP�"D�E]!�d ����d�Ӽ\�"|�Fn���y��M�B�<�)�SK	��!��C��(r ��=҆C�ɣ	��tb��ŕ]�ā��i��x>�B�	����z֍F�ԝ*vJ="8�B��&�f�藀�0{g�q{�LO �nB䉣9H-�`À4Q4i{��C�vSHB�	)�@�a��+�))�h�JB�ɬ[���eZ�S���Kbd@�Q�4�<�
C�Z�"~� �AR0�%��/^a�dH~�<�W��Fa���E�)I $��m�'x�h@D�L���S��y2 A$����1O�^��0�O��yb�M:?W��R��� !X0g�*�?�S�X�&�Nr1)0lO�,Q�B?�t(�A��X�H��`�'�8x������Iڴ$a��a6���TJ�X��ON�;~�(�'3P-�rm؞�a�Gշ����եQ�d��$#�(v\>�8R�8����O�h��DCxV�{G'�B_�(�� '��m8��#D����ŀ�=K^�S3��
8'���:LUd��?�~℀�m��Y�"@$����O@�Y�;!|@#&��_��PS�����S�? �D��e�2�H��3'�	� l�S�	\(ka���<w�q���;��L��%�1�P��C�����I��p%��>G��PSs�*����Q�3�̠I�� =Q6��������Gd�����T�D[�v"�9;�����h��P���r��'���B, .��1��V H��{���*�m��%�+b)��K�J�B�@��?��;�z��D�6"�XIb@���D���*&d���:��y˃��#PQ�����
v`��'
\,*Uň�?�0�8�q��)At�ݧ��@��.BYR�	�!�,zW�B�ɶ?]�d&L�R�Bc%.x�t�P�ЖOj�I�İT1����6=E���P�@�SnyrA��o�a��e�*X���n�3�=Q%��a���y&�B(cܮͳ���;/����S=/�t�t�<	���"��=6.��b�WBD��?Ѡ��<CI���F��.1�<(S��Sy�+��G�� ���=6M0l0o�}��]K��L5��#�Bv�KJ\9p�҅ ڊ]5��.�Ŵu؅�'R�ܲ�L4��4�M"}mR)O�: � 4�����=�0ts�� .Z��_�D���v��P�� WW����U.H/2�~���y��Z!�݃5�Rԉ0�	o��XS4O�=_�8#��x4��̍7F��kqŝC�$"[15�˓��iA/�rL@���Ӌ*U"�G}��7�fxi��Ky���d�<�s��?w���zp ׀!(�8f�:Eh\�;'���d%P��a�2�?���T�"�(a�B�LE" �ӥl?yG	�]�MBA�<��J�% hQ �IH�`�X����;C�,[ � �\�{�Ϟ6a%��Ud���Bjڦ�@!e/I�n��@�����"�U�"�C!#�Ze/~�\5��l��|��aP���2|*2�f�չ~$� �����p?a��P9��B�FH��$��7&Z?A&]�#ɔ#k�$�`H�{e��A�%>�J)z�(�<�6©`G� �ǀW�I \4b�ÃR�'A(�J�$��{
p��|�֮�Y���T��DOX��R+�Q ��˜���5���	n8�L:�g�8}�bBubq��ίf����>c4t4�cK�)Uw�S�3�K(Vst)S��Ӳ8�%s$�<.�����44<���-۲�Px�)�y۰,┉�>\J�qY1���ē}�������7�<yK��@�8����'G�8hh�(Ǉ�ڈ"P��gľ��	F�<`ƆS�\BP���c�Bʴ#kV�al<��UDĬi0�X T��E���d:$����2b�H�X1,Y.2��ȓ]�%	� �S��Aqa_�^v��'�FA8�GD�y�rQ��ɘ\�tD�bd��kp
c���>`�0���\�b�>��e�-X�v��!� ft]XSDX)�؊�'�JU�(]�"s�� �*�A*�8��Dߩd�KpD.�Ӭ�B`�g�Lp2 �yD>F��C�	�E���s�+ީ[ �֡k�@�I�Z�X�����!N$�q��"9����Ӯ�]Y0C�ɽBmJģS�P�Cæ�� �W$E�C�	$Ǥ���a��TY��˖T�C�I� ���3-������H�CWnC䉨;4�E"噬 ���Fǩi�ZC䉱C�y�4Ǉ�]��p��| C䉕q*��6ǜ�8�Je�L��`�C�<�,���g���u�O�-΄C�I/�T��v��AQ�"F�,��C�	*]>�3.X������Px�C�I�8�H�ʡ߱Ro`���� �yK@B�	 $�$H�U�ݤ$�6����2[�2B䉻#SZ�{��ދ<.(s�)j�^B�/�F����Z�Y.��D&�#�C�ɇm��Z¨�P��b��V(Z՞C�I�Kc��r�
[v���]/�C�	�WV�9{C@��()�HU�h�>C�	�/`��r����j%zɀ�.ōj�B��)�*�RlG,L5r 焪*B�ə3�BL��T�^�f%
� ?�C�B: ��d��Vp��0��q�C�	�6�Z����N^}*�M Z��B�4kΠ��E�J�&Vtʖ��� _�B�I�hR�����Cv��F�T&b�bB�	�Kb�<�� �iK�xR�U�@fB��	Ʉ� �V+��,�5��:��B�ɦ6C�$`AΫ^91�*k�rB�	+����m.7`]�5n�2V�TB�)� ��93�;U-����Ŕ!zG"O�I*���BNcR!�@�:�"O�#�^�$ �� ���@"O���l��M��їp�~yi��?D�4a�IѐH
Hz��Q�W70ɸ�.<D�$8q��.����%����M;D����  d��Į�8b�2�;D�8b�'Z�+x�{�c�1xMzӳ�;D�`xw���k��B�D=S�v88�-7D��{R���8�:�E�&m�Nw�2D�X�f�X�o���s��ܟ%�8���5D��e%O&F���[���<=X �Ԁ2D�ܱ`�Ԗ`�|�s�&[w��8���6D�T$$�?( ��rGby��u	H�o�<!Qi3���cBGq�l��!Zj�<����8�r���V �t�ҥ��S�<��bQ�q��yaH8rla��^e�<A���+A��%*�Z�nޝSŋ�{�<��a��L`8����E��Uc���w�<���QmŦ5��ܯ$��H
��	q�<y@ܓ+�C�KS�T���rf
Nn�<iŬ<��@��F�:�� A�<!2i �6����F5����Z�<�Gä��I�������U�<��	"}�f��H�3#]t��ĕX�<��f�0D�T�­�.W4�u��A�<�F )�����)J�w,T�Q��C�<����Hd��"	
9Egf���B�C�<��n,D�ȡ��9-���',�|�<�Ɓ$9-@�;Ё�Ų�U�y�<I��ۄx'��WjV� ��A�KR�<�́Q6�� Q�ߜH��rN�<q���:L:��#�5b�� �rA\m�<����&1�v)� ��L���FQ�<����=*�jw.
�7�Aȇ�I�<�C��=�����k�>2ڊ�� �\B��$h\t�A�+ ������8B��1"-����h���IE��"$�C�	4j��Z!˘hO���s��?X�B�/)�n1����L��-�b�UC��3<��ĺ5��Bt�q�d*�2��B�I�}�\���Z�o�DIh�/L�B�	!KMz��v�8]�<��p���6�B�	O螡8E�è:[����&G�G�bB�I!p3�p��Q;�&��q�b���"O��'ߵS��42�&'`h��'��Y�I�[o�I(gS�Ea���d����e�1B����n�Z؃#����D���H`�<����>�Bt���%�'P���CR�S�t���Hį��C����Fv+[�I�r�V�P�D1c���'@<��F��>�4�
n� ��0M�rg��P���wh<QQ�\�F>2�{S����b93���j��:Dc��2-yx�|<���_+v=���ۛs��x��I�],b�Gژv��pϓ#��qϓ�#����Gė�2��ȓ`��!(^��D� mސD��a%�L�P-�C��QY6n�_�O�I�DO�G���1��M�*��'����@[5\z��Q5DD��J�8�
�;X
�A�-OjL�b-�3}RjV�A�&�G��RX�H���_���x�R�m�e!�
�$�J)���ՎV �qF�E�k2�'��p���Y�3�~	Pw �iHJ��3�th��1jN@��'2��e�UZ7���u�m�D��'� x�7A�z�A���!l!��r�y��̠n$��Z�O�G�O���0G�5O��r��>��4�'�LC���.f��X��R�zpe���15;�Orm���Y�� �P�� j�{���6mA6iW"OJ���_24�,�@� ��[�e2�"O��a�+H�ȉ���t�
h��"O�|�Eeڥ[�T�S���!
��4"O�@���ͱ+�nTH&�A�&F	If"O�`��k��e����l�-7��#"OVa�ba+I�6M�3�Z�.�!�\�Y�����@ʆ���%L�>
�!�D�)Fb���F�O,���FL�/Gz!��цFTh���U:�e�W:DE!�d2~�:���"R�F�z	*Gʍ�`�!��-a;F�G��<�@�i
�T�!�C�u�~X)��0�Ji����p�!�P�hؐ�%�I�!�U����!�ą�L�lmʖ��80¨�b@٫O�!�䒯J&����C�F��h���<+]�*�����A�xT���(���c�/I("���D��5D(!�ӆ�d��� 7� 2R�ӢA�0y��A�<�H�M�=�|�<�)�X�	#�'V&/oę�/Y����S�[�O������%7�>�D���0�����	M�H.��>�dmU�'5�9��G�k̆��FPI�'���FH�=��[V@�Z��A�$t]#����@E��'`X �y
i�M��D�0��Q HI���DJ��ڬ;0� ##��ӈ�� ���ɂ�Ԙ]XzXh��ǈtl!�d��m�F]�F<T|`��Ԯ��}(i�&�Tu?�SCN�p:��#I~�>9��S7^���J�D�!*9�O��0D���@׫K�;����N�B����  wK2:����n;�I]�'	����ɡ
3�P��D,�D�E"��"�>� ���hP�Oo꽳Є��rAT��&GB�j�|�fG�@� z���y2��12|@�ag߼h��PtEY+���@�A��f��Ek��)]�d�����dJb�nѱ���J �NH��(�"�|c�h�<I��� ��E$Y��5
��@���d|&6�n�!X��vgj �O�|�r&��eyj���6S�� r��X����f��X��8��,�����=n�YA�Ad���`����Ö>��� �H�ܚ �F�@�����jDџXP+�;��&��tY�P4|L�6b�:'b��9Dn����i B�kr���E�����hO�Ր�-ǷY���ō0���_��M;� ��>�'2� �c���`20E��%�(aa
1���ʎ�R9bTK�.VV�:6�'b-����p
rĢӃ٦1�yb�a6}b'��Ii�}�d�-��ys���\pz o;l���]�Y�<����(��l l
es����!Z�$�a���K�ԁ�"ȭ@�4h���SH�!�D��}-���a���M�j��!���#(�fQ��b3�U���l�џ��p<�Ѡw��!�^.�`'ĭa�l���e�R�#~T�����i�f�@��f�<�Af\�J�H�&N˓3�Ѫ̡+�ҧ�4��"%�x`EdY,���(�*ek�pC�F�8� ���x��M�����jG6¶t�3����'n�u��'�3�������&7h�������9��t�	�J04��dS�
��`� K��Dx��ۓ%5*u��$�ܗ�X�Z�珼��'�^�B��i�r90c�M0��Ɂ��J�m��<"Ólb��%͎�� +pp"���\0:��oE�q}����Unzɸ�/_��{G�٬t�|�O��Ζ3ٸ��O�aA��mT��y .�+/��b�'>4Ո#�H�µ���� Jx6��'���goW�2|�gB�L�P3�'�b}�牕q�@)�B +��p�'�Mc��90�<�����) v�,��'�NhAmX �����#�����'C�Yp"R:so:,���Ȑ-��Ë�d�<=A
�Q��)��j�����*Ou��b'DD�!�$�C$T�@��#�\���	�jE����F��O?�ɢ��J&��;t^�5��� B�	j~����e�_�*�n͉tR���
Y�5�%ҁ��=Q�+@�).#��ĢH0^�K��o؞�HT��	t�����w��	3����-�D��eZ�T�>"p"O� �a��!^:-����Z4j������c�D�������#}����8C�B�d�Q5�X�+_�<����7{z��[�	ވS0�ZRڃ/�XM�g��?���9j	Q>˓v�{�Ye8�q vƀ(/ELՇȓ"�D���TLI2��m�)t��+��Ժ>�VU�Td�}�a{�iԕE�� �b� �pY�����p=)P��i;��F��M+��Q���vN˶{�BUZ�Kt�<�E �`��H���ǭ�~|BI�[�`:0	��A̮������CpV$�C�I;0E��"b��K!��A�b:��
%F�9�E��%J
(J�)G�q
��?O��|�'�
=S��r"�	Q�V�c��� �'�N=��F����AAA .>
H���T3;l�e@pJ���0>�2AP#9���2f��]c��ۑgT؞� ��1?���Kܼ����>�I�����p�݇ȓ4^��Rb��,oX46j�b��'��iI�l4@٬	��o�W�O��K�� rcB�7c�����'"ZY8D�,� 9�L��a4�SN<IR�ٗE�`:�
OH�����3���%I�2c����r�$ a��u.�PWMU�=ֹC7j˰:�2�H�O��4����	���	D�v����I;N%�XH1�(1�D��Ip�|0 '��:�ZqS�"O��PO�Ol���G+g��%���O�i����;4T-�L�b>!����4�r�S��I5<�J���/��,3�"O��a�炠]xZ��el ����>!�K�.��h�iK�7��H8�KK�i>��%3�@��G��5o�rp��)2�O�d����4r�v��f�v�
("%ぢ[	D��%��ao��P�K �P0�'��>	c���ׂڽ3�<�J���I^�>I�"P�2'���3�o.쑉�ؠB�:٦g�:�\�a�Y��$������d���Z��W��.�r�Tˇ�
�T=`�z%��F ��)��֎t�2�ғu2r,{��42h���m �s�(I�'��}�q�X$z��e��dIxNT��J<�D�>�������*6p$�4�]y�ԟxe���^):w�	��L�C¬����'L|m�ՠ#q�,P�ۧ�����8k:�e02g`|�MZA/�I��S�K�5�1���#��$�>��؅�8��xrF,x��ui����s��}�'���cw吐N����oO -���%d�&aP��,L:��䟬	J4�ɖ�R (?�呇Υ�Z�F���s�c@TH<i��S�{0���!ʃ�ov�Sa��K�'�0`B%���79�f�AAN �C^ֹ�
T��@9�"O.��Q'?X����^��ޔ�R�O8�Ѣd�>���h�����[S8]ju,?:�;�"O�5�AX�g=0t�r쟿R̫g"O�mӱlA�L��d߫Q�����"O�|ѳ�R�8�~ЁG��l�0z�"O��!1�D�ST��" Ë�x#R�#�"O�P��@�L,��c�x��m�"O�@��E�.��5��CR�z�>i�"O@ti���PV� J�dȐK�z�a7"O �BꁾT1rv�؎#ǆ��E"O|]{�/�+t�zTJ�P�oڼu�"O��6E�V�飲 :*����"O6]��	�llm���/3�:	۵"Ot��D�G���|ZRN����r2"O���" /Mo`iC�o�?	�HH��"O��!�J�|�<sD�/��qR�"O\����?W �i��CJ��$�b"O��A�+B*�r�hCBַBH���0"O��ygLz��t�eA�/����c"O����J��d(�ѱ ����Q�"OJtҀ �~*�*B�X40*�p��"O��5�Za�Š���\�H�y0"OD9;0��r��*�)��wvJy�"O�thÂ�B�ܥ�NK3z���"Oڰ���Ȉ9���$�˻%SLt�"O� ,��\���:rb�)%[�a��"O��ш<YD�	�t @�6�e1%"Or!HL[i�����YǶ%�G"O`豲�]�S0����ZF�Ti*q"OVb�D�;haڨ��$�|x:�["O��c5�Ax��y�i�gQ�$2�"O�$E��vi���\�l���
W:�y�P4n��K��FD���	M���'���j���y�V�=�t�8�y�f�z_�����-{�1����y�iف�~D�C¡�r�q ��y�W�tOtm ���	�x���,Ƃ�y��҂'��Y���u���b���yB� (RC��(a�š}+Z�7"�"�y�ȕ�4����B�-��i�ɇ��yb�V*w>X�	#�ɃT�~���ï�y�CK����rN �5{@���ޑ�y�L5l�d	Y7��*��؋VX8�y�,WQ��wm�8�ݪ�՘�y�#�D]˓�G9nڠ0eŨ�y⊄/e��Y��M��%: ��p?��֫�M[ރ�ؚh�R���k�q�P������t�j㟒�n��vJ]<�,wdP6�$0�>1Έ���O񟞝�W��rɪ����P�"| �D���t�x(��
����SA>��3G8a�DcÂ>�4T
��?r�ՉV�L�@	 ��0|
�S�P� ћ�M�7Gf) � �Pa<˓I��� �da��h�� "�WLNP{��S�ʸ'&�������O��	��E��LۗDW�P;����r����˶y��$�����������#J"�q�6���uZD�#ֻT^�9��O谀�g,w����	��T.��P���t�jt�_H�	�"[���) a~�Ş$��C.P�y�l	+%��I����?1�"7ʔ�ZRi�j�)�'��8�0�K`� A��n�z�lڑ'$}ap!!�Ԉ�M�ȟ�<�FD�R-��:���	w�i�Oo�B "��Y.s���`�a���g�S�@��:]x�Ĝ@ѬH����[�<�cZpc���#k�h�H�,\�<�..�q@
�Gt�eH�r�<#�Q)]��2&��>y ��xwL�q�<�D�R�d���D޻Hoȕ��c�<	&�V� f�ًW̏"dW^} Bg�D�<I�JT�9���H�!�8c��=(#@Hf�<�Ed����@�gV|@�+g�<�&�_;Gp�˔䑗7d8Laad^`�<�Q�̳�$�z�i�;+.:Xp�A�<q�ˆ�z��)7hȢ,������d�<�r�C�v�pk��Y�4�<�ӣ�g�<�Q�S�˼@��S���x�/�n�<I5�T�i�Xa���W�R��a	l�<�2�&g�l 8�O�=ޒEh��@�<��$��_��[�&�_�mB%�}�<� *�b����ɉ3]t`�F`�P�<�e��;���:|�p@"�u�<	���LB�l�`�	�3���
ŏu�<��iI*Ϻ%C�ĝ ��ga�o�<�Ȕ���e�v�PNZ���w�<	d.Y�uM�D0���d�@�Js�<��GK�E_(a����ZX"�HÜZ�<��W}�<�,�O��鱡� ]�<�ǫ	Y�Y9��37��Iq�\�< �N� d���'��=[`�rK[�<AP	L({�:��0��7|S\���FZ�<!֣F*n<��H�d��ܹ7��U�<� �QQ6vU�r�ÉS+,J��R�<�u��x�D�`E�� ������f�<���%�uK�l�����c�<�&�g�4�� �kW�1�QF�<� T��a�ŶG���u埽s+0mr�"O�i[g�E�D����S;z�aQ"O88��\D��b��8�0�"OT�:F
�>���ݫN����"O����I7�B@u��$4G���t"O:mS���<�h�A���nO:5�f*OzU1�(
@;�`ۤ�ƽjHг�':dE��l��x>��ƞ�7����'fҖ�i��h���v'�����w�<B@�|u)5;"}�%(��p�<��b�4h% !ڑ'�6$���
u�<���O=���W�Od&h�̘m�<1���?c���FIQ<WH(�CU�MR�<Y��"*F�Dˈ9D�4q��iH�<�P ��)}|��!�,����F�]�<��`d�r��V/D�k�̝z���R�<��)`=]�a���L@}2�BMu�<�塎�5+�i����Y�H8��t�<����8DR*�-k��y3�j�<!D�-��{��\@������Q�<	��=���#j��i�DdѠ�P�<ɧގDun�
�J��g0����%�R�<�b��2��u��M21�Ra[r�Q�<�6���`����C@	+�T �)�b�<I�fCS1���
�<��Y�1�H`�<���@,5W�y ���N�zL ���S�<y�	��"���*�Ǖ�
RmcQ)
S�<���H]�]�`� O�T���j�<	Pg���ѸP�Ғ60aDǟq�<i
;5�)���!<8Hj���m�<qg��K:(I��L�=��Q`�Oi�<Ic�x��FU���t�N�<y���	(�N��U���D�T���#P�<�#!Ciu�x����ơ���T�<��ٜ8�L��E����
(�0�CP�<D,]#oU���ޑ���w[f�<Y�HD�����R
N*��R$��a�<ٗ�W����bԇ+s��I���`�<���X(�]�H���`ΎA�<��S�AJӈ߼�er��@�<��M��\��"�:6�(����WX�<�`f�+P�`�ؑ�����pqo�W�<��ګ�@!��5b|���T�<� l�Ofj�s��٭jh 7�WF�<���ͧ����TMϦw�-t�ZC�<����4z� ����N�^��q!��v�<A����<�$����_�m��X�Ңp�<�Z6.r���͠H���#,�B�<ٴ�^�b��
ֈƲjŖ���"O��0Fe��rʇ▌<�Q�"O6��UI�?������>��)��"Ol�J�ZlY�����8��H �"OZ,�⣀�\�N�(�l�,r�JD"O�D���(Z�p��iU�l��I�"O��RW@�O��c
(F��3�"OD}�C6���*��%dX0D*�"O(]���WU,1�I�R~1��"O�I�����8�2<B�35��y1"Oڭ��@ʄ��Ps��*B!`"O���c�77J���)tbH�b"O�U0�lߴ�*a��a�#�PY��"O��t��6 ��fŚ(:~�Ja"O�e���HN>Y�4둲q8���"Op��b�If�t���DKa����"O� YBЊ>rWz�s!Ç�{DX�E"OD�"j͊'��dPȚ�b�*��v"O�l�����?dN����O'N��"O2e��ŋ,�9���[>'	��"O�{��ŗB>��
�'� �p��d"O�L�a$��4�p&�1%�DE�W"O\4
�mB4���FӖ-E"O��؄�:oA���Ճm��
�"O��cѬ˾4p�%ȋ?9Ȗ���"O�cOA��{(Fx��"g"O����Nݖ)G�t��-�t�F���"O��؇��C��}��P�$8��"ON��0!�"V~�dRDf�%0,�U"O�-"*�0�}3��V#C��j�"OXh�����$�/�buB�"Oz`�E\�u
��"����fX��"O�1���4x�"�Z�8�"OD�@��+o�D����K\�c"O���B'Y@fx�GB'zN���"O������5L��a&旱X����"O�=Z��*��(@$X$��	�"O&=�p�_	eNRa�D��X�R�Ac"OP����>/G�}�0Mǖ2΢�c�"O�y���Lt�h,�$d��)�P"O�x�ɒ"z��8�׭Ё)��I�"Oą"1���J@ 8`�FE��9�6"O�U���9i�ȠB(O���j�"O\�+�L')N��W*K���"Oz��&ٹ���y��۩Q�qH�"O�U��+�(=� Q�3���J�����"Op���U�,Ek��DnE��J�"O��@���h��,̪c��ѣ1"O�H�-�t���!�ԩ
��A�w"O�8����j�����ǉK�B�� "On��C(�?�����P���I�"O.�x��ىl��U#ťN6	�h�"O�,�%��Fh���c��0�U"O��[�-���EfN."g<) �"O�t������q����+��]�<Y1E?C�v�V%��E�xqy���\�<��ؓ=5���]��p�!��M�<��!��\����2� �u� đ.VI�<9I�Y�
�	0��W�Fa�a�}�<1I�+'��1����'/���N�P�<Q�GQ�E�@ҥ���(�8�FI�<A�l<B��yQ�㞳\�,�pgm�F�<� ��L�ʼ�vl_0z���7�k�<ٱ;ў%��Y*kЬ�!"�c�<�6�D�^\ش�����h@� X�<��sHZ�u&� ش�kb��P�<pET�]�(h{��H�iZ�0�M�<Q`��5�MI ˈ}�j׃���yrA�����ё!�l@*7���y���`����%�(|8�TM��y��
�O@�$�$�-v��8�#Ȁ�yR.��J��`d����H>�y"L�΄z�oЧn'XD�@.���y���m�H��F?�"l�@̊�yr!ؐS�i����l���Ó�yr�,.O�Y�B��&�����2�y��C<̬p�`�� �d��`L���y�F=O�|D �,U�nπ��`+�ybj
<
��T�kP����K5�yB�'N܌{�/ht��C�m�y
� �D��ڤg�FZ�%�&y�v�"OT%;&��"+�>�k��]�#����"O�\AE�2 ��@jJ�/�܀�"O|-��"D
M"� �G tz�5�T"O�(SӋ�0�8�8��͂^@��*�"OXPT$� ]älrdA?uA��y5"Or4��S!P`�q�����;��\h�"O� �b�с �Y�7�!czVu""O�{����B��ɂ��/vxH�"O� ���#�ly:�A.�����"Oty�D½Nζ)���0�J$"O|�	'X�x�Ѐ3���5:D`}zS"O���嘭�:ݘF)�+��Q�"OL,��-�,��QJVG����"OR�	�i߷=*fYjg�2Mm���"O
�Ӕ��o\�A�BO0T��v"O��j'��s� ����+U��uy�"O��[T*��@M�M""!��$W"O��ca꛱iKZP�� hq���'"O�uǅ�\R5�T�Ҹ���j�"O"���A$���e�	$�:�0#"O,2@I�7k3���o�4�:��"O�	����1^Qw�b�"O�� �GH
dx�M��o�d��"OvdP�,qb,�kGK'�s�"O M�瘃p=�|S�Gw�1�c"O������k��l҉\��ر""O���¤ЕB���T�b�HE"Of�C�F&)����b�L	'��b0"Ot=���D:'���	G,�<���(�"O�xPC'�� :f�
��޹�p"O��%��?S9�k#��:K��M�"OPp�\���D�eŽ'���p�"O���'Ѝ?u,��bQT[*�"O����V�DF��;��ՉK���$"O�	�Ć8F
�����B�X��"O�4'M�?_%�"�S�g0٠"O��&   ��   �  W  �  �  �)  "5  G@  (K  �V  �a  -m  2t  z}  ��  �  /�  x�  ��  ��  F�  ��  �  M�  ��  �  y�  ��  H�  ��  ��  U�  .�  ��   b 2 Q j% �, ]3 �9 �? �A  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e�!�S�)�Z%����� �Z��I`n!�ͷ�JP)���4�H���,\��Z��(�*�-�pZ��N���V��YQ!򤈧6��r�7Lޘ�զ�]�$�O(L��fÇ�0�˴E>]��(�q"OR��х�=~�6l�F���
ٚ�"Ö��hY)F^L��!I�l�H��'G�����MP��SR&K!J� �L4D��xÊU�l���ᠪ�D�2�ے�2D���J�p=����ސ!�&���#=D��I�b�".ū掛�6�b�kf�r�����d�%��$h&��n˰E+��/�!�d�K�"H�&�%���s�'\q!�DؙX�^,p*��y�V��Şo!��0��(g�̏R�j�y�JA�e?!�D�-Qv��o=u*@�#�\�m>���)��Y9�һ/�����>ސ�a�;D���rfʣv6<X0�ڏZ�z�B͹<���2Z���y��ӂ+X�2������0HX���$��}it�u�$��TAζI�!���!����?@�hLB����2f!��7/���O
�/nZ�:e,L+�!򄎺o�~}��	=\G��aB�!�d��=SdIH!/M�E2ne��@�2�!��
�Aj�dqE���p=na!�b�#Z!�D���pu�$*L@�� #Y!�D��b����#21v �6���?�!��A Q~�y���*"�<����� �!�ʒr�X�Q����0�_�:�!�Ē<_����eb�
1�L� #�ׄ{�!�dTJ�D�٢5�y�ī��!�$�@h����*ZQ�s�ǩ>p!�$Y2:�~���Mf�W*�3_!�d��7VB�7�ݾ�*4��)�K]!�� v��d	�A� X�������"O���!H_!5�*�j���2��PKv"O�D���C�C�~,H�k"H]p�"Oܥ�Fe؋�P$`ū�	*��1"O�xX����J�I$	�"O"�ғ%�tQ�����mt"O~�4FO8P�=��@��l�Z@"O ��҃_	2fD	����������"O>�%*��TD�٘AiN9Hy\Ŋt"O���S��� {��H����"O���!!E�U�E��lΤ��"O�})uaZv�����y��8"O����!?��fO���1�"O����W�8����
���0"O�`A��Ch��#gk�:k���R"OFԑ���l7����CŪa�Pې"OF�I����B/�aZa�R����s�"O���eN@��U;�Mi �;V"O�eσrf�Y��"�	��E"Oȹz�m_�c,�����v���"OL�e�R.��Xa��a��M�s"OصJa��4xa�H1U�uj""OT[�d�ڈy�'�L�е"OZ=�Ҭ�kz�׻8J��#�ŞH�Q�0 �6\0J�{��݁gC剷!���;0mH�P��9�T�v�C��.nڨ)�K�'6��	B��ހp��C�ɳRox��ᐝL4�)���[pO�B�I�JK&a�[q�8�h��U�C�B�ɘY�$��o���=�����Pi�C䉢t��Е�]Gv��G��&w�C�I�P�\�cG�<'"���Q��
%�`B䉥9M$ Cb���}��D��^�%�$B䉪s�y�1
Ǫz$�aE�δ�B�I!�lP8�(
2~�e�&!�'gNB�q�>�@�@�:��������-��C�I9;)�Lq6�&( �4����9`�B�ɳ>������"^��(sLA��C�ɍl(�MyG�AA��"� �,®C�	
�8�ka[2la0�0PA�C�	q仂��;�J��E�A(�4B�Im�v���(���9)��ս-5hC�	-`��j����P$O�w���7"OB�:m�n�
7m�E�~�V"OVcv��+��
s�U�/��� "O�[mS=$6N��Ӏy����"O4HI�_4��i���Z�5�"OB5	�D<Y�~�+1bP)'P�y��"O��;�@�g�I���2c4~�p�"O؅�%i�_ΰe&�Kw���"O���� �f ���e�4�h �"O��2�ݼvW��bqEF^�>U"q"O�� *��q������uF"���"O�ay�Ӓ%�z]���ָ<@�0�b"OdE�*�q��5�.��A����"O^�r�JT��Dؘ�F
s���"O$��̩U5�p���`ihm�&"ON���ǅ�gV�1�C�E�8�2��`"OH��e��?���Zf�� _�p0�"Ov����->Jq�&,|��{�"O~��h~>}�&f��?���J�"O�I��\�"z�%����0����"O�������|�&��d1�A"O���F�`K��S��u�ٻ"O� �`�@dO�n���sȬX�ԥ)�"O���Ejɩ�9�@̇�*�(��""O��ZLƜg3x4a$�.*�Di2"OFu��Ü0�����k�h����"OHq�q!2�� 	q��K�V�[b�'���'��'a�'�R�'���'�������$e�� r����"R�'D��'|��'"�'s�'���'J�8
I��H�Q������P&�'���'R��'���'���'���'��Y�mֽN^zE�!n[IL��Y��'���'�B�'���'HB�'F"�'�����ث�ByT�]q��P�'1"�'�R�'�B�'�2�'Z��'?�a��m�&9H���"b�*��V�'��'���'"�'���'���'ʈCV
S!� ղ��F3��e�1�'�B�'Z��'��'�R�'���'���r�K] ~oxH�������E�'�"�'pb�'�R�'y��'���'���9%�#I=��R�&U�\��T�'��'���'��'���'���'�h�`Ŏ*=[IҴ<'�F\h��'Ob�'0R�'���'M��'�R�'A.�R
�-nt�ٱJGy��Q�'���'���'���'%��'s��'��e;�`���^����]�(9��'�'���'OR�'���'"�'Xh�^�E�h�#	�9y����'��'�R�'x��'R�"uӀ���O�̂�h3��J��
'|��X��Iy��'*�)�3?�0�i�(�[��&r�J��0']�M�L��,���	��Y�?��<���UNu���l�h6�Q�*#tq���?at�I��M��OT��zL?-R��� 9��A��M�����=�IΟ��'��>���p	�0�&E�<6�0��ƚ�M����P���O,7=�ʤ2Ё6'x��qf�B��|�G��O��$e��ԧ�O
�i0�Dحf���k`l�![��L�v� P��m���k��=ͧ�?���Őv�(����~A���r���<a/O��O��lZ;H��c��z0k�r�vI�Y�����m��Fy�	��	�<٫O@���5T}�Ec�I1R���񂑟T��3�Pe��9擳��Y�88bkgY�53 �����*F��Cy�\���)��<�K�:���7�]:l��*$HB�<���io��b�O��nD��|����	���O#
��P�����<���?	��Mq2}0�4���a>us��l�X�3�Ϻ:7�"��N9|��sī5��<�'�?����?y��?᧤iV�e�
Ӵ�b��eª��D�����. ����I��$?��	�0V�C���qB��l��la4*Z}��'TB�|��TF��N�9�⮄�y~�� ��>h�@(�i��I�T���!3�OޓO�����ƅ4)��Y8T��.M����?���?���|j/O�oZӤ��I�Y>��`��L7z�Np9%�\ڨ��	��M�N>����	ϟ@�i��;����@�V�5 �s��8aw���F�m�~]*��!����O��a�nB�@ڝ{{����d���y�')B�'h2�'!r��"{�H@b �_�`��c^.kָ��?I��i[p��O%�#z��O�z0]K� ���N�W!P1�D1���O��4�|��i�<�G��L�ǌ��u����ǧqR�M0qLӌv��X�����4���D�O��I�K&�٤a�s���Bz����O<�:���%/�	ן8�Oz��;S�)�B�ăŏs�����O0��'���'yɧ�I@m��ҁkY�vZ襸B��Qx��q� ��7�1?�'cn�I}��@���)�?$��e�^1���I�t��柈�)��iy�b�2�x�)��~�~a�F�F0Jh��#�(�����O  oK����Iğt����I�l����1�Zt��C��<�ɍ-�mZ~~�D2 ���}
���!Z�L!b�3� A؆���<�-O����O,��Of�$�O˧"Լ�[%I�87����� >P��C�i� �(2�'���'I�O���b��n�f���6"شw��Z�_3u�V���O��O1��P4m|���1k�"�Jʻ J�<S�i��� R�����'@��%�엧�T�'j֝ST,�\K�3r��U�� ��'���'�\����4%�X1��?�&>�<���ZJ0%��"U*�$�h��@�>	���?�N>�Rm�-�=�cHń(�5�˃~~2��	���1�i.1����'Y�;�0�-�y��s�+��xr�'���'��џ$贩K�)%\��E��B2���l@��|۴b��4z+OhPnW�Ӽ��hJ�d+.DC�M��>9�"/Q�<I��?���[䬉�ٴ��䃽oN��k�O,��rd���s!�q D�|]���ٟ��I��8�Iٟ���]����H�xlL@fg�hy�Dd��Xzr�OJ���O���H�Ď5�i��!)z����Ã�]��<�'q��'�ɧ�O���PiE=^�4�@���<̐�;�T5U�����4CF�ĽP���7�$�<)Á	&�Ѓ��f��I�q͝'�?����?���?�'��U��������и���/�^��R���{�.�͟<
ش��'���?A��?t��=)bxA'!q�6���GW7f��Y��4���G�������O�� L�cY�e�T���D�'{аQ %<O��d�O��$�Ov�d�On�?�p�A��*���$k B��̕ݟ(�I���2�45�Χ�?馼i��'Z���e���'�D���"�*4H ���|��'(�O��r��i��i����ש F���fT	�N(Z�`\x��i�#I>�*OJ���O��D�O,�2vIV����Ү�n�	���O�d�<�%�i����X���b��$��3萴���*veZ�pW�����@f}R�'��O��1Me��	��9S���j�����4%�"�^	3`�~y�Oe���ɔo��'%���eh�5����j��U���'���'�����O��	��M;�JM�<~n�i鏐0���ф�F�!&\P���?�"�i��O�l�'���`�z�S��фH`����,l"�'��H�#�i�iݭR���?I�P���a@�_+Hݡ�J�26��Ų�g� �'���'�b�';R�'��(��(�LB,,�e��ݲ6SvLbشF� M�-O��d4�i�O�mz�uZ1���|�d�ѱZ~�ɐB�Y��x�	^�)� v�rUl�<�R
U�;|��׌�2;�a�cI[�<�C ¯���I]�I~y�OF2J�t��Ų�I;O�<��Ue���'���'��	#�M�E��'�?���?I�&�m�j 
c��!Mm4��5��/��'�Tꓽ?	��� ń()0�Q� �]r��	~���' H�T�0-�ի��������'���WNO�#B�z7#�*.��g�'�R�'b�'��>����T*�� �*Rv��v&��O�.i��'�M���#�?��5���4� �y��[�W�$�f��S���r9O<�$�O����R7-+?�lR�2����D#a`Դ���S{�.�X�G�:h��1N>q+O�)�Ov���O:�d�O�$���2��:���n�΅2�	�<Y��i����&^�l�IW��Ɵ$��G�xIt�"R�AG!�q*��-����O���3�󉅄Q��c�{���Jg��6n�Hp$hj�~\�'���p�e�b?�H>�*O��*nìI%V��Hj��Xv��O��d�O<���O�ɠ<y�iZ�3�'ƅ�sń�;��(�[6,g��#�'f^6M?����$�O���O��Ƀ-h����*�!���#g�&;�j6�-?9#(��@'��I;���߱e��I��a�����Bax��x����۟�����l�	˟�R�f�aQaU�/P.)� �H��?!��?A�ib|���O'�c�ܒO�S�Ą�تOۉ\a�MEL8�D�O@�4�l%c�nd�J�`��$�
K�a��L !A;8S̍�F���IZ�Iby��'K��'����a�T�r�f�o�Jh;D�
7ur��'6�I-�Mӵ���?����?,���`��3&� c/�%3mz�a%���	�Oz���O^�O��?�6����BM(�f)^V�Cakf 8�!t�@y�O*���IhK�'�ny㖈V1r��eڅbT8v�-���'�R�'��O8�	��M�e��b���0�A)@>H#DQ�N�:��?鐴ij�O@ �'��FU�1|�!�4C�GI�t�W�F�>���'YL8�t�i%���a:�S�O��1��%��Vpr��5�~h̓��$�O����O���O���|jRcT��j0X��X�J�Ɓ�*�>��임r�'�B�I���=)�j�C�ˀ�cΦ-�F�v�\���� $�b>����ͦ��Fa���垪>��)�c�P�~,�M_n�B�j���'���'�r�'9fq���W�ll����"�MSE�'���'��V�D��4GQ
�
���?��+F�;�.�L�2]a�ރ�hl��BB�>9���?YI>TcǺU�rpґ��7��,���TV~�#<P��au�i�1�r��'��
�3^~\hdM�T'��3�,
J��'���'�b���@�BM���)�-6W2<9Kw����411�A���?i��i6�O��C9�X)r� ��.3���R�yB�'���'V�aSe�i����?�:����O�d,p�׺eq��Wt��9��B�	Vy�O��'
��'Y"��)`h�Z�%Z\�\%�&��<��ɚ�M���?	���?�J~�-��HQ!��/u�l��������9�[����̟�$�b>UK��Ϲ3�M����RPi�FI�ToD~R��%0�����$�^LT��=���Z�"\}�d���O����Of�4�b�?�r�[>�?��+و)�|�"�OS1.�ȸ�k;�?c�i�O���'<r�'V�,��� �C�^��L"1OD�la<�Y��i���<�qàԟ������G�V�f�Yu�Ӱv�p�H����V��D�O���O��$�OJ�4��
\�������#�����@���������?���`>���!�M{J>9�� 	}��˧Ȝ5	��A��B����?	��|�����M�OLũ1`3?T�G�N���}���#8���'=�'�	ϟ@�������=!ة�GH�o�*Ѻ���v�����ß��'��7-O�2����Or��|*�Ȉ,��G!H97�2��'gn~⭣>����?�J>�O"�D���L�!�~�Z�e�o;����O:��0���i>�(�'��q%���w�%"�`4�Cm�5M�� v�Q�0��ߟ���ߟb>��'��7-B3������_�z�B͂0�<Qn�	�*�O��$��a�?a5[���	#�r qS'�:<�ؚ���П�#��F��a�u�S"���Ay
� EC�L�v�B�x�8Pպ�K�6O���?���?a��?���F�	M����R2�,��a] �
�o3L��֟���L�֟X����s�iK�H��&�11�,8�HA:�?����ŞZ���ڴ�yr�߷D��A$U5b��x�1�y"N�TPE�����$�O��d5M�̜3��-�T\����P��$�ON���O�כvO�Ua��'2*��m��L�dPI��A�k�T��'�I�>9���?N>Ivg�#���bAC�=�$�)��P~�$�H�����J��O����J���$-���bR�KZ��`���y/�o4~e�F�s:�J���1�"�q�`0���OR����?�;P.���9�F�Af�<I��̓�?���?����M��O�<C���1:��P畗a����`���B���I>�(O��O��$�O~���O� ��k��:pb�q�#�=⺬�֣�<�i�j���'z��';�OyR�Eݦ��a��0����!B�H���?�����S�'��)�AҗJS
�qD���-����a�L0-�.O��p��?���2�d�<�K�b<���g
ې���! <�?����?����?�'��D���E� ^ޟ�S%�L�_�������>~��
�\��\�ݴ��'�~듍?�*O�y#�J� ���Ə�-$��z�ů��6�)?�'+�3~�����&����+�"5�D�`��7Cˠ1`2B�<Y��?���?����?y��tOF�p0@� i&�|bq�]�l�R�'u"hӶ,��=���dæ]$����E
)*��ùVp@��X[���@�i>��6��-�'d�����D���k�"|oZ]�ץ�3%"����䓑�4�V���O��$�Pi@a�aЦi��{�Z`*����O|˓sy�&
�?4���'�2�O*�4k�s�\��4eW>qa6m�O�y��'Mr��?������|���Q
��p��$S�М�1��Ȳ0��g�~����ܴ��$��Q��':�'�$թ$a�6c�5Z�N�/����'�D7�@"��T���^Cd�!�/�1�ځtu�ɠ�M����>q����cl�3:��P�4���7�Q����?I�È4�M�O���?���V���b�20�,T�b�݊V�x�(�'R"�'#��'�R�'��S��v��C%ߘ+vޑoAռ�r��4@����?�����'�?qƲ�yG��K�@k C-T)xE�V�Y�b�':ɧ�OE\}I��ig�����90��A9�rq���6��d�4O�{�'%�' �i>��I<���:�	!�(� ௝�aن�����H��ߟ��'�.6MR+A���d�OT�D��Dw���R�	]�"xQ�lɶ^�Z�ؑ�O����O&�O<g��(`A@�-IT���0Ý�Ȃ gې|t͘��u��}b��R���8�(!�`�Z(� ���T�IƟ��I˟�F��'��ÄW	#p��;c �yi�|7�'t7�#qf�D�O
�oZ_�Ӽ� ��(T�~�QE'1���L��<A���dX��6�.?�QlJ?M�~�)�(h.JQ���7�|���j8J���L>�+O0���Oh���OL��OR��ӥ���ִ��k��4�z�,�<�ҵiè�0�Q���	Z��hh�̋�@X��ؔ��X$\=� @���O���9���%X(�����A��!"���,�f�P�}����'��`�D�k?�M>9-Oܴ��#��Y���Ճ�5+wVp��	�O����O���O��<�v�i(�M��''��r�LZG>Ҹ�q@�((I���D�'��7�'��1����O�˓Q�rg�V-JE����qs�¦���M�O�ͩr�Ĕ��U�;�i��^���n�ʜ:l�TIt\=O��d�O����O4���O��?���C�%q���:���@s0�����T�I�T�ݴ<����O��6�+���R�����;����h����Ox�d�O�I�(^�7�-?�����( l��r��u��j��6�	�?�A.���<����?a���?�ꛒ[٫s���gI�<��1�?�����æ�HhIȟ��	���Oǲi���-�d����I�����O��'Dr�'�ɧ��ԜD�@��٥FpxrE�/^AL�9E�'�mZp~�O�:M���{�� �@Ѡ[��2�h�'�܍��?��?Q�Ş������	7���$U�1 ���Vh^,��)�j��Iß$(ݴ��'4X듣?��8Q���XI�>y�AP�9�x�L��Q�޴��d��$�$�[�'5�˓,�J�
ub�!�桁�EWJ��M���$�O����O����O��d�|�&��ex7	�.T�%@0%�
u�f�[`���'����'5�6=�,��KM�y����@m@��L"!��O�b>�Q�]ӦYΓwZ~Q�	[� ���A�d"@�̓`��E��OdL>�-O���ONXTLR�����b̘�ft�(`p��O���O,�$�<��i@B|8&�'+�'�́����p$xEE �!D.�2��$�G}��'kb�|�o�q%�5�A�=y�hq�B�����D��V�z�ˤ�M?$f��T���!���O7>��0¢�:���`D�|����Oz�d�O�D'ڧ�?�^��!LU�(��D���F(�����	��CHv2�'��6M"�i�a��&�r4��S�m�)
��d3�
{�8��Ly��VU�V����0h�4"���&$� $���GY'~l�E2eݸR�*�r0o;�$�<����?a��?	���?!C�˘|��z��E�yV��9���⦹A��[�D������*�J�	`�b=Ah #�tkE�=�����Ii�)�s��+�!��=ʗ����A���q�'qR$��'�n?�I>�+ODI*E-+��$��-S�#�nшG�'�J7�k�N�$�M�Z  pe����	�R��&��C¦��?	P� �	ßl���#�&isQ$Z6<Z�BS��e0�ȁ����'��c�j�I~���{% �Z�	I+I`���#_:���?���?9��?Q����O-��U ��]�~$F��i�<	a�R���I�M�3�L�|2�K6�V�|��L�r܉`P�چ�D��ė5J[�'�����d\��V��`1ӦܞsQ�phFjʨr�t$�Ɩ*&�1W�OԓO�ʓ�?����?��8��@��a��O�R��T��&��(����?�.OZ�nZ�n,������@�	E��.��.7|����C�:e��	L��dDJ}��'k2�|ʟ�	G-�'`�b��l�\��}ʒ)� XԘ=�ǎ�:�i>esV�'2*�&����?}�����I�Q�ԎO������ßb>i�'�6MT�\^`J� 
�n��Y�G�5XU<�;�E�O��D�Ӧ�?�cT�x��%Y�0����Xs� 1D��|�r\���(������A�'�z@�"\ܧ>`��SC�=�X��F�I��|̓��$�O`�$�O����O��İ|b��� 洒C�L���U*�~���c�Vpb�'�b��t�'�X7=���XV/K�phƍ�$i� i�x#��O2��<��	��itl6�h��
Ub@TD�d�W(R	jf�+�p��@EA�{��f�~�Isy�O���	�iM���&��D3��kP#$���'FB�'����MS���?����y�J,9����L�5k�Bm�1�?��X�H�	͟x'� xA
��+�>����rs�!?)�M��8�`��4�O|L���?�1�X7 �2HH�B�B����N��?����?������ϟ|�
Z+R�lm�&��w:�Ej!���T�ܴQԤ���?��i��O�n�/e��,!3��#v�T��J[�3��D�O����OB=J�Jg�R�+�rFJ쟀��R��](j	Y��s@hQ
׷�䓙�4� ��O���O��$Y%涔+ ��


@ɀE���%^����4 �bH���?����'�?Y���/��s��	b6�����[#��۟�?�|���׺1R�"T�Z�G��$���=:ʨm�!����$/?�� ���ys
�O�ʓ+t�U�E'�&DX�x]R*��X���?Y���?���|",ODEl�1:�xH�I�n��2&�Y6'�~ex�ㄍC �X�I��M���ʸ>���?��6}*��Ɵ	����r!ÅaR	9Í5�M[�O<�I'��������4�w���D���v��e.�Qä���'���'���'���'����PG�X'�6��%㌃��D�ゼ<��)>�v���t�'&�6�*���.#�(p�V�ͬ�i��B�1O,���<Y�C߄�M��O���1�Śe�:x�f���s|ҧ�iL�q��hF��ON��?���?���>u��d�E/M�b�zg��mG��S���?Y.O��m�(	�N�����It��	։u�,��SEY�3B`őӠ�����p}��'�|ʟ��b���/5���A!��J��d�W��/A�M��qӀ��|�&��� &�|��gL�#P �r�U�{%΅��@Fԟ�������ӟb>]�'.�6�W�y�V�12'K�\�Ɓ�Q�aN�����O��Xʦ=&�l��;����O�=P��`�������`�+�Y%�?���?��`H۴����6�&⟖��/O^a '��B�b�EJ�_�ܡ>Ox˓�?q��?���?�����P�@lh	1A DO����aP�n�nUl�$�'�r��t�'�87=�`$pg��_ ysR�6X,4Y��O��D2�����7�b��$�X25 �p��H�H�2 %�v� �Q(��)���<a��?qb
��x�L5�kT&P�hcM��?Q���?����d���U�5S����Ɵ�@�,������g�0P��lNX��t3��̟��	q�	p (�y���0|-�PC��	�n�`��10�G�h�|� a�O�h���vd���u��f��e��Βc�t1�ȓs�Z��m��4\��jV�:�P�K��J��VD��'�^7-2�i��h-!Ѫ5�II��ɓ�w���I�<��(a��1mZc~Zw^�����O۲Ӆ!�:W�>u�jI*5trYA!(Ic�	jy��'���'��'��E�9�����NF	w���E�
3�I7�M���_����OΓ�����57��hv���DN���ʄ*`<�'o��'.ɧ�Oj�Q�N�0����f�ܥ(P��R_|��V��D!cM�|��6�D�<�BAQ�:(p�nL'q�ޜ���?)��?��?�'��$����C��՟	�mI�+��������j�F]џ�aش��'M
��?Y���?9f�qt��ŧ$w Q*W>{��)۴��dD�t�&�1�'��O���N��l��ʈ!sB�5*ƨ��y��'���'��'�"�i���FEz���L���S�*@(n����O8��Z�0�m>���
�M�N>��۷g�4u���\�|�v9�ri��䓼?���|څ���M��O.x��� ��E�lY�m*����+a$��ˏ�~�|�W������	۟���`�
��<XAn#D`��������	Hybn���A�	�OH�$�O�˧\ �e�Æ6]fy��+^:욙�'Q���?����S��N�R�6�RF�ՔP�.t�!��+K�4�+E��o�Ze��[��Ӏ>p2�|�Ƀ)�4�H0y�$�I�"�);T� ���8�Iߟ��)�Iy�cl��ͣ��]�'�)�QN,� �{�F��Z*��d�O(�nZe��T�����Ա�� ���h2M�=~%F���Omyb��N��v������'��bMy�ύ
?;`AÂ��8`5�Q �Ʌ��y�S���I韬�������$�O����H�%�x��_';h�B(zӀ�[���O���Ol����Jߦ�]�	�8Q����3�������a�Z��	��@$�b>=���J���ϓAߐ}J�)ӄ7rm�vH�'2s�ϓ5��M�Á�O@|*K>�+O�I�OJX(�FZ��x�4�&	v@�����O���O��$�<Ҳi�>y�U���� #���W�L�G�͛�O��T�T%�?1Z���I{�4��Y0ȑ:A�^h"C�S�&�*��'��e�D�F
v-�AR����˟TR��'�ؔ��G>Hzd��+�7���0��'���'��'��>q�I,B���EE�b`BAp�@�s˒�����M��
��?�F��F�4���O l]�|�#Ȑ�j���b;O��$�O��אo�B7�%?y�-\?d��IϾ{\���w��"{���q�"�$K���O>Y+O��O��D�Ov���ONUZ�O�:74�kG�P�%�D���&�<Y�i���t�'�"�'�O���<lvb����|�r!*EX�*u�듈?y���Ş*���zP�G����S�$���9�jU��M+&W� �E��-W��d'�d�<9p�Z�q�.lk�N�>E�r�81JP��?����?!���?ͧ����M�W����d���	�������8HÆ�{��ٴ��'xf��?)���?q�	�)V��
�	����hx��Y�p��z޴��ĕG�4}b�O)�O�%(Vg��xv�·Z�h=(��^'�yb�'���'���'4��	�N��¢䏿E���p��7E�6��O��D������r>	����MsO>���N�p��"7O��ܓ2d����?���|r�� 3�MC�Ob�[B`ҁ<����č;��4��@ȝr>���KAޒO8��|����?���-��{#!�6�D�񡂽u������?A(O�n�%��ß��I{��!�ek�|��\044E"w�'���{}r�'��O��D\~�p*F"+d���L�4��=@��G5�T����cy�O�LH�	B��'�Y	6��y�f��Db]�7��Q6�'�b�'\2���4�'%�dsCV���ݴ3^� f�F!F�\S���N{������?��'��V�'�I㟰��O~���yr)	S���b�R��������O�ёf�j����R���b+?I`��06$D�ZAK��QGx�'[�<q+OD���O����O��$�O.˧��}{uoћD��@C5*F!3��" �iW�ms��'���'1�O��Gg�󎑦r:���Oߖ��Ysf_q�X��O��O1��pJƄs�*�I,���lZ1�21�Ah^�0�x�Il��1��'���$�$���Ɇ�u!�D���`���Ss�J�/�axb$|�> 2w(�<��
�"���%�E;(��`3[\nŒ����>����?�I>Q�#��&��QQF/��C�~��n_e~��^(a[&�ճiA���H�'�R�Z��.����[���4��y�������[E���;��T
WBmvӀMI�H�O�����M�?������ W?��1��kl�	����ܟ�����⦩�uG��l���OUM��A�����1n�1#�q%�Ĕ']џ|���iS� BWk	�
k&���/?���i��0��V� ��a�'�<ySaH31;p�DК�p��[����ߟ�$�b>e��a��B�r��=y��Q�k���.�nZ=��䎺s���'o�'��I �ȩ"uA�h�,�0��.E6���Dʦ�# �Oş��l�s�Z�!2�ɂKS~43+����y�4��'Z���?i��?y�ˌsg��^9�P��U�j-�M��Of��Wo׮�:p�:�I���q���v�``
$(�9�>O�����kBͰ�e�:�>�Q��w��˓�?A�ie!�Ο��m�K�I,K�V4 aĝ�H�±h��;Z�F�&������Ӌ(عlZM~��^<1��i!ġ:c8�����KN>!������*�I�z;N)��U��R��v?�#<y½i���1��'-��'y��*G:�Li�M(~��tgκ\��N���ڟ��IT�)�� �mr�O^�`q�����ٽM H`�a�I�Q��J,O�	5�?�W8�$�+QZ\&��/�(;�Z��!��禥83�D=� ͓S��|D��K��H`�'.6�2����$�O0M�c��}�����?��)���O�����7*?y`�	z���iyIͦX���$��9k�M�s)W	�y2[�����<tS���&�567�0	� |�x	�޴.\���.O��>�S��M�;t'j}#�Y�`UД)���!2X�B��?N>�|:�8�M㛧� �s��Q=ˈ���"��dߖ���7O�ӳ�Z��~"�|]��	ßt�c� 4�|!�Gf�?E6������͟�������Fyk�T��#�O8�d�O��Pd� �hp� �Ap��s��;�ɘ����O��D �d���}bd�`�Y�CF	(s���)�2�
�Φm�M~�L����	3�]���R�Ď^�([�(�I�� ������y�O��o��E찰���t",�ӱM��'�"��O�%Hw�'�rLw�j�杫p��{��P�����ȏ0c��	џ4����c�,���)�'�((�c��YZ0��Y�p�І 5 �0�	�m�䓢�d�O��$�O�D�O
���>~q�a0	�/h�@� 5g�&=�˓d����!9�����'?Y�ɭ=t���ɓ�$ 8SA��_��(��O���O�O1����ҤE�T�����#b	%_c�7-�Ly��CX*������DB&,z���rjOdw�����9eP��$�O����O��4�f�ƛ'��(���5�a���+-�V4�#����p�r�4k�OP�D�O�Ǩ?�v<C���L��Jf�ִ%���	iӲ�ZӖ�@
�5�N~��;|M��YVܒP/�a�X	���?y��?���?!����Or� ȱDQ��$sA�զM��g�'Ib�'�<7��_��	�O�mnZi�IN�\�"�[�*�>�벎�CO�\%������擵ya�n�r~Zw�\aӦ�B'N*Dղs�ªĶ]h1f2l�B�	sy��'���'���WD�����`�p �1����s�'#��M�E��?	���?�)��){���=I��Uq�K��\x4R!?OJ��W}��'Fr�|ʟ�<!ԃ�.��"iڑ%��8t��o=�pk�J��+F6��|��M�O��N>�Cm�4H>h�BT�@s~�@ש�?1���?���?�|�.O��o�BB��W�K:�<ܸ1��j`x�RR�ڟ��I�M[L>ͧ7���:��@d��XF�q|�ɂ����� �I��8l�D~�(	9/�A�'��&��E�jl6�Il����;�̭DD�Y@��>՞] �	�)U�,��G�~DF��o� 
զp{��!
U2�y�(�6� �:e��%��R���ԁ�p�'�p=Q��Փx�hԹ��H6�Q)�Gͪ-�z�)D�%&�Q)$��$S�|z�.єl�8t�#�ԅ�.G���ґ:��	�*M�W��00 ؆8����b�G�Z��t�eh		������3btI4(H�C�����߈$�!��B�d2B�� ��H�AC	>�x`��$
(��l�ܟx�I�<�����d�<�d�&=S����A��(B�2/,�fM��VҖ|����O�L�����p#���oE10.�@��ܦQ��ҟ�̓K����O���?��'׮���ޯ6��s6���%����}2�Ak��'�R�'���;\:���N�va{��^6�k�p2sAn}P���IX�i����ʆ �p�2�V$|;��еb�>q���?A+O\��O��$�<��ҜJ;v�9��	�H��}H��8]���S�P�';�|��':�L)l�x���M�R�01bt���*,�e�'���ɟ��I�$�'�䐣�b>1�J�rh��M�d8N	GI`�J˓�?�H>��?�Q�S0�?��b��d��h'$��<B�i�hN3��I������\�'mL�)�~��d��e�R�0=@��@dڽ7�Bt�i""�|��'#�
�qO�"g��s$B��T�2�PB�i�R�'i�>]�1(�����l����1�84��!O*.+T�(BAP'�.$������ɄaXş�$�P�'D�ea0�>F:��`1,Z$y� �o�py�d�a!$7-�O���{��)]d}Zc `�C�o	G��h��hJ�u�n���4�?I�$�%Dx����I"��FϚ�&y�,�6��ߴN���p�ir�'-�T>�|y�!��M�����vMݡP/x19c�i;��Q��1��՟Xz�
4���s5�C$�̉4֋�Mk��?�'���:�\�ԗ'�B�O�A��[�`An��F�h(�4����č2�d�O��$�O:�d,%�������H��r��}+&inZ�<-��C�O,˓�?yN>��<��e��H��8p�L
:XR�U�'��y*�|r��5�4�?�*O� ��O�-P����<YNH�R�^�V�İ$���ퟄ%���u7f^�p�>��ΔlJ6��T��M�����O����O��v6F�j�5�t9��+e�T��׬cs��{U�,���'�(���4�'�qɑǛ�:] �b��D��n&��O���?i�A\�����O�x�E*�1*��<���9p:���mΦ��?����Ɔ�'�ű��q�^h�F�.	l�ٴ�?�����D�1�2�$>����?ט�C�&��qc�4!êai�* 8O�˓�?a����<��S�QأJ��;���Zsᘢ��t�'�r���� x@B�'�r�O��i�Y������BY��Vv�숚�lg�T���<ᐨs���'*�`���mҾX�<�8�J�P�im�(�����4�?Y��?��'n����$�]
0*�YE+�DxUAħ�X��6-�O4�$�O��O�3?ɐgӱP�dQ��@�.�����o����v�'Mb�'�yBR����	�Z�#O�/��T�1)	�lD����dWl��?i�']��{U���zu6Hr��B�t��ܴ�?�禇���dg����߫y�-ƕ[��� �: i�u'���w�;����@�'���+� �p�26 ,�S��֎|�$]�d�B����O���;����x�������Iʞ@���x�"O�|�%n�
.��?Y��?�*OҀ30���|��F]$cJFf�W�*T�A-H}r�'b�|bZ������o��a�z
s���@鱮9�'�P���I}/"Y�O
"n'[6���	�gDB�R�I�"\,6�.��şؕ'��<�N<Ӭ��Ur"��U�W��r�h�æ%��ky��'O*�`F_>���͟��s��9fo�0l�Ɖ����voT�O?�D�O�ʓ�x�DxZw���q��ְk�f ��Hז'�l
ߴ��D
�9�(1mڷ��)�O���S~2���BaF�17`�"!G��%���4���O��$�~�Sm�s�<,�!�΋K�䑙 �K���`�i.!z!cӮ���O���'��1�`��w��&aN c��^���4�?����?1H>����	�wI�P�"�(M���VE"���lӟL�����z���}yʟ��'Z��ւH8q�
�Y2�R��VJ2!�O�B�'U����:0�ԃDDL)��C��6M�O(�b�^V�i>Q��}�I;�����!~�W�7L76abs@;���O4��?��?�(O*y���!)�������m� r�����e+���O��+��<��=[��	��h���'�\�I7��oʟl&����\y"�'$l��ԟ����
Z}e�$�αaA@��i���'��O����<�aU�ɛG@W<&Ĉ�(�� (!��P�B�>���?���򄑑:Dl�O$R@W�,�, �a$S�0�o��5�6m�O�ʓ�?��?�ŮN�<�/��YH�N	� 3hq�p)kL�����٦i������'���X'j�~����?i�'-��a@lX2?Ǣ�gi�'5|
mz0V��������I%�$���?Ѹ���!~���G�P� ��!Q!e�˓j �5�iV"�'��O@��Ӻ��-E�
܂*E�U~r]Qi�¦��	П$�W�m���Jy����3$�pg��Eb`YSdO��f���D*6��O����O|���E}�V�|!!��,���t��v!҂����M+5F�<���?����O��C�5�\93#��vǌ�;�#� [��6��Op���O,��r�J[}S���	Q?A����A���FO�%s��Ѧ%&��pe��'�?����?idAM�;����"R��3�/ٛf�'��Ją�>�)O���<���kn�	};� �P�]&n�ց���TK}2���y�^���럈�	zy2�*ˤ���$J:�����ݦ:���K1#�>Y/Od��<Q��?��(�M���J�k0v-�̘G��Ap ��<�.O����Op��<y�iVs��� �]�PQ��� Y�l��,R���S���Iiy��'��'�h��'9���K�.C<`�CH��O@ v�>����?)���d�fy�d�O�KG:h��)���YƬ q��'�7�O���?����?16hT�<)H��P�c���v�z�
;8?:���z�D���O�˓T�,��V?a��ϟL��5����,�'O�z͟�A�&�a�O���ON��
�`��|����D�{f*�)3&�+���A�Ms)OjT���V��M��ɟ��I�?9�O������9�F�������(��'�囘�yb�|"�I�5n���J��@1.��e�hX�(Y��JåZ��6�O*��O
�	B[}�Y��Ô"�{����M�z���a�Mc��<yN>I����'@<����W�<���L�
�x��n�`���O��DD�:�"��'��П��s�/��$j��GD���'c剫.b$��|b���?i�A�"e�a�n>hI双(Z3"ٓu�i6B-Q�����O�ʓ�?��"Y8�q��$��,�&Kj���'j��'���'�"�'Y�^�Ps7�P2J|4��1P"�rd��Cٿ9�Ÿ�O���?)O���O>�$S�3��d" ���m��(�*�*�>aɲ�� �	����Iӟ��'�h0tgk>a#v)\.˺e ���� �f�����,O��<���?A�"t�ϓN���4ŕ�4�D�i@
��'Ø�QD�i��'5��'��I�)���;���DӔ=���%���J��ЮN��n��ؗ'���'�b�8���M��9NUز�2�ʩ�2���%���D�'�B(x��~���?��'0t�Xy�F� W��˷)Q�|�V�´X� �	����I�6���IQ��'��)�.`����և0��a���v��vS�#�(���M���?����R�X�֝�{��Y���� g�ڠ� ː1r�6m�Ov�dK/o��dNU��'�q����5��%Hu&,�@�؇
MBXE�i�����n�L���OT�d��r��'剠y�hI@O��Gr���q����Hݴ-;(��'N�IV���?A������D 6�A!"�8�֮:��f�'��'�$����2��Ob����0�5&\�5ޕ���!rdeҒ/k�ΒO<�r_V�ϟ��ꟈ	��Ǜyt��)��I���F��M[�ӂh.m��'n"�'�ɧ5F"�:,ބ��׮.\B�y�a�����^��D�<q��?Q����dӉi�܉c�\�R8FT���K�u'�X�U�BH�֟T��A��֟P����ʨE(;:���(a�'O�Xi����J�柼�	ܟ��'�½j%�b>ݳ��ާ;\{��C�Z�x�0��>���?�O>����?	����<ap�åy'r=�g%�W��&�;pV�	����I����'�R��w� �I�I�? ���g�<o��B`���y�&�i���|��'���Y�y�>�"I�	|�M	O���Q�R�Ц��I���'
~P���#�I�O��I�����RnA+ML ��`�F8��A$�D�I͟�@��ޟ $����R�	Yd`>$�8��
ڜL)�,l�vy"�Px�6�B���'z�h.?���9�d�Zr��:$�ƙ	��Aꦕ���X�Ff{�4$���}�cJЙh��-�E��j�j���e�����0���MS��?��������h��f ����R�G j��nZ-tN��q�	U�'�?Yê�4�=BFBïv�9�� ia�V�'���'����B,�����2���3S$n�4h�w&%1�m��??J|���?���~�td�.�5m� qs�ϓnfPx�i\�)˥nV�c����Q�i��r�EH�l����2<��h{��>y�l��?,O���O��d�<��+u���J�Q�z�(\�aeS:M%�����O�Ol���O��G`>&��Hg��-5��}@C�#Z�ĺ<����?���?���_�<��e<J�AЂ+V���e��.�5���i��'�|��'��Ik�7�S�8b�1�!�ȳ<�da ���u|������I⟬�'�z�q�~
�8bDً o�e#h%�$@m �l�i���'��O���>�ɖ!�����铢O�d��C�Z&?ٔ7��Ol���O��֗VC���O&�x��	�?\��ؐAX+8����ᕆNR�<$�0��ky�9�O���8B��m���,>�$�Y0GZB}��'�
�@��'���'���O��ߟ0e�"ҟy��m2CY�,M΄r�i~"_�����+�S�'+(!�່��EbE�?@��0B�i��``g�(���O�������>1A�J�x>�Q� E`��,1�Ƶ+�a��'�|�qJ��C3�pAg�*K9x{��v��D�O��$�9N���&���	ʟ��L4 y+�AFM'��*e	����>�p��v��?����?��-݃UE�I�O	���I�G-��t���'��EH�/�>/O`���<��[pI�
8&!�#�(t�%�u}�ሁ�y��'���'<B�'�剮+�
$�2o\�H&,���b��*�q)C�@��$�<�����O���O��oHKÀyP4!��h0��3�1O��D�O�$�<q��W�~L�IM*B:*����ZPpޭcg HD9��X���y��'|�'�8�+�'�t��� +'ؤ�T�_(����e�����OZ���O˓7�xxj�_?�i�Q�a��}��4�O+a��	���e�����<��?��t4"͓���2U�&���
�()а���)8# el�͟��Ivy"#A<M�p�'�?!���c&���a�A�]�j�e�	�#��I̟��I�h��j�Ȕ�yBԟp#qH�R^��W���h}� �i%�I�k9܈3�4�?i��?)�'��i�U��ޓ~h�A�7#ɪ��X@sGv���$�O2���7O����y�Ɂ:i|`�;Nۜh�u�A�Y��6�_�uj�7��O`�D�O�Ix}�[��㳇J0���c��U5y.2�*`J8�M�����<�.O�D8�����3q��zqM�6t��B��	�M���?��� x*8��]��' r�O������v����P�v�rL���i�B�'Qr&�,�yʟ��O��d^�
�"����O�^�J7K��f�<o�P��K���ī<������Ok�0l=T�Zs��
E�z]�aaθKț�'ܸU�'8R�'؆\[v�K���\��0X��(�@���Y��'��d���Q�;��H�0���j��X����a�3o˦8���V͌�,��0aq%
-<J���vt{�>ڄdA�rk� b�'��z�h�b�oЦCT>���';��7�bN�N:�aK���Ѝ3IN�Z�A�WJk�\�۱��3E�̴��u�\a��*0�h���L�+
ՈIZ^�m��H�����슰�d�1�i�,��A�'�b�'�V�S����D��ˆ+"��̑6��Zb#�!Kb� �VЅq	8���C�'av�)��ҩ|� �E���Fn8�Cǃ4]:�n�9HbL��!��>mU-���B�'�j,���?A��Ԯ@2K$�d��bȞb��UI��>�yr�'����.�2@�Q�ա�<:�B�a�q��'<!���P*4�+��¤&�t��'<��B�>����I����D�O����fq�f��{��o0�:5	.��͙e��k���O��u��,�v��+�j�Cs�+<t@ ��,ҢCH���� 7@4�PQ�"~��_����ΏN���& �h�}�eȝ՟4�IF~J~jI>QG�Hr�YgґB\q��	�^�<����@PH��fC4(� �14dv�'yx#=�Oc�# ��T�fe�租0)�(Af�'%��Yߌѐ��'j�'@�o�9��ޟ�� ��dH�y�3n3$v ��Y��?�tb�=	��ra	i-N�3ړ@dI�v
Fp�pQ���gɂ��s�'��I��B6�IS��QF{B�5���B�V,-�]�u�:�~b%��?���hOJ� @�����Lǂa9ă�=X��ȓp���PE��g\��13n��"�]� �)�.ObI
g�˦�"Ti���z�c�#��h��8%h�T�	����[{F��	֟�ɚIftP��!J�<��/F;�Su��[@<��U�!�Oी��Ӊ=;>�� �h��640<�%%�$~�4Q	6�O-���'�BjG)v+�0BЀ%�kb�/J,�'�'<�'�Ou�T��.�r�q���Q*ٔ��'(|leG� l�9	�)^�"Np!	�'p�6�O��]YL<Γ�?Y���雳-�`� .Q�zxN5�w(f��\E��O���O}!���A��	'�ʧ?q��n�;c�����G�1u�Fyb���L��p铀m���aF�P)4
�NK�)��<�2�ݟh�I��IA��J�Bq�uX� �$4"ī�*C����s��k$��|��!	G�q�l��b'�O�p$�����1���B,��v�"0�9�H��'I�U>�և�����ß�ke� JH!
�׺bi|ܹ�-�?�PȠ��?G��ӧ�)1��O�����`%@�j�>*]��[hޛE1$ ����S��?�'�ͻ]�����ŧ}�6U9��xؼ���?���?����'u�,Z��0D���]���!�W�y��'\�}��hUt���m�<Jm�����Y�O��Dz�P>Q�s��
8��2*� �,�����Yh<�Ifv�ȓ�EA�k�@n�<1���0۔P��"�x�aj��Hk�<��F�� KV��;�~�@Ck�<!�J́VsX(�FٍݢPxq m�<� דO=�ak�j�.������A�<��kU���8��/ۂ�6t�עA�<�o؝�F���f(>;�I6��O�<��!M��<PS���% 2<#��E�<9)�z�aa夋)!g���%�~�<!WkFa�R�R��x"\pJ��y�<�'޶ffhe�s$�#&~j�c���u�<�D���_� �H�A^}�mK2��k�<ɡ�_M*��e������g�<9�Q�_	.��g�}�^�P"��`�<��ØF2�\	�b׺o�n��&�c�<Ⴊ��\<�@ȶ#2��fDy�<�膴3O���%
1e��	[�%�@�<a�����!�&
�)r�H�1�I|�<��W����E��2L]c��u�<�Td	:C�jh���L�W��:P`Sp�<)���t���U�N9A��B�8D��4�U�c%�H�KVc��i��7D��F�ͷy�@t6�Ľc�}��6D��
���B�`Ӏ��kCH kR�0D�P��'N�1།ڲ���>��u�,D��
�m۴0�x#bk�Z-p�S�4D�����[6�l���l01�1D�Lj�`ƯAR���.�ͪ�N*D��E��&&ҭK���|��<P`)D�\������	C����`�(D� +R��<e��*��Z�_k.1{�%2D���g$��.��ٔ��W�ER`O,D����K�u�⼸4.E�Q�����%D�����$�P�e��d2�9��#D�<��/��,��XM7��d�7D�,��&]2f���I���א0zD�1D��R�L�_���^y6��(P.D�� G���WFE��}�䝣�� D��ӥ�FP"�L�&�zYQ��1D�g�øP{�S�	ŗ1h0�w�<D�  �Y��������g>D��8�H��*y���߿��=��;D�!���X�D�]@X���8D�$���G�%`����ܵ7��L��$6D�DK���=�Xd��,I�I�s !D�,�
L�y ��[j�xk����1D��0%e��#��\�qi�^��y�..D��S�	$��
a�
 kzY�Gc-D�� �L� e��f�x�z0K�(�F�y�"O,�c�.^�j=P�j��fKR�#W"OJ�sFW�7�z|Bđ�[3P�(V"O<�ZD�ڎܤ��b	Z/�}ȁ"O虂�fނ���⇺J>�D�"O��R���d�D3�A�-ބ5��"O&E�D�M�̠�r�����R"O�HQ�k��4� S��h\��A�"O�|���.Oo�H1�.��r+T]��"O@90w���C���E�V�,��HW"O�AE���Xy� t
= ��""O�2�B#]pp�W��Gj�B�"O��[DEK�<W�xA�Ą��	�`"O� ��N�"-\X�p�'�7}8��IE"OR���$�����'%P�X�s"O��J@A�u��8���,[蚲"O`���ŠK�"t��15���P�"Od��Q�PR���bĵ:~ؘbg"O�1Hʍk�����	e}I"Of��EH'[N�(�1�Ń~gbp5"O���,��d�H��B��6zKi�"O����$D +!��iA�*5�}s�"O:�a����ȝ��B�s)|m�e"O-i�g[�:�������9�*� ��'u)v���,y �h�($k��0Pg��îC㉗�l��틎J�����Y�Ejc��Bs�XZ}��7kWdt�~R�c�F1�[q*U�(�P�d��k�<i��μBX~��M!�D�*�c׆��$]�X`�(�޴&0fLF��Or�aH�3���x©A�d���w�'�YBFǭ<�����L�t��Um�;z��@�k�PZ�S%�1U֘�c�*��<�F��(��ѹ��_�Obd���.ZO�'0VD藁�0����g��z��pgM�^Y�y��%�0�C����8:F��Ҏ��$	B�90Sx���	�N�H�`�	���C	$|Kl��r�9R�Z��f�ȹZ a����WH�b�)����&xC|�/<�A+�c�F���I�Sq�C�23H,Ɂ'T�>H��阚�b�H-ȃ#]
*��H�E偨j�	���Ţ|�Ҥ���$[\��6!~�iR�N��2[k1.4�|��uB�(S���-�T�j�D�"측F(ͅwO��!a�߀f��j�ʟ9*�]z�L�<R��-h�\�B��Gx2*�9�H��E��1S��}{��� �OVu�cM c�"����
�f���l]�ArF$s$��)@$Q��B�t�n�3�E^/I�^�тD'\%�8��'�"�{��c��H���� 
�S	�P�6jR0k� �IG�@!|O"�y��O�$�I��5��w��v��pa�p!�Y��Fs�<�0��P�p�y$��4#�TU���Y�HS~l�
��g�L2�@L')Z���0)�z"��C�T�'[n�	e�\ '�����;(,��F��x؞��-tV`|��K�=Wa쥀5�[�`�ŉ��!Ɋ�8�DZ:8����@�x�������<a1�PMQ��q�T�I��H�')H̓	�I�!%8v�D�	�/W�H���8�b5�@�:2.�𖊘�V,��/9�ry��G=Y���$�#;֥X�mF�Y�<��j\�3�"2�oE�u�U����3-�v�P4c�v�I��ˬJ3�iL�S��
eVHk`e�73pn�8��L�8�!�dΊC֘��th��Y�P ��D��={b��o�����Z��H۷oު��rd��9��I��SpO�4��1q ��tT>���2\O�hE/�/c���BB�!<efΏ�yR���F��8t��C�!f�ɛ#X�)T����Sg8���D�RH[��0��
NQ��8�	�E�Yi`�ZTbA�vf�Y�V牅6@V\�G�/t������!t7G��l]�
OP0���
�����~S��q��| �@s6� ��� �3�Y}?����M�O.4�݆@oF���Įz
��@V�ڶD�C�	���Ȓ�1u����$
�d����>?��AY4����'�� !�&�S� ���Q��ލU0h�P��7}�ȡ��<��@0
k�{5���2m��ac��
!��{'���s
�(�N�9v���&��7��x��(:n}���6Gd�Lb��R-�OT�A���.��pa�-ȩ����ڑ#82}�� a��)(��ɨe��]�"B�I%FwD�;�B���9P$['0MZU`pO����A#᛿CŲt ׬%�)�;h,(�R/�-4�^�bIбOi�����	pS���b�*\h�⍙n μ��&�`�@�^瓻2�YP�RV��u��%�E;wEJ��쌬x���Sd �N8�\�G�!|��Vm� ��Ӈfݔ��4!:q
lxVm�=��L��I=�Ҡ��І�p<D/YN���%�E�,�E���t�':�M@
Θ��!�U�ljD�.O�y:c�L[�Z`�͜ZeR�3�l(4���˂�K
<��=Nh�ba�Y��Ò��<��}�h�`e�I�?�D���Oq�kL�:r��uK W<�X�J^�z5���!Mi���TK��A'T�|����<��ӂC>}�ȟj(�{"����B�4}��A�
�0?q���PI�q��8!�b�s� �8�h�O�QG�$&�Of<���xtd0�FG�z�B���>����f��d�3p;n���HW&c�t�K?�a�Y$�[�&�oj"�7D�h�M��&���*���/s�h�H��4�¯D)�>Y�'�Q��q���Ơ�a?�0m�98cF1�L_�Pޑ��@@i(<�6��8e Lt)�mN<6�m$!ְ>:R��ʥ>�ud� I1��ӕb�0��O�� X��Q�G�,�� �
�p<14F����y� �č&s�ay�ԑ/����\$ \�Ac6�-�O��[�!�;D��4��,�ԉ��x2iG1JQ�O  kì&�OL"\�c�C	y�a� %Q�n\)+	�'��h �)�h����(:p�y�'6��9��	~�2��E_�
�5�'(�Y;��Ҍ7.�h�'^h��'@$��2h"m"4��� ��
�'��a�k�L�������0	�'YBЃ�K�g����c�׌�LX��'�jth� ��G����T˼U��H��'�vܳ��+?�����	�v�:�;�'s"p����Xu���ғ{�0��'�R|��y�e[�d�	���@�'�0�hL��.P�ĠU.U��r�'�����Bgn"%ѓ#��6v����'��ٱN�4��H��(��@A�'D����(W�l�����&���'FH��0
_�S��@���ժ�6��'����nC�8�@�V�ɛ1B���'�>0�⤑� ��C5��#.���*�'��Y�"A(,TH���֨Z\���'�$�`Ӏפ�:�B���Td��'�4�����\Q8@��+�"T��'S���Β�cN�LC�拂L�hA��'SQ�@a�=J'�
s�K�71~�
�':�Ȇ�2$��!�'I"�H�'2�A w�ܐC�����U6%;b9��'�@�J�NS�jk�1y�M��4\��
�'� �C����jăP�'W�j
�'g ���+�. �H=�W��(a�	�'�葋D�O�Q g���
\8	�' ~��+\b�F��G ����	�'��T+���'�����	f �k	�'nE�c��$&�Q0g���	h	�'��-ʤOV?����s.W�5��'��Tq1ԙ�RdZc��&�����'(6a�QFH%�Hi �͉%K����'���q)�11������,J��	�'��L-UyXU��cX$E|��	�'G�U Q����MG?5S@T1w�
��y",E$�h�Z�>!X6h��^��y튔u�P�jV.I�A�6����y�BU�Z�FD��OA�@�F$��y�I�%j�4����A4N(���@��yB(՞R6<����,ɔx3'H5�y���LO"<�bY�ta<%�A�ަ�yb%H�PBC�7�N鱡
�y�ۯ$Z���bܾ�����ye�)2�+�(^&|Y�O�1�y�`��0��iWNQ'���E�y
� ��Jt?r�&,�'��v�<�9�"O�!(v���WV(5��cՈP��"O���ǦC �Uz�j��x��"ON��S!7 <(%��#yH���"O\ͪ�ǋXIP�E,}b�t27"O�a2ƪT(*��+� �c�0�"O�=��m�����f��`���"Oz�U�L z1���]�"O�5����9?QԜ�U�'|���B"O�xF�< I,̀��u��|AD"O�{Eɢ�"-%�E,(9�IQ"O��8cO�.x2a7F����"O������Ao�E!�[�5��ѣb"O�y0ց�%_������"O�܊6�
9CJ�3jG+z`ـ"O1�d�1m岁A1j�&-!j(9!"OD(�#JPA����"��>���"O8- tl�4��D�3BeV�pe"O�d*��%�a���	:,%p�"O2�KaL�<5Y��sa�@�&fm��"O0@�RMU�m!N��"m�����"O`����7KZ�c`�툅j�"O����B�j���u��2I����"O@8�1$��~�j�)4X�b"O���'ʐ���%1gI��<�nm"Or��FeO�uf2���P�@��9;`"O��B!�33�i�A\$/�8��"O�s�/�{fA�1����e"O�Q� *R&Z�hq��[��r"O`�VM�&*RXs$�s�r��"O�i�%j� rI0L���J���"O�0K7f�u�N�Ct#(咙" "OHxZ(K�� ���͒z��r�"Ob���T�"��W�c�H=�Q"O�=b�	�cp�˖ˍ�4����"O��qP
:V�~�j5�P�O�\93@"O�1�'�B�=���jBN��>�D̑�"O���W��J)P���-�: ����"OR�G��'��c-�tZ I"OHa��#
y���l
�,H�yQ"O��#�#�3�έ�UEP/W�xUB�"OF4h3��-O�t�:P�N�B��P"O�y��l�ZeD<R �G�nc�h�1"OA��τ-n�]j����뉷Z!��U��|���Ӊ����#,XI!���
�P��K,��ȱb�7/<!���!iEG/+��-�����!�DS�Y��[��
1�N�q�­{!�DL�Y�ث�Kɍ}����Gׇ8c!��K�ka�\i�l��e���	�G�!�d� �p�P�M'F����� 9�!�\�K<�ۇ�R3h����%Kp!�D<8H�(��ē�HH`��:)�!��5. j�RB�ҧ�\���ד�!򤙺Q�dQE�
$f��	�k�iy!�
M�q�7�]9W;D����n!��A&Dps��$��ݹ.ͳ|�!�$O�|b��P&�	gzt}C�'Rf�!�D֕]v�Р'a�e�b'��#)�!��>?��<{AkӥGd�qr��C�s�!�d6}�x##GV,Rg�4a�)L�|�!�D��U���y?[�-@i����.��$�(<��QS�i�J�E��~�f�aeȖ!"����Z/8��%��S�? �C���{�ac刟4| ��ږ"O��*��A�%�ɃtA�9� ��s"O:��W�x����ʤ�a"O�*�G�'�!����I��q�"O0ȃ�!�w
R���9�p@E"O��z`A̙m䬥y��٩@����r"O �����g�ʘ;q�ɯ�Ѕ��"Ov$	t�R��� ����;)��"OXUȳ��(����0�C��U�4"O�����.�=iE/�j���"O~�i���	8FLc'�f�Ur�"OlP�$��O��z`�	�d6f���"O��9��R� �P��5ΝX"Of��e#�
~�1��[N�q�"O�`��ePF����r��'^A^p�"OhM���a4,Çn�A)S�"O��'�s�ڶO�:��<h�"OV�C���|�<`�N]�'�X�3�"O Y"ԍ�a3T�*V�C�g�8�)�"O�8�c��e=����N� ��T"O>kl�Le¦�I	g(豈*O`($��6m\
��"O������+Z[��x�ϑ$tx�"O�$����[�LDh��X>	(5��"On�c���)vP��6I7�<�1"OB��h����u��;j��`Y�"O`�+	�3�4D���
�{zX8!"O*C�AYp�&L�9d��D!3"O6�R��~��`�� w^��y�"OjH���=9q�1e�w*�x��"OF�2bJ�%�A�A�S.���rR"O��3�O�>>ꔙٖbb�i��"O�| �b��u��(QA�4MС��"O"���F��3�H( �=�f ��"O�\�p"ܩ ����a��qj�!s"O�Q��퍗sq��i�a8&�C��y�,�-b��	�IӨe�P�YR�Ϯ�y���93���F@N3]JV=:B�
��{��\�S힤a7�U�x2
b��D{J|�V%
2�\��6(%���C���H�<y�&؀g$�����rb @�SG�<!@�ǲl�@�ړb��4��\z� x�<1�GG�K�%`R�Q�dZs��B��dZ����P��	�M�.��hO�>5�孕�@9�"�9cd��B� D�`��Z�A�Ԅ��KBD(K�I D�(ʥ*>\1�SB�14�T�D`?D����'5)h�+=#:�+DL!D�,iF�;@��3��Q�d��v�)D�l�Q�p�� ��n�=X0T�Y�2D��g�)J~��!�A(\:�X�"�<�����,���:�=0��9���z
B�I�6h���� =+��ǈ�	��C�ik=�H��aǆ'ˀ@�W>)`�C�I�^�!1-�I�Hqhq*Wf�C��{�ԭ $gR�
�*Y�P���C�I=όݸ�DӖkq�!Hc%O�lzC�I�+��bG^6�	��+�%�VC�	.��Q�㧅'bN\�m�X� C��'>d��ZE�W�20�Ş7SA�B�	(Z��u�[�U��d�"��9B�	�X��T7�
xH|���@Z�|�C�I�g�8�A��C�R�K�d�D��B��#>�x�s�� ~-��;��.C�B�)� �Rb�ǆ8�գ�KB��paQ�"O�%8t�:.��1d*� EK���%"On�����PR��Z5\AT�P"Of�HH�rx�0YD�CO���	S"O��d�=�٤EZ#�1�"Od�x��� #�N�j3�ڮ%8��q"OhDz�m�)��m2��?43���"O>�BaI�0W�����#��ku�Q�C"O�\ȵʓ�#���"N"	�4Q�"Ob,Ġ�#�`Ԫu��dú@�"Ob��q#�O�a�0�Z�e�����"O����S&\	R]���T�3
(h��"O�]ڃC�����@�-���"O؝"��
%(�X&��0�BL*�"O�QS++���Z���:�ܣb"O:��U��k�P��$FB&j���"OQ�0I�NN�UP�M�'�Ezv"O��Ч�$|�`A�Gϛ�ꪗ4�yr�IBd�hP0E*%�LMkYb���ȓcf�L3��!#x]��#�E��1�ȓ���W��G�=jD	�;�D���'�\�
ώ*��)[�W�	喍��'�>��	 (*X"�FI#|��%�':�81��B�Z����ӋX�Cs*���'�04ش�AJ���fީ�M��'� ���@�J���M|\���'vpD����Rچȑ���s�\T��'<�1�eD[�ބj�lŋnYt5C�'��$Z nC v���"5��;R`\ɍ�1��Oh�5�q$��)���D��D�\���jX�e;4�4N\ �
f��-5��ȓG�B��Aώ��*F���4��ȓy�^}��g�uw:�:�n�V�\�ȓ'P�T$l�la��)�S:Uz��HN�
��(JwKɎY����H�|�<��ԏ}��YaB��+܎������(���'�&�2A8�1{���k�GE%qx�=�ȓ��l�@��3����%☻%�Ն�3<B����ع`��	�E&]8�(%��)*�a� ��z$h͓a-S1]�$��=<>����Z:]#�p'LP.n����ȓ�-	A���N�hMˁ'��k����i��Y�#@<4�1���U�����ajy����E��IpW&V�8t�|�ȓ@�lp� #K������۠|y��l�t!d��:w �ؔjW1�J��ȓV�ҠH2� �h퀐х����ȇȓi�Q�#G��7T`���'O��P��#��XR7���-A,�PУ�	vR|�ȓ,4��E.V3~�h���d�m�ȓ.�)��H<Aen�A ��+��u��z�:A �� d�i!se��XJH�ȓ�$B/�1�2�k�$tt�ȓ��9u�ޔ6���Є&�m�A�ȓz����h�lp`�㛧ns�h���D�P��t��gD!ws����k�l-x�n��[�la1�͔C�ȓOϦY�g#ʏF�����h��Ї�3��J��A�w��4!���;U��C�I�oV�����UC�H��u�=��C䉯n8���SAs,�5@�:[�C�	�|������U�q� <��b�7s"�B�	�?4����P�U
����߹A�B�I7"b�),�W�&�cV��5`��C�)� *e1W�.p<5( ����b"OB��@M�B��!���	>Y�H�a"O���őD���3&�xaf"O i�Y� �����{��,��M]'�y��/��0�a�5� ����I(�yR�_�9�xI
@� ��+�d]-�y�D�N�����4-��������y�M?&�,���W�Π�D��	�y��Hc�����
KY2�#���y2/�X�
��K3 t9����y�O�?VM	e�Ƅ'���"P�Ў�y���"~���R*k²<;r�ˍ�y2 T-9Z��
�w������R��y�`�/b_欸c�L�\�x<Q�,�'�y�̕�2��QmՌUmB�8���y"cT1<�@c��Rݶ��g�Q"�y� ��w`$b�� =�隗&��y�˔=pU��p�e$�8�	 _�y2��(Ô�� �GYL)�K�y�fΠO:)�we>:�(t#���y�JS�y�����%:Dv��TkI��y�!��p������+�F�#t�Ƨ�y´�Y�`)�=zur��Y2a�����'-�ð�]J����@30��@��(�p��A
W�o�8
�-�q�2Ԇȓ
��;����x!C�,8�y��?lv=��LT�By0��*>�e��2�(�x��M `�@����&Jt���eߺ8�Єӱ^*��7(ݠ�6h�ȓtҤ��AC�^���f٤L1Z���a$![Ɗ�*�	Ǭ�O�H�ȓAnDУŭ�(\�Y�W��`l��K�x}zeE	�bV��1K΀:�H����l������LԻvp���^����v�$�R�kO��ꑇ�_J�	��1-%F���̚�!����ȓ6�`�Z�B�/�N(JaׅB$�ȓ^��9{#�Hk�����\�Cc2���I�<(T䗤R�RBn�$u�0�ȓ�hYH��3?�z�n�!`�,H��q! ���)H��(i�
���d��`>��х�]��Mz��]�Z�����4�1�S��:S��&��v�V�ȓ3]�.o&��"��r�.��ȓ`m�d�Po	�{X@a#@����v�T�*����K�"��j�-Td��ȓ8��͂W�Y=���ׇZ'
��ȓ!bD�@�-o�Yk�$F s$�ȓ���
�cJC�ݒ#e I����:�x;�	C5w�����k]�d��ȓu��}{s�>*�4�r�[���8�ȓA��!�U��w���q���BT��/u�	;⭅�=�ѠVh��@�����{���F�S�&��� [�f��3�2D��� KL�>z�XZ.E�Hp�0D���1�1^�-p� �??��Ɋ
-D�P� �G3 ��7��{�a�E'D�X� cAl���P��F$T>�q�0/'D�PR�R�C�@���AP9z��`��'D��; ���v�,`sN�3_�h��b&D�X�c��n�D`RCo���.��p�'D�������T�ڡI��m9��Kq�'D���!9#��!�lѦ*����'D��Nŏs7�m`P˔�dQ�p�w�!D�� ��Z�##�D sR�d���b"O���bD�FU��sI�h��-�$"O�hV%��e��\Q�f�4e��8Q&"O�� i��B��b�ʫ92�P�"OXI�3��'k�f�#��A<;)DI��"O�9�Ȇ�>���&���w�XC�"O����
J	S���,X�"O�iS�)�7� �C���X�d��"O��Pq
���L �,��M�ڭ�F"OP�4$`z�Y�E�g�V��v"O��8�.�x��u���Ʌ$�(y�u"O�����T���"�2���"O00Zd��
7�����Cx�|l�"O��k�� `��&Ĉ	Y��(j#"O�i�1�Ӓ~3Bd��!T/Oz8Y�e"Ox���*	+#� �	PA˂%kvY��"O�Aۑ�	p��Up��CPL�!�"O�y����f��@&$�4[ĠӤ"O��"�ׇ
o�u��0"��u"O�L�Aܤ*��Ն�.y6�I�W"O�M2`ܠa�`��%��(8)2�"O��*�ɑ��� �¤M+"ܐ�"O��P��֜ϸH����n�|pKV"Op�B���_��0�¡G����q"Oz�(�*�=q�>�	a��3W��2�"O.LIŜ?ik�����<Iؕ)W"Oy�r�=�b �0엑}5��(�"OX�	��"�P����˥G.*�I"O��"���ԡ�I�s>�Թ�"O�<5�ٞm�6��7��<1�����"O�t�ckR
�i��GD�.�ht!�"OB@� �N�)�
fC��rT3�"O�Q�D� 0E[��:��ݣ�H�"OR��EI\#��H�c��WC�5��"O:�Ӵ,�����wD�B�C "Ot!(B��5� @G&I�Z�90"O ���P-/Č ��E���%0�"O�бp�پL�r���FF?�b5��"O�A�fG�	y�U�&��q�-yu"Oz�В��Q�v�q��
�n�8�"ODI�Q	��s�h����v�lˡ"O0m1efăA[\�Tg�c�-�r"O�	�c c���F&�s�`�{`"Of��&�%
Zd��a#�#7�A"O���X�~JE�⡎4����"O�4��m�<~�@yu!���؈X�"OP��7��5EMdlk��Ca��1C"Oz@K��ď4�MK�ʈCF�h��"O����I�y=|��a#�&C�H��"O`� �\��=X��A��"�Y0"O���^�<a�&�:ch��2g"O�(UC�t��Y!��\-̵��"O2d�䝾=�Ri"��;'~�u!"O����N�T ხ��\_(={ "O&�� c	��Y2e�D5�:�"O$PSe\�i:�3w@[=*��"O�=Ȥ�@9R���}�aK�"O�mp��tx¸ -5V��0"O�T(W��,	ܕ�!�ן`� uq"O��A� �_�v|���
M��%0"O8��v��m�@\k�����=�u"O�0�0 ׆�Pa���{q"OYj�I�%�Pu�tn�^�h �"O"|�c�M�M�Nxr�����"O� Ι��mT�8Aƌ�d"G�(�� a"O8(83h�"xp�+��\�U��!;""O���*��hRH�e畉\Q�@"O*�sR �?Qy�Y�c,��Uq�Dʰ"O�,	1D2e�Qp���!fU�x*�"O*x�w ��hq �_�kVP�	e"O��P�%H)o��y3����[O�� �"O��Q卝L�0򭓖n?r�@5"O}�!�_2�$�f���$"Oh�E�< 	&��D�#ߠ��"O���	'���j3固�P��f"O2<�� �yg��pC8h�D}�Q"O\Q3�'=I"�9T�	�?����"O�]��7�����DSxn�<h�"Oة���*# �m3�֪`��"OP1��BԖx���H�gR~A8�"OH4��Ճq^r�y��=�R�	�"OX�JU7J�,���	J��yx�"O���T��5� �*�̠F�*�2"OF���ЄY9�a��&��=�$e:$"O�p�`ʍ�MD�Ă�e�H X�"O
m#�D�?AS�'vK���R"Ob	�UA��gR�X�̃�i:�k"Oz�RU�?$����6k�3���"O�@����
��� wl�&-�E �"O��C�eJ0*p�ʑ*��#�"O�e�Ef�L���<Q�h`�"O�]�p��YHn�h�'^;$��B�"O�\@�,�� ���OZ>�Y�"Ovq�w�N�^�T��;�T���"O���mE�]�XA���� �����"O�!�E��J@Sr�M9N�4 9B"O�)�&����r���7� u"ORA�C�	�Z�l��G 8��ܓV"O���.�1?fػ�ß����J�"O~M���(�`}+��������"O�| 5��er��N�A#�k�"O4��#i�)����ІȗVe�U{r�IW�p�B�2Z(�9� ���XN!�d�315�u��R�`@(9�A�n!�]̄����_�_1��;gÄnY!�dC!�&�b��7].�tQgB[�^v!�d'3�\�� f^#3+ ���HA!�J�p��T�C\z�&�Z�Q B!��G���s�.S�������W�!�Ĕo� q��+H5���� �g!�[�^r"��цL&���"� _!�D�Y�j���X�Z�0ٸԬҐq!�$g!0�e�!
�4|b���v6!�M 4�T1s�Ϟ|̌�ñe�U�!�$F �0��/��UjQ� d�"�!��;;ĸ�t��2 �us$Ĳp�!�T�+7$X"Ea�#R��0�1I�"�!�D� �8�¨Mt��(	�!�,E�8�ȒL
�9�U�Րo�!���`�#��v`
� '��u�!��ɠ
�R��6e�0��@�!�DN7q���CB��e��)�b��<w~!��&�ta��Ҧ2���Iu�
�t!�[�MpP��_�B����W�F!U!�'	~�z�*=C� �b0�F(!��`� �r��sA	h�!�$Ǒ/�I �@�6��Ÿ�I�\E!��:Bwf��,P�rvĬ��E=@.!�� `I�P�	�\\Q'F� ���"O�E�!�u���{�� \m�T)�"On���@;Q�lCUCJ>8pb�"OP��ܷ(��!�A`���x��ȓ[�H��_�#�� E'�1g��-�ȓj[ht�`]��̼C�P1Y�D��ȓ��*q �
z����(>�l�ȓ\mʸ�W�F�V�����un����*�ZD3��%h�Hy���h�hL�� ���"2�آL~�=�@��3��8��S��`@UJ� ��*��ܒ� ��`T��FA�d��<�w��}�l-��!G:�@�^�7�����Q�@$�ȓt�pC�H�BZ�P�`����b�<$M��.���c��Ofj�P$MOU�<1C@�F�@0��h�酆�M�<!�@�7q̙!!��SJ��#u�<B�FN���`��|�"�K�c�o�<��ʘy>$�� E֚1�=�S��P�<�v*κ}ߤA�#�^�D�sgXG�<�ŧջp�����a,nO��c�C�A�<���,��!B��#M�&M����D�<�T�,�,�%�X*à�q,�~�<�G%�9�VD�#l�!hspdp��[|�<�v��i���3��\�k5�0���w�<q��ӑ%n���{q�����i�<Q���&ݦ�X�dC�v�ri+�eo�<I�f��7oHI��%�m�PXS��An�<Q�ȑv�d�2��"|V�u��
�O�<A�F[D��0�nK�Fe��]�9����RJV�G�|�!`�݆�=J!�$׶(6W�6*|������~�=��}�I���9Y���6��2s.��ȓ)z���oҗ?0�P�/<?¹�ȓh�h\��
�}X@�����ȓuW(��(��l��lV��k[X��?)�Q��f
�C;�]�$�Q�cfvl��Az��� kִ���IӍx.���ȓE��!�i����P���F�l���ȓ:a$b���%��F-����upq(3���d4*s'N��@��&j*��B��K ��1��*�0��j�.�*�/�:vA�@��J�x��Մ�3m�� ��J�)�`�Y<��E�	~<�#�M"Ĵ)bF�ř>樁���a�<2�	�(?��&�C�� ��0�Ng�<ђ�ӻ=t0�!N�J��W*`�<)��" ��W��%Ռ�� �e�<A��3?�Ll����h�Кu*�I�<QslD��.EH�0�R��T�|�<9��(�
}� �o!��p��	x�<�K�K��8١�@�-2A�%�u�<q�ͅ*l�����,f�����L�<YҦ��r�:�#��6����j�P�<�T��"ml���H�0B��Tn^L�<QV� ��$�M21apԂg��]�<�Q���L�:ClZ-}�7��\���0=Y��WШ���	�Y�i�5ʔU�<���ȮI��jF�I�V�,�6��Q�<��횽%�A�BF�p�ș���i�<���ډCʸ�0�^���-D��e�<q�)�a�H�A��wp���g�G�<�rn�#��%��ɹ-5�`�c*\�<a��F�9F�%qg�U��Td�W��V���?�
�S�? ��%L��2�}��U;YyІ"O �5�,`ҤeaĆ��JH�y1�"OFM��+�,ڄ�hD埕1�0(��"O���¯�b�r��d��;w��|��"O����Y	*��@�����<�W"O̬h���9u�`tX����t���"Ol���Lá3�)�A�2yz��iP"O�87��	t�t3T��.Q@Š�"Oz," B��=+�`��ز��"O���Q�O>�He�\(pĄy`"O��4��J|���
T\�x9�"O^%Ʌ$A�3�
��"
��G �=�B"O~4x�oR�>�� �&�[,�f9�0"O�����XAP	����0��"O���4eI�w��Б�e�0�K�"O���J�]��4�v������w"OT2s
��E8*,�殈�#|�|ء"O�4����s�襰Vc'd�i�"OL	{�!FP���R��)��c�*Oƥ�c�&p�<ӕ�:t��W�<MS7xt0Q��+v�R�Яey��)ʧ%�� ��\D<RLk�8Ҧ��p���2IOZ�F%��$��md���ȓ0l��8�\��	�v�з����]������{w�G$ô����k��
������D��@^�%�d��ȓm	����[Ѥ���O b��0�ȓzLP!SPm�66�aCAS�6m`��[�u�"o��g��5�e �m���^h���TO�lq�'��H�ޡ��::x�B�C/i�T�HS��J��ȓd��D���7^}��fJ�D.t��KD.a��÷Zn���(�01�9�ȓLNX=3��[TZ�#B�(L����	�Δ�ר�?P�yZ�/G�I�%�ȓDf$��̜�)@z�`r��5cW���[fT�ga�I=ތ��*�Q}��ȓ"Ո0r�r!B�(��*m����Q�<��G^9��D8 I�&9��h����1ᐪ�
��\JcB� 5�@���6���!��q�a+`�OvbdE�ȓd�\�D+ϱX@���V v�ͅ�Od�`�hU�lp]��H�;����ȓWn���AI�
&A���N�Z`F���J�P���SU< ehqm^�>��܄�2&\Y�CB+C�T�����(�&��ȓ+]`v%�#$��#T�A2��e��x^e�nށ�h9S!�
#[B��	t�t�ϟN ��H�$HAE{��O�<�S�� �8jkC�4�q
�'@�����۷z�-�S�� �"�(
�'��p��
j��	��ӵ��@�'�� 3�D�n�|kBŝ"/�j�h�'	L`)s�gZP� b'\�Ld�
�'���Y��G�t�8`J�lI�i�(�	�'��Zf��\yP����ůn�p,��'N�{�>�,-�u�,�̵��'v�˓�3X"�L�e�Y;��M�'�^��CC/d���ѣ+� *tB�+�'�� 2��Ԣq`)
@Ύ�N����'�8D���d���۩M��T�	�'aY�E {x�����7�:���'nfI��*����X��]x48A�2�)��<q��u�Wȉ!��|��K��y
� �t*Ќ�y�Х;��9e�|�c�"O(�ԍB/"����"�)�'��'J�)�n�0y�#T�R�D�� V
KZiP
�'s,=	��υ�f$y�b�K��as	�'rН��!ڻx~��`K��r��<P	�'�}��痥=�:�cR"��}�&E
�'�Х`���<l� 2�A%}<�i	�'�>IJ��H��#v�B.=5nЁ�'I�-q���<� �p��h=�y(���)���&MK҉�`j�*x��L�y�`��3(�ȟ�p	��r��)�y2oT��DE!�(_Ic`'���y��`���ï�8>#�DSAl߶�y�e�iZ�)��oF 3Y8��0��yb��&�zر�B!)?��pM��y"@)A��C :	�N��w���yb�
�E�&��|������ym�+����f_�|��تC�8�yB�ƣY"��`�ـ{�JI���B2�yrKOj ac�ń*�b���L��<	��d� i�F�3���{=dyq�* j�!��3<�^aP5琙Q<L��h��D�!�A�ސ:��F<H���Q�S�B�!�N�_�z����X	�y�sJ�:r.!�$.e�fu�!��ॳ0	�?K!�D��h�Li�@B�N�h�'H�K�!��`��Ñ>�����9H!��֯p{�M�TbH9.�[�מ*[!�DZ�h���9Ê_�*�E���T=!�d	�����eۂ�UA��X !��]��i��^�le��@�L�"�'jB�'�$!��� (���8�ʍ$3):��'�z���>B����Ə�;��"�'���(��c�ʔ�6l�u�FT��'���A�BB���I��k��x�'8VY����"eV�r�Q�b�t0�'�Z� �L�:hze�$C�>[�'��UiB��f	�!��H��o�D!����xr+Z�M����oYD�$���!�?�y��>i�T�p��B5�:�Ý��yr��0q��R��� ����e��=�hO���I��GUѡ�K�;m�� ��
?�!�$�Lp�)5�\S�p�{�(+Z�!�dǓi�@]��G�!r�Bb�H�!����p/��Z���7*j��I��
n��'���'@ldP�*�)[Ɇ9r H��w()�
�'���a�/���A�`À}b�@�
�'��֍+<�ptc7C�5xa���	�'#ly���:Bͪx3��P�v{��!�'T�/����h�/n�n�Ɇ�S%�y��T�F���4�
���M���>��O�l� �B�j�X)� cܤ �� c�"O���B��7n����;H���F"O��Y��_�4�k���k��(�D"Oh�J�MO*l�d8���FZ<�#�"OʸYR(�p�8UA�&�ԩ.!�D�Fl��eEF�c�l��'�
��!�-pdiK�È�n�#3���!��<j:���˃?L�ʖ��)-!�G',�Q-��:80)xu�RL{!�$� 7��c�D�
�ı#�&B�h!��iN��`S;R���R�Æ�1�!��Z�\X���n�Qh�@اX4!򤋊�IW�,�\�� ��$kE!�� �葱΃�^�α����>Q��@H�"O�4��b[-1w��+E�Š
��yP"O*Ī�hS4��!�P�0qHh�"O�|� M�T��x:rm�m@�'"Or����ѶL�R��k�DN� �O�!�E#�1.��if���X�`<I�-D�:��#"�p� ł: (U/*D�؊T��=���ɳ�;6"�@��'D�(9�B1PD���M�7G����a+D��3�Q)8{�+�62ּ�R��'D�p)��F'��j��b��l���8D��!ǩ��	L�����3^��bc�,D�HS�/�x�8Ն��_�숥�)D�̢��N���m\F~�AC�"D��:�D���$k�m�-FbX���M-D�P�冢{'�}�g�pc*�)���O0B��.F�D�c6m�5o:m�a;e4B�I�4�h�����R�@ab%DM4R��B�I/	��4�!W+?ZAF��QzB�<*�r�Ҡ��n
6��f���C�I�gXf��#��'<�*��gN�5[,B�ɐ�0aГ���KQ�؇��W��C�I�dN��{�Ę����%e^B�I�u����'R��h",v-B�	�u�0��oO���$9�Ε�.#C�ɔ;;�����5&j>%��NkDC�I'�����?a	���b��B]~��0?��M�\Ni�"N	B���E�LM�<��+
(�(P�WƓ�xd� HN@�<ye_�'�-&P;A6�)�l�W�<�2/Z(a�܀-�"Y����	S�<�r�U/�}iƢ!WgP���#�L�<��� *f�����j2d�f�@]�<��?à�� �ZSN �s�[�<��jB�Y�vK���������Y�<�RdQ6>�T�I��T�v$[�<�0��?7�(��E&�� ���2�A�r�<����+gk�����u�`Z�[i�<��|r��C��3ZF�H���	K�<�vE X R��c�E�kQ���Q@�C����<��HB{�ؑ��O�=��UZ�Ĉd�<� �4n�}:CI�9fdIWn�\�<��+�v��r@5F[����^m�<�TL��8��<�2i5y���z��h�<�קR1#MH9�gF�I�-Z�B�\�<yw�ҁ3l ��˲^��e2�C@�<1f�QT���e��~w2�)ġB�<a�,p�j�Y�F��e��mA1L�C�'ax"�̽N[�q��X
�����ܱ�y�-[�,���Q(\��� %� �yB,ӭ|vԙ�sc-u�$�B����'�'td�R��?F�,m1�b�7~�4 z�'�ha@��%e���C�ւf�>�J�'\(B��'q��ꥄY�\)̅3�'[<��D�+���ɤQ�h.� َ�d1O����)jX��06h� i��:*O�Q���n�����W������?����II�v!�a-
�àa��ތbmT��5�L�H\���P�'MڧQV���6D��{c%�e���W�x�D���e2D���$�S�w¦L�GkU�rb�T�-D��Õ�3]��=���r��pyR,�O��c���ycS�2~��
}�̈́�ug0�(P�ҙ�,�����>�"���S�? V�+E�[��X��񉚞N�ܸ	���Q����Aҝ%�^T�w�.�lDV�'D�������A�g�%�08@'D��!&��
Tr�B�Y)H�l8�,$D�H  gG�C�a���}X���� D�ܳ��ƢU������&Ah�A0��2D�,��S�I�<�Aҥ՞QL&�H��2D�0�%f�#py�ȩ��V�w&�IQ�1D��:w�E7^�<�uÓYS)/D��[4G��J�R�WC�=3>X�k D�����H%�H��4�f`L[�>D�4�(�:Fu!ڂ�D*(*X�d=D�`���^>P���h�6H�F�i�<D� ���HwZk�A�6i�lu�.9D�,
V��P��P��C�W�^�s�3D�D�v�R4��舠�XKJ!q҅/D����R�s6���@![�P1�-D���tL�3~��*M6�BxR4�)��0|�`�&y��XcCa��~E��L�O�	[���@�6{'���#�H�j>A��9D��۔"����g�o��6D���p[�xa���wi��a�y��!D��y�j/�`��1%	%����"!D�h�����3�j��"B��&X���I,D�$Y�'�E|8�f%b� �s�h/D����#q&N�r�.Z5�#�+��;�Ol�$B�E��\����3e��kS"O�-C�g��Ke�=k���,���"O�0�ͥ7��,h �Z��8@"O��RbC��t���ōLR� L�"Od$�W#6{�>��&�<-�*5
G"O���G�X,UEAC�eR��d"OdH�C�d�&�� M8���"O�pT�L#~-���c#�GFJ1"Ot�����T�v�!�,+� �T"O.]1B���)Q�(��=O��љ��7LO:��vM�8�1�^O��@0�"O*<��E^��n aы�2{m�"OJd��%ѷt��
���� sE�7"Or�[��� n����J׎am�\:g"OD�Z���	mQ���QV��R "OD�pm�9x v���F��IӃ"O���A�7�
)��*M�H
��a��f�(�CH*'�u�C$τ<t�ᄃ6D��Q�����3��Fߴ4`�'D�z֢ʑ�� ��W6s4����+D�$*Шǅ7x~`@�cQ%aK�E���(D��P�H�S�y{�"<V��(D�ly��.��F���b] �$:D���Q�^��2)zO0E� �	�#D��Ձ�U�:���c:	��" �+D�+V�լȥ*�$^��[�'[l_!�[)�*��[J�[t��q�!�<=�ĸ�a�R�h�0�+!��?()P�mC����럖p�!�G<�`��iR�vHɉ�)��!�=z���h�aZ��S(ȸ
!�$�N��1p��?f	V�1�FA�D�!�$��_Ь��D��a�Ld�W�T:y�!�'vI�mkRaF�1���XP���B_��$ϻ\p�V�9C����(�B�I�/%��`BZ�3�jPca�]<d��B�I7R���0�ʱn@�3!J�M��C䉮+B�0ZQ
կf�"d��-�JC�)� �)���E�0L(p�U�4!���F"O�eK�!��X���$bH�~]�`"O�H�E B�D�г��Ji�p3"Or�22CS8�H�g\�uL���T�IV�O�̺5��.-���c��#(��	�'喕Q0�N䠲��~㞄*	�'dbt��
#-P0��aF��(���'O+E%I#/�>}�qcP��5��'�
(�f�Y/(N �ybĂ���	�'W�Q����aGP([%� X��'��,�M"�ժ��\:EN7��􈟺�y�ѼP� �%�
1��r�"O�<ᒠ��ben4@3�F�M���2�"O����V�yV�q�3K
1�&����Iz�i��H7X˰��2N� 7���A��<D�,�"B:�l{wGՁ:ut��g-D����z@��#�Ul�C0�*D�Z��%VY����"ξxZ� =D� j����C��E1��=jġ8r�7D���2N�%~�>��S-\���3D��b��Nts����I({w���0D�Шƌ���� �F�&!rD�&;D�x����6�h�Ǥ�=-jл�
5D���v�7bs���H�<��2�M3D��(W��|���0�φg���2ь�O�=E�E���B-XP P�Qɶɫ�@Z !��0 #'	1*�.�z!�ϫ�!��n&�	���_�tp")���!���!Y�D��C�r�� �c(��e�!�d��g��@[anK���y����6�!�ۯ0U�������j9+�ŒW�!��C��|ȡbP�}��ѧ�ߝJeRO�pr��!)9���� _���"Ot�i�Fĉe���d��<�:8��"O�4���S�u�6�P���"O Q�R��P�lc&�`~��Z2"O��2F܂$e�lC`GWbP�Z�"OaHo�0�hݩ¤B�-�.q��"O��s�G���$;1a�<�,ب�"Ob��$���X���Q�ZO&���"O�,��H}���2�oS�LX���"O�P��UZ ����:�����|��'�B\@&&��0��%I���k����'��䀶�Ҥ&x�0C�-;Z����'R��D�2%r��p���@?��`�'�Е0f  .�U��U�3K-a��x2(�5<:�`�
l���ْ�C��y����6آ����M�Z��R������<���~JfL�z�DX��qIA���	J��C䉰:�b�As��8�X���dG�ClB䉁7��{�	��I`!:c�O�+$�B�ɯ'�Qj���7�t�G�K�B䉖�2%s���|�+�?��B��;�>�'��e�PL�fjE�5Ȝ��7��'ړ��d�f00@�eGV -����a�'Xўh�<�����[Wp�+��L�*��A05NY�I@�0*n�;p��"%��Iw��%�6D�D���n���$�%t�	pc2D�����6 hQ�D�� 6��@�3D��S�1�U�����Ӏ&'D� 0UG�����@@%U���#!1D���c!V�"�P�j ��[[��R;D�@c�a
l�j=�g�Yw\�a&D�(��h�p&�%)�A��=H��O#D�� Tɳa"��b,Dqy��1h��:�"O�h���3�$\E��.s�9W"O24�1�	�O
���TK};l<͹w�d-LO�ð%��-ƌ��I{4���S"O#�o���� 6/�7:B����"O����%��z�Dŋ��_I2��P�"O�hզ�N��,H_�Y��"O<%�Rڬ���%�ػP)��"O�%��GC]&պ�]�4��E"O嚃͍�������X�~5�"O�{��Y�:xI�'��}["O�tb ��^�r��cz�E"O|,��g*b<����	`�]
&"O�񃀐9Hޮ�2v�H�A[fQ�!"Ob�����n#f�X1nZ�5>8eZs"Oҹ���8yI�yP���֌Y�"O�i1��66H<�Ԏ�$��py"O�% �� �H�R�e@hR3�'�,X �ŵk�.Pj�唘E��8h��6ړ�0|zS(�%3�PW��1U�H�Pr&]c�<�qȔ
dۚ@�DA{z5[�ƈ`�<�ԣ�*)YNl�A
�qfq�q`Y�<yE�;)&�;�/��q{�b"+TTx�l�'�p�H$Ƒ�d⒣�>$'*�q��)OP�4狣;0N�Br�<`׌��S"Ozl��cM%	�~(yt���a�Hu{��'w!�ę$�mxfb��bP��jGR#!�d]�Qdz���F�h��Q���d!�䝎r/�XSuר��  ë z_!��� IM�9�A�]4��1���9K�!�ǴlB�C��t��`a��;��'�ў�>�yaֳnr�"A��y:~�*��1D�`�G�=v�g�@Y��H��K1�	J��4��n����%����F*( �d�<D�dI�)/��qiߜ#�и���8D�0�� ",�I�.� q�<X�G8D��ش�yD
����0N��JA�!D���M<-���ã�+/��j�C$D�4�w�=@�9�o�4�XC��=D�hm�*?�bd�g�Z6s�r�2��;D�l�EBX���pT��P��:D��Ɂ���wf��5�Ў}��D�'&D�$Cq��`��,!g��;%�^TSB�&D�P����<:����E$(�V�
[�!�dS=� �	�o��E�N��7�ũVv!��Yjl��V���ܔ	$��0^!�d�Y��%�{|�<P��9 �!�$	6V�21q��Fs@$Sg�6^�!�ą�A@�D
я[�l����p�Z�!򄖥q " ��Dc#^DV��-5�!��I�H��Ś`9�I�F�֊u}!򤒋���X��F�D~t�s7I�'^!��ܫk0���Ĩ7NjI��甲XG!�Ea�����
J-	��B�A�^�{r�B�XB$�꒨�����E&�1�!�,Aā����de�$�e���!�ּG7���N�* R\�c�d i !�dF�<\�  
�
c������Tx�!��Va,��h�h2]��]�3�!��Q4�q��#���Q��;��yrቤ'@3Ҥ�8T��N%����1ړ߈�����/�=���GB�Md�%��Z�І�I�E��=�d�:0�ڷfI(00C�Ƀ;�	���=;q����fLgj�C�)� ��wo
߂�"��fH� S"O�y�%E���]c�cZw�xȉ�"O��Ko�J��F��J�ܕ{��'����qr lA�Dȏwm�ՑbcS�PsB�	��ȉ5	ʲX�k6���c�C��!xq��M=ei�(�wN�0+�RC�Ʌ_6L1����I�䂴�GN�B�	1���Pϕ�9P�Iy"�%s!򤋎|�.a�(ɶ`3�����Z�j!�؎W�بb��݈`��z���"��	_x���'O.�W��\H��D�[�n$��'�!8��n�) F,�Z�fUz�'����ьK�ZD:����Ov�e)�'\��
�֜�64��H�>��T
�'m:��Wi ��P��Kա7�^�y�'^J�7͐/��4ZŖ���X�'�-Z��U:^�"i+4�G�xR0Z��D*�XY�WGޯ��hx�G��z��+�"O���&�/��2'��Y�.�9�"O>�����n���5�����["O����A��9��]Cp�˓z���A"O���g,��{��p̂�h��"O���aF�	Exqx�íZ� ��"OB��3��3�x��L�8�
\��'Bў�'���O��Gk��("Pnԇ%p�X<D��p�E+m���EыQYX�Y�¬<��h5�m��=E���rK�ML8���s���h���D�d`
�V%�̈́�P[r�JGe��r"�y���\N���TZ6���ʕ\�x�A�<\� ��q�t�)AJؽ�F��B�e�=���ڭ�v�фc~Q�nXjUP��p�\L@�a�D�v
C<Ajr��Iן��	�P����,&�C�*�8=��C�ɰ}�,Y(�(���9yt�ڙ}�LB�I)�D�pԅ�2p��Ka/*Z:B�KY��z���9�Bl{e�L�n@B�ɴu�H���TT� �"��*ʓ�hOQ>9���C�}��s��X�#��mP@:D�,�G'�b��bEJ�`�!3�=D�� �K�*&��3�8��1"=D��Ǖ77:�Tz��7+*�����<D��[#��?P�x���뚸	:IH�<D��!s �fk|��AZ%98D/9D�T'+�:�Q���?���3զ!D�t����"�8t��	�|��,K�*>D��Q�F_:z%����a
yC��<D������A!ܱK5�:n��1%j D�\���,3��(�A�{�ʴ��A>D��
#�ݖ� 9P"cL�l�(;v�'D����_�o���!���>��� �%D���"E��^1P�#�>��+a�#D��;u�	,���j�
D�ߖtd�!D��`���&�����$�N��,!D����ʛ
˲��� 8x�2a1D?D�,ѢݙG�@���\3P�h��&�=D��"�C�P�@2Ě	f�hyE&D��!��@�/�&43���B~���0D�`���#(�J-���U�^<��g+D����Θ�C�(afkY�1f���v(D���L�g"�� �	~6H�I�a"D��c�!�u/t�p�ݫ/{||sd"?D�� 6�Z�@ʠ�)a�Me��#V%<D���@�d��`�V�Zn�LZA�8D�� ��%�	4�$�*�'
A�*�"OT��`N�<T��h�X1 �QW"Od��]�XE±��g7_�T��"O*��c�uP��[�fިu��Q��"O��g,�]����D��|��P�"OPa��lZ�$�@��é��<���`�"Oj����@$�^��O=x'�u"O�Ԁ��C�~�.�%F/l
��p"O�����%�J8 ƃ�t	�(v"O���d��$ g�4_�����"Od�3��-Uh52�J.�"�xg"OD@�Q.�4%z��땯р�V(9v"O4�4�)��#�V��@�j�"O$QPr�0K'NHH=��5�"O�4/�Z.H�Z$旭V�b0"O��؃b�t�2}��%��Y��D�V"O����N\ʪ4�2d@�s���(e"O�Pq�R���rc�C<WѤ� "O�s�G�|q,�hASh�4��'"OqjQ��M�p7�ʺ7�Pa˄�4D����ƞ�lA\�y1�T9lQs�-D� C�E�$M����`�1;aش�,D�\�����t4B��S�e��C7D�s#�Q�)��a�pG�(��	���8D�<���GeԔ��$�p��1�g�8D�G�ӹ܊���� q�*$D��)��QO�Ҍ+@�����f("D��w㇛FA<Y[�bA�?���f"D� (q�Bh�PКBܙZ������ D�\{�H57Heq��?>Ҁ�u#=D�P:�$R"N�Ƞ ��)��9��:D�t �b��v*�%�׸6���QS�9D��`0JQu@E��K@�M+� �FG6D�@�ā�:F� P!N�)Ԉ�zb'D����ťefT��Y#�X f#D���n�>���B�W�)�@��a"D��r��[�&哀L�r(,�à3D�4{%���X��KdfF21���(��&D�p�H#�^�X6�L�Qq�#D�l�d��c[By@�%��5$E)�)"D�(�5�BS�R�0�2��X-D��k��ٚ>~v��Aݱ3��XӨ'D��5Bڎ�^�K�M�n���r:D���C�y$���C.>ny�#D�t���@�(��X0�h��#D���LM�?#��B�k�4'ri�$�+D���N�-�^蚤�B���;Qe.D�t�3��m7��!�FP��Ԃ%�+D�X�V�	�Vi�̈́!/����EE+D���A	�.bv�̓ӎ'����K<D�T��LS2{eZ9�w��X��`��>D��2d�=��PSv�+@����A>D�p��n��\�U�V�7F����<D���2�zڬXP�U�FxܨE;D��r�	�mNey����P1rQC�9D�l���L}<t����M���y�7D�����٠���o��Uxy �4D��ғ��C���aW*��;} �Y��4D��y�k�J�Šd�Ǥ	!�r��1D�p�Ke��!A���%?a�+��+D�tӢ�.'k�5` ^�J���C��)D��i�B�LG	����Z�P�g�%D�ӑÖ	XሽC �Y�Pڴ@`/(D��`��N�+�9�a-�"n�yD�0D�� H��a\ w�,�فR +��Ye"O��ֆ�%2� ��#K�c��<
�"O�A�Ǯ���"}�Ynj�ٗ"O`%re��1rXx2ӭp+�p�"O�� u)W.T�iw/�I@��P"O�i�n�8~�lqe�I���� "Ov�)�^B�J1"07�
���"O�m������{F���̙�"O>	��e=D� ��`&�#��a	#"O`��FҷJ}��cB��T"O�	ӁN�:�|�3�q�:g"OJ��E	>1{p`�OF�Ma��Pv"Op���5� UiV�Z7���F"O��)We�H��H�]��P��"O@u�$M�!���*��>s;����"O��2VD�b�ɩ3��� *jAp�"O����>7��,�"�;|=��"O����,&ekDa3A� �ک��"O���%߿|�p�z�/į���4"O��{V�-b5�ġd�L�.�"h��"OVQ��k5o�튒B���l�8�"O� ��._�D����&g���"ONZ�A���	����զ�A"Oް�����ip0��%F�&(ܸ"O�����7wM���$\-K�"O���ǋKgf-R���=0
�[�"O�aYԈƵ=N H��
Ϟ�v"Oh�;!��
}��j�g�F�T]ا"ODՒ��9C��ȓ&N?����"Ob�i" ڗg�آ�G��H*��"O��@�A:���������7"O��@�CS>&�j1�F%;�3�"O�ٸ��
~T1��eͭNa�ٲ"O�Yb�A�?��إ���: �"O���#�Yɖ4�3J�o�����"O��Ӆ(]3�>Mrdi�R܈ar2"O������I�F�ˣ�4��"O���fU*@�2���g^<�F=�S"OZL���"��Pe�\`�~Y
�"O�u�NB�\��@!)N'c,1��"O<��QG��.�&9X!C�~�J`Z1"O $��#JH���r� �?�΀��"O���eC@: ��k-7'��(�'"O¹�������!��"=�PXg"OT����S�|��`�g눆c��͹�"O�hG�܅|=��<Z����"O6��K�
��H�,��<��C�"O�q����z��h�$�dc"OM�qH��45� c�B�Щ�u"O>8�SBH9*�BQ�5�$|�r"O$�׃؅w��}ca��F|U�"O&��N
-	��S��|�4s�"O�5x�év#�@0��(�a"O��I�$N�T �A�-%^ɲu"O~��d Y	11�hq��+/��(�"Of�"T�8���Z��/q�2]�"O,0ZQ�ԓdP��EΚ���`��"O਩b�.����է^ ��#�"O�I��$�1��Xs���C�"G"Ot�!L�4w�"��V#	)2����c"O��hr9n0F T��0g�:@�"Or�K5���r�
B�Ӳ~B`��"O�����t�1"�C�-9�tA�"Oġ��'@6A0��I �\ȹ�"O� H����G0'@B��E͔-Kv�*"OLlې�,���*0��s� H4"O*�R37(B6xqd��U��A��"O`M#��64�L��c�}�̉i�"Oli���	sش���B�1�r�j"O����Ù(�,���!�X@�"O}�5P�wZ �B�
@*XJ8�;�"O�H�6�J<6c0�V䉾T�d��"Ot �7fG�m��s��v��	�#"O�,��
:I�T�7�y�����"O y�`
��.�pY�dP�9ߨ`"O�����l�����K*���Q"O�Ӳ�F1k��:fg�ur����"O�ɸ���[���f��Z|�ܚ�"O<�� ʋ�v���2�?�"O�I�g�Ƭx�4
�$V�c�"O���()A�qZBd�<$WRP!"O�,"��͡�D��3�XUQ�R"O����D2(���)p�Ζ_�e�"O�i�tKC;!^��A��'���r"Ov��fi�%[�J�(�?Z�`)�"O�Y'�X�L�B#�9�,<��"OVŪ@M�9ѮU�Q�/M�����'���Y��SP�Lf�Z�)'�L�z�`E�2D� �˚�zTE#�e��j�� 1ړ�0|��b�'&��;���H�C@�c�<Iq�d4����6�c1jZ+w�C�I(�|��!���,��)�=ݞC�	�zL�٘���F$���s!��B�I)a�P���1����0:D�B�	`��t�"������9�FB�	�Y�3f'H��ڤX@ń� <b��F{��D���P
�P �CH=�8Y�ߋ�y"�B����Æ����z��A�Oh��D��a2^�i�B:vFd���a�!��U����V*�DA�9IkW�]�!�I����U��1�!@L�� �!��s��PY�̯|���p$j�%,!��n0��A�2s�H$#a�A1�!�� Ʀ
G�ʸ	��"�!��^�����IO�y}����d� u!�$��P����Ԗk^t�����rt!��ͯ9���ī��f��A#��#\!�$>�"i˅O[#�p0{�(W�X!�$ȧ����c\i:ĳ0&�KN!�d�\Dxj ,2-�^`��4H�!���=8����%�O�P��Q3$�/>�!򤖏#�����Y��]x�L7zv!�$^��("F���6|T)r�Ϋ]ܮ� �"OV�#�7xt4}h�ʣZ���"O�h�g�V�p�85hW�f�Z	��"O�q��ד;��a4��(VϬ�� "O�`i�e�6s���]{�(TYt"OP��犖��f�i�C$˔�:�(lOf���	�N�"b������"OtSl� :���h�^U����[����	Jsd�knR�)��U��oC���p?� ��;z����ܛx1rT�Ï�r���'�b<�OZ��� 
U�b���&(�Hs��>9K��j��iƨ?T�!h�D�,?�)r��Ç�!��
��m1���2$x����&�b�2�O�٠a�)^Z����Oؚ�U��4O΢=�'��O��)5��4qS	ֹ �*Y���>4���T'R4~j�ɒ��<��
k%?QN�Gx?� �xU?XN�S���s���"O��*�I�h� P��	q����"O�Ż�o�L�FIquÆ)��$!�"O�5#w���T1�DYD� d�xm�:O���� c��t��'�4�����Hܪz!�_��Y��:�v�+��o�!�
8P|�r�A^GH�٧���}��$:�I�T�?i�g/ �5^rP��$@>(h���R�7$��	��������k�5v<�����Dn����I-t�L]�-E����a��S}j��<Q�'ʛV�ԍY�2E���[��5'��9��C�	�$�9h����4�xƎ]�F�>1��I�6����k�,`i�̋!�D'�*���'ü:j	QǢ�]��y�I�	�����%t��Q�DW�$C�	l�A��TU��U�lӝ(��B��9��M0:���a �2��b�<�>a��$���/A�|�oB�SND4�TmY.I��D�>�6�{�KE+ZCD1!$oWGGqO6�I~�Ӻ��Op`�\�c�|�8���7e3 P0�"O��k�@�U�
er��N"�(�Q�I�HO^ʓVzV�Bƅ���\E��\�"����G���g��HV�!e Յ~�vAs�OF��t*��,(h��6��))"O�KD˒*$�$�2��U�u�	�"O�h�G��'hOԈp��� n,v"O>���Cզ2�� ?w �t�d"O��[��Nh�Y����,T�&IS3�'��ɧ
=�������zɈ�B�,x[�C�ɺ;3(ȋ��oPl!Q�@2��#=�$-1���0�P��1��0XK�E�z̆��D�'��i��̈́b�m�Ω&��P��!�S��?�Q�[�RIA�  ^��Y¢��g�$	���?E���5U�4�d- �u����N��(���c$�P�c?2:�]��#K0Hh.�4���+}��Ab�x�K��?��Q��Z��Px��-�ذ�&g���9�%	3�B$��f,�=S�E��iI���T�ȓi���c�^X��P#V��O@hx�ȓ34��vM�2^(I� 	N�]��e��mMV�u��$]��r�E׬F~���7�|�KQBB�]�d@��h����%�>������(B2sY%c%�̌t-������y� Sp��A����{o�$���'b�'߀�j�#]��d�)I�t��I�'����s������U�[���Ñ��hO?���7E�M��Nl"`p����<{6!�D����LIe�ߣ+D�B�&`�V&�K���kp�E�F1�m*p�y��d�����F{�Oc�OI��#6*�`�b0��.Sn�� "O�%ʲR�2���K����wT��F"Op�jW`P�H�p1Ε�c7�J"O|1��c�<���C�1%�������'�ay2�N�K���9a��p� �	ʨOzb�$�OuxX�v��wbH!�����HK�'� a(�"B-M�����J������'_a&��#����`� c/��ط��xR�'��#��!�f�EZJS�`R�'Y(�틥�������<�$���'���A7��I�ȉ��&�"91�̱
�'�~p��O8K�hY����8�d�Z��d,�T*^�[@$�W� ���n�&E��y�lP�UBҽ(Ӫ�c�%��vT�'�ў"}��+^�iJ"�S�
�FI8&N�r�<� z"�LҺ7V��BI��~�x�"O�h��@�_13��[9�Ē`"Ot������"5z�`J�8b�w"O�:c"/�½@ T/3����"O���Q�0�V(��ϕ�g�X�D"O� ů�#c�8�m�[�P$�G8O�=E�4��v����ƀM���C��y�o@.�-r�ҥ\��)�U��?�H���O���YZn�r��-S
��#l�6C/�M�ȓ;f�u�ƨ�2i�+��	�;B�X��^�["��W�.�R2��Lh�ȓE|���]'i	R@r����6�^؅ȓ]"H���gL��2�΂)�����?! ����	c�@
��O�7�^���p�ء��jo(� 	N!X�D���:L�A$ N�,��y��K�`�(�ȓ5:h+6�ܵz�0��ȕ�N�~��U�̝HA����+]~�� %�!D��� m�C��M�Gb�Pp$ؤ#+D�찰�3��� 莃e2pj"n#D���5eђd�496J˽�=�s@%D���&�9cX�[��ħE�h�T�$D�D���پt���c���W�e�n$D�x���T�q�4{"(�/;�
�/D�@"CE�2D�4qMA u��-D������.�p[��B/���S�a,D�z�o�K_԰���c����f(D�h��e;$ 8��Z�pw�'D�x(A$�;�TI����>��y`�8D�����
R!X�Q"�&^5�d.7D�|�U���ra"�� �0V�X!W�(D�TJ�fAg��RG!�B�z,Ba�3D��A��s�r�񧩏&;����'D��0�?ߖ� �L�]�>���$D�|�&���x)�K�4�8���'D��(�.�']rJI��#�H�S�%D��'�9[
��CUg�.2�@"O%D�8j6�N�cڪ|P��C�b��m$D�����>߄�	&��#�HGB"D�$;��Ǭ$2Phr�<qk�f%T�ԫqB��x�p�C�ռ��ԋg"Op�9!��1����FH�I��,H"O�`R��5G3�HX1f�`�l�H"Oi	�h%8�ޘ*�EO���(�MP'�Xm�S�'y�]�h�i�쁫��ޣy=��
�'z�br�;lM�Q*�K�i�ZPa�'ΊtQW�Ÿ���bq����D=�'��<���޵{��0��H�P �'�����IӧS8�p��.x#�"�'���J���$P���Չ�i�2�Y
�'%��e�	SX���ӵi�,`	�'��<�b��<�T`�ٝk2�h��'�����+i��%3��g&�4@�'_���̓�}��yjs�=\.�U��'��q�F	N>8̣�h-�K�'L
���IN�XU͕�';
1��'6ހa���/�TPQ�T��
�'Q��XGD˞<Z�\&�6 ]l8h�'���3�N}`z�C�����'MR��W39�|`b
�.s�,�
�'�D��͜2�9c�ǈ�r.Zd�
�',��V+xfTC��ʺb�L��	�'��p�ݲL��-@�E�Rh.���'`����s=$ V�"q?0�2��� yQ�́�-G`e�!O�F��LZ�"O�"d�FR�PC��+K���"O�0�7*
�g9�tӀ�bP��r"Od�k��޽.�v�ۥ�\�E��ز�*O2AK�j�g\ y�k�Lp��'a����m	�j��u��E�>H��,�
�'F����R 
,���b �J�"���'h�Q�B��f�D8�	�
88�c�'y�2�jY�S�\�K��M7l���*
�'���p����=�c�
+g�80
�'z�͛Ň�N0��b��	U5�s
�'�s��C#�p�'�Y.B���@
�'��]�W ��2�U)3����'b���%��! %�16����' @��P�w	��Q*�?"���'��Q�"ؿO:���ƨ ㈥��'�P����@<`k�5���|�h�'�`�F��aH�!@�Y0px����'���24G��<��+���3O���'���k�kݱּ�J᠊�z9渪
�'��t2���ch���BF䈐��'�6!����%��H# 
՜!6� ��'dZ����SfD��w��M�H�	�'��M¦Ȅ����` pM� ��'\����[:�y�WB���b�'/l�@��<y�����i��!�'$�pP�5�9'm
��(�'�D�aM.*R�pIv����"�'����F�L���y���Y�'4�(�<|!$��d"V�F.x8�'�D5�b�,&�g�:2�}��'#�|Z3�U�P�X��ǽz����'�,�т`��)q�dO�p�Z�2�'(y���u��m��%�1jNZ5��'*� �r��9#�Y��̑o�#�'qxD�"��k�H����b�
���'ff��3��J,���劔Zc( b�';�1aaT836-�b�[.�<ĩ�'���&�UW3�X+Rɚ?v
���'��km=b�����e1v�j���'=��!�ʊ*!B�: �<��[�'�	Y"�Ww�d��0b*)�ո�'�~D*���u2��շ
���'�ZBZ"N��a����a M���fF�=�a��	D ����[�nƤ4�3"��J�$��dƥ@�b�R��(j&�q�ܿ@��X�[)�щ
�'ov��ī[8C�ػF�K�t�6�qڴ�zqCG(��I00����N�/���k�KQ��Ol���"��=$!�$�*�<�A`��-mg5�"h˩i�BiS/�����P2*�剥Oc��G+GϠ�'KB� i�I�V=V�I��(��9�ۓ2h���AX:e����*�Q� Ph�/	�Iy@��]�8�`�}L�d�3���1��qÓ+&8� `�;�����jQ6`2Q���5)8��&eD�dM�C�?M���E6,*&��ץ��[J-Sv����\�
�ԍ˧e<���B��#aC���`s� �IL&|9��?>dxQ�'
���C�(�S�Ç���pC� μkV �FT��ꖅ^=2�B!+�m�r�<�rU�6�"��r�O9m��t#�$� -eV]bS��.������ȶO��&%4�,ɸ��N�n��d;�h>U���5"qD��ň4f\Ԣd.�F���"��0&xyb�A>Lx�}��M�.EX��EL�M�&�($��+�Ԉ��0][�XᤌR@CFl�28�Z�?�n˂����*�J�� �%��OH���!�U% �L��i���Ĕ�m�8�E�Z�Y�J�a��BY���s�"ZƮ��U�@,=0ߓ�
�@�'��|��K�JI�/(U
P��br�d�l� ���²�����P�g�}��s@�-(,YZ�;fþ��w��u����Ad��1$�܄Ɠ=v0��١�|p@gY`C���0gÀ
��9R
Fr{��I��
y,� O�����$�Fl�Á��v��Y������I�B�(~qX)���?��U��a�+y~D0׈�V�? ��[�ĕ��I����b�d�P�FH?q�F\�a
�Y��	6E��K�Q��O$��Qe
�ڐj�9+n"UHP�-�D9)k,u�ĨCZXɑ&�)�x��"�����S ���+ģ��W'.PD㓑&��6-�u�l��w*�$��=�&��t�g��'<� h�P*NiD á�~�P�#� �3��t�F�ĀSA����U��Q�3'��2�Ε4�9��&4���Ù-, H����%��(���

5��� U�x*��*
�8x��8�#Y�/Z͗'�����BD�e��yIr!;a<HB����ŢT�'"1����W�vybq/�	����qB!:�%)G��N $;aH�-�<�OY�����0^�q���	�O4:m �%��x��$Y'mk�1O�,Ag��
n�����C�qX�KH�s�⭘�8��PA48�8	�I��Y̠L��"Ot���� ?Ԭ;���*n6�K��׮z��1�sAL�ft�&�B�`�җ���"�y�s��:2�і'Š�HgFO��yBLs�̑���^j+�@��%>1���H'��n��͙b
�iW��+Cl��r�¹��d �h((H:���;�xe��KT�cKa{r��[`���If�H��r��g�䉐���u��(��	.�x!�	�
z���$�:�ڭ�	�(�d܂�I�r�O<a����r&�;�n��W�рu�1�n^����#E� l�hT'G!��\*F�i�1��j�2��D��"̭B��؇e��vlBNrTe0pbܪ�(���Mnt��֦��CS֙�����!��^~��$D�9'�
m�bV-A��ѵY8@@��cn7o,~�B�۟�#=	s�1A�d0P��"�nxU�d؟X�D�)d�z�2S�3�Xam\�����P,0JRH��kX���j�T��(S�'��f�2AXV�.��r^�c�Ĝb2���T!�~��@V.9�<QJ����ȁ�^�<9�
�+o�T()RR/,��!���DXy�$�L���G�Z fD�F�$/TY�x=)�<�����Ő�y���,�&��{��0JUU��y�1���d�sϟR�Θ&?�X����%��͠�gԡ�"r�C3�\ДIHcpYp�U�x	���O$[��@�AV�;	�B���	�`�K!��ޟ)���	�@T(�����yz���'5���v[�L�8�
��|����	�'�t��4dۧ;Wb�M͌E>��P�y�G;��@q��&����"'��A��,�dC�>R �	`�c��s���93hޟ3��3%�;�	�Q>˓V� #�V,A�̏:��Նȓ��D����qt.��d��R�Tȅȓ|� EA�"ǩj���Ʀ 5V�9��P}�]��'E�4�0��8@��Ȅȓ:d������6 I��X�j\�-ڬ���^~M�A���q ��c�V =	 ����0��c�}���S&�)��`$ �*4��9[Lr%QT��NR����2e�pG����x5�ؘͦ���M�N ��/:�hp��>B��Fy2�N!L�JD��l��Q��Hz��>kvhp�bː,�y�*2P 4�⍷a���HB���v1+U�A2 ,�|�J�>E��'�R}�"�٪R�P� �P���3�'�̠9d�G%+R�� ��3Lթ�C�pL�R�� �z��d�`�`�����Jcd����4>��{�8f���oV�v �i�J-q�� 5�4���+[.�y�H�'� [�(ѥq�*�b�oI���'��1��ǐ� I*�E��M�>dt�� �c$6��sB��y��ݠL�@@��h���S�'��%�TኆwZ��'M�>�	�1��4�G)`)��#H
\�NB�i��b�k�l�ؑb]3G\��c�!�ORt�6M�#�!c��u��jA;(����JJ�4�nх�ɻ2���������^���ui���>�Z	��������2u�%c�$ٗ7�DE�?�҆)7|�!��)�'9m���!�]"Aw�}�Qʆ7!]JT��A�� �Qomb6���A��`6'۟?����|��9O`M��[��@t٧C�Ȩ�6"O M�!�2=�X�� �H!6�O���A����0>��/Z"PI��q#Ձ mZ��ay�<�g̶G�%(�`��,L̤�FH|�<� 6](Fm�!�J��*�vB���I+�2U8V�S>B��QbaW�M��AIv�O�D�zC䉶6��C����F��UPD썠W~m�!C
��h$�"~ΓfH�Y�l̿��y���?hu���ȓ)M��B��/V����5xL����,E���ZŁэ�a{��+Pe*=�D��n���wkK���=Q����~���Y��n���X��`����`{���{�!�x�������O��[5�Ϡ /�O��!�`0�����)؏H� � P*�P�΁´�D8b!��M��h���H�,Τ�ՏܗCD�I`�5^����O��}��?Ĥ��E�i)�t���J�8���7zb,�Ӂ�gFL툃:���I"8����:�a{R��r4���;��U(�m���=��	^�7Ѣ�!�mӀ,8�oӥl$��R��ڜyb��*�"O�i3��+>�0�F�dg� �A�Č�b?�:����H�: ���9�Ց���o0pK�"O�8����Bd�աۘxX�����[��u�*���S��y���4{�Dh�6)�#Z�1kB���y�nئY�#TL"9�9�A�>�~rH��[bm��	$uD5�U��^ ���º'�B䉁f�Nm���6 a�}x5�#V�jB�Ʌ�����T= �� 8tgL��rB䉺���Sa��T���!��B�I�h��+���>|r1�
�#K8C�T�8���  k�(�i� #4:C��#)S���p�����*�M�9<Q�B�ɪN�ƅ�$e��I�Hx��$bB��w����ANI:/�D��gg��TC�I� �˰h@�$mTY�w��G�C�Ƀj�܃F4@*�:�E�5:C�I7!<H�#X���V ��v��*F�4D��s�H�4 -^5���� y [D/,D��;�8C0iCv�Z7,Q�CL+D�T��O%bRt�DK=r��ԢS�)D�гfPK�<��)�+��Щ#)D��Tgˎ^���
�E���x�ᴧ(D�Ĳ�&��Rk���Âw��;�  D���4��{�2����!zH�� ��!D���D]U	|�p�߼_�\�"D�dx�I���1`�,]5?���Fj!D��2�n)`�4`���yA҄��G0D����/D.�@�4j��^,B�K�*/D�P0�-�bx�LYEH\�0�*O<m Ӊ]�A$P��"�h�3�"O���_�/	�xR
@�Jv"O�a�G6*��h6�ϴp����f"Ox	JV���_}l�G���B���P"O���Aƃh��P�$�P�/�$��"Ob��"O5b�zh�6�W9+�.:T"O"�be��"�^l��
�k�L��c"O��z���<�0�Wc�O��L�"O���G"�:,�@�J�B�(��"O��i��ٕ1���P��� ���"O^�"h�0�̹�󅋾8�ܳ6"O>���#����B�͛̌\��"O����H��9iR�(
o��"O��%�[�:\�E!U����"O�p��	Y�9�S�M��E�0"O{^�8�6�W'~����pj�*V�!�䉓L��h�rχ� ֤��eU�!�$M�?:^�t$�P��My��֘N�!�$ύ���`6��k��=�@�!�$_::2d!V(��4��mӢ��0]�!�d2m�b��26����A��P!�� �t�̓��X�.��0�T��"Oސ�t��~*X��f-��7�����"O� c�m��<5�<H����Z���s"O�9#�KB�t�\�5N��9̈D� "O���K�6x�����#.�N��"Op��$(�kBbm+P�¡T��| "O��)fN_�ր`#���Z �,�E"On9���E�O��d�cŲ\�@��"OȘҰ�&F�(B������´"O����̃M[��z��74�"�ʵ"O�)@��/���B�A�f���W"Oxl��H���-4Qv�z"O��	#'�!c?��+Zhx��"O����o��
��5ӖH�?m�8�T"O������(h���b�JI)h�"O*B�Lݙ;^1#6�9M\p��'8�5�� j��%��������'/~�ǂѿK$.��2�nb�2�'�D���G�N�z��N������'�z�AR�ͻ� y�1�T2m��'z��%��&�\���כ���r�'����!+�8{��H��q���'n�Q����hʜ��c�&]�`��
�'���b�-(��L��'Dd;L��	�' ^	 ���o���"`]	μ�I	�'J����I?�9���6��X��'q��3�,�,%:�Q��Q�pT�
�'��ȵLà0��8"ȇ�a�
�'!.�ˤ���qc���Dԫe�fM�	�'�\���E���ޠ�����Y���'�p��֬_�a�z���ĉ�)pj��
�'�P*�h�;��M��j�� ����'�٢D
zJI�.�<�
�'֖0S�$־ d`��.���'r�)�(]2"m'�y> l��'�V��Q@n�z�ӝ����'���b�F��(�02D	����'Q�|2EmU,|�~�xRň.he����'��L	GgW,b��#8N�E�	�'�6YT��?9��`�2�2	�'@B����3F�P�J��7u,=��'�����(DI{ץG��t��'Drx�%gN�Y�����eɷ�)�'��@�g�J10��E�U&hM\���'���3�*���s��6o�H���'*��(G@I��0��&ܗ_)�\�
�'+�]�F��Ecn@1�$H�FO�5��'���dΝG�p�[�4o�Б!O���DV=h܎���.7Pq�m�a��B�x������<X�Vd���ϔ$H2��Ic��*D)�-}��DA
�'���D�M�u��P�Q ��LߒѠ���V-s<*�@���"1�tb>u�0dMq�����=P@8��6D� 16��5!@�u14�έ0WdxjC�O�L#��Fi��:3�<E�td�!r"H�$��Q{婧�2\���Z�u��qP���23�X�J5����P������M�)�P��$�z�(��I��h+�n�s�}��˔���'!C~�.�2P��r�J�b ���-i��Ot�@e��Z"�*�e+��%��ɸ0t9��@u�
�!f�����T�3j�0�(xå͐?�C�I� �޹�wƚ6G� �u�!.T����zo�A#����[a��`�T���O��*S��Bz �Y��H�%%	�|�ց�#����?��@�7�H��'��P �Z
9|��Tk�5jw�	Y¬Qw����]�H�@��O��H�F��-�����M?S����A#�n�v�ʱOH�f�#��[_>\�oG�o 4�i� ��sh�`Ԇ�8 �
T�&�ÞB�"`܄�)� `�K��ۦlB($q�\G����"�O2u#�a�m�(����c��-��-�6 �0�6J�^a9&�Ok�,P�+ �`)���
�GL�8+�'ʪ�9�Œ-��s�a����+�L�0�R$���dNIrpo��Gƾ��;���xI�λ}��x	���eG���n�
�ȑ����p#�QK#e[7\8+����`��z��8cŁ3$���a�X����-�=Y��$f�lA�e�ٙb�Q��/Ȇ!�Q�hBn��d�xq���e�a�o	#��	�.B"�&P�i���Y
$@�4C&��bC5�X���؏z�h�D��?M�dr#�>(G���',�CҎԃth��6�����x��ӦG>���_�"��P(Q�`��M�3`�,�\;�y��1�4�HE��)�|����T�{�Hp�
�V��t�b(���Nթ��1�>�p-O ���Ġ2���dxܑ�C���U�*LIu�#|O�hkU�C�Q�0�\r�"��8c�A��D>i a�j�+�F��>M��4A���BG�		'��l3�R��˱��-U����Պ�;B���Ě6�bW�Ђ^����'A�$PA�I)Cl�]�T����Dt��S0�c�U�t͛��@#�,u�X�|H�k�'P�}xq�N1V7��J�w5�E��FQ,n����P��>�8�'mr]��ņ����y�`�C�Hw�ֆ<RlD�K�$�����Ε���%��O�lCE�ʁ����F�]�	4���'&н�0 �8d��\;�� �x��aw��2,�T�`��F�\P���s-y��'�ZQB4HݙJ� �� Jם*�n��B%�� ����(��5�X���T/8R��(p1��lB��SPl�P!�0D��C"O,�B�ex�y�ÊtR2ى�A�".n�{�ٓ2(�G��
$ ��9�,I�'-P04z%E�E5-&=��"O�Ոs�V�� r�(�i�AK%���;�j�;�L!��|�P��Q��	>ғs����
�w]��yRa�'^i���+�iI��Μ9�|�"��z�
�q��=���)0ϵ.f��K/pm�\ �R�`Ԓ�JU�Fz�џ�!A�8N��a+�j���S�`.�13�E6��58t)/6�B��+k�q��kM�B]XA�F�<)�ZgS�\�!��2��#���"B�� .3W��UEEQ�<)t 9iI %A��� 3HQ0���D�����O�� jB NU���qO@���Y�a�@P�� iVd*�OB��#F�/^X�u �>V ��`�l�0@�h<�"��\X������ã�C�Z
$��V;J��$�/`1��X3��m-��;�L�)q�X���E�*K�4��ȓ%��]K�ƅw��dc�B��x�<D�ܙ@��pP����T/�D�ǆ�)�X�I"h!��
�tb�*�%P�r������UF��Y7�dS*�(��I8sR��9�V(1V邳�H1a>DB�ɍ9Pdx��ƕ�7e��;F)�N�4B�		N����H�فE0�6B�	����H�.�1A�a�_�W�B�	<U��dkvL�_CL1��Zm��C�ɩ��HS6�ؤ-���[Ac�B��C�$"f�]�r��E��z�-�N�C�ɴI�~в�ǡ���#�e�&;6xB�/K�h��a.J�t���:EE�W��C�	�_��H�¾�R��7����<�+��^��#~�В!�V��鏢&ZRhAu�r�<9Uj��b$�Ux�D��<�r���-S�~�����S��yR*3}5}cWN��@&x=@����yb�V7�����!T=�N�)E�_�?y��٪L]��4lO��t��&�R5�@c�</>�����'6�гB���oZ4����c��5# ��a��Rr:B�I7jZn����ڰ�Sˀ���8�уhؠ��S�v�B��#���ag�(y�B䉃X��Aa�C�*X�āC�C#w�-����<6P�J��G��'��}Y� �`�����5zL��'D�pnc����8BW2p��6�p0��f}�|��$�M�����dU&
��@B"�@�{BM .&xHt�Ԧ�9v.�cӢ���D�4C�M@�l!D�<"dㄟ#�x3��7>�%I�2���%L�HB4�>F�>e��T�As4���HL���y��N2D��r�A0@���	���z��0�� �+�+��\�)��<� ��!�˥/�����%h�q86"O�RjD Tv +&ӦzVT)�O �ʐCر�0>��j�i"H����� Y� ��X�<��˅6=6��q@�' �R�[ �T�<A�i�2 ��a��� iq0�`�Ek�'`^�R�)�r�O��`�6UXZ� ׎
�:����5D� �Ɛ	%r��ui;F�`BW�� #ub�b�i�)��<�b��s��=Y�+�.�M��&�_�<C��<�8�qa �` hˏ��T�#*@2� ��'q��{���'Di޵r���&)1
�����` � u�6�s �A��bHlE�O�co!�S)Oh�q�Ɖ�T�p˕T+1E�O��R�&	�T�ޘ��I�=F3��[�f�pB��)dχ6 !���+@�ڡ��	�(��5oڧ$r��w�E�]��O�}�"
q�1͖^>�#���>�
��ȓ'���(�2$�Ĝ��S�fN���I0V�#"8_3a{���6p���0!_2]՘E[v�ٝ��=�MY�`M��9��r�r�� BϾd��k�j�)��)� "O�b�[#_�0$��ՎY��P�s����{ 1h��7�H�X�Z�b� 9���2
t��"O¼�LJ$n)��@��ޤS�mѠL�(ĮP¶b+��s���EK�t.`���W���k�B)D�(\�m�4�`7 Y�nc��ẟhK���� �a|�lX�sT��6nP�&pbR/Ĺ�y�䋜8�`bT/Z�O�h|�q�y��6�~��d(�p��	�y�,��"�v;�Z�7��]&W)�yrn�8���Yk�? �z��㔶�y�Ő�3G�@��+$p�@�7	�6�yB	�b͆a�1�\ 3��B�W>�ybdȞ=t���Ȅ=j�n��"mL �y§Ҿ?�P����	�1i<JI���yB�+%��b��*�2ak�N�%�yb`ȧ������#��s3�]��y���^���ƒH� ��D�y�O�:Y�-��bN�͚����7�y�J7�xu�G ;	�\�NZ��yb�LiC������:ܩ�g��y�ִ3���u��xB�y���6�yr(Y�b�,s'����*
2�y,Z2di���e�>z��9:��D�y���6k���ؕM*��` )	�y���"��1�6/��@	����
�y��zS�`f��*�8-ʐ`ݴ�y�+��̸a8E$�5-���� I5�y�*A{���2�V
&8@���@�y���*8̺D�`''�Vъ�g��yB�2b*�ف���d:hSwj
��y��61�� B�6��.��y�
T���V��q/�E;_p�B�'�hJ��T� /I�Q[',VB䉁ZK� ���D���a�Z3�r%�E�ͱP��DT� ��\�Q�&�i�"M��"�!�d#|Z |�4*/n���"�!/!�DQ�&������+v�%q�A�=)!��0;E"c�	LjJ��3 N�Z&!�	5z�>�K�'O=L�U�����!�]�9D��#ݑ'/��fO< �!��Z%T�"��� >\S-��Z�!���ykw)�K��M ���0t��cJ$}Rn�b���Ԉ�?i��I ;��@��g��]��


f�I=�(xO�z���x��OK�A��B2[�
t���?T�~�д�_z. �5� �l���K�:O�>)��	w�Z���D[7|ժ�s%�H>S6�x��E�lO�q�G�Z��M�wʃF>!�f�+A��0ѥ��?hl�fnV�rit��J��M��!A��Ɇ�3� 6!wF�A��T���Y,z��ʷO��rf&t�	Y���ɲ�I)|���;�'xȢ�pA;%Ǧ��U�UNR�i��<O��SbLZ�X�\Q�4�F�OPB��q��0�XP��\6��D�ۉ��u�ʅem<��EAÈ�?E�ܴ{>tE奙�(���1��o)���c�Q_�M#�����	u�L>���4u,Ɋ�͋	7�$��Q
�	&� ��G���0h`������g�$l�ȓU�l�Ȧ�D��嫂�+>h������&��O  �L�=����]ud�-)���8e\�Pw��ʲ 'D�H��T�/7�ɘЅY>j������:D�pz���7K4Ւt�[�]c<Aѥ7D���������D8vĤ����?D��SA͗�Pp*0mz���'(D�� ����m�a,�Jh��!D��#�%"���9a�o�L:��>D��3AM�[K��1�	Řwx@�w�<D��P��\=:��°�z}�D�-D�12M�b�@-I�A�V4��C��&D���@�4�ܕ��_��J��W�>D�����-B˜]s���'U��y�O0D���F.�	q��P5č*:��%�H0D����pMr&+Ѩ{��Y�A�/D�$y��K�t@��2PIJ+v�`sM1D�h���]7~�"���d�eP�u�/D��`�ʆ�<��d��0ߪ��1D����k��ܨ'�Y�;p�h��':D����)�"Q�zaC1�K,
I�ѡ6D����ڢ����#�ĝlD�`Š:D�|��&d��ģH*���q�#D��!!�=���+&d�*zˤ�{$#D��⑮Xsޚ �[�n����R!6D���Ƭ��('fx��@0��r�>D�� /��t��l��g�
n�	�#�/D��x􀐹v��y��*#K��!���,D��#&K�H�� ���Ȳ�)�&D��p��[�4`�@�Ʃ�1'�����?D��ԡ�x
�Ycl\�VCĥӐ@*D��(�F���ڔ f������(D�|�%��8x`���»:q��U�!D���q-J�F��eƁ)���� D����a\�j�����V�i�̊�<D��h5 ��=�4!��OхJ��P��	/D�\��5F�x����(<s||{t�+D�8i�I	b��PB0�B�	�$!4�/D�x�Qұ[���[�ܘ:26�3�a.D��
�@O=g(T�(/����>#B�	�.�X�i�Ǧᒓo�B��<9��
g�GNr����NP�^� C�ɟ;Kxࠇ-X��������N�2C䉢;nP�0v,�|.�8��6� C�	W���L�@
�聒陫K��B��ܕ2ER�x��)�Ǔ�J{V\��'0�����X�0J��G8Z��h�'�f�Q�E�Y_� p�ϋcU[�'_�8�deәSX�����p�T@�'<|�3���|LJ6g����]�'��@HYD!�]8�E�t^���'� ܸ�c�;���
J9I	�'\�O�nƴ� ��Μ�
��':$�����F�"���48��'�J��-9沴���ؒW�����'<����@l����gJͽV��1	�'�>�鳅��n;���^�]�k�'e��1Ѓ1n�`8�j�b������ ������0`����Ϳ},9�"Obm����)M�1#�ܩY&p��"OBл���}��y�-��F�x��"O@�4�Ξ*o����V�i�&��f"OJP��)5�Y�A+��*"0s�"O���5�]�t�X�� �$P�"Or�1#��4Y	��ƅ�h���"O���!eH�\�m�����^��t"Oօ g.^ O��Bf��s���0�"O�0FI� J��"��j$Q�"OP��eEáY�^�W,�_(�"OBe*���W��̂��_0#q�;B"Oa�#�+���@�D�>hHԸ�"O*����H6�t��ӂ&^v�"O�Y:4�	�l}\̩��A�\��4�	�'�d��vɐ�%�@�U������'�К�OF���]iE ��}�X0��'�H${��E� �։�t�DD`����'��YS�� |�Qa'HєB�X�'w2T�$K�K�t�ٷ-$.{
]��'1�x4d��Z�L� dU*�͐�'��tu,�?"�`�OV�I��'
��㑋	%���#��׮	Ծ�0�'T�����Z>Mn(	R≓��ͨ�'�ZТ7���7�ЊffGxQ�=��'C�L;q�T�uP�B�Aښm��I"�'|6yiv��>np.Qc��_s�,
�'�}צ�sbd�H�ᗄ^��dq
�'C� y�A��k����q�G�&fr� 
�'\P�pQE�&v�~}��K�-�ĺ�'���a퐺Zr�=9�<��
�' l*D�96��� L�K�!k
�'5
{�K��A�N�ʠ�@�J�`� 	�'S�e�5��`�Ҳ�ЬH4N�C�'�v9�Ǹ��lR�NT>���'z����-�ڰ���جJH�q�'���g�=#��%ƜB�Y�'s���`��&�����#7*��A�
�'�D\hG*�;5&�q0�*�;VD�
�'��s&� �2��{�SX�@
�'��;b*�0m���� b?/l@!
�'<� �%lб'Ɣ�Wb�F�X�y
�')a��d��u.l�f�g��Y	�'r���fЭf���P��8`��'���2&O�4i�:4�E�O�)%���
�'<I�C��
���DØ�!s��R
�'%����ͅ6x�+������	�'��ݠD�7>�p��l��	t�1
�'��@��O̠
��*~���:	�'U��At��z:�M�"íG��Q��'�R�;aA�5P{�<�F�B���:�'�\�$N��M5j�3�]5��'���Q��P*������?70��
�'�ڌQw Q�BX	S6A	>a��d��'�P�b���&�����BH^H�c�'�vE�Uٵr<�DHBI]�Np��'���y�Lk���1'V#�x9�'/x�9�D%U��ZAX	PB@�'�F�ڦ&Ę=5Ь�᠞�p�����'4LQ�@�)��)�1��/��Eq�'�~h��&[;M9 ��g��t��	�'��<{S,z���%�̈́�\	�'���bD
N�	���JuC� |$���'*�kG�П�L�!U��&T��[��� <���E�1���	�34O�T��"OD��� ��"�a���h��i�c"O��z&�ً2���q��94��J�"O �E��5 �p`C�P��Is"OPh�UdZ�IW0����	uo>�Y�"On�+6b�270����[�5
�"O6�Є��d��H��8Xl̄3c"O0�{G
�s]tPkQH�@S���!"O�H��ɸ3��µ��	I���5"O+𬙧Y���S�d3�"�"O|	�S�L�.郆]b�{@"O9oL!c� �V�D>���"O4$(��Y�1	�b�MJaq"OT�R�����R�� =|��y�0"O�=��Y�!B|	�dS�#~�H��"O��G��b�|Y $��4Z��9�"OH����X��t#�3e"Tag"O��xQ�UWJ����#:��i��"O��� �x�D*~︹��"O\鹃��/.�ĺb�E�U��p��"O
�����o�w�^��%�+D�PqVJ21$�M�&ON�N����%D��XB��)z��� QF_0P"�#�'D��B�e�,4.��v�޷x��4Ag�$D��Rs�O� ��u�d��L�����>D� єc�8<�j% %G�HB��f.<D�@�烍gdL��fm
9E���I6D��j��ų)�J�i>v�I�� D��g�V�`��pI�dg1F�t�>D�LpE���`Z=�g��2�(]�d?D���Q]0Qx�|𷎛�1��r@�>D��;R��$C�
WN���Vʕ:�yO1S2�p@�J��TjF��=�yҮ�+!�fT�� F�D��e���y�$˥i*)i3�<HHd���y�ˋr��D
�79�:�l��y��_0f��Yx6�^'"��!e���y҆܇-��H�ɂ 6�p#7�M�y��̈hy���K
�B�xC�!�y"�ۚ-,P���NXM�Ty!�8�y�M�3,`�!F�\�M��x�s@��y� +�e�ԋ�RG���O	��y�#7�(����0L����eK4�y���0��jC4E��9xp�]��y�ʛ-R�9��ó	j�����&�yR�@'*��2*�K0t#����yңA��
�a�������I!�Q�y��ˊ4�N=�&�Æ48Q���y���C�A���щ��yR��mȨ���B�9�"������y2&�'J�h'aB�'�HS�>�y�*^QjℌN1mK� ��yB�$��#�I��=���PE��y����b�(I�l�KJ���@�I2�yBeށ`�h����΁�����ׯ�y�IH� i�Ο���$`�.�+�yr�M	db\�,����7�^��y�썲��hr��\b����y�ǖK1�(���H�<��F�ێ�y�� -�,\P�(�f�ӖȜ��yr�P�?b���TF�%(ż�Q��iH�Q��Rg��I��䗠0Z���e%�܁�.���!�O�{�4m��j3,STB h����EϜw����S�? �a���r�RP)^&�8@"O`LQ��רih��sURs�"O�p�F�S�2תA����5;��k"OF�8��ϲ2�p�iU�L'wFA��"O��p���>)t,B�k@�]+���"O�a��5�f�b�
�;���"O��o�;��L����i��-�u"O�A��9̤��� 3"rPy�"O���S�K+r�Ta
�a�4CIA"Op���B4
P6z$�Շ"��eI6"OT�S�'�9zp�j��6Oa
i� "Oz�w�OoL�A�̟6��p��"Oxqj��> �Ir��l� 8��"O� �����b#�ܛ� %"O�ሆ�"�(���o�
ai$"O`x1B��D���P��6lZ`���"O���"B��~U�)�cC��Ii��6"O�j%
   ��   �  l  �    �*  �5  _A  YM  �X  d  �m  mt  �}  F�  ��  ؒ  "�  e�  ��  �  ��  �  =�  ��  �  _�  ��  ��  )�  ��  j�  
�  [�  + � � n  �( 0 U6 �< 3B  Ĵ���	����Zv)C�'ll\�0"O@��!�գvk�b��z\6�qe"Ol�** !$���Z'�� |d��"O
`�(�;���8���-0��1%"Oj4��ND^[��"3/9�0|H�"OB���H��*�ʞRy=a"O�味V�!X��!&F�:J�$���"O,��a
���C�Ą�M�"O,$3%o�-���p���+Ն�:1"O��ݢ1����`���y14]2��i�<�6��{_���c�H�`�fX�$Kn�<��A̼VI�xR[�)�Ć�pඤ�ȓA5��('nߡ4�� �)˩%� ���,��r�؊b#`T�eT09���ȓ!�b��g��}�8�F��-? �ȓ
K|m�ș�VṔ���2�%�ȓ"R�X�j�4JN�1�˘X�i����̹	_�jZ��1!g��zܶ��ȓgil,*�J�
j�Ne��i�J%b���f	�(U��:���G��$Y^م�~r�� S�%T"���k\�jx�ȓ|4�1�îJb��@ӵ�ݩn�V��/[`�"�v4�R�!ʎ<��M�ȓ`:��z�ؚh�J�Z��$HY:	��H��p�m�C1��!��B:��0��EnjZA V;9����J[
2���	��4'J�EA�IVW&��~�(aZ��ӹ�>� o�Y�|�ȓ�f�A�
Ο7�H��M�$�����mޠP����/���ANXo*�ȓTv�����{ ��-7�*h��I��sB�8�8���3����ȓNe*M�悡;������X�o��!�ȓ'lj�#F�m�+R&;�|��2)n�C��0S4���T:
b���:�0!��e֊��)��ͷV��,�ȓ0�&�8#���� ع�L�����;�P�AFd���,w�6d��r�EQ�( �gVlɦ�M,H��,DP���|�I	$G#\���ȓ"�)���E�B	yt&B�^�LɅ�4�� ��eëF�ڙ��n��R�p�ȓp`@}bŇ�=�$�AUN��P����L��p���_�a�)�Y�!��-��u�5���o}�`iF�@A�p ��F�\�0��[���IF/5���k>bTؖ�;K'DT`�^��@��fnV���Y�b�lI��	����ȓ,nٛ��Ć3���kC��8�m�ȓ'� I ���x<=���޳{��	��6��(� N�����
�y2<��ȓx;6q��I�
=  yG�O�,�!�ȓW�>���.؜ɰB��;�����`9"�ˁl�$@��- G��D�ȓ���zF"� ~\�`%�[�ل�E�1�N�;f��P7�.
�T̈́�4 ��QS�[@��o�|h���h�c�A�,@�X*1�֧jN���"�q��� ��Hp%����ȓ]�9+���.E��T�qA:!Θ�ȓ<d���jF�,�*x�d(�9w�Ňȓg�\x�b��/k��<8�ɔ�(��U��Q^��ç�	)��c���d�6�ȓ��-	q �Gp�p�ԭPpGx��S�? ��KG��"����(���sa"OTEq������ �+�+?�2�R�"O��.ܮHְL؃h�2��""Ob�iU�Dt�Z�p��Ը�<Ej"OF�qSƏ��EXQ��'��Y��"O�|c����B�d�c�8X	c"OP��&�\ �za�H�A�P��%"O.��%kְڲ,�+v����"O:  dZ�@β��R=��IrT"O�- �Z\tu�[�輑�"O�×@ RJ���#qRaF"Oz�8�䞐%�L�FnM�blt�i�"O�q�t��|M�j�,�/S&0�"O$�& r�<�J�%kX@x1"O�88Ga��\H&�+�j. ��m�"O�U[�N��`��'��x�t���"Ol�Bp�^*���������Q��"O��E"ěI�d]�@�8n��Zs"O�%�R�U1pС�6�D,�Bzr"O���6�ۖ%�vP0���m���R "O�	�3	�07�Ơ�`"�p����"O�Y����e�@-B�%���q4"O�pZ�=E� �:���?���C"O �g�-d ��IR�Ҁ]�$}��"O�Ѓ�DQT~�Ċ`��"�m��"Oj��&��!U��p�ʽB:Jr"On����&�jE�C' 	v�BE"O�,I�	�(�  H�O^%b^e" "O|h
ĄG�I�&�: ު(�&"O��	DB��g�R%Ң�¹b�̅!e"O8�H��I*Hă�%�it"L�B"O�邵LF�T�"}��ł�e8C�"O���q�˴K;�����\�fz>� "Oy㕋ͻ5�i8��ݮ$`4%#6"Ox�[cG��0��(��&xz�D �"O��;2�"$"�Z�Ub�с"O�t'$ǔk�����O�؉�"O�U��v=z��cB�1�C"O�8����N��ч��؉!"O��6���w�@zU(�?}ʴAS�"O~Ab�ޑYp�yQG٣A�Bbf"O�Ya��=!l���Ɔ�b�V��!"O�!)��Y�fx���eE\z0	J�"O>��pg�0Z�2=�C�A�Hy��'���^8�'HZ�L@t{v��Y�!���m��h�U��{B����M��>�џ F�$�3mJBd"`����:��V�y���%vd0�U{N���c�҈O����N���1��3~�\�QWM�l�<Ia��V�8�a�KŮ8�B�gK�d���=�҈�!U����@ޔ#	�a��Qhx��'ʴ���W�Bg����(�vD�d��/D�@c��уo�0܈�`ʺh��E��"O�7M;�-,����.J��%K̰F�Ʉ�t������;kX���N/Mc�E�u��8�S�O�(���,Ui�"չ*���'��4�B�'4v����[�&u����'Px�+��Qe�I+��O�T�`I�K<��O�c�b?my@A�R�)���E� j�KQ�+D���!��pF(���$_�3��
�`.��C�&3lXG|BV�@ZF$ߕ1F�)�fA�Xt �(�,.�����{�B��c�	Fik@�)Z�l��Ɠ&D(���L�j,�p�6"$p`Dx2�|��)E:�A�'M���H�n�)�!�� �3VdL-0����Mִ6>`��f�|��)�ӾBA��S�ل��7�� >M��'a}���H����h_1V�Q1f��y�dޯ<y�Lj��C�82��+W��y��νf�z�����@x�"��O�"�c	V�f��TB���`�~��6J�x�<!re��t�0��LC#J� ��ʂ|�<� _kl~�B�L[��"����{�''xF�D��V����,�/xrL;P�]��y2��/��\�b�?#��(�$���y❟P&����7�$5�K��,itH��&PņȓW��E(bw�h�&D߽k����ȓ}�J$��
(f�Y��NR9��d��1�`� @�]����B�E�x}��c��:4��B�*��$g�,B1���0,O��	Y��,�(����n1>0;��P�=��B�I�_&�`��E����FMλ�˓�hOQ>�I`� {����H� *H�#w�0D� 1d±'qX�s�ݔGs�p��P��HO?牡a�\�s EM
S.rpB���'�����)}�I]�~e����%���z�ϔ��MS�'ya~2��d���Ɂ�Z�r�(H�#����p?Y�OpP��O̔r��ࠥD��l��"OZ��� 
�z��4Y�k�UG�����	\�O��LX�MBF�$U�E �$%xl��'2l���Z#\/$�u�Q�zqj�'" hcT�Bn�4b�*9�	�'���Y��ǡP145ڳ/԰AR���'�6�#m7sv�Y���q�T1Q�'�8�;��
4N�(���زle��P
�'� auE��HP\��4�X���)�'�*}�c-N0H����3W�}�B0��'�aA�E�%
�lI#(NL�l���'6�j������KU5C�~�X�'���	� ;K&X2��-�U2
�'���6�	�@:l���Ɣ6k�
�'K6bT�=iqx�����2�'�H�����%���k�ǌ�ѴM��'9��:

34&�؄Gւz4���'��|�PI�ؘ`$�%p����
�'԰	
W��6�1d+B/4`�Z
�'����"�đa>���SƁ�g���	�'�LC��"r�6}�BK	sy�
�'�حe�Y'y5��[�)\:��	�'�&I�Sˉ5�0�Q�ٱ���J�'�\ԩf��T3�C҆�5
P
�'�FEpơ�de��	%*�0�B0��'?��S�:,p
�ZT��2*9��'��=x�#S�(��*b�x�
�'?�h�Dh�d4��cM��7"O��Ƈ��[,P��P�Q�|$���"O�yt� 4,��s�P�Qb��8�"Ov H��B�U&8��"_�2I��1"O`��I��N=��@�*1,��2"O䱹��ʙq���p�o�.`D6I3s"O���w"�u��:Ί%dpB""O�Yh���7>⌻���w콻�"ON��D�:M%��sթ��8.9��"O�ɱ�ː$W�� �S�L���:�"O��3��a�jXn��=���"O��a�ܷ}J�0���K<b2�i"5"O"�b����b��
c@�À"O�@��˽>�=9��3��8u"O:dk�Oˍ_ņ�C��L�ƌ��"O� ⠲�уr��a#׷Ԭ��"O��;3 ��T]F�� �#f���K"O��qD^�2��(��Y����"O����W#44�%��B �X���y�"Oh��l�D��cDIҔB�"�i7�'�b�'���'R�'s��'���'���6�{��85n�S��%���'�B�'�B�'V��'���'�b�'�V�z	-74�H�ƩV�l�`�ä�'���'���'��'��'���'����L�#n�F�u�>�>����'��'w�'FR�'��'�B�'�4�z@��CG���r���H�˵�'~��',��'wR�'��'��'p�ؑ��µw@,�(�B��H�6M���'��'s��'�b�'R�'�R�'u0�+�'�`���2��.K2����'*��'b�'5��'�R�'���'_��Z�/�@�di�S�$Y/�Q ��'���'eb�'�B�'�b�'��'��� g/����ن�޷g�aXV�'���':��'#�'2r�'c��'Z��L Oņ.>B�#�Y1�?���?���?��?���?���?�6K#+/��#���}8I�Cc�?I���?	���?)��?���?���?9��ک]QE2�8rǄ��F7�?!���?���?����?���?Y��?Q�-�T�x�D�J�i��� �ѷ�?����?��?���?�Sh���'\R!K)cP�i�rHP�3�b1s��ʁ-[�ʓ�?�-O1��Ʉ�M#0��̢�`�K�!N
Jo��'\�6�0�i>�	��4�5H��n�@c�Ӡ���@@Cӟ��ɕ$x�na~b6���a��ë%(���$h~H`U�L1OJ�$�<���N8za�٣��^�h�4c�8qz�n�"~b���r���yGK?OĪ�{�n���(?q�P�	័����	��+��6w�8��B�x�bc��-��-i�tϓ6g�Ok�����'ժ�Щͦ���;f�-dPѠ�'��	X򉵞M�1 �A�*�@���'*Y� uY��S�8 ��"��>���?�'����^�l%�E6��,�5	B�!���?Q���'C���|R���O��8�`�P�C�V�``� �K%p_6�.O�˓�?E��'�f�c�EC(>���@�֠I.2��'�6-F��I��M���O�dS礉

Y��a�K�>C��y0�'��'�"��^śV����'j��M�)�`�6�"'|���Ay��&�Д��D�',��'^��'�Q�bD4J �*@�?4VZT� �ڴPv�����?����䧣?�a��_�b�ءC��e��I��0J�ɶ�M[Q�'މ��O.H%�W#�=y�A�L�c�*BU(%�R�S��!��H�V�b/^�Iwy�h�A[�0w�փ|��ATH�r�'�B�'�ON��M�0B��?��.؀٘1`�F�⡰U��!�?�B�i8�O`�'-�7���qٴm�jX�'��5\��S
�4�> �0����M��O�H�ؽ�����wz\Ţp�L�#pV�ꖤ6�`P�'��'s��'@��'J�H�x�G��`C�([P�A�O��X���O��$�O��nZ����'(�7�(�d�$����%��-.�`���� 5�v�&�@��48���Op ����iU�	,X�Au�Ň^b.��7���w����n�U���]��Uy�OeB�'@�"��B@sTZ�'�y��xr�'b�I1�M�g
��?!���?,���	r��{�6���"�2�DU�Ҕ�8[�O�\o��M���xʟTА���
�Dh��T�sE�*��7?����T�l@�i>9��'̀�&� j�jڅ<;(��3��]Tdh�����(��ٟt��џb>�'��6��>���Nаw�諥a�
"��-�s��O�$�����?a�_��Qܴ$HVk�e�B��,�tΛ�88K��ii�6��5866?i���M����,��g7D8b7�׬2�ك��yT���I�t�I՟���ɟ��O���U��lL
$��Ѿ�
�p��kӪ�����O����O
�����Rʦ睪i{��Q�C�0j�h��0$��޴}��#��	�!z�6�i�X�W$X@�����e�E��m�fl�$ d��[T"˟V�	]y�O�b'�|$8ѷ-ԔF�<a��f�*AR�'�"�']���M��#�?����?I�*L�x4�Q�~D�*�����'p���?y����A�1]�A`�JU��P��B~�
�>-��{�9�O=���I;j
B��!��Љ�E<;������� _"r�'�r�'^R��̟Xb����MSTb��~�ʤ��	��(ڴA��(���?�i��O�� �͑��- Sٲ7�J	,��I�M�"�i��7��L7M$?�u�Q�H�I}ݱxC�_Is������#IL8#��%�d�<�'�?��?���?Y拎�n��ז� �ЩKd�ʂg�˓?
�d]�Vb�'����'�� 	�& ��[L@��1	����?��aI���Ozj�p#H�u��K�ɔ<Rk^�ؐ�¦o��8��Oм��	�?	Dc3���<�f�>Fs�I�e��0+��PA���?����?���?�'���ɑ f����{C�U�RQzg�>ROhe�� ��49�4��'V듍?��zN��-�7E^�� ʒSB	 ��ŷvY&�
'�i��	���1ۖ�O�q���� :$�"���b82�(Z�K��`�#=O �$�O"���O���<�|�5��:^#:��A���A��\���$�O�a�IA ��OP�mr�Ʉ73Y�����3PN,UY\pK<�s�i0V7=����Q�r�l�o&�?���*fe��]���V=nC0��+����4���D�O����]nm���  ��;b��l�*���O�����M.���'A�U>Ź���x�x���'f5bH�<?�A_���I��p�O<�OM�tk�,Mlw��t�,y��P��K�V���2�����4� %��@�O����$�s'&���bR��VA��O����O*��O1�X˓	&�&�**x������4����&�2Y�����'[Ҧ|����H�O� n�%4�>����'/��P���ϛ��YP۴T��#��5���������!-���~��!9(����d�R�YP�_�<�+O<�D�O��$�O����Ob�'=�PUT��&�M�� K4`� �1�i0�����'�B�'x�O�҃i��/x�8U�Z6.0�
&G�  �I�y�N>%?ɺ&L��)�|�����6p������`^�m̓lji����O�N>�/O�I�O���٧G�����h8g��O���O����<���i(z�H�'"�'Q������{�)K/�w��|y ��[}��'OB�|�K�T�>dH���`���+�b�����:E��]A��ՂpZ1��Yi��uZ����15#��� �ǟu�*]��A�2����O��O��8ڧ�?9D5g�x��� &  P�N
��?i��i��1ɤ�'�"o����M�b\A�d��l"�є�S�K�������	ٟ�P�%�ɦ��'f4e�����?}��
��)g���A�D��;5��H��'��i>%��ϟ��	Ο�ɻ=9� ;�M j蜠7gҸ}��T�' 6�Q������O��$'�9O����ǁ7A����� ޡ { Y� ��F}��'1��"��).5jġ�W�5��s�ýbj�v��x���{yĀ&�'�4�&���'��8��R������y
�(��'~��'u����U���۴���F�ꁙ��0$g*�����7<b�Γv4���F}2�'�R�}�r��V�A���7rRv�#l"@�8��`Ӯ���1���j����w2$�E��q�X���b�k���ʚ'�"�'��'��'����'M���4x2�N6@d�Ǆ�O���Or$n��.���'1B6�'��9A�pkD�U:�!X":�1��<��禉���|b5%)�M��O��d֒
dl�r��Ϛh
���Gj��!0P=��Mx��OT��|z��?���]�(��m�s��#�dR)Y����?�(O�Mo��q,��ǟ���l�����t�@�p/X|��M���$p}�q�To�7��S�$�Ò^��ǌה\rJ���V�>���n<�x1�O���'�?�bf.��ЈKUjm��;j��lki�w>��O��d�OL��	�<q6�iSv=�vf��(�nXc,և�ză3���ldr�'�:7M>�	���d���5{1/�,a]���rP&xbI��M��i4*�w�i���/`�h���OD�m�4 ɥj�"_�7��;���̓��D�O`���ON�D�O���|�v�r���Q�Ɖ,/h�HdFܖO'�F�>���'������'ܔ6=�l��m�Wޔ���JEU��!�C���M��4!����OĬ{v�i��JCp\�2���m�<����� zf�d�*)�>���r[*�O8��|�����BpG^� <ʂ%�'w
�)���?��?�*O�l�0N��I՟��I!��;���O"<�dT,w��?�@W� ����	L<1��/��	C��%v�>��N\~"��K���c��טO����i�t�'�d�i���w�@t�Ι<��BP�'��'���'��>��I�SN4l��=#��+��
S|��I3�M��g���ɦ�?�;`z����6ud8f'����?i�dw�f͂8�����,�3��@e�$��C�P�G8~D��Q���%�H�����'�b�'X��'g`�SA��l�*=h�eۍJ�p%*�W� *�4{��Pj,O0�d9���OP}��^����Z��L� !"ѣ�l}��'v�)1��i��l�׫^�8�${ l�.s��)Al�~b�	�@�#�'���'�X�'8|�f"����rR�˞.`��'��'E����P�<pشj�֍��^�X��c����t�P$c�t��r�v�$VL}��'(��'�����`tÑh�; �3�ɏN��f��4�'q����)���	볮K f�Ƭ¶éT��s�<O��D�O�$�O����O��?	�T�QW$��30IW7����[���������ٴ�bu,O^�l�\�IBh"�h��� /J��z�2B~%1L<AѴiK7=��j�x�*�"��E��Z$3b��R�ŕ�
$`p ���,,�����䓭�4���d�O2�$�x`����G�!P�(�AfC�
�V���O�˓(5��	Z�0��'y�Q>�(�FZ�9b����^>d�RyC�k2?��Z����٦��K>�O�Z�
���DaA�Z�}�Zy0D���P9�hh1����4�B��,�`�Oր� D�0��+���"�TX��O4���O6���O1�J˓p�V��X����!�͝����Q�W�I]�(��'��m~�f�4�.O�6�W�@���l�Q)�)�6� �m��M#%i� �M��OV�
���K?� NjC`�z�����Ԇ7 ���5Od��?1��?!���?�����	U�@� jPe�w�R}�^*
�nZ�wS��������j�s��*������GA���`��f:(K� �?�,���O��Җ�i��M�h�^��E͇�[�"���B/Q��8u�^���h.�OT��|���yi�m���VjP����Z��"�I���?���?�(O"em��8�Z��'�N�|DZ⣝�B���ä���.��O��'$z6̓��$%��@���*�Hd+��`�D�0?���G!� Z�iE���'/�>��D�?�� ���܉�H0J���A�n��?1���?i��?Y��i�O
U���Z9�ny��H�?o�X96��O4�nڊ";Y�	ߟ@�ٴ���y��G#��E�D�ܝ��㵩�y��H��I�9����e�'���%��?�0��O�R� �U��P8���Ni��'���8����	����	
7�x�{����Qx�zcO<i>M�'��6mn���D�O���:�ӗZz�Љ3cͳ)8V��6��	�|(�,O��D�O �O�O+l�`$ӥr���P�&B���IԈӛ�u�I�|y�፼D�2���%��'��+�P|�V�W�4� �ɂD �$�'jr�'0�Of�I�MC����?���J(W�(pE�a�������?���i��OD��'b�7M¦��ٴ#�`$���ǥy���렁ۇ|��E���MC�O�a$�-�J��D�wx~P��K�4
��g�ŲB�p��' R�'|��'b�Q�b>	�"��
e1G/.S~6h��+YП(�I՟��4Ut�!�O�7M>�dL>L`��e � /��4Z��Cv���'� �����,�\|o�I~&�0J>�s��V���9�Glېr��\;ե�������|�U�������Iџl�5NX� ,P�"�`-a�N�w�����	jyBgv���5,�<����ɟ	r���P�,�H��R��O01�'r�ip�O�
\`�u�M�|>�nK̼����X�a�$X�18?�'k�������4��%ūn��9���� C��p���?9���?��S�'��$Hצ�[���\V�� �*�ۢ�V��4����'6�8�	�����OV}�BC�#v⵨7�73�d��o�O$ oZ�Df.�o{~Y;�^��SX���J�(�����#�\@ACC�}W�D�<y��?���?����?!/���C��	Pn�홤�&xaj���韈Z���O*��O���(�$��~W�Y5&�����)ٺ���a�b�'�ɧ�Op-��i���� Aʉ�^lJ�#񇋎(���	�9�������O���|��fr��a����pY�8٧kD���1����?���?))O�l��C)�P�Iȟ����Cm�1a��j�ygڪ]���?�7R�l�	蟸%��c�b�7T��e�uZ�,?!2����(�z�`Eņ�"�$D��?��e�5N�h�D���0����?9���?Q���?i����Of(j�d�
q���M܍'�������OT�m�f��������1ݴ���yG-��6v�]����:��l5J���yb�|��4oڽ�MC6Y��M��O�9����&�?�pyUH�s�E�P��,A0p�O���|����?����?��dd���I�eJd�	�ř��.�s,OilZ4��4�	����q�S�(co:~v��bI��@8��ܕ���[覵:�4
����Ox�C��А[��AˀoW�ࠪ�C�p�
]A�O"��POf1��4��'6�I �z`�Q% ��0ϛ��R]��蟔��ԟ��i>1�'�6�K�Z���I&@��`p`Z���Љ#�T����d�¦U�?1fR�İ�4cS��sӴ�ɀ�W�H�j	��A�����A#n��6�,?�� "C��i7���ߍe逑W|f��\M�%0�(y���Ɵ���ş��I֟��S'��JF�!#�Z�p��Wb1�?!���?i5�if�T*W��pߴ��0G��;�Ř�H��ĸ(CS�x��'��OV`��u�i�ɘ#0�9�F.�=k9t9I`.�2޶0�V��j��C�S�Vy�O6B�'t�L<f���9B%�A,P����M���'m�4�McuaW3���O8�'>`Z�rT��!��eK� �Q�~��'W6듑?����S���:b��x��� ���s�$(�@�"�bɺ9�H(*�O��?TL<�D_�+w����,Z�<�lIɳ+F$A��D�O���O��<�U�i�B-!�lۉb��@�A�	]@ k���R��'A�6�"�	��D�On��;O�,��J�+�*��v��O(�D�37x6M/?���Y>AB&��+�4�ӬDu\��㊧T٠�fK�y2W���	֟���П��ӟ@�O�(��b)-7��SA��9�Ν���hӜ����<�����'�?a���y�9OѾ0ã��Z�n���-��z�'Nɧ�O-�a"�i*�d�(fhJ�ń0@�������JO󤁦|Zh+�n��Od��|R�(�L#��-s��j��V�BRP����?1��?�(O�ao��5�V��	ğ��I�j�M[��A4)G|�;���_�<�?y!Y�L�Iԟ�'��+�-W3V��I�,�?M��XǦ(?���S�'H1�Όf�'&B�����?�B�-'� *tf�e��8cC@���?���?����?ш���O�U@�� 3���
�c��i�J���I�O�Loچf�t��	�0�ٴ���y�+�n�M	GdA�+� �2)���~r�'
�6Nr��=�&�|��p��B�F�i	w�? �`"���=R!t�Y5�O�K��i5E*�D�<ͧ�?i��?����?9�H��n�xU
�f^����t��9��dΦeR���D�����&?A��;P� �[�!�6���
do��f>��b,O��d�O��O�O���	�kC[�dk�Tt�b��D�"_,6HSZ�܋тӖ[�� {�IVyB��;@\�(��
�-YD�]	 0RL�'���'$�Og前�Mcq�Q��?�6���T�a�U�h5�]������?)R�i)�O d�'6�i��7��]��� R(Xђ FM�W�X���zӴ�7�6�/����>���1����l5x�ȏ7[�,�Iߟ��Iʟ�������L��Jg><Iv�vOv4R�c��o1\5�,O���Lۦ�b4�1�5�i`�'�D8F�%�"�_�y��p�.�D�O�6=�4� �fr�v�vJ�aπ�(rZ� ��]E�\�ŅД��$G��䓗�4�&�D�Ol����a���oB�$��G�J�
���O��PP��$U�w���'W�^>R���n��PSr��6g�q��0?	dV�����8&����0�Cݧ+�p�CF��D�	�,ԉ_V��B�OFI~�O���	���'u$�!�� C�|�9!	Ȅ(L��R�'���'�R���O����M{c�)qM�p��R�|&"	ё�G�G������?��i8�O��'o�7-����˧g��x�\�qß#p�DmZ�MSiJ=�Ms�O��+��Ε��I?-�򎁧ɐ�C�ۖMntP��o�l�'Z2�'�R�'�B�'哟o3��R
�9K ����_J��xܴ_���?����'�?1��y7��>^�C4� \n(3�h��Zs.7˟$�b>I�g����͓[6�THg���
��L��슺CeV�Γvv�q�)�O��sN>a(O��$�OTd�(�FZa�eǤ�qa��O�$�O��$�<i2�i�����'n��'��S����O�V%��EZ�b�"|�5��^Oyb�'��V:��ԚW��ua"@�
*x\\J	�d���9��T����;&�b>=�a�'���	�D뒯�!_�,�S�׸W|Ѕ��������h�IP�O]Rj�-�P�)0
$)���zՋ�����VH 6%�<�w�i��O�΋�H����jKL pA�)۹T��d�Ov�Cצ�YD�[ϦM�'�H�Ԭ��?yb����xWn�{�@��O�H���$�T����'B�'���'�>���O�Pd�gDZ^ɶ\����4�.$����?)����OO���%ʂ�6�m��bZ0rXb�@���>���im��d6��	ȬE̎]�gB�?$�xUA�+��y��iX�lԵ{�d˓^���.s�/�~�	sy�kSx��́�#'���'��U���'R�'^�O��ɿ�M�ш�*�?�dM��TZ��Ve�[�*rfKZ��?�g�i��ODi�'6�7�	�PoZ�wp�����.�T���X�>�BmX�e���}�'I��-S������'����	�iP��B��
305�5��<���?���?����?9���U�~��IK'�����
�	O�;yR�'	�pӘ��d7�������'����,A�`���NC�5��Ɍ�ē�v�~Ө�i 
*N6�x����Fhꆇ�/o��EA0g���7L!lw���c��`y��'���'�"���yS��CU�����#�)N�!�2�'u剴�Mː����?���?�,��99�c
�`�@�!��H�L��D����O���O��O��8X���a��D�5��;�݁2Zv��+	�tĮ8ZC�7?�'K���/��
����O-],��C/�6TZ��P���?)��?Q�Ş��������a)��PB��/v���v��$���̟��4��'����?��%��Ti���r�yA"Q<�?Y�S��q�ڴ��$�/U�i������9	z5V
	E��(���R�b��by��'?��'���'T�S>��F���D�Ppx3JL4~�~`���M�p\
�?���?IO~���r��wl2��♭L ��Q����0L���'�B�|������)��F<OJ�XC&�z��@"�C
+p��2Ofy �JI��?�!���<ͧ�?Q(T�`*Qp����d�/ɝ�?Y���?����$̦�)�ˏ̟��Iߟ(��ǌ��0L#DO�=��9*0��s��m)���L�I]�!T�d8P�Ƅ-�����нxF�Z�Q�CF�N?���|���O��9�e�,�Xĥ�u
6%	�.E=Dռ�����?����?���h����F�-xjA�M�:蒍��DK2Ext�DOŦ��A"��l�ɘ�M���w��ZB�v�<�1+H�b�A�'t��'��6�P3B%�7�2?��[���)Ԓh2)Y���iX������>w�ց�N>�,O�	�O���O��D�OB��	�g6��� IC>��)�<���i�	��'�B�'���y��$<x̸0P�@�s����P���듺?Y��Z����OZ,�z1慠Y���v��,iN�i�ˋ^4b�OԜ��B��?Ć>���<����S���P���d����/���?����?i���?ͧ���T�51��ƟTZ�J.Bx�zs��ҥ�(�$���?�EX�d��՟@��F~��bA5m����@�<�e��ԦU�'\�����?q�}B�;U�PP��#�h��S��.�����?q���?���?a����O�0q�u,G3_��HH��ڳr� x�D�'�r�'P7���)���oM�&�|�n՘^`�ag	N �Ey��ąm�R�O���d��ɞ3^�7m(?Y��Zo�? Z s��*��H��H�-�@q�K1�?A!�+���<ͧ�?����?��կz�ZQ,B(n"
����T��?�����D���VΗ��X�	��ؔO�l܁��V�Y�4�!D� =��4��O ��'��'�ɧ��9gLr����\�aŜ�*��ЬID���d�&���H����ӶH2L�s�Ij)Q���79�<2� ��ThT�Iʟ0������i>Q`+H�8	�'7-ЍI��q1P)I9H�����,� ��j�O��� �=�I`y�OW\˓�M��m�~2�P�$���S�o�ٛ�+a��E0�x�L�Iԟ�KPjX/|���-??�'��%s߄����M`����M��<!/O4���O��D�O����O�'	҂,��9?�hd8E�ŵm3\��"�i��*��'�r�'��y��c��[nJ�"*Z�-��}B2�?z\��IΦe�I>%?�7�����I�<UmF v�3�������S����!�O �I>�(O��Ot��p
Q'Ze�}��@���[7+�ON�d�OV�$�<i׼io�uC��'>"�''�Y�ө,f ��щQf�d�E�dFU}��'��1�d�,<U$�p �_�zz^e��Q9'i�I�J��ӧB��rKlc>����'Nl)�I�Lu��C�@�(5)�1�=���	�0�Iӟ\��v�O������0q�4���F�s����by��)���O`��[���?�;4�]�W���r�!@:w�y��?��c�fʅ7=�����%�:��t��:NF��Q��
8�L!�OB>]��8%�H�����'���'�R�'p�Y$"6z���J�n�r)�T����46�p����?������<�3Ā.H,�XA��*bm��Eo������<��S�'u����ʜ�|�BlR���9Ӷ=˦hW�����')�-z�����|�\�h��K7P��L�o��=]�$k��K������t�I���xyr�1^����O�sA�5a-�Q�AC�� �C�O��ot�N�����MCV�'��&�͞Z�x�W�F�R��H[�aS���M˷�i&�ɆM�nlZC�O��5$?���%�&�˗��w��Q�XM.V���@�	�������	d��JDP��i_~��#W)7������?A����c���D�'QZ6�&�?|! =P�)�(x�0I���x�'����4y���O�����i�	/~DB�[⭎�ueLQʅd�5+�Mڡ�;%��Te�zy�O�b�'�R"��X��=qo�3V��j�
L0R�'�剸�MCl ��?���?!-��4і�
�0��ayv�R��n ���� ��On%mZ0�M���xʟ�չR"MTO�͒s%��m�@4�r�_�u%�E�Ad�,3��i>��$�'r&�|��S	{:���S)$=��������	�\�I̟b>�'՜7M_�q�z��b�Q��s��;k���1t��O�������?�_���۴Y$e	!mҴ
��`9G
�e'�):��i%�7MN&B >7m0?	1�Ŵ����(���]�>�̜�e�@	(�"���_��ybX���������ꟴ�	��OE��0�aEf�$a���9u�JmC�@`Ӷ�(���O��D�O�����dQ��� V|(Q�ȄOJ���!9����I��l�L<�|�c� 8�M;�'P�[h���u�i>l�8�'��I�K��P���|R_���۟(a���{�|�+��OG��P����I�x�I_y�t�*URՇ�O����O�Q e	��E�*�9���Z�f��s+8��9���ۦը�4j�'� ��o@�4�*�`M�cf-y�O�i�Pd�������ڏ�?Y+�O"<�"�UT�P9$�Ҹ\�pCv��O"���OP���O\�}���D�8�!OԺM��չ[�R�N�+���^W����	�p��4���y��*+~�y���e���tD��y�x��umZ�M��:�MK�O��$ɋ)��e�׊~/¥#Tǂ�)1Չ��/�uA�EҦz�)�ɖY����[NO|�ʖ�	�8��qT���;4敁5&�U�� r��+E� e˴�Z��*�� ==}d 37��9R��}��O�q�f[Ҥ���'��	�K����,{�e(_�&���[�h��p��{IN��ꁪt��u�	S���[Vg"K�vx*��\9��0SC�=0|����m� ��U��	A,b �P%A4 q:v��WQ6]��F�+$`���y�p-�����y1S	E`�
4�Ŋ�s{z=S�l
줬�ui�>�
H������':�P���䍂w�А��' [	��ֈ\��M[���?vf�B.�l�<�~j���r���a"�'P�����N���J+�ȟ�������	�?Ŕ'��SP����m�i̊h�7mդ/���޴���k�b�n�S�O��W�ѐ���	�	r48��2��Vʰ6M�O4�$�O����
�O��ĳ|���~Rj_�l0�IIѯW�L�n�{P*�1.Zb�\y�i���'�?���?����!wT`P��[��zp�t����'��A��S��Ӭ�Z��%���5D,��N_�c���R�"ӸYJ�M�'ׂ�b�*H��D�O����O0�]~M�g+/G�p��q���Ҭt�_pI�Q[�̔'~�|��'���I������6->(��T@�h��|�'�'�	�P��O�킕F��|�X@�+īYV�my�4����O�O����O�ic�*����J�Z��i� ^	OOZAh�i�>Y���?�����dD8����O���'� �ң�J�1"T��43��7��OR�Ov���O25�F�Ot-i�Y��+�BªT���:��]�� �Ss�f��d�O4ʓO$n0Q?y�I���	|�B*�|-|�	'�Y?�2�8I<9��?i�j�'>�iT�lơ�������O��]�FS��Bcȳ�M���?���:�_��8� ^}�� ֚Z YV���(l�d�i�B�'��Qː�'k�A�O��'���ȳ&�<[U��6
j��V�	�M;�EH�	��&�'�r�'��m�>	-O�5����� �)r�]o"t�3
���A��
�`����O��wxHy:�FőkP�p�i���j7��O��$�OjD�m}�V��	M?1� ʎy���I��>X����J�"Ơ,?)� W>/��O���'e�p^Y)�IY�I��E
G� H6�Oi�'�Ku}BQ���_�i�MB�L� 5'�􊅭�R���)��>A�f�����?���?�-O�H�A����43���f� c ͊80�ح�'�����<'�D����,�^֤����̂wT�i�.�$�x�h�O2у�>O����O���<�*�'}6�i�� �T JcI�C�1!%�
�($�FT�d��a�	ڟ`�I;V��L�W���@0�	lJ��0��r� �'~��'�2P�X�2h������O����H6�^��GӾy��������	C�I˟�	`�=��.˙mC=��ܱ�FD�խ���ퟔ�'-V%[��~
��?���<g��ɒ)�?.1Px�$�@<K�d�IƘxB�'��Q�P2�ٵ��D�?]����@bD��/P,U�6]k�Jo�B�*�ԭꂹi�R�'��O�6����� y$�鑄	�z�)�#������ at*�N����O$X��5�ҭI��	�F��=GֱjشA�0T��i�2�'���O�&���D��||�@:fg_�?e U��n#(3�$l�Zκ��Id��P��O�� �0���e+��w�>�C���f���o�����Iǟ�Yw)�	���|����~�]��ܘh��Kk^����\��M�����!I�s����|�	�L �"�<h(���5	�gV��4�?tNN�c����$�'��'Ƚ�'�K�_^�%p�'b8���"�$�O�ʓ�?A��?q*O��eق��t��j[(<<5EKR}g@ $�|�����$�x��u'�G:p?00I�f/v��lA��K<�M+����D�O����O�ʓ5_fp�P0�4!)�+bؤKS흗2]<@i�^���Iʟ�%������'O"	��B��`D�9C�\�3�D�{��7�$�O���?��$P
��i�OR@��ҩ-1�LC�9M�q�N��Q�?����U�2�'&}�t#	�${�M�;02�!޴�?)O���ߔ4�<ʧ�?�����1��(x��w�$�h�#��?�<-&�L�	Xy"���O��.������5>�'�O&x�	�8�- ����̟����?��u��ݡD�y�Q�3&D�lm�4%m�f�'�	�kZ"<%>���!ҡnɤ)�U� I	r��k�@��O&�d�O8���2�S��!R���-٥���!54h�`*#]��3B�Fx���[�:�Pt�V�A�Tyʄ(��>�h�l�ğX�	؟|y�$_Myʟ<�' �A"拃D�^� )�'+Ì`�o%�|�O�B�'���?C��H{'�BE�"P�*J�S(�7m�O�X��D�i>��Iџ��'�̔�B�"`���Pw��s3��H��,ʓ�?�(O*���O���<!�V1G�����|M��j�!	��3s�x�'SB�'|�	��H��E�Rб#'��������gT�PoZ��h�'b�'M��P���Sz�	Ŧ��m�,F��a'�ɦ������?1���?)��@_٠�m�1H���ʰr��P�(����Z�H����l�I_y�܏V&��4����p��U"�莔cꅳEgO���I�ؕ'z��'^�8��'���vP a�nv��x1�I�i�%nZßD�'N�ă�p:�S�|�	�?��')~fQ�/M6)��y��d�O����O�i�$�]�1O�S59K�hYRE\?a $BCM��l ���?�D�X��?����?���/O�ɞj��Yb'�sMjMږ][H�F�'J"OF�W$L\��y��J]��D�W�ؐ&�Je��*�6�MۀAبL��V�'X��'k��>�4�V��E�#>���#JnpDQ����Y��I���INy����O�P賎�=u�W�Wfgx�#���1�	���	t-&Ė���$}r�Uw7ܭ����l���თ	ئb��c�'B(��'�?����?a�D0d���5f/gL4б�nܛ��'+��e#�>�.O����<����FdR�]�m����(�L��ǯ��qF�'�������?��Iߟ��'#���$�	�c���ҁ���\��AAP��:O*�����Orʓ�?i���?YF�P�j�l�Eꁜ�^�b�-Ƃs j]��?)���?���?9-O������|� ɏ�.��=�ʙ/h�.��tn���ٕ'�BX��������	 <d��i��
�.ŏ�F@R�gЂ}�;]x�<��T���?I(O�A	`��'�R�A���l ���DI	h,�R��l�R�$�<i��?A��0s�\ϓ�?A�'2֡��@�.+���1�N�r��۴�?���$��?�q�Op��'����ˎL~ ���*w���"��لX����?I���?)�a�h��O��Sj+��ˋEZ�`���)C�j6M�<�v�C����'!�'J����>�;eO>h
Gh��zt�{��&��l�ǟh��}����9�S�` d��i�Lâ|�3�Х~7-Q���`n������d����d�<�!�#/�t)i&���agR�ɃRW�&��yr�'�IW�'�?���Q'v�I��)������)
1<��'|��'mh�H��>�+O�$��� $H�$�u��9�U�V>�a"��i��'K� �U��yʟ�)�O��A�JF�=+f�A�(���A�h*�]m���t3�A�-����<�����Okl�F�d�ᥢƽ2���hW�_�m2�	�z�2���d�	���ɟ��'=��в9F$�x�P�Ӧ~;b5�Q�_�-�&����O���?����?�cf��_�NhK��K�tY�
݃@�U̓��D�O����O˓9�J9H�>��0�L�$Yh6XS�ĳ$~��(��iQ����h�'P2�'�BBƈ�y��3��1
=f<P	�D�X>��2't����?�)O�Q1��QG�t�'�a@m�p����
ݚLS�k�j�ĳ<���?����A̓�?1�'vẶBZ��(����%Dhjٴ�?����d��)��P�O�R�'����t�.�s��Z�X�*&�R�E,꓌?����?�`~"[���&-Ќ����)������B�Zb�lZZy���l6��O����O�IJM}ZwR�0�!l�E��8{�	�Q*��ش�?i�q�|Γ���Oڤa!�P=^<Tt;��Oz���شQ�^Z�i���')2�O�x���D
;X̽)2i�1+�T
&,#'�i�m��'�2[������Qo�l[��T�;e
񈠇�0E<53�i~b�'"l�5f�XO �d�O�Ʌ#��l��Ĉ�rD���">nd7�=��ߘt
�?�I����	�6�k���N��ڧI�S��7��On�3e*IV�	؟X�	V�i�E#����`dT-��m��)�Aͨ>)Bi^��?�/Ot���O���<� �îK��0��֖+K�%��A7C��z�xb�'S�|r�'RbkQ)���+&j�-X.���l��;��Q�'��	���I韄�'�\���i>�+ �Տ9b��Ap��"��%b%f�>9��?�N>1���?3!�<�ԪΔeM����a�-i8Fbqmۿ2��I̟��	Ο��'���c'�IY@U����l�e �H�hЕ!�(�n���&�T��럖�e��0}�� 'lj߀G�D<�����<��f�'��X�PAc� ���'�?��'�5%]�V��Xȴde���Q�x��'�R�X'< �|���a�q������S�?>�u� �i0�	���شB���@�S��I2)��)# �R�HaFJ����6�'�W��yғ|�����S+�Z�L��u��	�q��/�M{�f̀:ț��'C��''��h9��Sd�q�F^��jb�΂�5����4f��ϓ�䓣�Oe����:kl�i� p*��r5�S�{��6�O����OvL	g�_��ʟh��C?��
[S蜓b�H�k9`Ő���]�tK �9J>���?���l����N��&�a�
��1���?���
�<�A���OT�Okl�"S����N�yt�Q��`��I�-�����Ty�'R�'R�'m撌��^�&k���CbM(E�
���'0��|��'1�Z`��d�pAL�Z$�X�0�31k^U2��'�I��h����T�'�l 3�u>��5�T�<��tU/ܐ-��B��0��Or�O����O�,�g=O�	�^g� ��G-J~T`�R}��'B�'��Ir�Y�M|bB$�H��="�ΰj��+��ۑB���'u�'��'����'c�O����F�[Q�2p+I0N�:�nZ�d�Ity2��4Jfv���d��<�2�k�"6�������e�xE��B`�I����I�[!6�IQ��Bڳ�B�^ARԋa�Ltaڱc��Q�'�=��bs���O(�O�0�dR���@ԜPߞdr��U8���oޟ��I	Z¹��W�S�']8\X��fA�)�8*RMʹ4C��nZ�/+؈2�4�?Y���?I�'-��'j��Zf��|��F\)����"Z�[�7���,��6��0����\Z�+�,x��QJ�?ݢ@���M���?���Vq���d�O��	4vV-!��[�`�����fQ$6-*�d�u�H$>���˟���GR�y1��50��0�n�j��4Cش�?q���X�'j��'%ɧ5& نQ��Y��Z�犍RV%������$��Ĵ<i��?�����d :Y�x�vg��~��q�s�.B"�Q��WW���@E{�'ώ�x���2X Rh:A�'K��D9���qGP�������I@y2�̫c2����1�L�YI3�">���?��$�O�� �e�O�1b��-�1 L
�W�N�+�e�N}b�'L�'��ɚ����H|�E+\2<:X0j�&�V��q�,�9���	ΟL�wm柤�O�(��J�>�mR
�-^P�`�i��'���'���X�'|��'�2�O��]"q�.J�b�y��h�^miw�9�D�O.��Q�UvPA+��T?}���G��jIA6��>Nz��.e�ʓ T��i���'���O{z��{�K\�)��YmZ����Kr�[@���?y�g�	 �� �TC�H V��A��>�7M�>n�B���O:�d�O��i�Oz�$�|�$��0L0-�%��.$8���3&��*�oD�I(�y����O0�́;eN2ѩ�Z�]�@�V���e�I�\�	�[�� �O2˓�?��':x�8���}m�@�[�r��}��SG��?���?�q� �r3Vp�S�H�i�"I`�"�F�'��-`�³>a*O���<i������ �A��@+[^�ᥪ]}2�.�y��'���'b"�'��	�����3d�FcbI�r��jĂ�7���<y�����O����O��� �D��w�|1�^4)�h�FJ_�<i/O����O����<e =��I�8�6]�eVUr`��t�VR�,�	iyB�'���'Chi����pb1×1_~�3F�O'R�2��4V��I����	gy�`��u.n�'�?i1��+�)�7C_N0�+�@Y�&I���'��	ɟ0�	ڟd�cf����S?q���'"!��3�	^�?����Zئ��	�ė']$��~����?i��c�T�;�dM�Wo���e��l���"Z�������?$�Ik��'X�I^�
t��ϗ�e�"�祟�~y��S�x��X��M+���?������U��ݙxe�eZ!�j)�u�+}".T6�id2�'Luӟ'����<���4��*�>�"L���S�%<�Mka���b�F�'��'��ԃ�>	/O8U!)�."��xy��B������㦕
3�r�@��py"���O���+\�\]�i�1GO�$T$`j�fۦ���������u@ܬ{�O�˓�?��'�(�X�m�/���F ��hպ�4�?�-O���<O�S7n�����ٰ ��hɄ̒*$��Qc��Jy���Ʀ���y�dџ\�-ÆJ=H�f${Gcѿ�p=UO����d�B�Crn�(�J�c]Rx(��ɔ@Yڣ"��x�܈����(l��y���7>�ihWH�wu���-E�9� $��L�تfG��r�zz��Ń��pB����5;�F��F��S( ����
����U�ȂT'L}���\�B' PY��(s���iU��"+$=�� [ޟ���	>c�����ḑR��a�ɸE����V�d�bX�a�� s���$���O�Q+(�:]�� @�AG;wz��H��'�p�����?	+ON�Q�ה1<���/۱w��{�2Oz�D�O��"|Rdb m�D��Ɵ��If!^~<���i���Pk�x���
[�
 ��' �	4u�:*�Ob��|J��7�?Q�$ c�F}�ՄW>s��Ś�'Q5�?1��T�5z�OV�~Ra��>�O���Z<� E*�(,��c�*�h4l�'|�h�4�X�k�(�Kg'�~q�H&b�Jd�
��V�Zp���O���e�'������pъ������$A`pM;�E?D�����[�vI�"�_�'[b�0e8O%Ez���E� <��J\:�%PE�ʏ|/~��?���M�@=+&"�"�?9��?Y�Ӽۢ+ް�prS�\j<x3n��ܢ9�Ө' ��@��ʌҊ�L>���>M��т�'�3]`��:�n��?�@��w�-�1G����}&�P��aɝi_���'V�5V-����ɟ�'4l�b��|�����3[X.4!�F��N@uB���*�!�D�+�vT;��H�1܊jB�
 ��I.�HO��dy�+ީz7p}�TV��*��ǈ7��A���9H[B�'N�'5r��՟����|��k��vhBԉ�ljP���*`���c%H���>�
?��K�	[3R��8�0K��k��Մ�E�^���E�E����1�E���
�̞�:R�����'B�'�bU�l��f��A'�9�P.�@���k�ȳ^��x���"e2W3�B1��%���<��R���'*Y�$��>���s�Ru� z�`�C픭H�RD��?��Y��?�����h��m�H�� ��?y���sָig %:��XM����,%T�-��J6��-	 $8�4@G.7�o�685bh;�o<^TL=�'O�����}���'b��M�>���@�gz�!-g�c���	Ix���@|;|h	�.ћY�L�r�' ����4z&҈����G�v�y�Dȉ)�����dB?@e��nZ��l��q�4��|��L�	��!�5&"y��싫w��'��z�d�0�1O�3?ᄡҪJ��S�m�8�B�[�,�w�d��(�1�{����C'}���"[�<ɂYI�G��I�	y4�D�Of�����F����Έ�)A^�//��z2��O���D,i���R�Q)a�3c�kax�j7�ZyF	s�]*	�dIp�	Mh0	���i���'A�Y�}�U6�'X��'��w���K�U*Z�n塃��/��h���'�DR��7�|��M������I�-j�x3h�G�b�O�ma`n����,�X�@d@�)X��Ѐm�2����?���* �S�gy2�'�̅{�c��B��[ ��~�8�O�ba�Θ3� Y���ڋ/G<{S���I������<�Q�K�p�jB3dAp�S�<�"��
'����ȆT�ݸ�ΆK�<Q)^"x$��XD/S�'�T���Yo�<Yd%�>-Y,Hق�_�=<fĂ$�_T�<9�R�X��1;f���`Tl����O�<�Y������TQJ�+�͐bDB�	 +��	K�j�6/�F��ի1J&B�:"T�R�h�.<04,?\|�C�)� �燁(:i���ݙ,��lQ�"O����X�,/L)@�)-Sy�Ԓ�"Oj��B�{u2�9R*QkR~�#S"Ov�X���A@��iSM�T
v"O~5{¨o*������ .NM��"OxXy0o݋9�t���nǜt9�"Oik$��$e�"Y��#}��(�"O�{��T2a �/HB���0"O,mX!a�2,��[E���Q�n��1"Oj5�bc�2
�bE�D
~l9��"O|-1��^�I��|AK��Z`n$��"O�����v�Q�d��Ze���p"O`D�F��
y�SSB�+c��(�2"Ofaz�i��SB��⧈9�։bq"O�h�Ⓐ 7�ՂT'�I	��Y'"O"8 3C�)@<�X�=�,<P�"O Ak�	ͱT!���f��v�@�"OС�s`��bR��0Bnѽ_�n5Ȥ"OH�8�!8/��):q,�?Q�(�P�"O`pYe!ݓq�	��b�"OԔ،X��� �U�g���A"O��)J-e�����V�tU8xچ"O\x�#-�!O�,\���N�d�qf"O�L9TH�z�,����J t�"J�"O�l6D�(�`��(pZ�"O�<�a���i��ٲLjx0�"OB`Q'��<Ml(� P�E�FP�Ѡ"Oj}z��4U�&��E�S<�j�"O�|�!@\M�d�c��ܶ_ Ը!�"O�,���S�@fe���^�zܑ��"O�b��H�#|��ū8	]s�"Ot�25j�r5"$`�;8	 �җ"Ol��&z��!����0�%�&"O��Hq���g}� dK�Lc�r�"O�Q�� ��P�
�s�@BH�X�"O� #�i�����?9`���s"O��9��	�]��m<���"O��p"�:a�"=�?C5���&"O0rq��r�^Dr�G�,mn�b�"O�1�2NOS> J�̏E6���"O�����>���v�U�T�йZ�"O�Q����y�dݢD�ď��i��"Od�#�H�yrTq�V
|ða��"O��f
��m��V�Y�y�>M(f�'��9�VA8�O�\�oV=2�j�B��H���MSG�'3���@*�<��$�R�Y��}�(��q�T�<�r��[�:ՃكM�DT[�ij��n*� 5��8�@�����m��"����i�C�	70�Lа�,R)0B��ǅS�T+QCC�O��h����.������ļq����w�J�6h!�$S3rK��q�-�F颡� O32������Ϝ[8��	��6d"�XD@L�{�&��A��s��A��6^:��1����&І���-i�L5�9k�6D���Fx�V\*�#0$�a�e�u�ڌA?�%�am]e�<��A�d��M2�iT�z*`,�V��b�<��m��F��HN̏=�� !0��_�<��;���u��$h�����W�<��͙	N���$�1+��HG!�S�<��4���D;^�"�8�ϜG�<11���'�p�6�ڛ*�xE�!F@o�<���B=
�]$ac��tB%�i�<�qo��E�=�E�IfZ���Fh�<ё"؈_���+���b�zm�1Wy�<� ����Y�-� �1Z�Rk�"O.$�>E��Rv��)3����"O�;e�ƱV��쀆F�
i�����I�W�~<G�4⏯Z�Xe�pΑ*RD	���y����(����e�1�"�bQ�'�~2e�+�O�>%�5 ۝x�k�D�0H �$D��@�AI�RA��*�E��B�H��7}Ҍ� -�a{B�B4S%�4C�v"��wK��p?�R��M�B�ɰ3B�ł��ۀ7&�����i�<��
Z4p��8�I�0�[�?�Qز����ԭ<y\�[�I(jֆ B���s!��χM�"1XuG�O��Y�˙r�!�D�^��%�Z/�6ԩe��	R|!��I�B(����q��A��40c!�D#����0� RA�ظ���)"`!��b�N���!Į&�֔�'ǱT`!�$2� ���\0whdX�&� ;�!�S+x@p�"��$s��� ��1
�!�� Jר�3?�P�Q��,�!�$�Z_�p��̊Bt����Ʒ�!��[�2����I��&�WOC��O�ԑ
�T{��	1��N���與�Ix≐x��	��̊ 5���2��;���rQ�`(<����9I"�4�$�uƺ$r3EF�#���'��5� +�����҅��	�$��fL�B"B䉩c謍�3�΋O�A:#�̜HZ4�8���?��� �s�A�F�����p�Ap�ۂUk�u!g�\�X!� �Cl%����>�4X�6��ZP �	�v L�{��J�A4�l�[�l$GzZgd���\�`�@�Fϣ9�l��$�#A�V�A����� P"�E����;�d)��0aZuHDj��F���ڄJ��͏i-��P���s� $��R���3L �U�]�T�����J	Jy�O]V�k�� 0֊�À-O�UX����'�h��� ֖Ol�)����.�2���
�`l��N�\l�a�,O1�2���gxލ��	�wm:����'fȱbf.$4�<K�M
=����$뎄7O�ܱԯ�O~�A�=I�ջg�O�_I�hC�o��O��2V����|�+��ORܦ̘U�'|�)��_&\�͚QI^#��	�n�;�^��e��-kr���ŀ� Ahк��+v�����2�n�qҊ�#Zi։� Hw��'�ֈ�@(7~��)��V9g-=�I<��&�𳒨T�t���@��P��C�	�`w6���%<((�)%�.r�7�ބ:�� {Š�Af�A�m���T����=Z�G瀧E�P��"O��ق�.2�X�[%(X�MD�d��mH�� Í�
���@H�0��9.$�Od)���ܖ:�$pz  Ѥ6n8%yW�'��Qv��aT��o ͖u� �<m�f��RI�:pv�dI�O�����ɎL�b��c�!?đ��(��"\Dz�C�y�FQ���ݟ�b��ެ��nO���ӄ.�o��i�M
<4b(u	˓G��	��N�48��Q���O��׆�'���#v�M�t�q��'eXY�A�K>f����0w����_��!r�]�4}���v�\m�(�D]�R�֮#"��H<� �č�.E��I��-��ъX@��$�*዇$y�Ē$�(�b �QGR�R>xh�gBQꚠ�D"����K�^��8��c��p�Pٰ�A���ԉ�蛞{F�c �-k��O���� ��g�MJ�HQJ�~�!�Sh��Pæt����4U!�����p=��_��lY�m�g�ܽ-?�f��*�i�0�И]n�Z3e�\��qK?�@1nۖ� ��΂s���B�8?@��dS�Egn\���E0������"2+�iP5c��t�� u�^5"���&t��΀-?8R��E�?�)�a@^���p�ij�Sc�D���߾>��(�*͐O:IcU&E�a��e���������(�e��-2|�6KB�FhP�j�ߪҸ'��>�	693�%�#9� ��±	��a�7KN2[�"�х ����ĂґI>��$h|�18�#�*g������3��	����pB�'��xR�͘�=�l�b�)�)��� R$*�ɴ-}d+̓2-F|�Cc��Q峟 *%�W
y�����L+#N���7,O�B���Ɯ1`!B%����˔#��=R��QY��k���;>L�3��U������6[���3�I{��fF���ɆEOsd���0� ���3䖅�4��A�f�8$�M�,���=�Ɔ�K��T��@G2$��T���XŦ�Xf��|ܓ/�>��2�	#5��:�rp��\,| Z�c�M�W& W������(r?�S�g�? �Qv�@�O0��jQ�� ��v;O�����p>�PD��Z�3�˂�Mu� ʤ���O�ĉJ���_�IU��Q�O�tXr,�T�]�d�j؁��I)�"xAqfɳm� ����	�$�Sk<4�����%��|�lG�YcbIº�x\��ط<A���q�xД'���>K��x1rf>f:)�s���d����4o�����\�.���J΢,��D�x@��3$*�4u��I�$��I<ЋKI�I�dE�%8�@��7��.�b(�3N�'r�N0���S7z�.扲{c| ��k�>t����PKbc�T���p�Ac!lJ%pt���KT�l����� VB�ESO�X8Dt��"0Ҷ��@ׯdjM�ҥ���) 'e�[�tO��J�$r����׆$��w|�La��\@p.�y 	,A&(i�O����n#K��i���H�����D��:1�X�m+M2KP�(�p��F��j}�'t�RD"�_j�ֈ#�J�l�@�wh��[��EhEÑҴ8���>�(u��p�F�H-h9p�J�6'���{��	�p�K+�l�rp�R9p�p��+�X `ώ�cVJ�����~�Y��)�e��&� �($��rR,d�e��c���̓R�҈(#�R�f�l2r�O�fA ��'��0���	� N����p�B�n����3Y��;��X/w��`���&|O�):�_.xP�Q"bިq�)����#	�������BK�/P�H�#�f�P($>�N�u1�9�E��{e��I���
TE��Ը�|��E�5[تM �!�/v�&�����Q�d]����4P�"�����N?�`Sc���l�����fG�Y��K@�&#�]@S&�p<)��-%��O���ҟd��$J�n���b��g��H��F�T.� 3��G|	��¯Yn%�?�r��&\�p� c�qӰ��%�Dq�D��A9�y"I�.Yb�`z�G�������8�5��۫~T�Y a���WOʰ���M�}༼�C�'�J4򮖶XH��CN�)X� �yBF�EР1b��\�@/jh9��D;��4�$����]�)�2M��&�'󮈉0O0��ªT�c��X3�Nu-ֽ��Y
k$Zd�<��I*+�Z�>1T+<<y�,ʐ%I�/yp�V,Cj�<qw&�
~�4�#��]E��+g�[(w����'Dr��BB2k�n� A�Ԓ<�Fu��'�<Y�����.��J�0]�p���'��mq6�	H�d=�h��Sqb�I	�'޲�YrfE�[����ܲP�r���'ܞ<H�j]� Y����
CHRQ��'����щ��ff#Zd��'M&�"F�L�+H~<��B�n���9�'�0���/�~99��o�މ��'��t��b]+/���B��0W8Pq3
�'�(�`�D^n��k@�ش?_�<*
�'D������i�BՉ�� �.�|{�'M�d�mЂp3S͒p"���'^R�#G��%�f0m�+��'���P$G��fH� G(E������'L���J�h�sdB� /.�A�'�I	����t���Ə�.]\���'��j���h�`�`��o^h4)�'�b��aFL�H�KƋ�6mZ��+�'
�(�f�`C��S����z-�*�'��h0f��:4�1��8%kZ���'�ʌ�u��=����V�Q�$<��
�'!r����͆?R1�5`D�l@�S�'zZ�9 ��-M�ޠ�����D��'�J���-����u�3 �Ih�'p�FKQ�w�K�'�ԙ�ԣLd�<����$�+f "t���4�`�<����#R�Af�A�4�!`bR_�<у+םŜ�#��6�"E��#�W�<��%C3H�8��`IV����'�]K�<9!���:��A��q�s�C�<AB��#M��P�.p��W�	k�<9Q	~N���fh��7�RT�v�}�<ҫ�|,�D�^����z�<�3
�i_�7��������=�y���3HA����̓�©r��ydҔT�Dqs��@1 ms����y�ɓ�cf@�����8�ZQb��_-�y
� ����OX�Z��h�C�]nD�"O��8�c�?q���˵�W�lqY"O><�#��R�@����S�ؤ��"O���V![��y�j	�v�n	Ȗ"O�(��04S�L�*��_8왉3"O�}9$�K�=㞰C"):��bU"Oj�f��
�`5���U�!1�t��"O�LYe�%&$Pr�_�B)��"O|�@Ӊ��7{�T��*X
cޥj"O�3��%tքu��L_6^� q�"O���C��)�t�kq��#
4�P��"O����$O�M����3�ʠ[�u;�"OL��Ӏ�7E�Bqju ۼ�*�[�"O�-
G`PR��(��,p��A"O���#j��S|@t�ٶZTE`r"O&��ER�� qd�ŽtG�s�"O���KG)M@fAQT�M
��!+$"O,�+��Q�����D��asz��V"OX�ńW!9N�kE� �mU��p�"O�2��@���a�"B;Hi�w"On�ԥ�}��t��;H/��	�"O��թa2�͚p��;=2�"O�,���-|H=�@.ɀ|a��1�"O�0B�DM�p����,�� �6�)�"OB�I��`R>$��CC�8���"O����P1�FD��i�02y��0"O�q �R#O���F�_;nC��z�"O�aAG(��0�a �Y�مĈ�!�D Ht�mH��� ��D�b�!�d�K� �m!H�tiHr�ǯ<�!� �`���Ҿ|�K	}&

�'{4]��O�2�2��A�x�k�{"�)�) *Ľ�d���n�M2�ժ/!�$FS���@KX�a�O@�&p!�$�72�尕f�3�*�s�.?�!�W)y�,�fђ/��Iʳ�Ý
�!���<����P���=�0�H(!�$�4+:�p)��^�[�ɲ��%�!�䘳g#���G��hid1�UD�!��R�u�� �AѬnKpQ���G�!�>��HUNǄr���P�L}�!�d֬4&4��aO�s�*��1BB5r�!�
�m�Pm��ްG���r��/u�!�dM b{���HW��*��ua 
6�!�$V�i�6D�+44~�G��T!���ej��cg��s,L� RU	!��B
 t�Cfb�#O.P���)�!��E����Iۋ��A�K�Rx!�dZ�(	^`�5"�	:pJ	�R�ns!�V�sI�	�R�_���Q@�\�!�dش?o�!�uc8AJ����s�!�S�x�6Q8R�a� �!��N"c�@�4�E.�P��㎺5�!�$�z�$ ������%b��"N!�ī��j#��a# k� F!�D�s�0� c�+s�>p�*8D�!�dQ�T�
T�g.)��Q
7/ċu�!��jFJ��b=r����soˮ]!�$ʗ=����4�%h�x�Ig�]�d�!�$]#"=�j���|��H�f.�;t�!�E�93DAD��+�dp�Vo�4�!��V{��E2LG�]���r�!�$�,��)`�
+v�jVM3�!��ȼl9r�R a��+j���A͠8�!�� :���M�^\�����<��xD"O� �!��[�EcV���W��;P"O��H������ȷ!_2�,Yy�"O
 �W��R�d����]��<p"O� ���Ň'�ĵ���;1��h��"ONa�`��� %��Γ�0� �"Oh�	9����͒�
)�V"Ov؂�Xq(��Y*�*�ZDh3"Oy��ȏ%
h�y2u��y��"O�U�'BG�v���a.ܽT�x�҅"O�$�7�B.X�ZSM ?~��P�Q"OBX��#�i����
�.��á"OIr�\6'<� �!� &xҜSG"O:3*ˑ{R^yQ��
_ �c�"O���E�Q�;9T�{EF�D��b�"O��A�������,�ر;�"O��j�)���0ؙ&��G�0���"O��j�AL�KB�]��fQ�m�f}�S"O.u�5�˜u\ %`�#Z����Q"O�Mۇ��9kƪ(�VŒ9|4 0�"O�<��O�d�(�k� ӥJ��a�"Ol�j����:M���_?u^��"O֬� œ�("�c������b"O��˗��K_�`�¦Af}�"Or��i9���I�P)�"O�	�����$��	B*_��(��"O��kE�,�9���E��90v"OZ���8Z:����ܖqm�@;�"OP9�ƀ��$��pӂ�P?]�'1Oܹ�Uɚo�z��b�J�5�zLc�"O-k]	�D[���� � @�Qo�<���o5���kR�3���c�RD�<��LH2�f=R�=I�{� �|�<i�]+]��т�P��s�PA�<�N��g�f�K -	5d�����Ts�<�%���1��)���ԭj��$H�b�n�<���խQ
���j\�v��h�<�ҁBI�i���t��4� �Og�<�v��
JM$�1�6E�⴨Lj�<!t!�YJu�c��/:�@��rI�c�<�ǚ3�������+���weM��y�,C����C�0�C!��L��!�'���p���Q�D)�l��9��
�'��x�N�
&
�"aM3�ܽa
�'��p�\la"�S5�Q�<K�:	�'�"�PR�
�5{J��w�<<�)��'���z���dЀS �W�aBj]:�'��ZS��K
8�i"eҠ1�E"�'E���Uj!b�d���W�
0��'ؒ@���N@	��$D�5�'`�d�.�ds�%����H�
�'�pK���$pr�l)� 
�Ȍ��'�`	�e��v�IѠ�Y[j��P�'��0� �E�a1��B�&ݓ�'>�i�i�+a�-Q��1��c�'���� �PAAu���!)��p�'�����F�����c>��L8	�'2��%�MI䤭����@�a��ONA*g��9�)����)����I����xe��E1JXQ��ɞ�3ux)��"O���)0븴a�)Ćig�"O� ���������H�
�r��"O(P`�T�M������7�Z�hg"OF� R�@�q��m7�5!�l��"O� ���/%��"�ӧiu�0�"O4���a�#+��t� N�d$M�w"O��3GB�Y�h@��K;L�A�"OL��#���$���Z6�ϙ#/�S`�w�O�ک���Nq@$4���b�͓�'エ��DY�,X��R�eR)Yش���'D`4[�hޖ81l4F��a�IB�'4�M��<r���
��M��(��d=<O�Q[�Q��0d�C�U���tK`"OF���[���4Dx����6"O��)���V5@�اC�2�r ��"OxA�bɁ�.�q	U�w�Xq��"Ox5t.ۀoE�PS�҂3��;�"O~D�Sj�v���Qf� T�X��A"O.�q��Ωh&�t1�!J.g��;�"O�̱�B�aT�a���vi��!�"O���F�/*�&��'E?EQę�s"O�u�Cě�%�j��!�)���"O|��iЂ;��A��R�^!�%��"O6M����9��h��N�C�T�@"Oܐ�W�4%�����R�MVx3�"O(xhp�8R�ޔR%cڷH�,�"O�I;�6M�FTC��+^!��"O�<�� P'hn� 8r�T�L�,��"O���!�.u׺k����8(�"Ot�	"O�=:�I�NB3E�)��"O E��K�X�����зd�XW"O֠�q�=�H�Qp�1U00���"Oh�I*m�-b���q�"Op�y�%Tv���_�Eg�0�"O,B@@�>x��a�� [8��A"O�xHԡ�y��	!͕&i� �C""O���JYW��ݻF�:׊<�T"Ox)9�f��z��Ig$J�h2�i�"O�H���E
D��Z���5tS�<�g"O<�����bߚMЗ��`.��"O��1��¦
 ��`��A�ٰS"O8����
I� �@�J6o!�j"Ot}�c�"�� Dٵo#$pjP"OP��Q��.]`�e��Us��+e"O�8�J22����_)s���d"Od��ɗ+l�4���ɀw��a"O�y��/�*x���
C��h^̰�"O�I���̫I�@�JsHL0i�"O��!��� �s�(yJL`#"O�A�5.g$ͫb/Əc7���1"O0��5 ҵOQa0f��&FT�t"O���B�� �a��m
&s
,�"O�� 'i�Epʙ�W�d����"O�����	�Z��GG���%AB"O�('R�B�2�Θy��1"Ob���j�?kzB0�]�B��U��"O���1�H� ^�q*��I�q@�"O�h��m�1n�L��gM�:.�\��"O,�@Q'@�n{*�S�B^�4IYf"O���G�[ 01P�i���'�(y�"OԽ�B΁u�H%���W�&��"O8|c�B�;qt����bW�h�\]�"O,�넢�X|x(w��*O �!r"Ox�Ӂ�
�~�\��KF(~�d��"O�M7H��.x�|IK� g`��p"O���geN�8�0}2FI����B�"OE�Ї�5SrыPg˘?�4��"O��F�W����(�:y�"O� 00x��D�Y�p���o���"O��� 1�B��D	���8��"O�0��7m���[��K�w�L-�"O\ɑ! 7c�P �(Ȥڠ�§"Od���fՕZhm��;[�(rf"O�L*ĉ�!Ar�+���2>˦4C�"O�bd�Y�X�*�˦!EW4�5"O�!���/yj����,E�|;"OR,@�%� 򎨈ǯ�-(4��kF"OL! ����Y����$�>6%�`��"O(`C!�j��yBP�ʤK�"O���O�X�g��`e���b"O򩢠e:/X-���;e(HD�"OJԫE�և[ː��tjW�n�@dc!"OX�����&��4$��5�P��d"O���A:4��Q&U��k2"O,��� ��jt�viW DU��"ODpU@�8O�	h�'��4��V"OjM�'�}��s���^�b�"O.T�Wŗ3f|���r����&��"O<i� �Q���d��,@�J�H�"O����>����3�ݎ+�Ҕ�"OX�"A���3�V�sD��e�,���"O�y
td\�!Ҁ��s�U�2��a9�"O�K�#ΟKs+����J=ZA"OP8p�H��B�s����j��܁�"Oh�(�c˫'ʐ�;�/ǼL����"ONq�T��.+=h,�2����x� "O��p@�mSx�+��k����"O8�
D�%aa�0� �I�pU��"ORQsU��O5�H�ot���"O��wi��v>fhDއ/�"�#�"O|!c���ug�9�Vc#S���Q"O�KEǈ?�\�g�P�����"O.P��i�
Uy�)��.5�D�ʔ"O`ݡ��-CP�e�^�t��F"O* k� �1�<k��I�s|��b"O����+��`A�����R�]��r�"O2	ȃ�T<
�L�f��.\����6"O�aQ����dP�&b��P͌��B"O`��'�S�%)x���@˶�����"Ott���2�H�v��:���:G"OԐ*�a���pH}�����"O�0`�����XM'��*�&�"a"O����Ns��eJ���0�"O(,Q ���zg��M�>T�T���'��T��eg,|C�
�5��)�'�H��'M}\Ĉ�`� S�'IN��, 8U���3N��h��'�<��0��:Y�h ��{�H9��'��\s�H�^���J�Gވo���'���3�̙�`B���� ;}�&=�'�8��f��P��b#]X�г�'�v]�@Ɣ�9[�C� 
B��e��'b9�uF�^��#��ʺ3�|D��'8�t1�58Y�	T>NL�*�'=���$J"9Ne�:�m@�'8Pd�'���ޙ�o.��X�	�'�J-�G�9Uk&�P���	Tr���'yLx����d!X(�t��O�����'3p5�4# \o�*E\����)�''��S��P�Of:��X$:�t���'0�D�5!���0D�(4��#�'����B��eMFh�ƈ0������ �i9�R6s�(y�� �!XH9�B"O��x��<"�$pe%Ԏ-g�<�#"O�q2aC��l���+��L�8S|`��"O:�!�]�O��� �˃#Y�Ԁ"O.5zqԗ�j�y��ِSK��z"O�� �_��-��)�
H� u"O,����	}7��3/W�>�6�B"O��N��8)��kB��DF���"ObW?2_�` A�J�4��G�z�<	�n����'��;5�)��Xr�<��^w���B呐a\���Fd�u�<i6L�?Eh�ͰR�T�Jy��x�<d�40�H�^#cԍ˔�s�<��M�1u� ��Lo;���*p�<��
	�rq�+}$�p�3,�h�<aǂ�>�x]���Y�=���U�M�<�� ��:������>ro�P���m�<��ȓ$K�\XD�͔b����P@�^�<I����`��"̔�� F�@�<�DΛ�|��Q�ČV�H7�!h
@�<�%.�@���@�]�1Pv�*U�z�<����+�>���0n!��)�s�<����(X�*m� ZWF���,�x�<�Ъ6n8v��'eֵ1̬!!3g^�<�E�bzm�%�q���X��Y[�<����r{",�@�I*$��(c���X�<����S�T9�@c��j_J��Q�<���E��f9 �Z�]wL��S�M�<1%̀�A�� 2Ꟊu=䤚�CWF�<��F��SA��j��B�0gv@�A�<1���J}��Y��?V���I�{�<�J�98\�XE��/<jЄ+���t�<��l��
�,0sF$@.O��!;� n�<1��],pʤp�(�x�B��s.h�<Y��X�� B�ɉ�A޲�ӪN�<��� fF:tZr��2Qp�"0��c�<��+�)5��C�ȲQ��e�Bd[�<$]�W���{�eI.:e�Q���Z�<�b��8C�0�kC��(,*�٣�*_�<9`㜩��b��T?�cE��|�<!�#��2#��)�`��т� QC^R�<�' P�h؉$�K���,`Re�Q�<�h�Qffس%Bߢ�VPy�N�<�"�[�2��Vc�mx��d�K�<I�M�"6�h��s#ҁF�:HGI�<Q�Mg>s�N��1
�/�D�<�r-�\1�!��Kр[ ��Cv�FE�<q�@�9i�$B��d�C�n!�d[+b��������U��b�B$!�J�&Y�� �)1�v!���Q�b!�M�v��I��)PIn� ����
!�D��/��T��N�2AT�: !�ē�cF��gKN[�������[�!�Ă
{6��Ha
��qxp1(��B_!�dվs<Vܫ2L+(T�ȓ��Էe!�dR
*� �����rhX#��-	p!�d))W.-�3`�6r� ���(��kt!�d�`�6MÁ�]��QJ{!�DV-,�8qs#.�Kwx�����N]!�:G���Ae�@fA��BQ2y�!�Dι.S�X����G&��(�ԘF!�D���ܙ2�$��?���[�@� 3I!�dޠ_m��!�8Y��E��T�e�!��B@.`�KC=�� C�oJ �!�� ��(�E�&LH<K�苗u?���"O�A�3B�f�|q��L)_�����"O(,�V�3�5����+�N�8"O\��!��J��8�ǂ�K�&�X�"O�YB��)U�� r�h�Sg"O@�1�����ٻS&�i�<�I�"O���#K�-@���䔒f��U"Ov�y��������,_� ���	h��AE��
s��i抠Y\HPgB2D��Z��Q'"��c�G�5\� �-D�X%kF��
��D8f0���0D�@���,�Z�A.D8k��-�7�0D��i@�[�z��ZăĚy�^Q{Rb3D��1��Hj@��B(Ƞ1,>�K'�>|O�b�h�VD��+ܮ=a��E�U:�vd2D�8+��S"���2�ȫaN14�@�դ�$�!3S�*mj�i���V�<р�Ǒ�> �!Û%e��Aa���@���?a
Ó$�)YF�V�Z���$Ǥ9���ȓJ�ʈ蓬_ĖVI�jOn�>,�ȓV��cD?7��k�a�)ș��	����<��D�	N����/
�W�v�q*�R�<9�%�7��B�a���ڼ����t�<y�@��	&i"�B˚w�TBL�<Q�Ô�_��Daq��iz��{Ј�D��0=)&�B�����s��*�4�Z��u�<�+�)n�H4� �Q9֬�g��E�<9���ܾ����9vh��u�L�<��KZ�g?�Ir��E�~H��_I�<)��I�e����  ��Z%��F�<1a#� �����b-2�2��RF�<&�W�m�H�s4�X�a�z�!EJ�m�<��� Q&��'VI��%���s�<���M�hh[�d[��&U:Q+Ti�<)B�ɏd�L|
�h�
?���!��N�<Q��l�(���2��E��kDG�<�".��r`q�w��*h�(8��@�<��%�
�0��)��\�A��	@�<�A�0:b�Y�eɋ)W�Z����U�<�U�<UaL�"d�H������*�|�<9Rl�JL�����`�� 1�O�<��Dp�':6#���.G�<��G#/�dP6�N>a:a�s�E�<!���E�|�Ⅱ�7g���hG�[~�<��O5V�R���ּj�b�pB�o�<I�ᐒI�\�#�I9mb�Hxf��P�'wa���[f�N�ХAQi�JԈ�']3�yb��l�F���Ë�[� 0��.�y�Ǒ�?S>�V�W0X���۷�׮��O��d?�'>��3����/�p��,��ȓE�����r�@:���w4-&�h�'�ў�%.Xҙ�#�T8`��1�T���r�0C�Ɋ:W����Q{ohd����q��C�I�Qd���� &4ĺ0�J�{�C��,6���(CK�
W(��g̛}�B��NY��Sjҍ&"�YG"�A�v�?i����8,߂}`v�ړl�:��7G��bO� ����F8H��1g]�EKg��(LO�x����L��V-��2�:g�|R�'=fi@�@��8�<� �&�<�^8��'��IC�����y{�	C�k����'�(�YBΐ-~�Yc�NJ�d�T���'jD �^&#���� O����'?fA�0���x���?uh����x
� �x1���rc���#&R���h��	I����F�1=��bSMɓa\6�����<�
�T��4�#X�$�0Ĥ� {|ȇȓB($� B\l�>L(GBӘް���.���B��}��M�"� �:͇�|�"8�Ð�L=�ER#qM��I�����*�m��BK�Q=��G�n�<y�B�)#��1�IZ�@��a!�E�	z�ГW�S�EҜ0�b F��(�C�2D�`��,��I��i�tB�S���"q@1D����)��2�}�%��yz:!���0D�be��/����I$fN �kh0D��zPo�
i����2�@�[�,�d#�SܧZ���#�/ȁe�D��s�E,I7���e�'��� CѠo�<P:BCO�x��$���<1
�`T�T-i0�P�Y�t��e�2D��XW덓Q:��@��7~�Z�B	5D����,%k���%�	�z�Npa�3D�$��m˳"�@�!P�m�6H�2�1D�� f[�zpa����l���*.D�|��K�<&�EZ��-	�&�X�)-D�l`�Y6=b���IPK�.��C@*D��*e@�,h��8u�� J4A��)D�T�3G�<�G@|��lXb(D��1U"�8�R�;���FjaKW%D�HHP�O�J����нFONIA��6D�tXЃS�3��5�̎;���S5	3��b���2���>O���en!'?$��@/D���I��lDr����JD��p	e�?D�XZ��S���D���[4�~����<D��J#���\1��t��4w���db>D��tb�zaD,�4��24���) D�`BR�Of@�@fˊr��(D�8[��oR�yT��'*��aG��O�˓�� �'F
t�����@��Z��yՋ_�<�5̀�N?r���˳x���5 �D�<1q�/x�6Y+�h0|����-vyR�'Z�� �ϑ*u���kA�2XD���'|UJ˝�Vђ��al� 5�L p�'c�	i��V9w�Nj�B#`���'�p� #Fܡa�:�PR�ݾYP$I�(Op�=E�T�N6:������E[��1�y����t@"��@}�h��h�"�y�M�0X(��Ve T�i�����y�&C�	!4�b7̱7 ځ����0�y�!� P�zD�yʆD���C��y�� ��vՉ�I s�4��`�&�yBmR�hl���%h{H�a���yrϝ>+A��V(����!��,�ylH�ݼ,RT'�6A��A��*��x"瓺5����
��q |[���a�!򤌶%nv�a5I�9N������%z-!�$ɃR��!	�@Ď(�Y�1�"#!�I34���j\�D��b�Ԃ!�$ήjNxa��q�l��*0 ��}2������YB���F@�A�@�"02D�8��+Ia�������[��a�1D���uK�,'�i���P�%� )!c�OC�I<+2�R��J9J�� X�6�4C�	1y��$�B r�������w��C��.�����T�Vǖ��" �4��C��%v���)��$bĈR��;цC�I)�Nh0�E-l�,���E�6C�	5W��� e	b��8���&x}$�=��g�? H�0���JI�%
s��5d��[q"O(�w��KD���w��W^4�f"O��Bc�s�RTyХ6r@��9t"O��b���.e8c�!BRp+�"Oʌ�H+4U��C[d�ib�"ONTYѠK�?��*�C˿A���"O�ȁ���	PeBq����\��h����OJ��i��ͩD`�jV:D���}�s�Ʋ5h���"J3]i����|�	sV/��Q*j(q�S�Zl)�ȓ0|L�15�� �@�kڳ=6����X�hպ2�C&v1PW1\�m�ȓ1�F���<;��iVɞ,y�z�ȓ5���u*F)sfx � П~�f1��O�n���@\��i7Z�ȡ�ȓM��!j�:R�^�N�Au�B�	m\��@�� d��^B�	#T�~(h��J�p��-A�O$D�XB�	_��9Q� ��)0򌎔hF B��=Q��4$N�^k�a��ћp<B�	�p�
�KT��\}��ԚCU�C�#Xa2iۢ�#�%+�g0Z{�C�ɂ�Ȱ�d/H�аR���*~C䉜2_����a��J�dPQN��(�@C��$
��4@b�	"=�B5��..�PB�		��}jե�9PIX=2�nҀ/�vB�I51|���3�ـ^�.�Z1IP$-�@B�I+�4��CK!?��ÔM�>!"B�	2H�p��ٗZ6! �h�#1 B��&0K����O�-[�%A�+ՎZ�C�	F*R���O��F���R+N�"˼C�	�R�����ڏp`j�cTg��#��C�ɐHS�e���B�sF�l{��-'�C�	�;�Ju��ʎ�vkusF 'a�C�	�V� �	©K`�m��Zz�B�I<O��f$�J�t�g��.x�C�ɵsJF����~�����Q��C�Iz� �eh�NI�kC�C�	������my
���l[4f��C�Io�8�ɓ����V$U%7n�C��6y�yX D
�b�\�&�ؓ��C�%v��鱃H*r=�\z�(R�?�dC�2�]9��ݬq�&���$r�`C䉔*h2=I��E�� \��Z�L �C�	�|9�(ۗd��pŪR�AC*C䉴sk�U0S.ڔM�f���fQ}� C�I>W�^��3oUB�����B�3H��q��@u(0N �AB��C�pp�n��"x$iu�>_��C�t< ���OV!c�["lnC�	>[� � �܄S�bh3s�WY�HC�	�}� }�S�[�a�}C�	1c�^�r��ŀyX��ec��b�C�	�R=����]n�H�J��Q,�C�ɢW~�ɋ@
���ܡ�dH:3fC�ɭJ�&�"��M�]>�6Ǌ�P)���ȓą�y�l�paE_}�y`��i�<R�� �N·f�����B�m�<��)G[��)�I�P�؈q���b�<i6���1�mB��(R�X�AIJ�<�ʋ� �X)7c@+ K�H�T��Py��)�'=#����!��Ru蔊�A_<?N���@WP`B��C�0-S�\U�NC�I�u��i���4!h�;����ʓ�0?� ~!��(�%^6| p�I�Q��pBf"OfMy%�ȼ>�t�S��0��z"O��:Á��z�V�i��[�S�v�R"OȉZ%��%'���GMC=�p�Ȳ"Oh9Ica($Z4��C,�Lu6��G"O��T��
��1����!}�}`"Ol��U���r4�,�4̇
M|��D^�(��Ie���c�&Ƭf�ha�L�7��B�%j�C��2�F�F�1�B�I>P  �����).��<6�C�I=P������}/DHi�G��C䉣[ 8I���ٻUq0��i�KN$B��5XE�3��L@�2��s<C�ɃH�F�R�0C��Ea�Ҏ]=��3��s�*��j~V�b[;�h�c0D�xr�(OV���Ё��>�����9D�#��߱-�DŨ�-X�(	�F�+D��(��6s!��,<F:4��.*D�8�Sn��{@��'����[��(D�Lаm)`
�(�sH�<@��*6L*D��f�CL���36�R�j2�k��(D��+f��*V��VfO#�՘�$D��$�({|���fA�q��9���=D�`K���2�@@�HK�����"(<D�����sPb�܍p�l��5L4D�D8&G˸T2Q����di�W�3��������pe	6n&�! ���H�P�p�"O:jFD�5��('`������e"O�|y�NKs �Բ���p(2a"Ol�QG# ��ya�mR2y��	�B"O�X�I�Z���cW���v����d"O�r��˕�lb#)�8~��@�c"OPD�Ƀ$P$��N�O�}q�g�� c���=pU�(��4D�$��%��g �b >=j�J D���� $oH��i�'�\�
	r�!"D�<��/��� "�
?�� b3$D���횄CN$,s�JV�;��-D���1�� tt�����/&df�9D� �s#�<k��a����Y�8k1��O�=E���X)b���1nP�r��U�C�͚P�!�d;��	�#}�x�1H��!�dA=8��i�YZS��&�0"�!򤏷��L�g ��4�+���!�$ټ3���E!�5<�D0 A�!���>3�aH�	��>rB��2@�!򄌐4v��;���]���Ѡ֗o�!�dɏS�� �E9MW�	)��ć_�!�Č�-��E��L	�wT���#@�c�!�d\�f�u�#%F7P� Ȑ'_�u!�d\�Ojz��S�=oS����Gd!�Y�3��Lh�"��y>�q1a�ǼUm!��D� 
��72Lr��FN��!�L)}KRdp4�߻4,��3&�9�!�$�F-P5r�LV<{�y6��Y�!�Dһ �@��Q�}d�,[񉄼t�!�X�Ggv�	Q���z���G�X0u!�M,\34�µ:���# �COO!�dJ1
F�)�c.V/�f�A#��B9!�D��m�����M�8Ϣ	�G��3T!�$\�o��C�@ue�]"���,K��IV�����d�4eV.�����La��P�bN=%�!��)�d9�g»4h����]-:i!��D�s�RE�M��h�<��j�lg!�� ,��d�Rv�PGN?N�P��"O>uQ�N�5M~�˒˛�g�(��"O �2��&\�$�Q
W)Z�d�c�d>�"���- ,�X�s�R�
�j���=�O<�|��ݻ#F��=0���J&0u�ɖ'�R�D4�OH�u�� b")�`�$ޒ��ȓi`H��	jٛ�ۖJ�d��M�����ϩe��ICJ�G	 <��&�P	��G��q���U�fP�ȓf�l��k�^��{��U9QT(�ȓn�� ����IelţHG�D��i����<�2w&�<�IV6�Y৊����'ў�>��qb��l\X#��^Y,���*D��"(�)� �ITK�E@	�F&D��T��{�&��-'N�$�c�A&D������a�
{�`�6�#D�x�RA�����:3K*BffMJ�#D���B�p+d�@��J�8E(�� 4���#I't�F�b���;�|H���TA��hO�'M��$u�M��jY)Cm}N�,�ȓ#����U M�)<�F$3Q ��ȓo����YMA�O���؄ȓ90\j� ��Q-N���N�)4�N��ȓ\�z�!�-T?HCf�E�@�*<��@�N��Fäs��g��#C��ȗ'��y��� ʄ>�"��֋�4O���ڧ�8ړ�0|*!�J�)�j)���R�D�1�Wj�<��F��[_d\q �Ъ;���s ah�<1eLQ+7 �W�=y褩�j�y�<�"��!po1ր KB��F��a���^�YT�ˠi�XYB�N�3j�D��m�Z���nԙ��T����u�nG{����O��  �N��A
H @,������㟌'���'��	�P<LY@c)F3(���,�h�C�	[�.�H竓f�3�	ӂ֒C䉸�V)���BQ��B�N�qՈC䉬�f�� |�X!��N�U�&B�I$*�P4a��6K�� v����B�ɷ�V�	v�T�;2|<�V �1O����d-?��퉿ZFS�%C�6�@.CP��x̓V0�1N�%�̱0��O;���ȓmL\�V.Â/:�d0�ȝ[L�ȅ�W:BxAN�3g�z��'( �&�ȓLtđ�tÈ n1���f�-zJ@���R8��k_%����pe �����J�p|Z��7L��KP�N(����p�:� S� U���/��o+Έ��Iq�	�<9%��/8plh劜 \�`DjQa����<���0�XX� �\2n\޴��Z\�<q3,4�d�����&2����
[X�<�1"'ju�%�Te�o¶�{�bAS�<��o��'�a)',Wޔ��6CMO�<io[Y�xI���<2��|�'�q�<9�AHR��ك.�Ժ&2|Oc�$ �Λ%N�v���(B�:��<D�����>b��˵,I5ڬi��/D���r�H�g���k3��'��\��)D�dcr��"t�j����!c�X��
'D��B��;�B��� Oc����O6�=E���9-FM0ŉ�WP��H1!�$��-�0�dDA�R>���J�:!�DΈ^��5k�b
��i!�V!��F��8:�j��n��Ȁ@Ȓ2�!�d�:�����SV �do7�!�� J�ɖ�?s��4�f
0K��{�"O�u��f�$A�Z$�Q�G{0b�H��'��$�,�^�� �5� ��*M!�'!� h��/J��$��?e@�{2��(qKt��l:G�:�$�k��O�QG.�?}�B)  ς&鋇�y��X�4!�t!���RQ���y�C�Ρ�ψ� of�Ч(_�y�/���B��Ǹ�T9Р�6���0>�Q�X#MͰ-�MF��#Xq�<A�D�
�褓��ԿX*�8ʂF�Eh<�a�����4���-��NJ>�?��'����!��	*$��P
�ZZ�'���I�C�?�f�s4�D�ʙ��'�d���O����sу*᮰��'c�h���ݘ ��Pm�'tD袅f�
�@��@*��\���'��,{Wd�	K�Ɓ;�1]�ΌI
�'������d��){���
R�f=)
�'p����הs	(����6+&D�	�'4lP��_��Z���ʛ4�h���'��]�`��>}��Ua�
�'J*d��'�$�YS�Io�9р��$�vy�'��a�ւ_)/�r�����]Zl��' � ���DA���W.�t��'�R!*�;(�ܐ�s��E�(!�'J��1�@��IX�"��-�P*�'|)�A�ѻ&y�tA���!*^u��'1BE�3D�8G��daR4sމ �'��S� B��e"תL��l�i�'�x���1*��iF��pY!�'qv�ߖ8On�ϛ�����'� 2�Ì/b�X��,J�h	�'����lI�.BDE �Nmp�'�8��d�96^h�O�dH}�'��\i�Yv[����G��[�
aS�'��+S�B���y�b��L����'�����;)�>���FAڤ$�'1^MsI�}TB�� �
9�P]
�'J�kV얀-
�� �Gٞ<�����'�� ���~�����,,b*,��'�-�U��H������\*V����'�����_b���a����X�Q[	�'_|����,/IF�i����HT	��'��#+��~#����c�/D�<��'��uiQ,'V�"�Q`�I�D�v�'���#Ц�t-rm`�Րjtb�z�'R������$C��0BgJ�0*&���'��j$��hw��HVB�,�b�;�'���p�"t�.�A��KVz���'|�ݘp���!sU���;�b` �'�Ԥ� ڮ-�^5�Л2J���'�" P�E�H�����+H�X�
�'��D;�J�a�I[sl��!��C�'۞h�cNW�vQ�D�£F9m�,Vh�<�t���z���)� s0��w�<�*H�@-�y�p��1��DjČv�<yV݁T������%ʽ٥
�m�<Q��*@��}bبs^ͨЈu�<���� ��Q��k�Lc��v�<�#�>A8�����U)�0s���\�<AV*1A�`��!�S9wn��a�S�<�i�L:~�8ס��e�&=ǈO�<A�	�=@ �c�N�8x��KG�<� �d��<#��Ћ�KC\ft��"O"���aܛ)"�$B���3S,(�1"O2���a?��T����T&�ԩ3"O�#�G�<ٲX��	�Wop��"O@�&铞Z��4;C�{1l�K"OD�N�D�ΥHt�Ӑ0=&�	3"O�Q*�Q�I���yA�^^d��"OV�j%c]�M��<q�&�
u"O袵 �'���Q�ڞn��"O�5{1�P�m���r3�ެp���T"O�d��M/�Z�Bs���M��#A"O!y�E6E�`Q�R�M$Q�Q��"Or���lH2<�)� �{ކ2!�d��4�X5�L1IӖ����!�^�\��ŖW(:�¦�.[]!��˦u� @����0�Q6E��h6!�$�3(�#g�X:�$Y� �S�{�!�;�=8`�P���T�ŋ?�!�d�[�~d �f�� !��'!�$ܽHv�,;h�>���˔��!�%�f��c�.]��|�s	��!�$��8J�P1�m��M��H�!�D�$Y�oa����0l�(�!�,d������ܤ��kճf�!�$P)Mb`�2GjSfU� ���Z�!��I�����BaԜh"e��,r9!�d@�^���k  Y�"�Z k�.�Py���
qH��pb��.ܖ�tϟ��y2�S,;�F��-J7�H<��!@,�yȳ[;�=1A(ap$+�A���y��Ѝt,tx#JńA�nȚ$`���y"��l1ށ�!�M�D�#�F�y2 E%,����G�.yR�ҹ�y"��	̜�3PaS$G��"ULW�y"�� �n���ڶ�ȵ�$ȓ6�yr%�]׀��P�~1pY���k��'܌ ��T7:⌹'��l��'G�a�'�'��#��ie�l#	�'ʈDid�[l����-�)a��u��'R����U)4<:� GÑ�Mظ�@�'�J1�c�wr��7K׮|[�]��'OH�(�gZ%<�m�F�Иe���
�')��2#.�8OϤ-QE��G�`1�'HT��D�\�ذ��3/gH��	�'��� q7�|Т�y��@:
�'�}IWl��J �D�a�|��y�	�'���EȄ9j���^p�!G�+�y��e���8�bǚ@*�:C#'�y2��%P��%��d2����F��yƆs� ��h�)��J��y���!)���0�˨'��a�%��y"��4��蠎T� w�$�W��yA�)}��!EX�'��Z��*�y�H�	��,�u(Z�|T�+��y""ÿT,RE���D�~�:�͍�y�ʒ*d:�aq�[�p�,����y���W�L��A���f�8���4�y���:3�h5��h��kuD�{�!��y�aη=l��pMܵ[U<b"�Ύ�yҁNTP>��D��+j��e0���y2B@"M�,��K��X��B2�\�yb'܁'�8�N��N|9�cN��y(����ۤi̽��QQGو�y���2|YRA�:'�Dh��7�y
� $�����'f���ǨT�T�c�"OPP�q�^2U��g�(X�$yAa"O���/a>�sEl�1�&ѻ"Ot܋F��d���0��  :HY��"OX�y�O}s�{p�Q�7Z"ȓ�"D�8��qK����0����h D��3`��=i޸��&<�����-,D�T�'�,���d�s�$��i7D�+7�Z�7��E��gŊ"��`*�4D�Љ���*b��1�s�O}z���#1D��#�B�in4���G�.&�x���,D���!����()9� L���8��4D�"���0U�D"U����h	0�&1D���W�8�x�1F�-���!#D��z
V:��ɖ%�4Xp�!D��3@�X+Q#F�	G��?��Ш�(4D��q���T(8TI�%�5��l��1D�1A��)��K��rp8c
:D����ǰ$Z�U���\_�b����"D��B'N�u�tY��L�Wdut�3D�P�� \
:��-�m�)��$�g�/D�p@�ME��Ҍc�#��)pc�,D� bi����AU����Ń�&0D�(��E�Mè�5k�쉂�#4D�<k��Rgv���Q�f�q;�! D�|�e�ة4���A���9Rx��Y��2D��2�G�?n��A�u�A$�
p`0D���$OƧh�8�d� \ ѱD).D�P�Fl�%� G��(V�aKP�*D���w��Y���4dK�[<9���#D��{p)K	@��/	$f�-Af�"D��p������p���?D�@��_!�Z�CI��Z���7�(D�x�4!�PYH���H7�LJA�%D�ȘċP!][`4��e�*�|��!.D��¥���m�&�s4��
/0>���+D�|��Θ����<t~�Q�gl(D��8�@��"�(T���"��9C�$D�̋�(��}!�X� U�^�����"D�8*��!u��Y�w�����s�,D�ذ��Q
q���È�$uo�x���(D���g-��;t�8�0�؅k�z�dM'D�`�J�a�����!0H�&��R'(D��慘Db9O��sϺ H&'D�p�≈�E�Н��B��ZÎ<Q�@&D���'�jϖmSb$��]'�%D��Ks��T �Q��L3ADd�4�9D��hU���Q�lx�EfJ�B3`�6D�@�B�h����H�����*D�x+���1b(Ї�G�wT�Bw�;D�� �\"�@Л���'`��J`�5D����)�yjHZ��&=����H4D��A�K�Z�ቱr枈���'D�P`N�}��eS�G�w�V��QK&D�\r���e�03��V:i!@��#A#D�����ĆV��J�	4'?fHYci+D�Тר ��ꄃ��6О�Ą)D�L�Q�Q�Y�N�;��1O�&��4	&D�L��20j�!��K"3y�a��'D�\:�b�
w�t+��=�)cv(2D�H8C�^�YZ�� �
q��:�#/D��z2O*$��a���"GKL�B!��u&�P��R>kָ��ޚq�!�X�f����jH�}cĀ:�钼ja!�� �*��*U��E���U^��K�"O���B�� "p`q�dC�[I���C"O��ؕ	��t�z�@��.G�J�"O��q3k7`v��YPI��B�6PR�"O �i�.͆�45�TFV#�X8""O2��r�ɲ��S [�Mn��2"O��� ��(#�����Vc��"O�ä��&1���	����jZĩ�@"O����*�J��lQ�P&]�R��D"O���VU%!�`s�k�)�53�"O�<�ˇ�[^�����"y� w"O�T�p���AL!�׋ l�̠t"O�t���f���D�H#-gDHj"O����͊@Rt=it��KJ��#P"O��T�X�|�l8*Ё���Qj"O����HO�)��==�R���"O:I� �_oB -K�I��9"O����лL��[ψz
����"O���#j��$�C�H�������"O\�c׃6�@��({�����"O.� �ؒx8�Q�ץ����#"OD(�u �+p̬
�.\&�h��R"O
��။b���.���"O�(�ֈT*����2�=9a"O����F�`,�dae�(pY�"O� �'�c���8"��zIz"OبQ�'�;0V��cW�в�"Ox x�$��D.�S!�#@���A"O
Q���_�.͖|�Bţ2
�@ؑ"O$�#i�RE�5��%]<(��"Oڨ����s@6 �۲a?2��"Op4��섂g�>=B m�(���"Op�t	k�}�#ɅLJ&�"O�-:dF�M�:��G�l�����"O�͸���-�H��u���f��5"O��)EE�)���K�L@�}���a"O����'z1h��Ui�D��"O>��G/��P��bG�U*���"O*}3��<��\;���:P�vY�"O���bʇ�N��s���C.�#7"O0	k�)�m�X�&�D�b��1"OR͉������H���/b�Y�R"O����O:���;�d�B&�9��"OҸi�䘹qV�e��"
�`�r`{�"OjLc�!�r�αC�'w�HE�2"Od ��ٻ$��� �"*j��"O�ƨ�X����v.0
�B���"O�iCtAܡ�pنL392a�"O:y  ��B��M���?/T��T"O��E�ׯ<Ԝ!��"~�4�"O00"+O0l�d�sD�R�x��0�F"Od�K _�a��Qg��P}���"O�@�7 Ai�X�q$F��KI���"O�-�Qk%��u���9}T�E"�"O~�v/ϲo*p-���śO���"O����ũ0�t),��>�DIc"O8��d��oTMjRᅕeq����"OX�:vƏ�;s����l
�@�s"O�p�ۣ6��0p��Lb���1"Or}�d�Q8Y�h�)H��j�j"O@�K!�ܱ�H>#�`Q��"OX8����fE��T
'�PH�"OU'):mΝ�@'.LȀ#�"O�80��S8y�a���1=�� �"O� ��Y�D�}"��#OF.oo�ib�"O0l�'�d�u+2�M)~(�s�"O���0b[�����W���#"Oܽ����*R�fu	p�#�0���"O�p[�j8b(Œ���.���C"O��cvm��ڐ�S�T�_���!�"O��,�yZ��!D�Z��&Y�YE!�ċ�"	�5�7j˟q�X���D�NF!�$+E�4��b?���L�Z!�D޳5�� C�cU5@%Xq
�E	�g�!�@&V�<r Ο=-$^d��-R�!��>�2���Q������� �!�.�� y֦��!��[f
!M�!�d�T�՘��8%پ������!�Ƃp�6��P��s^�œS&""�!���hq�W�U�fE�`�P+�[B!򤖂L"a@u�$DZ�B�L�t�!�K�1{�(���"p6>�Flp!�[�f�z(b�-F��j˓6�!�W��Q�炌+&G��z�O�5g�!�֨�<xJS�!<�QX��J�Pz!�R%8��IPfN(BL���QeP+T!�$�_����G휛47���!�[ejT���L��)З&\!��ܷCL09xt�A�zQ$�����A�!�D��;�(h�vF؟G3����T�!��O�#Zب:����!��Q�;܊�B׭W�/�d�� ΜO!�d�)H���6���^�T�jD*�X�!�	:'@�Cg��m�Z�`P��s�!�d��	�fų�ݻ�ۢ�I�S?!���p�Ќ���^\2�G%'!�$R�$$��敊/�P�!��=!!�\���7s�&A�
�!��\��Q;���\�V�@�$�!򤗔7#�((R��p�
�M���!�VRSnI���(�v��#zs!򄅈&H�3$Xx���cKX�}h!�� �3?�zuL��2���32��%%S!��N�j�R�������Z�ak!�V� ۘ��G %`����X3�!�dםG�Qsɛ����:C��!��"����L�m�Mj	��'�^Q��GA,�z<c�P�w��)�'|� �sf��dh��d�6p�l\�'����g��y�L�7���o3����'�h �S�J�Nk:L$k����'m|�J歁:��4z�b	=\�VA�
�'W�40q��#��XQ�¿Z�<�	�'e����ۻBΒ����[�KZ��'��3'YՊE��)�0@B<Y�'�p�	A�˔i(��B�72��
�'�;�W�e�0#4��>�$D�
�'��H�R��}�a��@j��'
H�����b��`��_�@�'��8��իU�8@3u`%QnX@�'��9i���~�܄@�X��3	�'���R��L8�����_M��'�>9�я����BMι\Ez���'X��S6N�g��A����T�<@�'kRʍ� �|�Ǡ�a ^li�'gv� �� ܉P��^p]Q�'�����ͤ]َ�y7%��^��4r�'3����nK�Y��[�0P������ �Ƀ&��;�������U��!�"O���qEY7S�2h�wո�X q`"O�Ȓ���#+^8��Ѷ�j���"O���-�=*=���Y+g�<���"O|�bw��<4
4ٸU���"OL��� 13e��*�fOQ�$ x�"O�5*q�� *0�Љu�#���"O4���5�����A
�1�
�9�"Oz��,[.[�<!��A4Y[NѨ"O:�A,�L5(w��^>�Y�""O����5,�*|h�+Iİ=�@"O��KՇ�a*ڹ��ᇷ0X��8�"O�[����w|RѺ�Ƃ�cQ����"ON`j@-�.O7:Hs���	� YB"O��1�%��.���ʁR�J�#"O�YTc�)���!Iߝr�l ��"O.0��nH�&[8(���:xtm	t"O���a�fv|5a��̪y6=:b"Ole��3%q��s��a>�a�"O: ��i�,�}Q%��)]�*�a�"O����N��/K޵�6aV�~�Dy�"O��b��
�#ľ=;��_+�0 ��"O*Y�s��[E���2���9c��9c"O�}��^�v�Եz2�_u��"O�����T�n�� �$Y4qH"O��i�gX��A�T T5y1��u"O|5�RnG%I�� � -�� "O�@JA��$H��H����Z+�բ0"O:<cC�P%-^m#� ��_j�jV"O��P �77��|Am��u����"OJ�	'U�E~hYU��(4�d4bb"O2��1ƈ}�p̸BH��.��#"O����䁡!�.�2r�[>ƀ�R�"O�$#rD�
l�Hmh@k�7��`"OBcVCH5]��8���U�J��i�"O��г�6�z���fyN8a�"O$����D!a�.�[�茋'���p�"Oji�um��O�@�AA����y�g��H,rH �ݣM�-��͠�'7&=�f�_60���eEd�
A��'�Xl)5��O ԍ�s�èh�|�
�'$�d(��Gi�X��
�a6�Ѫ
�'�0"��Kw�D���X�-��	��'?:=��AD�^�r�K��dI��'#��~�r���ԓ]~d#�'FhB�G'CU���`��+ �
�'tLH� ��Y�6 �	͌`j
�'D��H1�I�g��2Æ�T���'����ϙ5�����Y�K�����'�jܺ��!��L�B��Z��p�'FZ���#OlFHZ�H
F�����'l$�A�i��x����Ky��:�yr�D'§>" ��Cۉ�ūg�\����ȓm�la�gJL$xU�"h\9t����Ik��X�[g���	��M�6F��!��E��$5��̾8�ֹx�HO�1�����Ɋ ��#a#�LD�\��/?�C�I,�Ĵ���t��X�0��Y*�4�Ɠ��ɳh��Nkr���j>Q^EEz"�~�2#��I�`p΃? $ҩ��C�ȟ@���LJ=:f��pݣՇC���%��F{���G��RW�X�c
��M "�֖�y⃃5E� E!p��;h�<�J�唼�yB� v���!$%cq�0��-���x"� �d+��U���WK-?��i""O6�[���2�<����F8���'�qO07M�U�������}B�Ǳp!�ė�y�q��A"H�Rt���U�D���p<�TG�}J�`��I*i$^�bGO�<�Ul������F������ͦ��\��T�C�9Lb:|�#�Z{�Ι��B$(aS��y�J6Č3$����O�����WaFX8m���.P(��I�y��I5Y�`���Ŏ|,L>���,D�hE���2�F	kwS%I��  *?I-O�=�O"�}f�!bvbL��	,,6պ	�'wz��NK*r��-�ˌ* �Ε��)��<A�.�� ��e�h�T�`�J�Rh<�S�zv���̐A�
ۀM��yb�֟r*䃔�� ?Y>a�U,�yB[�[lČjwi&nrlō�y���'�4TQ$(ԃc��9s'�ԏ�y�$7mʂ���
.n���6��y��$Za!1$�aȾ��i��y�ו��,*v��Dx�xhV��+�y��ߝ+������O���ڐ뀵�y��)�"EjY���XBY>���E|����nL]�����?��Q2�iO�L(���J�҃@�=���@�"�h��q�ȓ@#͓7Aչ$<0Р�	�8��gs�՛3�3yފ5�7��L8�\��� �#�	�|�xu !)ƀ/Z`p��Ӫ�֮ip���M[�;C�`��"O���� �����3$X�e"O�#$H����$���L��ԉ�"OT�8�A�^���)c���bź��Q"O*)r�O�@ň!c� b��bG�'ZqO�`��"�&Z\S#E19�c "O,�i���o�R��E<�(��'e�l��h]9hZ�����\�ժ%K2D��x5F�֢�q���[��)��/���O�c�$�S���'[, �Bǥ��eظ��V�9j0��ȓ���t���``8"(�2+`֨Dz�a*�g?�Fۭ=F�Ԁ�Pg r(���M�<I�	��vq�u�bJv����<i�ˌ<_��H6B�r14�����f�'	ў�'<N:��h$ɫņ��S*����#��K��ʞ!�b)[Gl@�s���'~ў֝O�v��ňۑ&6p[fUQ1�ȓ.��Y`*��Ԩzri۹IJ��>Q����d�Z$�P�GN"BѺ �׆'�B�ɳq� %�C�	o�R��4&�(~w*#<QN>Y�BE�,B�L��O�a�8��A��O��=�O{4�'fDT�N��)�T��tp
�'�Ј+��л���ƈ[99�z0���$�O?�	�t���!� r�1�U-N
!�������O�t���� @{I�S�g b"BE@�'{����ß@�Z�V�� �R�N��(j��+D��Bv��X��p:�GN�q�Еs2E���'��	�EFx�OZ5��,�4Z�=1���yNra���$%�S��d�'0yF,2тŬ4����J�3�O��j��	��ZH4A���3.ё�,D��:��S�S�#�Nu`����-]�ȓ
�ZD��Z�ԐV �ڬ��	�EQ�"~BU�y=��aB�H��2�Q?�yb)Q�3R&�R�m��9�L�"aP�!�� �O����v�(�A��00̠�#F�M�R���@�zM���#5����������ް?� H��g�"����a�+��qȵ"O��Ǭ��iq����͕.�n��!"Oޘ��_�д��@�w}<$@F"O�0��@I� ��#�)l����4O�����|��,`W�,K��#P�I�3�|2�x2�)ФS��J��$���I��y����$�1��~��ur-K#��'�2H!�)擓L�:-35IJ�ab���ҧ@<MrB�ɉ^lu���'ߨ!
Ь]�b�`����O�p+��ֆ�&9X�ɟ�� X1d"OL�X�� U�5��ɛ+ ܌ 2"�OD<��I7-���I��4���6��J��u�����O�8I�F��"��d��'�����'3Q��Y�H�/����C��^9�(����	5)0� ��� *t����
 �Tt��d�<Qam��b2�,0k�=?EN�5A G�<Y���ޒ-�@�L%N7�Ie�@B�<QE%(~H�Q@�H�6?�ڕ��Y�<�Td��5d,a�=�$�4�GҦ��>	�����D:��Iu�+�I2!y=!�D@Lhū$lN6�"�C�į!%!�dԴ�Xu�7b�;�Lئ*Zm!�/
��z�ʑ�+R�P�GA*!�R�(��-:1f�h�����ו5�!��a��� �CХmMP��".�!���p�}(rS٢T��� �!���|tA��*��1v�H;����p�!��	 ��7@��_^�phe ĹHo�'4�|�!�VmNࢰ��	W2>��B.��<�J<)�'b%��Px,
��T��(�Ac	�'����H�L�\�ST���S8`ד��'�h!��!�&e"ǤJ,a�^��'n���d]!l�@M�A�-I.��I<ъ��i��*g���0/�i`��� �O1I'!�D�U�8<����'.�бKr��)!�$��v= ��g�E��q�@�_��ay��	n_��R��>g���w
ś!APC�I5Ti�w���+
a7LB�o�B�I�S�@�a�E��@�`��$Za�X�'��*'O9`NW�Y��m,��&K�Q�l�'�ιH�K>O�� �!l��1�
�'�\�0P������ԎfȨ���6�!�َ`�x��� �$��=��ԩQ�ay�����'�V�ꤡ�/�IXV˔l0rE��y��'�&$j�$�31�-1a �#|�p�+N<!��)��-�L<��&��q������3OzLC�ɴb���MK����&	4��B��<16Z�׮� h؋��N�3E�B�ɿ���[cmP6PZ��Z��� �B�Ɏ] N�����LX(�c�3'�C��UA��(W�~hc�5�B�	�_�JQڤDr� ��n�h��B��#~}J���4{�
��&R+~+�B��(�ȃ%S&f��9c'�O�(�B�I�,�)9s�NH����m[�żB�	I8�}`d���2�z �W�/�HC�I:/e1�c�>[ũ&i��&PC䉄0��$��0(��^3�B�I��N���#�?$9LX�
C	 9hB�I�0�r�3�7|� <(''=2B�	�$���0D�_;zoJ��el��B�/_�n�9���;�����؊ ߊB�ILm�}�G�(��Hb ��X�\B�	2p�fx�]T,�[]���C"O� >����0,=(p��o�>D^�P"Op���iL��ܸW�_�gf�\*v"O��{���=3zR�jF/�!nUzLx@"O���!S�H��%��/\�aD�T�"O=��%u!P��ŧ\�^4���"O|��aO@h��LA�C(m�&��"O �3T�Y�G2��D'5��Ȓ"O6�@qK��vs
	fĒ�"Ǧd�W"OR�����Q�QrEDR"v����"O��GEZ?3'Ĩ`$�Y�b��p�"O.4"G@3Pm&A�u���P�<�Q$"O�Hre�iMn岠 \	T��"O����k�t
�I0 �,r��4��"O8y���LwN���`�N=#a"ODaqB ]�D�`aQ�[�e]4w"OLI ��H)�Z2gvL(�"OH�e�9�`y[���%W��"O����N�r-�L�F����Vu��"O�h��ֽ�+��_��(Ƣ���y��"٠�X�"�<5�2A c�,�yfF|�i�o�' �%2�J�>�yrU�Vި]�ǎ�$��D.2�y�%�QQ�����W��r�x�Bž�yB*t�ƅ�	Z� ��e�2K��y�À X�����E�8X2l��%R	�y�����=��KD-9�r�8�y�.�<IQE(�w&( B�5�y��	 9��F!�	m�prëɣ�y��D�_�֡@Wa��\cN3Ջ�2�y��gW��w�-T��L�d���y�!!*��$PP+PTQ�������yR�	�
�AV�H[̵�N�"�y�� ��T�Kw琇HH�m �H��yb�Θ|?���e��'C�b��� ^��y¦ŋ.�F0@��2�[S�ӆ�y�� �/�@h��3Y�>E���yR��+k�nA�կ�*R�n��g��yr�T�1?�ukB��,[��N �yR`�>� ���Yڀ`�B��y�֍�r�9��\[��<�#f@��y���y�d��ᮔ9 ��@�r#2�y�G�1CK> �5�L/���#힙�y��Ȣ	
0���� :�2�	%���y¨]�x�.H�@�<+�A:��[ �y��
�E[��e
x|��O�y�n� K��
p�ٌO>iH�I3�yb�N M�x|���܊rj�$[6n��y�n�9MG�p�FH�h�<HAԤ��y��x)�u�K�ZWt\ca���y�+�/q����V�X�F٨�BD蕷�y����D�T=�4BN�<9R����	��y��2:��hV"�)7�-���^�y�'-T��L�7�F	�^ŀ%V��y��=$w	�JdTU�d�J��yb��L =y�C�f��M$�y�A��Rb؍k��)2L��
ó�y� �YzEŤ��H�dy����y��p�����C&T��Uj��y2�M�<���jRD<�"1+�����yB-�v���`�Z |p�Dʃ�y��=,�xeh˃T���H
�.�y��� ���%j)BZ,=�r�9�y���w��4X7ʕ(?��a��V�6�8�k'+)�$ּ�(��	��`��o�3e��p��ǉ�
��B�)� �QY4Kv�&�I3Ì�P߾P�ʙ�G���IG���p>Q��	"��[pc��E�p�"�E�dx��K �]F�~����<	A��q���b� �0����g�<�6cZb������9zF$�@G�y�I9|V��;j5�]E�$�N:�P("����@���E�yA�8l;<\&��N�'��6A���#�������?�'䦔�3�DAE��y��Z4$����'~�옷d�f��r��0�:�z��
�|GX�Y�)W8,a|�ϖ�P<��z�L��	}���[7��<i��@�q !�&6�y�$��~
��h�.¼������y��M3	�~,�g̓�,`H��m�4��-dD�Cw-D6h�$���I�i��m�����l<�&*a!���s���Fǲg����'b��U���؀mU�Ɉt�BH��O三�	�8�N����E�,*���"Of�ې�C����K�+�Dƾ<��D��!�p>��ȗFز	�Q��
r؀��"PS������7"���'��`As��K{��#�W#%D��d�&@崽Ps�A(�-�#D�̩��L !w�	�Em��a�,phdg>D���eB��H/Fu a5�FL��>D��i!��;m�ɦaۯ�X\�0D�0q7h�=Zg*e%Rd��.D�@A�%)��`���`2l��*/D��)�햎g��(�qAO|I@-ҒJ/D�y��d�"�;��p�.Iiċ,D�ܫ��@V���!���>����B+D��A�,�nL͸��.m��p��?D��a�D��r9i���m'n=s (/D�(h��o�֬�2&�1ug qI,D�tK`"��K�I�7KS�4�	sD7D�0 c���p�aۢ��>t��XB2D�L2Rѥ2�� "CE�i�T�ђ�0�9��F6/���9�1f I0hlт�(-a~2�T�j���H�0m�8	�ث�0<	m���m@�Eɠ��d�&!LM���/�Ц�7*�!�D��_�Z���y�B�K�ΉL��	>a�3��E9 >m����F�d�QG@9������F�0C䉝w�*�T,�#��8���T���)wj��~D�YN�RT���{b�N ^�d�!奂�E�UPAT��?q4�XsZt����x�r�R��Z�|=��'�~r賗m'�O�	�e�X�tU@������	�`n8`��A��C` 0T?)uh ��(x2�@Ә�(P�bm/D���V�.Eu�%ʦnКj*h��l�<)���Gg����BZ0&/��}�v�˴��ad�ۏt��"��'OBD��1��H/��B��|s���E�F)9�'�a��:�'w5��
H�8�iԡ}m���Ug1���eڈ�T+˩���0���0����fݤ()���z�z�zk�y-*hG�J�a��'�׬�(ݪ��A�d�/��O��4�G�����;��:�|�p��D�\�.T�J� �O�U00��%m�f���!V1{X��� 8}�Iíf�������{" �('eXDa#J�)2��e����ͩ1�p�t�֔6vڢ}rs�N*!�H
v�~sz�)PdU���Q%L�Ї�I�K00��H��� �P��D���L�,iT��C�>d�QI�& pY�b�DR�C׼���5�����8�*j���_������"�H�����F�ސ�B��*3d R�.�)I�d,S���/�X��iHй U	5�s���u��7,Ҍ[b�G9\�z��1��z�Ґ�.��p���z��� I'�aX���<\.ibBi��+��E�� p��C'HD$�3����@ǭRNTi����^�V��'�@%e#K�p��O�	ڡK�l��JD�{�&]	dOI��|���b��e�d��C� ���<H��@ S|y�D"5+��'��ٓL���4*W;D���iБj�IЯ���?�3����F���
�dA���ٌqL�٨Tl�p�� �6�c��[a�*q�$�ĭQʒ�Ek=ZQ ���&OH�
�<O2�a��G��<����n��-�G'����aa�NP`�'��u:��\�b&>����T"�@{�L��D��e�"­��:��
f��1�ד':R�Sr��������7����'lL�b�ƪE����O�ӣrkxUc�g�� aa��\'{TuC3ƌ�r����"O����H�|!�X��Ɗ jܼag<��
 hٶ(A����}v.yI�i�4;��`�KX�j���@>:h�Xa䂁=��`!AM�/��� �&��x
��t��C��0	d�u V��yRÞ�/�$����8��Ye��0�y��וT�|`�O�D���(7���y"/[�o����V�8��=���Q��yrDV�&^vI�[+˒�����yBF?�� A��¯|�Be��m�"�y� :]��$;ĬH(>��kB�~rgY!gG���I_� �P�L�(Z$s�
�*]���T%�@���O.!�����E6dm�Un?,Ĩ�Q"OԅhP������按/g�dr���LNh��3� ���H�d-"%�Wf�va�S��;|�Lq�"O���� Q:S�� ʃD¤~zD 
�+�s��b~� �q^ B���`ީ	� �,�>a�6��`����<D���g�ν cHq�G�U0i}�y҇.�O��+�f�$y�V�.O���@T��9S�y�lA�`��H��,K:Ok��X7�T�p=���o2�W�=٘%l�4�^q
_'Q)Ṇd	0\ �W��1�R�ܘP��0Z� #,O�Y����� �NLp��3*T�)%��Y�)����dMK8��ɣ=F�A���٩KߦL���+nZ4��B[(��l�B�?B���Z���҂C=Lm����Eؘ����A,'(�s�0O� q䍙Y����"C<N�'m���]�g����#n�_& �aJG�
��B�I/-��d�!ުK"S�^�'/T��KϦS���0���s�"E/,��Lz5�_(H([�gy��
G�����)�J�H����p=�A�ʽ,��!��ߟ�s��2zP軔�?�ĉ�*�>62���ļN$�C�ܙ3�����ҍusp ɢ&�>d��Z3lA�9fqOp�1���0�d���'��-s ��et�i���8:,�B� k�n�ۧ-R�b1�C���!A���Yƒ��q�t�ZV�@�y��� l	 �8�	W**gsD�agX͆ R�Ic�L���y���R�2�ⳎB�r9T�kG�O>��?�ू�S� %�ݝ7U�p8g��i�Jt��AU|���e��vtl���D&)��]�6W�p(7g� j��	?�f��&mܢTa�yҰ�x@#?I�ƶk���OF��3(}�v3�'#$�!��|�xɧ�1gv$�@�bW\��ǋ�W�'�`PM���Z(��a?}X��'����^��'��% � ^
g2L�/@(ZY�)� ��*h�m�v����
K�}�tE�$�/��?ّ�Ң�*-�D�]݄�;��sy�$�OjQcV/��R�`��tȅ'NC0��a�5d�)b�<��xC�L�^���U�؅���9�'`Y""������*樂;� m!��S���XJ�Iܬg�<�3A��s�61Z1*̤���OY�9��H�<�P�$$�Ȉ	�@�*ky��Y��c�'b\bl��n��',��4�ǃ<�H�S퍤@
��k��0az0���A%9��`Z4����h��$��Pa�eV/]j�1��bS�:��-�t�2s���ӧ��&�#*:9�s.�* ǂDqZ -�����4:uM�T�(HR2)�R<q���Dn\h0 BL�a��Z`�$)C���LK�B�Y��ɏ	��	�>ļ@�Oܶ)P��3 _p����W�2�����i�֠��vXzժ�жE��#�8I�f)����$T��x1X/�����XIr�҉��O����6�`�Xv�� �e`��	�o$��G��rܧHn4�i%lª3����R'��IV� ��A#[����U�'�v�q6fX�� ��غw��� a�<�6L�
b����'w���8�nƠk�в)��z�*,�!@�u��R֡��xBGG]t��"��?����To?�hO,��Q�b�D5���,I�<�+�#|��a�$���ybg��<@�@��e��z裰V��?�#���Z�X���'}��)��n�>u	��ʍ!�Ҵ@fk^*Q�<C�ɐ4	��5��F��s�h���(q��ug�q��ɀ�����EP%%v���>d$��$�	FZ�↊�)�T
q�U/|����5f9�yB�ļ<��3!�!��]ZuÆ$�yn`��E<b��,dcB�Gz�!`�' �A�M�@QZ��O�5%h��'6�����"VP�zG�ע.�,�a�'��p�/��`tDJe�ÿ"�J�J
�'��H)�ӭ��!��⑩�dQ��'�LЁE&u^h�H˯	�I���� ��q�lP'� Ա㠀 /Q�,��"O�,�BňU�5 ���.7���8"O�ȳD#{�]P�aY�����"O:t��iL�L%tp��6d.��b"O��yc��!¤i�䟙l@���5"O4�㇁+h (#b$Y��Ar"O (��N�{<�a��лRED��"O:t��)�"YrP�s)�$9f|Cd"O�A��0d �ԫD�����"O������=�j麵	L�|�)5"O`�pĂX�C�|�g��!.�5��"O�H���z��3�h�Puږ"O �N����Ջ�fb��("O�����Ҟ=���A%�;Pz���"Oꑡ7G�(���#RO��9BLٱ�"O>]��̞!Y��}(��0sf����"O ���Q�|s�5ɥ�ϕnЄ��"O�	��G�/Or�	x3Ν�%�0�4"Oz4�G��������h���"O(�3ˀ�B%���o�4B�Yk�"OJ$Xweǩ��Q��/����@"O�<���ڢ{8��m�4@��@�"O�5� �1��4�j��!�12$"O.���ճi�6m!���%*���"Oj� ��\ARtj��ފ<�����"O�����ΚMXvǛ�K����g"O��!�GUV�x�L��y}F��"O��RW#(_���NڣnNY��"O|����':��hi�cD�m�<(8"OB�[�c��1�ec�ǚL�fIc�"O�5�ro L%�5��d�&OBt	!!"O�P'��!�t��@7F>��"O�m+2��[��eK���8m�a4"O���*�l�(A{%`�4 �Q�F"O�����ƾ?B~� EE;7��m0p"O`��L�4R��} �.��r��Yڑ"O���Z�pM�h����2e�,�A�"O
��%h��K®EKp/O�	��	�"O�1*�	�(t�0��̰4|\��"O��2э��̉s��2 b"OlaH�	:~�@��u��UKly�T"O橊���0o��Y6`P�F>��"On��T�ز0	�D
� ��6 �٠"O�E��B��F)�q�);B���"Op�"~'� +�&A,����W"O"hz�aZ8DI�yB��W�E��`�Q"Ov	Ri� )���wiޑAqV�
"O̝�u�]� ����iە}cx�w"Oδ���>y�J��"�Ό/W0�"p"O����R�7��]���nб�$"O�`�WE��B�в~�{�"O�`V�U�xԈ ꔆC�daXE�"O�-�-̩T���KކF����"O��F|����k��R��`��"Oحzu!C�4��hk�H^�v�-z"O�1�C�a��U�Q|�4�d"O`�s�Y�RL���ry��{�3�y��\�R��U�o]�D#�/ȷ�yB�A;�%�f���Z��)��͛��y�L�dז8�0M��Dy񠘁�y�j��8U�����J"A�H�������y��D�UAC��[  B�y���&V���Ѣ�"D��v-ݴ�ybhY:Ѧp� i��H�5`���y
� �U:�ų����"������"O��§\)J��̉�Ռ(�@0��"OF�Zv��D�DA�3��m�&���)��de�%����<��� �>Ɯd0B K'!d���@]�<���Aj`�����A�,��פ��i����@F�{)���D�uC�����-4f"��ĄĮXi�yҊX,7a,��D��Yh��Pd2��¥�����"�5<!�@�a�py#c�H�2 �>�'
�P��@ <y0��J���0��6��A�r���^C�I2�`P�I��l-k�a�t�*N@���ʓ<S�eʌ�L����oͨ|�A���.Ȝ`*4��q7g�^��0���w�f��I�ut�񓕌J����ɱ�R�p�ղSRԕ��:�v��D�3PX̥c )W��r�I�i
��z�*�)���1���
t<C�	$���fk@�GD"�'K� �ԓO&�����a"qL!�'R�b���a++Z<��%�s�1�ȓb_(`��d�G��8�Q 8
��e§M���'�D��>�f��)	�x��
�bJ1����S�<�`P����B :H�(�^��cpI��b<��$0O��	�*]�����o��z`�z׼:�:�s_��*t͑�:�e"T�[>��Y���1D��w���bd�=s�)�49���b-D��A7I 	:��]p���5�-ڱ�(D��#ǋ٪I�
d��H�@��s�3T�h�W�5(D��)���?�m+"O̼��o�� IJa�\+QZP�s"O ���$�=)#��R��/���"Op%I�Iʛ\�tTD�6
n��S"O���@��0�����a��]��R�"OlD��a�9�H��n �9=Ds"O��@bb�oV�@u��*^p%��"O���A�KU��-9�J��qLTLh�"On�P����3�R���"OX}�R�G	 �H����o�R�z�"O�- ������c�z=©;�"ON����
P�Vl�vጘ@6��
O���2�ZH�X&�x���Ԧ
�
�(���Ğ�0?ٱG�;U��� �<5�>`��dM^��r��ԅ
���A^yB��;�����/s4��j��y"��+pm"4,h��b6��DKe�'��a�k-y�1q��Y�OE]S���;�� $=w�:u�
�'/��v��,}����.5bl��#E	u0��C�'}�m�#�#�ϸ'6&$�������҈-Md=��x3(�"��� ����X.�~�)�B^�i�	,���L��t0Ҥ֊O����eKH<5�G�a��_' 1SwC�.$��`�O�>���C̆Jji�`�I�C���`�'V����Ҏ>n�ӧ+�p��-O���M�8��%
��h���� M��+�7���k��׃SOhTz�f�F<���i�N܊�
��,r���� $!*Y���Ot��Lܖ	��4o#dQc�� W�ɘuVb���K�Fč� Z0Z���dLwPl�[E��-��9�&a�BG�D��@;V ���)��o���ʤ��	>fڱ��!�,M)�2��R� Z�p��ɰ6�Ě�*�m� `I(�(���b�D�vab&eI�\�4�� �j�ʓQ�0A u�:�����5Z�!�N�R���T)��e��ɻK`Px�.�$~���F�*T�0V�<��JD�>�%����~����ɐ}�N܇���KPpe�S������Ë�;}�ͪL�,1���p�*!�UI�.z�%H� �1b��S �_�(�2m�BJG]�Tts��Qr��,{p�^�0iB��!A��\rD%���H&K���z����UU}q�x�Իimʬ��"�s�x1F.�S\嫵D �#�
-�0��-7�y���U���bŋ
2��q��k�;��_�v,R6��'=Z�{�-�~-��>���1��8 E�g*�0<%�tP�J�<�D%�^���-}�O���Pc̩l{� A� /�z��r��T1�ܑu�5��:��7�O^�������i�Ȑ]R�p��FUz�$Ѡ2���d�(p��,H�"�4"�	��H����W���h�f�$���c�Ȁp�����NT��� �9'o�mP��d(�w&��네�u�j=��A�+M��e`w2O�iW�WA��<�F�[?֘t���
!�>��C��N�'� @#r��$/*�'>q���	0;M��v��g���#���A��1(�V(דh6A{�(�u�&I�O]45(��'E�q�T��=v�Ф�O�:inV�#�@mӺ˖띘h���H�B�f��m�q"O�[����`@�`8ӆ�1�D�B�j,����;My�5%� ~[�L����8����=�HyC��I�&Q�I	s�^�{V���x�^$h��६��B��)a,ٛ�y�R�cDV9ٔ�W	��������y�CG(e��h0���v�@K� �yd� )Y��NH�{�@B D�y�@�w!0����՟B�2B �y�)!D�`�L� j����nY��y��/[3P-Ja�"Ow��[#�ǈ�~�*�
�}��I�O��p�q���IY2'V�q�����!:�Ș�f��OR��4�T:�SLޔ�V���"O֤��Y�p�s�kÃ�������Q>s���q��3�H��e��I�	���kc��1M�P�R@"O���й\FLй�kP�ٞH�� 	+��D�]~�!�g}"�$5ض ��#���
ݶ�y"մE�.����J���f�Ew�REs���������/lOv-RA�E(x�La���� ���:F�'CPu�aɰ;����i�VYH&ay�Be([8��J��o�<�+�eH�Y�Vd�=�:��_ܓ�V53�nZ�~9S��i";e�����MLr���	�q�!�d��R��`f`��7��� �ǹH��Pe�p����<)GI#�gy� S㥉N!}��\�@��5s �ȓ(L���#��!^��鐠nC�!�
H��D�:.,����a{��ʚ/��Ȱ��e,H!9�S�p=Q�	WB��\f�D�)'��*#��3�tp�҈ÿk�!򄆔-gT��*W"�EHD�G��qO ,
�C��Y2�d1����>�ٰo��e�<�t��	6�!��D�+v� ��kBA��ybd�<d�D��2g�0��d��>�'�.�	���]�����+��s@���I&�*����Ј`�m�g��9X�hi���?�F!]�Aya}R�C�(G�P���3�R���O�r4h 8`�8�>�Am�#?!�M#5M��]4�	T�1D��+%�����w��/Nˀ��Տ��0��\<h2peJ�>E�D��=x4�
	%%r��+�J�/�y�Ć�~1(��U!Z�w��(����ɴ?�$b�'�9�ax��ҏdwVPYci^E�X"�B���p?A��݁M3�ի
N:�\Xb��z�`���?	��䨓�%.➢}���{�� (�	OPX��Dg�'�R���+�8��d�|�ው�X�ih@&�*&�0hcǄk~��LWI2�q��'��D�#(\J�8c'Խ `s�'�]����>���O�O ��(�?1����׃�%��x�e�����AUKH<AT��t������i\!���WT�dE(ڬO��(�&�� nY��R�'S�אVt�'��.�5�GjӤIa�~")�]DTD�3���䨛�qG ��"�Q:�@����t�9W�>)��� 8�҅)���u��0� ҂Rʹ"?i� *4 H������.M��O5w�d� ���HI剬=��5�C�;4Iay��L�;D~� �H3Ҫ��,���#|N�@��{ʟls�Ō�4O�yC�\0������9C����
���x"�׌!hv��&ت3�aIcCD��hOVе#��������n�)v߀Y�i�)z,��ҏ��y"$�2���p�,\�XA�BD��?)���:�Ѻ�-}���̘+Qn�(8M;�C�I&s�}x6!ފJ�u��7I% ��$���c����<)$���vbe`�7v��ȑ��c���x���S���h���h��/�Zl�4"O�`P��k}�T�f�˼~	�
"OVr@�[��$%`��D�\���"O@�����`�N��'��|��e2�"O� ��a�	��?��l: $�.`;�E:�"O��ID�?�H�ټ  %��"O6DYd#VL��ĺ:�z�0�"OzĈ�� ���Ugj��~8�8�"O��8 )?s��Y�靍Z�0�"O�p�S
¬|�I�d��eWd)�!"O�d��e	$n����
14p��"OX�〨X5[D�Z'_�(�p"O֤�J�,S/T�U0j� �HU"Ob��7�ՠ)O��H��D����g"O�y��#�峂�}���"OzY��Hwo0Hz��6�F���"ONճ�U�C�P�i��)z�b�"O,�j��D5��yx���%�� X"O�����r��M���I�T�e��"O���߭j� PjÞ?���6"O�Xȅ П?h8��#�1�����2D�$��F4@`$�:�
]q)��˦o"D�ā��G�'�:���f_26h)�C�6D�0�fփ���yF��<I�d�{��7D��'ޯG7:4h��N2'Up���7D�P��� D���u`��`�4��4D�̨���
a��iHP�UJ��5D��������i���[�L��5D��P�F�B߾�y�h�$^𺨢0�'D�8BB�U�*�1PJ�M��9�*%D� �f��l.$�9&뇒SZuWo D��"f�K�Qql�8�(�� D�\�$� i�!��� 8��$J1D3D������(
�`Cp�+�l4PgJ2D�p��E�}��]ʰ�.��](��:D�L��B��7����A"g��� =D���j�}>�X�Cޗ\���%D��Q�!!��ܢ|�b� �%D�|B"čE����	�� l��/D��Y���T�f�P�g6�cCb-D�|*!��:'Lժ7�0$Zi�`@6D�|�Ѝ߸����4,/z8(�!D�����`l���m�z^�l��*Oj�T�X�$�� �d�BB(�J���A?�7%9�23�=`��Z�J�"ǆ�G%�$;�J��Y�u��O8"��Ov�q+Tc�!�x
p�˨]��I�tG[7B4d�	 _D��mf���JF�RS�Ǘ5x�j�%U�QTt�t4O|xQ�G�!V[P�B e%���{�� �x{<��UCN'l�Tk�R������dst�sy�dE�r��b�� �S~�����ԝ�uh��V�1O֙�eH��ֈ����M}�R�ـdU"ʶ�FG�5��"˴�
V�T>Y����}�b�3�� 8���0�fֆU���&�OŁ6F�7�4����p>���	�k�t���ݠ6mJ��PLzӚ8if� y4�Ħ)�~��Ė�8���e�<��P�Ri�cH2}���S��S�$(��0|�5ŕ>_�r�B��Ԏ+�\E�r`�,_R^���	'?��ŀ��0|
�L��0(��ލF���:`�� ȶ��.9�e��%����A�EaZ��)�	g3a;!�U3����ZQb�x&#Q6�y"� ����Oi��A'��v�%���5���'�2�C�'͸�3@��v�^R�`�Wc�]�'!>I�W��p�
�c��D�fӂ1��'xp���:p�@�;�eUc����'s4���!��3Z�P��/W6-�
�'��ꀮ�-2��;"�9QZ�C
�'y�I�u
�/��(�`��}_�@0
�'�b��f2��#�-KnHJ��	�'��1b���-���kE��btȌ9	�'Vhl��W�	��XC�O�9Z$NmX	�'0�����2gr�mB���V�i	�'�v0P�I�|����Q�BрeR	��� �<;��5Ұ�Y���	+�"O]�$�,Z��r ��=H��	v"O������WR-�uH ~��y�"O�i��@� hU��Z�ƻb��"O��� �Ao0Y!4��<���("O���ģ�<d����v @�h���bS"O�@�Х0Z���C@�
z���5"O�<��Ʉ*�Xӧ��	WRԺ"OPA�>\7�a�e�a�
"O��Iң�;-\����o��k�xCw"ORd�r���4hC�d�4K���W"O�
E���a9z�af	�
L���"O�I�VKS�^X�S���juF 8�"O�ɲ@��9�4!���<3p�8RP"O2sODո�#a@�'XP�i�"O\��cGG� ۠t���~Gr!*B"O�=��A9n�Yю
4;��"On�K�',��X�RmIXu1$"O&5��˞?I�x
�m��c��T"O�)��)H�8��?P� �"O�I�w,Hmz0�L�����@4"O�\07�ƍJҜق���%W���{�"O��Ǝ�H ��IҢ��z�"O8�{��M����(="�II�"O�	��nYW"�8��!`�a5"O�T��C���0Iɨ5�8�q6"O:��5i
�V��ã"�g�
��""O�12'��B�� �	
/x$��"O���1��l@�	F��XB>Ԋ�"O���GbF*<��P�4�',Ј�D"O�=��Iܩv���T ݯ3����"ON0���� @����%��%�Zt��"Ozԫ����Z��E�P�r���x"OXH���@o	��z�C�x���&"O��Kp����HСc8."}��"Od1S�Л[�D�0�&Y�l�0"O����g_�x�P�+��?.�&��"O��B��z_�$Z��$T ��"OR��J�`�t$� %j!�m�A"O��Xp"�2^�|���	��Jf��U"O��X$��F&plPի4e�q�"OBh#eCT?\bP�5k-�R���"ON�"�'m�>���)�/�h�"O -��D
�t\z=S�̏W���r�"O0��E*�f�nlHWF�>ht��f"O@5{p�W��L�V�Z'pTZ�h2"O�:��V*i6N�xw.�>NDP��"O���5)�ᖔY#��*(J��4"O����L	D�P�[4C�H��u�`"O�ٓ )�.J�s֠ܘQ�A2"O[�#��\z(�P�!�?`*�,#"O>��%�
-:bu����r'd�ˑ"O�S�Ɍ�tf�����ڽ }d9�3"O���cN�R�]h�d�~a�u�"O��9��� <
����W��Br"O�e�hY�N t3��.x����"O^�yf�I�
�\�㎃aM�eZ�"O�P��f2L�j�ƁP�|/�ey�"O.\zaD	�<`$�іAM4٫4"O,�C��}"y+�)ѹ56x��6"OzicgE�Y<ʔSA�A�x0��
G"O�=���*/)�w�_�m+��"O�e�ǋ��EH�	ƥ@��t�1"O����" ��H
NVR��"O� 2�R/�3~�f��w��Z<���"O��
��Xk���n(�D�d"O�Tat�B�J��a�!��L,��"Oҍ�l��^�[m�8W^4$� "O�ɣ$��[��]y�,X�[U��I3"O؁$O�3>U��m>�{"OVHТ.H�T���H�I��(b=�c"O�����75�� *�g^{�͈a"OJL;�NRm�n�����\�\�"O6�ӓ@�Ns�MqLP�f@@!�&"O�T�W�]��� 	�jX[0����"OH��1JB�v� �JB�f����$D���(�q�>y�a��/j@ެ: #!D�\5+� l�6$���f}�,Kg� D�`��5�� sG�}���q1�#D�l���Ɖ��Yfi
�`�t�@#D� �WE�S���{dJ-�<q�s$!D� �D�C�D��)K��L5/�&-���1D����ƐN�h5����s����%�<D�����M�p�"�V���)sPI(D��p�D�%�X��5�S�F&�!K6�%D�8Hp�&ZbQ$ͅ/���{é D�K��6>�N���a�Ru���*D����(e��4 T�]΄@��$D��[wI �^H��X4`�2y\l�9 �8D��Z�#� q��}���fiv\r��5D�x�r'����ΗZ�ЬS��2C�'%:����ll\X�m�&ZqC�I�u��(�SeGjL��qA�t�C�I
O1(�ۤ���F(ॊQS��B䉊7bpz%k�Lt-����(ժB�1�X��Q�\Ob���A��B�I��xUk�#&y���sF� )�LB�I�b�P���ߢdG�-k��?z"B�	�=2��#r�ʳ̲1ʅ�N�O�B䉐'6�	��̫OmV�ۤ/�(_�C��.7�����:��pN���C�I�u�v-��m�5^�L�1�2��C�	'!��@���7m���ҡO[��C�I�]�< Ť;B���`�j��B�I�Y�ؐ��a�Yp���ɟ�m��B�I�M2���&YSd0 #GQa �B�Ɉa�$,bd��4*�Ϛ iNC�Ij*p)P��];���Fo�E� C�I0zP౉�ꌺH�$Yy�CE�w��B�I4V��9$	_<\4e�掂&�B�	�{�,��Cb�=�,�a�Y�DC�I�I.����H��`�ћ�.ˎt�zB�)x���@d z�؍k�/�RB�I2�̔
�J�*b�="����B�	<.��Ah���/X%���-b�dB�	�ppc#E sLN��r#�}�4B��V�t��# d�@��	�kB�B�I>Q@�j���s>�50��bT�C�I�#DP���CF�!P�N����C�ɃPp����aĞ��@GV��C�ɐzn6���a�&L�Z���&m~��ē8�Ni��!�6�`dl�6=J!�1,/�Ty���z���rj��B!�0N�h5!CD}ad�D�j��"O�����%jrذ��̓!���X�"O��pCn��Ա*�HP�oh�Y�"O|`P��5R��ɡG�9P�e��"OL�yR͇q�L�[�#ϙ�� ��"O� 8����H�YܪPJ�M���hA!"O��u+�%%�Y�P��y�|�c0"O<�sPiZ��BX#�KJ?�\]9�"O2��6,�m���
��!٦���"O�e��<o��]���D��� ��"OdЈ!�. 솠�qA�?P@�"O�S3��:L2�5'��#��"O��l@p��� άm��]@"O�P��n�CW%Rq�Θ1�z�R "O�(���i��@�֯;�pm
""O�Hj����{@;�N׺$�"Of��)MR��� x�r42t"O�����ݏ	����ڑu��`�D"O=�qM2Q���A=���)�"O�$�L_O�X!r.�����$"O pz���",i�Mѕ��q���۷"Or@2AlV9}����kB�4�,�"O�M!���i<XRK�jl=��"Ol�0D�1;������ԳUpR څ"O0}���� ��C)	~�3�"O�M���, �Ve�����+:X��"O�A��ִr�4��c̔�c�F���"O.P˓C�-��@��r�\J�"O ]CF�)^���jG���n���� "O2�Q2O-7Ѧ@
�IU(uxLD�"O�U� 'H�8T�D �̧8L�0��"O�1�WƗ��L��W6=�JЋ�"O�Qq�ج�X�Θ!�(��"OR���j2V���!d��"O0a:��e�@alí@
��*�"O| �c��F�l�p�
!�Ayu"Op��N�j��*pJS,o���b�"Oܨ;�ßS�@)f� Q߲ �"OPuiфY�F�PR�^�=�.	�F"OJY9�"b�P�o�1p����"O���P���]xte��`B<��L�"O0��e� �(i���	R���۲"O˰F�<Ay�R���C��X"O��ql :e´�����N���3"O��*�M�k,
( e'�� ��؉�"O�ȄON�TU�5BF�R#< 0�"O=�SB�e &u;���+QK"O��aw��	Sh�����b���"OJ}���H�g�T�Z��ެ�"Oh���@ �`��Ş�5���"OTy�OȽ%&�q)�I�#��PJ�"O�E |H�uڕ" `�.��3"O� �d	!1�T����Q6D�R @'"O����+�\,��Q�_��)�#"O�5��ۄso�iPSA�ZHڝ�4"O��RA	ň �O�>P2���"O2�S7�ڈ ��oкxY{�"O�Z�j���D<+�-N��Ȋ"O� ��6<�&��76�l ��"O`���!ǯGʄa�mO�A,x��"O�q싾8w~0�e�O(�+ "O���g��\@�q�eBc���"O�m2    �